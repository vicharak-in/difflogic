module logic_network (    input wire [399:0] x,
    output wire [59:0] y
);
      wire [549:0] layer0_out;
      wire [549:0] layer1_out;
      wire [549:0] layer2_out;
      wire [549:0] layer3_out;
      wire [549:0] layer4_out;
      wire [549:0] layer5_out;
    assign layer0_out[0] = 1'b1;
    assign layer0_out[1] = ~x[60];
    assign layer0_out[2] = x[394] | x[395];
    assign layer0_out[3] = x[71] | x[72];
    assign layer0_out[4] = x[3] | x[4];
    assign layer0_out[5] = ~(x[261] | x[262]);
    assign layer0_out[6] = x[293] | x[294];
    assign layer0_out[7] = 1'b0;
    assign layer0_out[8] = x[165] | x[166];
    assign layer0_out[9] = ~(x[309] | x[310]);
    assign layer0_out[10] = ~(x[235] | x[236]);
    assign layer0_out[11] = 1'b1;
    assign layer0_out[12] = x[325] | x[326];
    assign layer0_out[13] = ~x[178];
    assign layer0_out[14] = x[145] | x[146];
    assign layer0_out[15] = 1'b1;
    assign layer0_out[16] = x[286] | x[287];
    assign layer0_out[17] = x[73] | x[75];
    assign layer0_out[18] = ~(x[1] | x[3]);
    assign layer0_out[19] = ~x[32];
    assign layer0_out[20] = x[308] | x[309];
    assign layer0_out[21] = x[355];
    assign layer0_out[22] = x[297];
    assign layer0_out[23] = x[289];
    assign layer0_out[24] = 1'b0;
    assign layer0_out[25] = 1'b1;
    assign layer0_out[26] = 1'b0;
    assign layer0_out[27] = x[56];
    assign layer0_out[28] = 1'b0;
    assign layer0_out[29] = 1'b1;
    assign layer0_out[30] = x[23];
    assign layer0_out[31] = 1'b1;
    assign layer0_out[32] = 1'b0;
    assign layer0_out[33] = x[317];
    assign layer0_out[34] = x[344] | x[345];
    assign layer0_out[35] = 1'b0;
    assign layer0_out[36] = x[91] & ~x[89];
    assign layer0_out[37] = ~(x[93] | x[94]);
    assign layer0_out[38] = 1'b0;
    assign layer0_out[39] = x[364] | x[365];
    assign layer0_out[40] = 1'b0;
    assign layer0_out[41] = ~(x[67] & x[68]);
    assign layer0_out[42] = x[175] | x[176];
    assign layer0_out[43] = x[184] | x[185];
    assign layer0_out[44] = x[321] | x[322];
    assign layer0_out[45] = x[171] | x[172];
    assign layer0_out[46] = x[240] & x[241];
    assign layer0_out[47] = x[41] | x[42];
    assign layer0_out[48] = x[245] | x[246];
    assign layer0_out[49] = x[132] | x[133];
    assign layer0_out[50] = 1'b1;
    assign layer0_out[51] = x[241] | x[242];
    assign layer0_out[52] = ~(x[130] | x[132]);
    assign layer0_out[53] = 1'b0;
    assign layer0_out[54] = ~(x[18] | x[20]);
    assign layer0_out[55] = ~(x[350] | x[351]);
    assign layer0_out[56] = 1'b1;
    assign layer0_out[57] = x[327] & x[328];
    assign layer0_out[58] = ~(x[249] | x[250]);
    assign layer0_out[59] = ~x[232];
    assign layer0_out[60] = 1'b1;
    assign layer0_out[61] = 1'b0;
    assign layer0_out[62] = x[98];
    assign layer0_out[63] = x[18] | x[19];
    assign layer0_out[64] = x[31];
    assign layer0_out[65] = x[43] | x[45];
    assign layer0_out[66] = x[147] | x[148];
    assign layer0_out[67] = x[105] | x[107];
    assign layer0_out[68] = ~x[186];
    assign layer0_out[69] = x[150];
    assign layer0_out[70] = x[96] | x[97];
    assign layer0_out[71] = ~(x[85] & x[87]);
    assign layer0_out[72] = ~(x[234] | x[235]);
    assign layer0_out[73] = x[158] | x[159];
    assign layer0_out[74] = 1'b0;
    assign layer0_out[75] = 1'b0;
    assign layer0_out[76] = ~(x[68] & x[70]);
    assign layer0_out[77] = ~(x[303] | x[304]);
    assign layer0_out[78] = ~(x[118] & x[120]);
    assign layer0_out[79] = 1'b0;
    assign layer0_out[80] = ~x[35] | x[34];
    assign layer0_out[81] = ~(x[214] | x[215]);
    assign layer0_out[82] = ~x[86] | x[88];
    assign layer0_out[83] = ~(x[359] & x[360]);
    assign layer0_out[84] = ~(x[218] | x[219]);
    assign layer0_out[85] = 1'b1;
    assign layer0_out[86] = x[83] | x[84];
    assign layer0_out[87] = ~x[106];
    assign layer0_out[88] = x[25];
    assign layer0_out[89] = 1'b1;
    assign layer0_out[90] = ~(x[26] | x[28]);
    assign layer0_out[91] = x[227];
    assign layer0_out[92] = 1'b1;
    assign layer0_out[93] = ~x[352];
    assign layer0_out[94] = x[230] | x[231];
    assign layer0_out[95] = x[36] | x[38];
    assign layer0_out[96] = x[322] | x[323];
    assign layer0_out[97] = x[0] | x[1];
    assign layer0_out[98] = ~x[192];
    assign layer0_out[99] = ~(x[126] | x[127]);
    assign layer0_out[100] = x[73] | x[74];
    assign layer0_out[101] = x[45] & ~x[47];
    assign layer0_out[102] = x[114] | x[116];
    assign layer0_out[103] = x[315] | x[316];
    assign layer0_out[104] = ~(x[154] | x[155]);
    assign layer0_out[105] = x[273] | x[274];
    assign layer0_out[106] = x[24] | x[25];
    assign layer0_out[107] = ~x[114];
    assign layer0_out[108] = ~x[37];
    assign layer0_out[109] = x[336] | x[337];
    assign layer0_out[110] = x[48] & x[50];
    assign layer0_out[111] = x[135] | x[136];
    assign layer0_out[112] = 1'b1;
    assign layer0_out[113] = x[52] | x[53];
    assign layer0_out[114] = ~(x[163] | x[164]);
    assign layer0_out[115] = ~x[263];
    assign layer0_out[116] = x[107] | x[108];
    assign layer0_out[117] = ~(x[224] | x[225]);
    assign layer0_out[118] = x[253];
    assign layer0_out[119] = x[295] | x[296];
    assign layer0_out[120] = ~(x[393] | x[394]);
    assign layer0_out[121] = ~x[4];
    assign layer0_out[122] = ~(x[8] | x[9]);
    assign layer0_out[123] = x[112] | x[114];
    assign layer0_out[124] = ~(x[256] | x[257]);
    assign layer0_out[125] = 1'b0;
    assign layer0_out[126] = x[126] & ~x[128];
    assign layer0_out[127] = x[209] | x[210];
    assign layer0_out[128] = 1'b0;
    assign layer0_out[129] = x[356] & ~x[355];
    assign layer0_out[130] = x[79];
    assign layer0_out[131] = x[119];
    assign layer0_out[132] = 1'b1;
    assign layer0_out[133] = ~(x[118] | x[119]);
    assign layer0_out[134] = ~(x[79] | x[81]);
    assign layer0_out[135] = ~(x[39] | x[41]);
    assign layer0_out[136] = 1'b0;
    assign layer0_out[137] = x[72] & x[74];
    assign layer0_out[138] = x[281];
    assign layer0_out[139] = x[55];
    assign layer0_out[140] = x[75] | x[76];
    assign layer0_out[141] = x[257] | x[258];
    assign layer0_out[142] = x[130];
    assign layer0_out[143] = x[161];
    assign layer0_out[144] = x[33];
    assign layer0_out[145] = x[330] | x[331];
    assign layer0_out[146] = 1'b1;
    assign layer0_out[147] = ~x[194];
    assign layer0_out[148] = ~x[223];
    assign layer0_out[149] = x[49] & x[51];
    assign layer0_out[150] = ~x[62];
    assign layer0_out[151] = x[173] | x[174];
    assign layer0_out[152] = ~(x[208] | x[209]);
    assign layer0_out[153] = x[51];
    assign layer0_out[154] = 1'b0;
    assign layer0_out[155] = x[144];
    assign layer0_out[156] = x[312] & x[313];
    assign layer0_out[157] = 1'b1;
    assign layer0_out[158] = ~x[48];
    assign layer0_out[159] = ~(x[82] | x[84]);
    assign layer0_out[160] = ~x[133];
    assign layer0_out[161] = x[223] | x[224];
    assign layer0_out[162] = 1'b0;
    assign layer0_out[163] = 1'b0;
    assign layer0_out[164] = 1'b0;
    assign layer0_out[165] = ~(x[57] | x[58]);
    assign layer0_out[166] = ~(x[390] | x[391]);
    assign layer0_out[167] = x[139] & x[141];
    assign layer0_out[168] = x[60];
    assign layer0_out[169] = x[1] | x[2];
    assign layer0_out[170] = x[110] | x[111];
    assign layer0_out[171] = x[42] | x[44];
    assign layer0_out[172] = x[38] | x[40];
    assign layer0_out[173] = x[20] & ~x[19];
    assign layer0_out[174] = ~x[21];
    assign layer0_out[175] = x[70];
    assign layer0_out[176] = x[287] | x[288];
    assign layer0_out[177] = ~(x[215] | x[216]);
    assign layer0_out[178] = x[168];
    assign layer0_out[179] = x[76] | x[78];
    assign layer0_out[180] = x[17] & ~x[16];
    assign layer0_out[181] = ~(x[23] | x[24]);
    assign layer0_out[182] = x[290];
    assign layer0_out[183] = ~(x[231] | x[232]);
    assign layer0_out[184] = ~(x[236] | x[237]);
    assign layer0_out[185] = 1'b1;
    assign layer0_out[186] = 1'b1;
    assign layer0_out[187] = ~(x[91] & x[93]);
    assign layer0_out[188] = ~(x[124] | x[126]);
    assign layer0_out[189] = x[141] | x[142];
    assign layer0_out[190] = 1'b0;
    assign layer0_out[191] = ~(x[133] | x[135]);
    assign layer0_out[192] = x[74] | x[76];
    assign layer0_out[193] = 1'b0;
    assign layer0_out[194] = 1'b1;
    assign layer0_out[195] = x[148];
    assign layer0_out[196] = x[190] | x[191];
    assign layer0_out[197] = x[32] | x[33];
    assign layer0_out[198] = x[255] | x[256];
    assign layer0_out[199] = x[25] | x[26];
    assign layer0_out[200] = 1'b0;
    assign layer0_out[201] = 1'b0;
    assign layer0_out[202] = 1'b1;
    assign layer0_out[203] = x[138];
    assign layer0_out[204] = ~(x[212] | x[213]);
    assign layer0_out[205] = x[48] | x[49];
    assign layer0_out[206] = x[193] | x[194];
    assign layer0_out[207] = ~x[30];
    assign layer0_out[208] = ~(x[80] | x[81]);
    assign layer0_out[209] = ~x[328];
    assign layer0_out[210] = x[339] | x[340];
    assign layer0_out[211] = ~(x[104] | x[105]);
    assign layer0_out[212] = 1'b1;
    assign layer0_out[213] = 1'b1;
    assign layer0_out[214] = x[297] | x[298];
    assign layer0_out[215] = 1'b1;
    assign layer0_out[216] = 1'b1;
    assign layer0_out[217] = ~(x[181] | x[182]);
    assign layer0_out[218] = ~(x[5] | x[7]);
    assign layer0_out[219] = x[160] & ~x[161];
    assign layer0_out[220] = 1'b1;
    assign layer0_out[221] = ~x[159];
    assign layer0_out[222] = ~x[380] | x[379];
    assign layer0_out[223] = ~x[323];
    assign layer0_out[224] = x[298] | x[299];
    assign layer0_out[225] = x[31] | x[32];
    assign layer0_out[226] = ~(x[182] | x[183]);
    assign layer0_out[227] = x[111] & x[112];
    assign layer0_out[228] = 1'b0;
    assign layer0_out[229] = ~x[87] | x[89];
    assign layer0_out[230] = x[313] | x[314];
    assign layer0_out[231] = x[125] | x[127];
    assign layer0_out[232] = ~(x[124] | x[125]);
    assign layer0_out[233] = x[227] | x[228];
    assign layer0_out[234] = x[84] | x[86];
    assign layer0_out[235] = ~x[275];
    assign layer0_out[236] = ~(x[81] | x[82]);
    assign layer0_out[237] = ~(x[149] | x[150]);
    assign layer0_out[238] = 1'b1;
    assign layer0_out[239] = ~x[28];
    assign layer0_out[240] = ~x[28] | x[29];
    assign layer0_out[241] = x[228] | x[229];
    assign layer0_out[242] = x[96] | x[98];
    assign layer0_out[243] = ~(x[12] | x[13]);
    assign layer0_out[244] = ~x[273];
    assign layer0_out[245] = x[47] | x[49];
    assign layer0_out[246] = x[382] | x[383];
    assign layer0_out[247] = x[371] | x[372];
    assign layer0_out[248] = x[56] & ~x[55];
    assign layer0_out[249] = ~(x[247] | x[248]);
    assign layer0_out[250] = x[17] | x[19];
    assign layer0_out[251] = x[94] | x[95];
    assign layer0_out[252] = x[225] | x[226];
    assign layer0_out[253] = x[237] | x[238];
    assign layer0_out[254] = ~(x[106] | x[108]);
    assign layer0_out[255] = ~(x[229] | x[230]);
    assign layer0_out[256] = 1'b0;
    assign layer0_out[257] = 1'b1;
    assign layer0_out[258] = ~(x[136] | x[137]);
    assign layer0_out[259] = x[125] | x[126];
    assign layer0_out[260] = x[105] | x[106];
    assign layer0_out[261] = 1'b1;
    assign layer0_out[262] = ~(x[103] | x[105]);
    assign layer0_out[263] = x[112] | x[113];
    assign layer0_out[264] = 1'b0;
    assign layer0_out[265] = ~(x[282] | x[283]);
    assign layer0_out[266] = ~x[357] | x[356];
    assign layer0_out[267] = x[174] & ~x[175];
    assign layer0_out[268] = x[220];
    assign layer0_out[269] = 1'b1;
    assign layer0_out[270] = ~(x[358] | x[359]);
    assign layer0_out[271] = 1'b1;
    assign layer0_out[272] = ~x[63] | x[65];
    assign layer0_out[273] = 1'b1;
    assign layer0_out[274] = 1'b1;
    assign layer0_out[275] = ~x[389];
    assign layer0_out[276] = 1'b0;
    assign layer0_out[277] = x[100];
    assign layer0_out[278] = ~(x[72] & x[73]);
    assign layer0_out[279] = x[46];
    assign layer0_out[280] = 1'b0;
    assign layer0_out[281] = ~x[43];
    assign layer0_out[282] = ~(x[101] | x[102]);
    assign layer0_out[283] = ~(x[134] | x[135]);
    assign layer0_out[284] = ~(x[197] | x[198]);
    assign layer0_out[285] = x[284] & ~x[283];
    assign layer0_out[286] = ~(x[242] | x[243]);
    assign layer0_out[287] = 1'b0;
    assign layer0_out[288] = ~(x[148] | x[149]);
    assign layer0_out[289] = 1'b0;
    assign layer0_out[290] = x[16] & ~x[15];
    assign layer0_out[291] = ~x[374];
    assign layer0_out[292] = x[137] | x[138];
    assign layer0_out[293] = x[291] & x[292];
    assign layer0_out[294] = ~(x[334] & x[335]);
    assign layer0_out[295] = 1'b1;
    assign layer0_out[296] = x[244] | x[245];
    assign layer0_out[297] = ~(x[22] | x[24]);
    assign layer0_out[298] = ~(x[102] | x[103]);
    assign layer0_out[299] = x[166] | x[167];
    assign layer0_out[300] = 1'b1;
    assign layer0_out[301] = ~(x[347] & x[348]);
    assign layer0_out[302] = x[141] | x[143];
    assign layer0_out[303] = x[29] & x[31];
    assign layer0_out[304] = x[96];
    assign layer0_out[305] = x[276] | x[277];
    assign layer0_out[306] = 1'b1;
    assign layer0_out[307] = ~(x[79] | x[80]);
    assign layer0_out[308] = 1'b0;
    assign layer0_out[309] = x[142] | x[144];
    assign layer0_out[310] = x[61];
    assign layer0_out[311] = x[11] | x[13];
    assign layer0_out[312] = 1'b1;
    assign layer0_out[313] = ~(x[301] | x[302]);
    assign layer0_out[314] = ~x[299];
    assign layer0_out[315] = ~(x[220] | x[221]);
    assign layer0_out[316] = ~(x[22] | x[23]);
    assign layer0_out[317] = ~(x[381] | x[382]);
    assign layer0_out[318] = ~(x[341] | x[342]);
    assign layer0_out[319] = x[137] | x[139];
    assign layer0_out[320] = ~(x[127] | x[128]);
    assign layer0_out[321] = ~(x[50] | x[51]);
    assign layer0_out[322] = 1'b1;
    assign layer0_out[323] = 1'b0;
    assign layer0_out[324] = ~(x[71] | x[73]);
    assign layer0_out[325] = 1'b0;
    assign layer0_out[326] = ~x[54];
    assign layer0_out[327] = ~(x[102] | x[104]);
    assign layer0_out[328] = ~x[81] | x[83];
    assign layer0_out[329] = 1'b1;
    assign layer0_out[330] = 1'b1;
    assign layer0_out[331] = ~x[350];
    assign layer0_out[332] = x[156] | x[157];
    assign layer0_out[333] = x[285] | x[286];
    assign layer0_out[334] = 1'b0;
    assign layer0_out[335] = x[140] | x[142];
    assign layer0_out[336] = ~(x[353] | x[354]);
    assign layer0_out[337] = x[132] | x[134];
    assign layer0_out[338] = x[78] | x[79];
    assign layer0_out[339] = ~x[173] | x[172];
    assign layer0_out[340] = x[187] | x[188];
    assign layer0_out[341] = ~x[62];
    assign layer0_out[342] = ~(x[110] & x[112]);
    assign layer0_out[343] = 1'b0;
    assign layer0_out[344] = ~(x[142] | x[143]);
    assign layer0_out[345] = ~(x[88] | x[89]);
    assign layer0_out[346] = x[331] | x[332];
    assign layer0_out[347] = x[50];
    assign layer0_out[348] = ~(x[85] | x[86]);
    assign layer0_out[349] = x[108] | x[110];
    assign layer0_out[350] = x[91] & x[92];
    assign layer0_out[351] = ~x[340];
    assign layer0_out[352] = x[136] | x[138];
    assign layer0_out[353] = x[64];
    assign layer0_out[354] = ~(x[317] | x[318]);
    assign layer0_out[355] = ~(x[97] | x[99]);
    assign layer0_out[356] = ~x[270];
    assign layer0_out[357] = ~x[346];
    assign layer0_out[358] = x[246];
    assign layer0_out[359] = x[120] & ~x[121];
    assign layer0_out[360] = ~(x[100] & x[102]);
    assign layer0_out[361] = ~(x[57] | x[59]);
    assign layer0_out[362] = ~x[147] | x[145];
    assign layer0_out[363] = x[44];
    assign layer0_out[364] = ~(x[178] | x[179]);
    assign layer0_out[365] = ~(x[115] | x[117]);
    assign layer0_out[366] = ~(x[263] | x[264]);
    assign layer0_out[367] = 1'b0;
    assign layer0_out[368] = 1'b1;
    assign layer0_out[369] = x[144] | x[146];
    assign layer0_out[370] = 1'b1;
    assign layer0_out[371] = x[278] | x[279];
    assign layer0_out[372] = x[87];
    assign layer0_out[373] = x[251];
    assign layer0_out[374] = x[176] | x[177];
    assign layer0_out[375] = x[149] & ~x[147];
    assign layer0_out[376] = 1'b0;
    assign layer0_out[377] = ~(x[60] | x[61]);
    assign layer0_out[378] = 1'b1;
    assign layer0_out[379] = x[123] | x[124];
    assign layer0_out[380] = ~(x[75] | x[77]);
    assign layer0_out[381] = x[36];
    assign layer0_out[382] = ~(x[107] & x[109]);
    assign layer0_out[383] = x[305] & ~x[306];
    assign layer0_out[384] = x[67];
    assign layer0_out[385] = ~x[22];
    assign layer0_out[386] = ~x[8];
    assign layer0_out[387] = ~x[23] | x[25];
    assign layer0_out[388] = ~(x[29] | x[30]);
    assign layer0_out[389] = 1'b0;
    assign layer0_out[390] = x[151] | x[152];
    assign layer0_out[391] = x[128];
    assign layer0_out[392] = x[338];
    assign layer0_out[393] = x[248] | x[249];
    assign layer0_out[394] = ~(x[69] & x[70]);
    assign layer0_out[395] = 1'b0;
    assign layer0_out[396] = x[311];
    assign layer0_out[397] = ~(x[204] | x[205]);
    assign layer0_out[398] = 1'b0;
    assign layer0_out[399] = 1'b0;
    assign layer0_out[400] = ~x[30];
    assign layer0_out[401] = 1'b1;
    assign layer0_out[402] = ~(x[368] | x[369]);
    assign layer0_out[403] = ~(x[157] | x[158]);
    assign layer0_out[404] = 1'b1;
    assign layer0_out[405] = 1'b0;
    assign layer0_out[406] = x[335] | x[336];
    assign layer0_out[407] = ~(x[134] | x[136]);
    assign layer0_out[408] = 1'b1;
    assign layer0_out[409] = x[77] | x[78];
    assign layer0_out[410] = ~(x[202] & x[203]);
    assign layer0_out[411] = ~(x[66] | x[67]);
    assign layer0_out[412] = ~x[397];
    assign layer0_out[413] = x[5] & ~x[6];
    assign layer0_out[414] = x[281] | x[282];
    assign layer0_out[415] = 1'b0;
    assign layer0_out[416] = x[122] | x[124];
    assign layer0_out[417] = 1'b1;
    assign layer0_out[418] = 1'b0;
    assign layer0_out[419] = 1'b0;
    assign layer0_out[420] = 1'b1;
    assign layer0_out[421] = x[180] | x[181];
    assign layer0_out[422] = ~x[61] | x[63];
    assign layer0_out[423] = ~(x[307] | x[308]);
    assign layer0_out[424] = x[398] | x[399];
    assign layer0_out[425] = ~x[38];
    assign layer0_out[426] = 1'b1;
    assign layer0_out[427] = x[320] | x[321];
    assign layer0_out[428] = 1'b1;
    assign layer0_out[429] = x[244];
    assign layer0_out[430] = ~(x[95] | x[97]);
    assign layer0_out[431] = ~(x[275] | x[276]);
    assign layer0_out[432] = ~(x[266] | x[267]);
    assign layer0_out[433] = 1'b1;
    assign layer0_out[434] = x[210] | x[211];
    assign layer0_out[435] = ~(x[302] | x[303]);
    assign layer0_out[436] = x[200];
    assign layer0_out[437] = ~x[179] | x[180];
    assign layer0_out[438] = x[362] | x[363];
    assign layer0_out[439] = x[146] | x[148];
    assign layer0_out[440] = ~(x[93] | x[95]);
    assign layer0_out[441] = ~(x[387] & x[388]);
    assign layer0_out[442] = x[304] | x[305];
    assign layer0_out[443] = ~(x[144] | x[145]);
    assign layer0_out[444] = ~(x[65] | x[66]);
    assign layer0_out[445] = 1'b1;
    assign layer0_out[446] = x[65] | x[67];
    assign layer0_out[447] = x[117] | x[118];
    assign layer0_out[448] = x[240];
    assign layer0_out[449] = ~(x[123] | x[125]);
    assign layer0_out[450] = 1'b1;
    assign layer0_out[451] = ~(x[357] | x[358]);
    assign layer0_out[452] = ~(x[127] | x[129]);
    assign layer0_out[453] = ~x[164];
    assign layer0_out[454] = 1'b1;
    assign layer0_out[455] = ~(x[196] | x[197]);
    assign layer0_out[456] = x[319];
    assign layer0_out[457] = x[183] & ~x[184];
    assign layer0_out[458] = ~(x[198] | x[199]);
    assign layer0_out[459] = ~(x[200] | x[201]);
    assign layer0_out[460] = x[9];
    assign layer0_out[461] = ~(x[345] | x[346]);
    assign layer0_out[462] = 1'b0;
    assign layer0_out[463] = x[6] | x[7];
    assign layer0_out[464] = x[38];
    assign layer0_out[465] = x[342];
    assign layer0_out[466] = x[264] | x[265];
    assign layer0_out[467] = 1'b1;
    assign layer0_out[468] = ~x[380];
    assign layer0_out[469] = x[94] & ~x[92];
    assign layer0_out[470] = ~(x[152] | x[153]);
    assign layer0_out[471] = x[389] | x[390];
    assign layer0_out[472] = ~(x[74] | x[75]);
    assign layer0_out[473] = ~(x[279] ^ x[280]);
    assign layer0_out[474] = ~(x[133] | x[134]);
    assign layer0_out[475] = 1'b1;
    assign layer0_out[476] = x[30] | x[31];
    assign layer0_out[477] = 1'b0;
    assign layer0_out[478] = ~(x[113] ^ x[115]);
    assign layer0_out[479] = ~x[40] | x[41];
    assign layer0_out[480] = ~(x[260] | x[261]);
    assign layer0_out[481] = x[314];
    assign layer0_out[482] = x[156];
    assign layer0_out[483] = x[361];
    assign layer0_out[484] = x[150];
    assign layer0_out[485] = 1'b1;
    assign layer0_out[486] = x[277] | x[278];
    assign layer0_out[487] = x[153] | x[154];
    assign layer0_out[488] = ~(x[216] | x[217]);
    assign layer0_out[489] = x[343] | x[344];
    assign layer0_out[490] = x[40] & ~x[39];
    assign layer0_out[491] = ~(x[44] | x[46]);
    assign layer0_out[492] = ~(x[104] | x[106]);
    assign layer0_out[493] = x[189];
    assign layer0_out[494] = x[191] | x[192];
    assign layer0_out[495] = x[19];
    assign layer0_out[496] = x[50] & x[52];
    assign layer0_out[497] = ~(x[185] | x[186]);
    assign layer0_out[498] = 1'b0;
    assign layer0_out[499] = ~(x[265] | x[266]);
    assign layer0_out[500] = ~(x[221] | x[222]);
    assign layer0_out[501] = ~(x[116] | x[118]);
    assign layer0_out[502] = 1'b0;
    assign layer0_out[503] = 1'b1;
    assign layer0_out[504] = ~(x[55] ^ x[57]);
    assign layer0_out[505] = x[271] | x[272];
    assign layer0_out[506] = ~x[8];
    assign layer0_out[507] = ~x[37];
    assign layer0_out[508] = ~(x[115] | x[116]);
    assign layer0_out[509] = ~(x[20] | x[22]);
    assign layer0_out[510] = x[188] | x[189];
    assign layer0_out[511] = 1'b0;
    assign layer0_out[512] = x[8] | x[10];
    assign layer0_out[513] = ~(x[90] | x[91]);
    assign layer0_out[514] = x[41] | x[43];
    assign layer0_out[515] = ~(x[238] | x[239]);
    assign layer0_out[516] = x[393] & ~x[392];
    assign layer0_out[517] = ~x[2];
    assign layer0_out[518] = ~x[367];
    assign layer0_out[519] = ~(x[122] | x[123]);
    assign layer0_out[520] = ~x[214];
    assign layer0_out[521] = 1'b1;
    assign layer0_out[522] = x[2];
    assign layer0_out[523] = 1'b1;
    assign layer0_out[524] = x[88] | x[90];
    assign layer0_out[525] = x[121] & ~x[123];
    assign layer0_out[526] = ~(x[324] | x[325]);
    assign layer0_out[527] = ~x[151];
    assign layer0_out[528] = ~x[131];
    assign layer0_out[529] = ~(x[83] | x[85]);
    assign layer0_out[530] = x[205];
    assign layer0_out[531] = x[143] | x[145];
    assign layer0_out[532] = ~(x[63] | x[64]);
    assign layer0_out[533] = ~(x[66] | x[68]);
    assign layer0_out[534] = x[99];
    assign layer0_out[535] = 1'b0;
    assign layer0_out[536] = 1'b0;
    assign layer0_out[537] = ~(x[94] | x[96]);
    assign layer0_out[538] = 1'b0;
    assign layer0_out[539] = 1'b0;
    assign layer0_out[540] = x[397] | x[398];
    assign layer0_out[541] = x[169] | x[170];
    assign layer0_out[542] = x[162] | x[163];
    assign layer0_out[543] = 1'b0;
    assign layer0_out[544] = x[201] | x[202];
    assign layer0_out[545] = x[267] | x[268];
    assign layer0_out[546] = 1'b1;
    assign layer0_out[547] = ~(x[135] | x[137]);
    assign layer0_out[548] = x[170] | x[171];
    assign layer0_out[549] = x[103] | x[104];
    assign layer1_out[0] = ~layer0_out[344];
    assign layer1_out[1] = layer0_out[487] & layer0_out[488];
    assign layer1_out[2] = ~layer0_out[286] | layer0_out[285];
    assign layer1_out[3] = layer0_out[177];
    assign layer1_out[4] = 1'b0;
    assign layer1_out[5] = ~layer0_out[431];
    assign layer1_out[6] = layer0_out[292];
    assign layer1_out[7] = layer0_out[249];
    assign layer1_out[8] = layer0_out[114];
    assign layer1_out[9] = layer0_out[196];
    assign layer1_out[10] = ~layer0_out[520] | layer0_out[519];
    assign layer1_out[11] = layer0_out[39];
    assign layer1_out[12] = ~layer0_out[54];
    assign layer1_out[13] = ~layer0_out[165];
    assign layer1_out[14] = layer0_out[493];
    assign layer1_out[15] = layer0_out[84] | layer0_out[85];
    assign layer1_out[16] = ~layer0_out[87] | layer0_out[86];
    assign layer1_out[17] = ~layer0_out[117] | layer0_out[118];
    assign layer1_out[18] = layer0_out[379] & ~layer0_out[378];
    assign layer1_out[19] = layer0_out[531];
    assign layer1_out[20] = 1'b0;
    assign layer1_out[21] = 1'b1;
    assign layer1_out[22] = 1'b1;
    assign layer1_out[23] = ~layer0_out[441] | layer0_out[442];
    assign layer1_out[24] = layer0_out[12];
    assign layer1_out[25] = layer0_out[102] & ~layer0_out[103];
    assign layer1_out[26] = 1'b0;
    assign layer1_out[27] = ~(layer0_out[250] ^ layer0_out[251]);
    assign layer1_out[28] = ~layer0_out[512] | layer0_out[513];
    assign layer1_out[29] = 1'b1;
    assign layer1_out[30] = ~layer0_out[151];
    assign layer1_out[31] = layer0_out[296];
    assign layer1_out[32] = ~layer0_out[491] | layer0_out[490];
    assign layer1_out[33] = layer0_out[348];
    assign layer1_out[34] = layer0_out[83];
    assign layer1_out[35] = layer0_out[204];
    assign layer1_out[36] = layer0_out[549];
    assign layer1_out[37] = layer0_out[66] | layer0_out[67];
    assign layer1_out[38] = ~(layer0_out[213] & layer0_out[214]);
    assign layer1_out[39] = layer0_out[303] | layer0_out[304];
    assign layer1_out[40] = layer0_out[67];
    assign layer1_out[41] = ~layer0_out[99];
    assign layer1_out[42] = layer0_out[191] & ~layer0_out[192];
    assign layer1_out[43] = layer0_out[73];
    assign layer1_out[44] = layer0_out[449] & ~layer0_out[448];
    assign layer1_out[45] = 1'b0;
    assign layer1_out[46] = 1'b1;
    assign layer1_out[47] = 1'b0;
    assign layer1_out[48] = ~layer0_out[307];
    assign layer1_out[49] = layer0_out[418] & layer0_out[419];
    assign layer1_out[50] = layer0_out[206];
    assign layer1_out[51] = ~layer0_out[145] | layer0_out[144];
    assign layer1_out[52] = ~layer0_out[508];
    assign layer1_out[53] = layer0_out[491] & layer0_out[492];
    assign layer1_out[54] = 1'b1;
    assign layer1_out[55] = layer0_out[453] & ~layer0_out[452];
    assign layer1_out[56] = ~layer0_out[327];
    assign layer1_out[57] = layer0_out[421];
    assign layer1_out[58] = 1'b1;
    assign layer1_out[59] = layer0_out[78] | layer0_out[79];
    assign layer1_out[60] = ~layer0_out[499];
    assign layer1_out[61] = ~(layer0_out[184] | layer0_out[185]);
    assign layer1_out[62] = layer0_out[299];
    assign layer1_out[63] = ~(layer0_out[423] & layer0_out[424]);
    assign layer1_out[64] = ~(layer0_out[210] | layer0_out[211]);
    assign layer1_out[65] = ~(layer0_out[458] | layer0_out[459]);
    assign layer1_out[66] = ~(layer0_out[524] | layer0_out[525]);
    assign layer1_out[67] = ~(layer0_out[515] | layer0_out[516]);
    assign layer1_out[68] = 1'b1;
    assign layer1_out[69] = layer0_out[276] & ~layer0_out[275];
    assign layer1_out[70] = layer0_out[95];
    assign layer1_out[71] = ~layer0_out[366];
    assign layer1_out[72] = ~layer0_out[124];
    assign layer1_out[73] = 1'b1;
    assign layer1_out[74] = layer0_out[506] | layer0_out[507];
    assign layer1_out[75] = layer0_out[317] & layer0_out[318];
    assign layer1_out[76] = ~layer0_out[52];
    assign layer1_out[77] = layer0_out[265];
    assign layer1_out[78] = layer0_out[159] & layer0_out[160];
    assign layer1_out[79] = layer0_out[524];
    assign layer1_out[80] = layer0_out[161];
    assign layer1_out[81] = ~layer0_out[23];
    assign layer1_out[82] = layer0_out[201] & ~layer0_out[202];
    assign layer1_out[83] = ~(layer0_out[7] | layer0_out[8]);
    assign layer1_out[84] = ~(layer0_out[243] & layer0_out[244]);
    assign layer1_out[85] = layer0_out[402];
    assign layer1_out[86] = 1'b1;
    assign layer1_out[87] = layer0_out[88];
    assign layer1_out[88] = ~layer0_out[545];
    assign layer1_out[89] = layer0_out[107] ^ layer0_out[108];
    assign layer1_out[90] = ~layer0_out[299];
    assign layer1_out[91] = ~(layer0_out[98] | layer0_out[99]);
    assign layer1_out[92] = 1'b1;
    assign layer1_out[93] = ~(layer0_out[328] | layer0_out[329]);
    assign layer1_out[94] = layer0_out[400];
    assign layer1_out[95] = 1'b0;
    assign layer1_out[96] = layer0_out[416];
    assign layer1_out[97] = ~(layer0_out[412] | layer0_out[413]);
    assign layer1_out[98] = layer0_out[356] & ~layer0_out[357];
    assign layer1_out[99] = layer0_out[518];
    assign layer1_out[100] = ~layer0_out[301];
    assign layer1_out[101] = layer0_out[188] & ~layer0_out[189];
    assign layer1_out[102] = layer0_out[532] & layer0_out[533];
    assign layer1_out[103] = ~layer0_out[403];
    assign layer1_out[104] = 1'b0;
    assign layer1_out[105] = layer0_out[117];
    assign layer1_out[106] = layer0_out[320] & ~layer0_out[321];
    assign layer1_out[107] = layer0_out[347];
    assign layer1_out[108] = layer0_out[232];
    assign layer1_out[109] = ~layer0_out[54] | layer0_out[55];
    assign layer1_out[110] = layer0_out[542];
    assign layer1_out[111] = layer0_out[522];
    assign layer1_out[112] = 1'b1;
    assign layer1_out[113] = layer0_out[393];
    assign layer1_out[114] = layer0_out[35] & layer0_out[36];
    assign layer1_out[115] = ~layer0_out[32] | layer0_out[31];
    assign layer1_out[116] = 1'b1;
    assign layer1_out[117] = ~layer0_out[373] | layer0_out[372];
    assign layer1_out[118] = ~(layer0_out[134] & layer0_out[135]);
    assign layer1_out[119] = ~layer0_out[461] | layer0_out[460];
    assign layer1_out[120] = 1'b1;
    assign layer1_out[121] = ~layer0_out[284];
    assign layer1_out[122] = ~(layer0_out[374] & layer0_out[375]);
    assign layer1_out[123] = ~(layer0_out[115] & layer0_out[116]);
    assign layer1_out[124] = ~layer0_out[343] | layer0_out[344];
    assign layer1_out[125] = layer0_out[148] | layer0_out[149];
    assign layer1_out[126] = 1'b1;
    assign layer1_out[127] = 1'b1;
    assign layer1_out[128] = layer0_out[479] | layer0_out[480];
    assign layer1_out[129] = ~layer0_out[39];
    assign layer1_out[130] = layer0_out[81] & ~layer0_out[82];
    assign layer1_out[131] = layer0_out[149];
    assign layer1_out[132] = layer0_out[130] & ~layer0_out[129];
    assign layer1_out[133] = layer0_out[353] & layer0_out[354];
    assign layer1_out[134] = ~(layer0_out[218] | layer0_out[219]);
    assign layer1_out[135] = layer0_out[181];
    assign layer1_out[136] = ~layer0_out[187];
    assign layer1_out[137] = layer0_out[530] | layer0_out[531];
    assign layer1_out[138] = ~layer0_out[14] | layer0_out[13];
    assign layer1_out[139] = layer0_out[109];
    assign layer1_out[140] = ~layer0_out[290] | layer0_out[291];
    assign layer1_out[141] = ~layer0_out[18] | layer0_out[19];
    assign layer1_out[142] = layer0_out[340];
    assign layer1_out[143] = ~layer0_out[320];
    assign layer1_out[144] = 1'b1;
    assign layer1_out[145] = ~layer0_out[178];
    assign layer1_out[146] = ~layer0_out[333] | layer0_out[334];
    assign layer1_out[147] = layer0_out[150] & layer0_out[151];
    assign layer1_out[148] = ~(layer0_out[262] & layer0_out[263]);
    assign layer1_out[149] = layer0_out[174] & ~layer0_out[173];
    assign layer1_out[150] = ~layer0_out[191];
    assign layer1_out[151] = ~layer0_out[407];
    assign layer1_out[152] = 1'b0;
    assign layer1_out[153] = ~layer0_out[390];
    assign layer1_out[154] = ~layer0_out[5] | layer0_out[6];
    assign layer1_out[155] = layer0_out[381] & layer0_out[382];
    assign layer1_out[156] = ~layer0_out[197] | layer0_out[196];
    assign layer1_out[157] = layer0_out[139] | layer0_out[140];
    assign layer1_out[158] = ~layer0_out[49];
    assign layer1_out[159] = 1'b0;
    assign layer1_out[160] = layer0_out[200] & layer0_out[201];
    assign layer1_out[161] = layer0_out[374] & ~layer0_out[373];
    assign layer1_out[162] = layer0_out[415] | layer0_out[416];
    assign layer1_out[163] = layer0_out[30];
    assign layer1_out[164] = layer0_out[148] & ~layer0_out[147];
    assign layer1_out[165] = layer0_out[221] & ~layer0_out[222];
    assign layer1_out[166] = ~layer0_out[182];
    assign layer1_out[167] = 1'b1;
    assign layer1_out[168] = ~layer0_out[309] | layer0_out[308];
    assign layer1_out[169] = layer0_out[258];
    assign layer1_out[170] = layer0_out[105] | layer0_out[106];
    assign layer1_out[171] = layer0_out[195];
    assign layer1_out[172] = layer0_out[363] & ~layer0_out[362];
    assign layer1_out[173] = 1'b1;
    assign layer1_out[174] = 1'b1;
    assign layer1_out[175] = 1'b1;
    assign layer1_out[176] = ~layer0_out[288];
    assign layer1_out[177] = layer0_out[429];
    assign layer1_out[178] = layer0_out[101] | layer0_out[102];
    assign layer1_out[179] = 1'b0;
    assign layer1_out[180] = layer0_out[166] | layer0_out[167];
    assign layer1_out[181] = 1'b1;
    assign layer1_out[182] = ~layer0_out[127] | layer0_out[126];
    assign layer1_out[183] = ~layer0_out[456];
    assign layer1_out[184] = ~layer0_out[254];
    assign layer1_out[185] = layer0_out[342] | layer0_out[343];
    assign layer1_out[186] = layer0_out[305];
    assign layer1_out[187] = layer0_out[321] & ~layer0_out[322];
    assign layer1_out[188] = ~(layer0_out[527] & layer0_out[528]);
    assign layer1_out[189] = layer0_out[20] & ~layer0_out[21];
    assign layer1_out[190] = ~layer0_out[113];
    assign layer1_out[191] = layer0_out[106] & ~layer0_out[107];
    assign layer1_out[192] = ~(layer0_out[385] & layer0_out[386]);
    assign layer1_out[193] = ~layer0_out[414];
    assign layer1_out[194] = ~(layer0_out[411] & layer0_out[412]);
    assign layer1_out[195] = ~layer0_out[337];
    assign layer1_out[196] = 1'b1;
    assign layer1_out[197] = ~layer0_out[313];
    assign layer1_out[198] = ~layer0_out[80];
    assign layer1_out[199] = ~layer0_out[400];
    assign layer1_out[200] = layer0_out[363] ^ layer0_out[364];
    assign layer1_out[201] = layer0_out[113];
    assign layer1_out[202] = layer0_out[356];
    assign layer1_out[203] = layer0_out[504] & layer0_out[505];
    assign layer1_out[204] = layer0_out[475] & ~layer0_out[476];
    assign layer1_out[205] = layer0_out[535] & layer0_out[536];
    assign layer1_out[206] = layer0_out[503];
    assign layer1_out[207] = layer0_out[318] | layer0_out[319];
    assign layer1_out[208] = ~layer0_out[418] | layer0_out[417];
    assign layer1_out[209] = layer0_out[369];
    assign layer1_out[210] = layer0_out[244] | layer0_out[245];
    assign layer1_out[211] = ~layer0_out[69] | layer0_out[70];
    assign layer1_out[212] = layer0_out[488] & ~layer0_out[489];
    assign layer1_out[213] = ~layer0_out[188];
    assign layer1_out[214] = ~layer0_out[72];
    assign layer1_out[215] = ~layer0_out[241];
    assign layer1_out[216] = ~layer0_out[168] | layer0_out[167];
    assign layer1_out[217] = layer0_out[156] | layer0_out[157];
    assign layer1_out[218] = 1'b0;
    assign layer1_out[219] = layer0_out[33] | layer0_out[34];
    assign layer1_out[220] = layer0_out[269] & ~layer0_out[270];
    assign layer1_out[221] = 1'b1;
    assign layer1_out[222] = ~layer0_out[288] | layer0_out[289];
    assign layer1_out[223] = 1'b1;
    assign layer1_out[224] = ~layer0_out[72] | layer0_out[73];
    assign layer1_out[225] = 1'b1;
    assign layer1_out[226] = layer0_out[1] & layer0_out[2];
    assign layer1_out[227] = ~layer0_out[377] | layer0_out[376];
    assign layer1_out[228] = ~layer0_out[336];
    assign layer1_out[229] = ~layer0_out[242];
    assign layer1_out[230] = layer0_out[448];
    assign layer1_out[231] = ~layer0_out[427];
    assign layer1_out[232] = ~layer0_out[96];
    assign layer1_out[233] = ~(layer0_out[118] | layer0_out[119]);
    assign layer1_out[234] = ~layer0_out[125];
    assign layer1_out[235] = ~layer0_out[155] | layer0_out[156];
    assign layer1_out[236] = layer0_out[542];
    assign layer1_out[237] = ~(layer0_out[337] | layer0_out[338]);
    assign layer1_out[238] = ~layer0_out[153];
    assign layer1_out[239] = ~layer0_out[165];
    assign layer1_out[240] = layer0_out[443] & layer0_out[444];
    assign layer1_out[241] = 1'b1;
    assign layer1_out[242] = layer0_out[258] & layer0_out[259];
    assign layer1_out[243] = layer0_out[309];
    assign layer1_out[244] = layer0_out[339] & ~layer0_out[338];
    assign layer1_out[245] = ~layer0_out[529];
    assign layer1_out[246] = ~(layer0_out[366] & layer0_out[367]);
    assign layer1_out[247] = layer0_out[315];
    assign layer1_out[248] = layer0_out[437] & ~layer0_out[436];
    assign layer1_out[249] = layer0_out[450] | layer0_out[451];
    assign layer1_out[250] = layer0_out[355];
    assign layer1_out[251] = layer0_out[388];
    assign layer1_out[252] = layer0_out[279] & ~layer0_out[280];
    assign layer1_out[253] = ~layer0_out[217];
    assign layer1_out[254] = ~(layer0_out[137] | layer0_out[138]);
    assign layer1_out[255] = ~layer0_out[45];
    assign layer1_out[256] = 1'b0;
    assign layer1_out[257] = layer0_out[47] & ~layer0_out[46];
    assign layer1_out[258] = layer0_out[210];
    assign layer1_out[259] = 1'b0;
    assign layer1_out[260] = layer0_out[173];
    assign layer1_out[261] = ~layer0_out[298] | layer0_out[297];
    assign layer1_out[262] = layer0_out[455] & ~layer0_out[456];
    assign layer1_out[263] = layer0_out[233] & layer0_out[234];
    assign layer1_out[264] = ~(layer0_out[543] | layer0_out[544]);
    assign layer1_out[265] = 1'b0;
    assign layer1_out[266] = 1'b1;
    assign layer1_out[267] = layer0_out[57] & layer0_out[58];
    assign layer1_out[268] = layer0_out[192] | layer0_out[193];
    assign layer1_out[269] = layer0_out[425];
    assign layer1_out[270] = layer0_out[207];
    assign layer1_out[271] = ~(layer0_out[516] & layer0_out[517]);
    assign layer1_out[272] = layer0_out[5] & ~layer0_out[4];
    assign layer1_out[273] = 1'b1;
    assign layer1_out[274] = 1'b0;
    assign layer1_out[275] = ~layer0_out[375];
    assign layer1_out[276] = ~layer0_out[493];
    assign layer1_out[277] = layer0_out[28];
    assign layer1_out[278] = layer0_out[419] & ~layer0_out[420];
    assign layer1_out[279] = ~(layer0_out[96] | layer0_out[97]);
    assign layer1_out[280] = 1'b0;
    assign layer1_out[281] = layer0_out[406];
    assign layer1_out[282] = ~layer0_out[437] | layer0_out[438];
    assign layer1_out[283] = layer0_out[477] & ~layer0_out[478];
    assign layer1_out[284] = layer0_out[59];
    assign layer1_out[285] = ~layer0_out[331];
    assign layer1_out[286] = layer0_out[348] & layer0_out[349];
    assign layer1_out[287] = layer0_out[183] & ~layer0_out[184];
    assign layer1_out[288] = ~(layer0_out[235] & layer0_out[236]);
    assign layer1_out[289] = 1'b1;
    assign layer1_out[290] = ~(layer0_out[446] | layer0_out[447]);
    assign layer1_out[291] = ~layer0_out[466];
    assign layer1_out[292] = ~(layer0_out[467] | layer0_out[468]);
    assign layer1_out[293] = layer0_out[445];
    assign layer1_out[294] = layer0_out[259];
    assign layer1_out[295] = layer0_out[380] & ~layer0_out[381];
    assign layer1_out[296] = 1'b1;
    assign layer1_out[297] = 1'b1;
    assign layer1_out[298] = ~layer0_out[14];
    assign layer1_out[299] = layer0_out[40] & layer0_out[41];
    assign layer1_out[300] = layer0_out[267] & layer0_out[268];
    assign layer1_out[301] = layer0_out[121] & ~layer0_out[120];
    assign layer1_out[302] = layer0_out[262];
    assign layer1_out[303] = layer0_out[484] | layer0_out[485];
    assign layer1_out[304] = 1'b1;
    assign layer1_out[305] = layer0_out[93] & layer0_out[94];
    assign layer1_out[306] = ~(layer0_out[478] & layer0_out[479]);
    assign layer1_out[307] = 1'b0;
    assign layer1_out[308] = layer0_out[131];
    assign layer1_out[309] = ~layer0_out[512];
    assign layer1_out[310] = 1'b0;
    assign layer1_out[311] = ~layer0_out[22] | layer0_out[21];
    assign layer1_out[312] = ~layer0_out[391] | layer0_out[392];
    assign layer1_out[313] = layer0_out[407] & ~layer0_out[406];
    assign layer1_out[314] = ~layer0_out[443] | layer0_out[442];
    assign layer1_out[315] = 1'b0;
    assign layer1_out[316] = ~(layer0_out[370] & layer0_out[371]);
    assign layer1_out[317] = 1'b0;
    assign layer1_out[318] = ~(layer0_out[429] | layer0_out[430]);
    assign layer1_out[319] = ~(layer0_out[171] | layer0_out[172]);
    assign layer1_out[320] = ~layer0_out[302];
    assign layer1_out[321] = ~layer0_out[449];
    assign layer1_out[322] = 1'b0;
    assign layer1_out[323] = layer0_out[135] | layer0_out[136];
    assign layer1_out[324] = ~layer0_out[540];
    assign layer1_out[325] = layer0_out[311] & ~layer0_out[310];
    assign layer1_out[326] = layer0_out[489];
    assign layer1_out[327] = layer0_out[69] & ~layer0_out[68];
    assign layer1_out[328] = ~(layer0_out[499] & layer0_out[500]);
    assign layer1_out[329] = ~layer0_out[217];
    assign layer1_out[330] = 1'b0;
    assign layer1_out[331] = layer0_out[206] & layer0_out[207];
    assign layer1_out[332] = ~(layer0_out[234] & layer0_out[235]);
    assign layer1_out[333] = 1'b1;
    assign layer1_out[334] = ~layer0_out[239];
    assign layer1_out[335] = layer0_out[476];
    assign layer1_out[336] = ~layer0_out[24] | layer0_out[25];
    assign layer1_out[337] = 1'b1;
    assign layer1_out[338] = ~layer0_out[527] | layer0_out[526];
    assign layer1_out[339] = layer0_out[481] & ~layer0_out[480];
    assign layer1_out[340] = layer0_out[143] & layer0_out[144];
    assign layer1_out[341] = layer0_out[463];
    assign layer1_out[342] = ~layer0_out[547];
    assign layer1_out[343] = ~(layer0_out[50] ^ layer0_out[51]);
    assign layer1_out[344] = layer0_out[510];
    assign layer1_out[345] = ~(layer0_out[329] | layer0_out[330]);
    assign layer1_out[346] = ~layer0_out[461];
    assign layer1_out[347] = layer0_out[162] & layer0_out[163];
    assign layer1_out[348] = ~layer0_out[111];
    assign layer1_out[349] = 1'b1;
    assign layer1_out[350] = layer0_out[340];
    assign layer1_out[351] = ~layer0_out[294] | layer0_out[293];
    assign layer1_out[352] = ~(layer0_out[62] | layer0_out[63]);
    assign layer1_out[353] = layer0_out[482];
    assign layer1_out[354] = layer0_out[205] & ~layer0_out[204];
    assign layer1_out[355] = layer0_out[97] & layer0_out[98];
    assign layer1_out[356] = ~layer0_out[6] | layer0_out[7];
    assign layer1_out[357] = ~layer0_out[214];
    assign layer1_out[358] = layer0_out[358];
    assign layer1_out[359] = ~layer0_out[547] | layer0_out[548];
    assign layer1_out[360] = ~layer0_out[246] | layer0_out[247];
    assign layer1_out[361] = ~(layer0_out[3] & layer0_out[4]);
    assign layer1_out[362] = layer0_out[335];
    assign layer1_out[363] = layer0_out[109];
    assign layer1_out[364] = ~layer0_out[249] | layer0_out[248];
    assign layer1_out[365] = ~layer0_out[283];
    assign layer1_out[366] = layer0_out[441] & ~layer0_out[440];
    assign layer1_out[367] = 1'b1;
    assign layer1_out[368] = layer0_out[119] & layer0_out[120];
    assign layer1_out[369] = ~layer0_out[255];
    assign layer1_out[370] = ~layer0_out[34];
    assign layer1_out[371] = layer0_out[267];
    assign layer1_out[372] = layer0_out[358];
    assign layer1_out[373] = layer0_out[19] & layer0_out[20];
    assign layer1_out[374] = layer0_out[501];
    assign layer1_out[375] = ~layer0_out[323] | layer0_out[322];
    assign layer1_out[376] = 1'b1;
    assign layer1_out[377] = 1'b1;
    assign layer1_out[378] = layer0_out[396] & ~layer0_out[397];
    assign layer1_out[379] = ~layer0_out[470];
    assign layer1_out[380] = layer0_out[471] & ~layer0_out[472];
    assign layer1_out[381] = ~layer0_out[3] | layer0_out[2];
    assign layer1_out[382] = ~(layer0_out[198] | layer0_out[199]);
    assign layer1_out[383] = layer0_out[236];
    assign layer1_out[384] = 1'b0;
    assign layer1_out[385] = layer0_out[414];
    assign layer1_out[386] = 1'b0;
    assign layer1_out[387] = layer0_out[469];
    assign layer1_out[388] = layer0_out[213] & ~layer0_out[212];
    assign layer1_out[389] = ~layer0_out[277];
    assign layer1_out[390] = ~layer0_out[545] | layer0_out[544];
    assign layer1_out[391] = ~layer0_out[255] | layer0_out[254];
    assign layer1_out[392] = layer0_out[324];
    assign layer1_out[393] = layer0_out[409] & layer0_out[410];
    assign layer1_out[394] = 1'b0;
    assign layer1_out[395] = layer0_out[388];
    assign layer1_out[396] = layer0_out[291] | layer0_out[292];
    assign layer1_out[397] = layer0_out[434] & layer0_out[435];
    assign layer1_out[398] = ~layer0_out[367] | layer0_out[368];
    assign layer1_out[399] = layer0_out[351] & ~layer0_out[352];
    assign layer1_out[400] = layer0_out[65] & layer0_out[66];
    assign layer1_out[401] = ~layer0_out[177];
    assign layer1_out[402] = 1'b0;
    assign layer1_out[403] = ~(layer0_out[83] ^ layer0_out[84]);
    assign layer1_out[404] = layer0_out[55];
    assign layer1_out[405] = ~layer0_out[394];
    assign layer1_out[406] = ~layer0_out[232] | layer0_out[231];
    assign layer1_out[407] = 1'b0;
    assign layer1_out[408] = ~layer0_out[496] | layer0_out[497];
    assign layer1_out[409] = layer0_out[453];
    assign layer1_out[410] = ~(layer0_out[100] & layer0_out[101]);
    assign layer1_out[411] = ~(layer0_out[36] | layer0_out[37]);
    assign layer1_out[412] = ~layer0_out[230];
    assign layer1_out[413] = layer0_out[16];
    assign layer1_out[414] = 1'b0;
    assign layer1_out[415] = layer0_out[526] & ~layer0_out[525];
    assign layer1_out[416] = layer0_out[56];
    assign layer1_out[417] = layer0_out[459];
    assign layer1_out[418] = ~(layer0_out[422] & layer0_out[423]);
    assign layer1_out[419] = ~layer0_out[219];
    assign layer1_out[420] = ~layer0_out[77] | layer0_out[76];
    assign layer1_out[421] = 1'b1;
    assign layer1_out[422] = 1'b1;
    assign layer1_out[423] = layer0_out[231];
    assign layer1_out[424] = layer0_out[42] & layer0_out[43];
    assign layer1_out[425] = layer0_out[260];
    assign layer1_out[426] = layer0_out[315] & layer0_out[316];
    assign layer1_out[427] = 1'b0;
    assign layer1_out[428] = ~layer0_out[435];
    assign layer1_out[429] = layer0_out[534];
    assign layer1_out[430] = layer0_out[275];
    assign layer1_out[431] = layer0_out[303];
    assign layer1_out[432] = ~(layer0_out[189] & layer0_out[190]);
    assign layer1_out[433] = ~layer0_out[494];
    assign layer1_out[434] = 1'b0;
    assign layer1_out[435] = ~layer0_out[390];
    assign layer1_out[436] = ~(layer0_out[37] & layer0_out[38]);
    assign layer1_out[437] = ~layer0_out[181];
    assign layer1_out[438] = layer0_out[377];
    assign layer1_out[439] = ~layer0_out[220] | layer0_out[221];
    assign layer1_out[440] = layer0_out[252] | layer0_out[253];
    assign layer1_out[441] = layer0_out[397] & layer0_out[398];
    assign layer1_out[442] = ~(layer0_out[163] & layer0_out[164]);
    assign layer1_out[443] = ~(layer0_out[141] & layer0_out[142]);
    assign layer1_out[444] = layer0_out[421];
    assign layer1_out[445] = layer0_out[314];
    assign layer1_out[446] = ~(layer0_out[509] & layer0_out[510]);
    assign layer1_out[447] = layer0_out[507] | layer0_out[508];
    assign layer1_out[448] = 1'b1;
    assign layer1_out[449] = 1'b0;
    assign layer1_out[450] = layer0_out[176];
    assign layer1_out[451] = layer0_out[383];
    assign layer1_out[452] = 1'b0;
    assign layer1_out[453] = layer0_out[501];
    assign layer1_out[454] = layer0_out[80] | layer0_out[81];
    assign layer1_out[455] = layer0_out[470] & ~layer0_out[469];
    assign layer1_out[456] = ~layer0_out[537];
    assign layer1_out[457] = layer0_out[333];
    assign layer1_out[458] = ~(layer0_out[103] | layer0_out[104]);
    assign layer1_out[459] = layer0_out[270];
    assign layer1_out[460] = layer0_out[256] | layer0_out[257];
    assign layer1_out[461] = layer0_out[91] & ~layer0_out[90];
    assign layer1_out[462] = ~(layer0_out[465] | layer0_out[466]);
    assign layer1_out[463] = layer0_out[45] & ~layer0_out[46];
    assign layer1_out[464] = layer0_out[211];
    assign layer1_out[465] = layer0_out[142] & ~layer0_out[143];
    assign layer1_out[466] = ~layer0_out[265];
    assign layer1_out[467] = 1'b1;
    assign layer1_out[468] = layer0_out[439];
    assign layer1_out[469] = layer0_out[128];
    assign layer1_out[470] = 1'b0;
    assign layer1_out[471] = layer0_out[379];
    assign layer1_out[472] = ~layer0_out[474];
    assign layer1_out[473] = ~(layer0_out[170] & layer0_out[171]);
    assign layer1_out[474] = ~layer0_out[341] | layer0_out[342];
    assign layer1_out[475] = ~layer0_out[199];
    assign layer1_out[476] = ~layer0_out[222] | layer0_out[223];
    assign layer1_out[477] = layer0_out[517] & ~layer0_out[518];
    assign layer1_out[478] = layer0_out[10] & ~layer0_out[9];
    assign layer1_out[479] = 1'b1;
    assign layer1_out[480] = layer0_out[505];
    assign layer1_out[481] = ~layer0_out[365];
    assign layer1_out[482] = 1'b1;
    assign layer1_out[483] = layer0_out[43] | layer0_out[44];
    assign layer1_out[484] = ~(layer0_out[486] ^ layer0_out[487]);
    assign layer1_out[485] = ~(layer0_out[495] | layer0_out[496]);
    assign layer1_out[486] = layer0_out[464] & ~layer0_out[465];
    assign layer1_out[487] = layer0_out[240] & ~layer0_out[239];
    assign layer1_out[488] = layer0_out[12];
    assign layer1_out[489] = layer0_out[454] & ~layer0_out[455];
    assign layer1_out[490] = ~layer0_out[440];
    assign layer1_out[491] = layer0_out[70];
    assign layer1_out[492] = 1'b0;
    assign layer1_out[493] = ~(layer0_out[316] | layer0_out[317]);
    assign layer1_out[494] = ~(layer0_out[224] | layer0_out[225]);
    assign layer1_out[495] = layer0_out[272] | layer0_out[273];
    assign layer1_out[496] = ~layer0_out[16];
    assign layer1_out[497] = ~(layer0_out[168] ^ layer0_out[169]);
    assign layer1_out[498] = ~layer0_out[203];
    assign layer1_out[499] = layer0_out[283] & layer0_out[284];
    assign layer1_out[500] = layer0_out[514] & ~layer0_out[515];
    assign layer1_out[501] = 1'b0;
    assign layer1_out[502] = ~layer0_out[361];
    assign layer1_out[503] = layer0_out[268] & layer0_out[269];
    assign layer1_out[504] = 1'b0;
    assign layer1_out[505] = layer0_out[289] | layer0_out[290];
    assign layer1_out[506] = layer0_out[62];
    assign layer1_out[507] = layer0_out[541];
    assign layer1_out[508] = ~layer0_out[241];
    assign layer1_out[509] = ~layer0_out[127];
    assign layer1_out[510] = 1'b0;
    assign layer1_out[511] = layer0_out[484];
    assign layer1_out[512] = layer0_out[473] & ~layer0_out[474];
    assign layer1_out[513] = layer0_out[306] | layer0_out[307];
    assign layer1_out[514] = ~layer0_out[393];
    assign layer1_out[515] = ~layer0_out[432];
    assign layer1_out[516] = layer0_out[197] & layer0_out[198];
    assign layer1_out[517] = ~layer0_out[77];
    assign layer1_out[518] = ~layer0_out[282] | layer0_out[281];
    assign layer1_out[519] = ~layer0_out[311];
    assign layer1_out[520] = ~layer0_out[486];
    assign layer1_out[521] = layer0_out[326];
    assign layer1_out[522] = 1'b0;
    assign layer1_out[523] = layer0_out[345] & ~layer0_out[346];
    assign layer1_out[524] = layer0_out[351] & ~layer0_out[350];
    assign layer1_out[525] = ~(layer0_out[208] | layer0_out[209]);
    assign layer1_out[526] = layer0_out[497];
    assign layer1_out[527] = 1'b0;
    assign layer1_out[528] = layer0_out[8] | layer0_out[9];
    assign layer1_out[529] = 1'b0;
    assign layer1_out[530] = 1'b0;
    assign layer1_out[531] = layer0_out[179];
    assign layer1_out[532] = ~layer0_out[158];
    assign layer1_out[533] = ~layer0_out[451] | layer0_out[452];
    assign layer1_out[534] = layer0_out[383] | layer0_out[384];
    assign layer1_out[535] = layer0_out[386] & ~layer0_out[387];
    assign layer1_out[536] = ~(layer0_out[0] & layer0_out[2]);
    assign layer1_out[537] = layer0_out[41] & ~layer0_out[42];
    assign layer1_out[538] = ~(layer0_out[513] | layer0_out[514]);
    assign layer1_out[539] = ~layer0_out[193] | layer0_out[194];
    assign layer1_out[540] = ~layer0_out[226];
    assign layer1_out[541] = layer0_out[123];
    assign layer1_out[542] = layer0_out[121] | layer0_out[122];
    assign layer1_out[543] = 1'b0;
    assign layer1_out[544] = ~(layer0_out[294] | layer0_out[295]);
    assign layer1_out[545] = layer0_out[174] & ~layer0_out[175];
    assign layer1_out[546] = ~layer0_out[64];
    assign layer1_out[547] = layer0_out[245];
    assign layer1_out[548] = ~layer0_out[133];
    assign layer1_out[549] = 1'b1;
    assign layer2_out[0] = ~layer1_out[512];
    assign layer2_out[1] = ~(layer1_out[126] | layer1_out[127]);
    assign layer2_out[2] = layer1_out[103];
    assign layer2_out[3] = ~layer1_out[24] | layer1_out[25];
    assign layer2_out[4] = ~layer1_out[342];
    assign layer2_out[5] = layer1_out[326];
    assign layer2_out[6] = layer1_out[230];
    assign layer2_out[7] = ~(layer1_out[214] | layer1_out[215]);
    assign layer2_out[8] = layer1_out[308] & ~layer1_out[307];
    assign layer2_out[9] = layer1_out[158] & ~layer1_out[157];
    assign layer2_out[10] = layer1_out[195];
    assign layer2_out[11] = layer1_out[99];
    assign layer2_out[12] = 1'b1;
    assign layer2_out[13] = ~layer1_out[119];
    assign layer2_out[14] = ~layer1_out[83];
    assign layer2_out[15] = layer1_out[58] | layer1_out[59];
    assign layer2_out[16] = ~(layer1_out[488] & layer1_out[489]);
    assign layer2_out[17] = layer1_out[284] & layer1_out[285];
    assign layer2_out[18] = layer1_out[493] | layer1_out[494];
    assign layer2_out[19] = layer1_out[290] & layer1_out[291];
    assign layer2_out[20] = layer1_out[67] & ~layer1_out[68];
    assign layer2_out[21] = ~layer1_out[139];
    assign layer2_out[22] = ~layer1_out[399] | layer1_out[400];
    assign layer2_out[23] = ~layer1_out[27];
    assign layer2_out[24] = 1'b0;
    assign layer2_out[25] = ~layer1_out[60];
    assign layer2_out[26] = layer1_out[378];
    assign layer2_out[27] = ~layer1_out[10] | layer1_out[9];
    assign layer2_out[28] = 1'b1;
    assign layer2_out[29] = ~layer1_out[145];
    assign layer2_out[30] = layer1_out[324];
    assign layer2_out[31] = ~layer1_out[85];
    assign layer2_out[32] = ~layer1_out[463];
    assign layer2_out[33] = ~(layer1_out[74] & layer1_out[75]);
    assign layer2_out[34] = layer1_out[398];
    assign layer2_out[35] = layer1_out[361];
    assign layer2_out[36] = ~layer1_out[30];
    assign layer2_out[37] = ~(layer1_out[204] & layer1_out[205]);
    assign layer2_out[38] = layer1_out[545];
    assign layer2_out[39] = ~layer1_out[487];
    assign layer2_out[40] = layer1_out[245];
    assign layer2_out[41] = ~(layer1_out[228] & layer1_out[229]);
    assign layer2_out[42] = ~layer1_out[451] | layer1_out[452];
    assign layer2_out[43] = ~layer1_out[235] | layer1_out[236];
    assign layer2_out[44] = ~layer1_out[207];
    assign layer2_out[45] = layer1_out[464];
    assign layer2_out[46] = layer1_out[400];
    assign layer2_out[47] = 1'b0;
    assign layer2_out[48] = layer1_out[412];
    assign layer2_out[49] = layer1_out[387] & ~layer1_out[386];
    assign layer2_out[50] = ~(layer1_out[489] & layer1_out[490]);
    assign layer2_out[51] = ~layer1_out[279];
    assign layer2_out[52] = layer1_out[307] & ~layer1_out[306];
    assign layer2_out[53] = ~layer1_out[509];
    assign layer2_out[54] = layer1_out[171];
    assign layer2_out[55] = layer1_out[385];
    assign layer2_out[56] = layer1_out[116];
    assign layer2_out[57] = layer1_out[352] & ~layer1_out[353];
    assign layer2_out[58] = layer1_out[145];
    assign layer2_out[59] = ~(layer1_out[119] & layer1_out[120]);
    assign layer2_out[60] = ~(layer1_out[32] & layer1_out[33]);
    assign layer2_out[61] = ~(layer1_out[528] | layer1_out[529]);
    assign layer2_out[62] = layer1_out[404];
    assign layer2_out[63] = ~layer1_out[515];
    assign layer2_out[64] = 1'b1;
    assign layer2_out[65] = ~layer1_out[232];
    assign layer2_out[66] = ~(layer1_out[508] & layer1_out[509]);
    assign layer2_out[67] = layer1_out[423] | layer1_out[424];
    assign layer2_out[68] = 1'b0;
    assign layer2_out[69] = 1'b0;
    assign layer2_out[70] = ~layer1_out[286];
    assign layer2_out[71] = ~layer1_out[398];
    assign layer2_out[72] = ~(layer1_out[152] & layer1_out[153]);
    assign layer2_out[73] = layer1_out[321];
    assign layer2_out[74] = layer1_out[146] & layer1_out[147];
    assign layer2_out[75] = layer1_out[331];
    assign layer2_out[76] = layer1_out[534];
    assign layer2_out[77] = layer1_out[450];
    assign layer2_out[78] = layer1_out[418];
    assign layer2_out[79] = layer1_out[467] & ~layer1_out[468];
    assign layer2_out[80] = layer1_out[540];
    assign layer2_out[81] = ~layer1_out[271] | layer1_out[272];
    assign layer2_out[82] = ~(layer1_out[159] & layer1_out[160]);
    assign layer2_out[83] = layer1_out[344];
    assign layer2_out[84] = layer1_out[113];
    assign layer2_out[85] = ~layer1_out[197];
    assign layer2_out[86] = ~(layer1_out[461] | layer1_out[462]);
    assign layer2_out[87] = layer1_out[88];
    assign layer2_out[88] = layer1_out[71] | layer1_out[72];
    assign layer2_out[89] = layer1_out[190];
    assign layer2_out[90] = ~layer1_out[110] | layer1_out[111];
    assign layer2_out[91] = layer1_out[185] | layer1_out[186];
    assign layer2_out[92] = layer1_out[255];
    assign layer2_out[93] = ~layer1_out[506];
    assign layer2_out[94] = layer1_out[438] & ~layer1_out[437];
    assign layer2_out[95] = ~layer1_out[188];
    assign layer2_out[96] = ~(layer1_out[430] & layer1_out[431]);
    assign layer2_out[97] = ~layer1_out[86];
    assign layer2_out[98] = ~layer1_out[137];
    assign layer2_out[99] = ~layer1_out[311] | layer1_out[312];
    assign layer2_out[100] = ~(layer1_out[268] & layer1_out[269]);
    assign layer2_out[101] = ~layer1_out[20] | layer1_out[21];
    assign layer2_out[102] = ~layer1_out[500];
    assign layer2_out[103] = layer1_out[369];
    assign layer2_out[104] = layer1_out[111];
    assign layer2_out[105] = layer1_out[359];
    assign layer2_out[106] = 1'b1;
    assign layer2_out[107] = layer1_out[17] ^ layer1_out[18];
    assign layer2_out[108] = 1'b1;
    assign layer2_out[109] = ~layer1_out[77] | layer1_out[78];
    assign layer2_out[110] = ~layer1_out[410] | layer1_out[411];
    assign layer2_out[111] = ~(layer1_out[322] | layer1_out[323]);
    assign layer2_out[112] = layer1_out[92];
    assign layer2_out[113] = ~layer1_out[319] | layer1_out[318];
    assign layer2_out[114] = 1'b0;
    assign layer2_out[115] = ~(layer1_out[545] & layer1_out[546]);
    assign layer2_out[116] = 1'b0;
    assign layer2_out[117] = layer1_out[57] & layer1_out[58];
    assign layer2_out[118] = layer1_out[213];
    assign layer2_out[119] = layer1_out[409] & ~layer1_out[410];
    assign layer2_out[120] = ~(layer1_out[394] & layer1_out[395]);
    assign layer2_out[121] = layer1_out[87];
    assign layer2_out[122] = ~layer1_out[71];
    assign layer2_out[123] = layer1_out[44];
    assign layer2_out[124] = ~layer1_out[143];
    assign layer2_out[125] = layer1_out[193];
    assign layer2_out[126] = 1'b1;
    assign layer2_out[127] = layer1_out[439] & ~layer1_out[440];
    assign layer2_out[128] = layer1_out[205] & ~layer1_out[206];
    assign layer2_out[129] = layer1_out[532] & layer1_out[533];
    assign layer2_out[130] = layer1_out[504] & ~layer1_out[505];
    assign layer2_out[131] = layer1_out[356];
    assign layer2_out[132] = layer1_out[536] & ~layer1_out[535];
    assign layer2_out[133] = ~layer1_out[135] | layer1_out[134];
    assign layer2_out[134] = layer1_out[409];
    assign layer2_out[135] = layer1_out[497] & ~layer1_out[498];
    assign layer2_out[136] = layer1_out[314];
    assign layer2_out[137] = ~(layer1_out[526] | layer1_out[527]);
    assign layer2_out[138] = layer1_out[215] & layer1_out[216];
    assign layer2_out[139] = layer1_out[14];
    assign layer2_out[140] = ~layer1_out[183];
    assign layer2_out[141] = ~layer1_out[445] | layer1_out[444];
    assign layer2_out[142] = layer1_out[419] & layer1_out[420];
    assign layer2_out[143] = ~layer1_out[140] | layer1_out[141];
    assign layer2_out[144] = ~(layer1_out[360] | layer1_out[361]);
    assign layer2_out[145] = layer1_out[518] & ~layer1_out[517];
    assign layer2_out[146] = 1'b0;
    assign layer2_out[147] = layer1_out[417];
    assign layer2_out[148] = layer1_out[209] & layer1_out[210];
    assign layer2_out[149] = layer1_out[310] & ~layer1_out[311];
    assign layer2_out[150] = layer1_out[339] & ~layer1_out[340];
    assign layer2_out[151] = layer1_out[276];
    assign layer2_out[152] = ~layer1_out[320] | layer1_out[319];
    assign layer2_out[153] = layer1_out[435];
    assign layer2_out[154] = ~layer1_out[519] | layer1_out[518];
    assign layer2_out[155] = layer1_out[101];
    assign layer2_out[156] = layer1_out[238] & ~layer1_out[237];
    assign layer2_out[157] = ~layer1_out[350] | layer1_out[351];
    assign layer2_out[158] = layer1_out[268] & ~layer1_out[267];
    assign layer2_out[159] = 1'b1;
    assign layer2_out[160] = 1'b1;
    assign layer2_out[161] = ~layer1_out[19];
    assign layer2_out[162] = layer1_out[468];
    assign layer2_out[163] = layer1_out[48] & layer1_out[49];
    assign layer2_out[164] = ~layer1_out[138];
    assign layer2_out[165] = ~layer1_out[350];
    assign layer2_out[166] = ~layer1_out[202] | layer1_out[203];
    assign layer2_out[167] = layer1_out[351];
    assign layer2_out[168] = layer1_out[77];
    assign layer2_out[169] = ~(layer1_out[370] | layer1_out[371]);
    assign layer2_out[170] = ~(layer1_out[82] & layer1_out[83]);
    assign layer2_out[171] = ~layer1_out[295] | layer1_out[294];
    assign layer2_out[172] = layer1_out[148] & ~layer1_out[147];
    assign layer2_out[173] = ~layer1_out[190] | layer1_out[191];
    assign layer2_out[174] = ~layer1_out[395] | layer1_out[396];
    assign layer2_out[175] = layer1_out[507];
    assign layer2_out[176] = ~(layer1_out[353] | layer1_out[354]);
    assign layer2_out[177] = ~layer1_out[62];
    assign layer2_out[178] = layer1_out[533];
    assign layer2_out[179] = layer1_out[392] & ~layer1_out[393];
    assign layer2_out[180] = layer1_out[131] | layer1_out[132];
    assign layer2_out[181] = layer1_out[367];
    assign layer2_out[182] = layer1_out[441] & ~layer1_out[442];
    assign layer2_out[183] = layer1_out[39] & ~layer1_out[40];
    assign layer2_out[184] = 1'b0;
    assign layer2_out[185] = ~(layer1_out[173] | layer1_out[174]);
    assign layer2_out[186] = layer1_out[333] & ~layer1_out[332];
    assign layer2_out[187] = ~layer1_out[542] | layer1_out[541];
    assign layer2_out[188] = 1'b0;
    assign layer2_out[189] = ~layer1_out[343];
    assign layer2_out[190] = layer1_out[19];
    assign layer2_out[191] = layer1_out[96];
    assign layer2_out[192] = ~layer1_out[248];
    assign layer2_out[193] = layer1_out[471];
    assign layer2_out[194] = layer1_out[294];
    assign layer2_out[195] = layer1_out[290];
    assign layer2_out[196] = layer1_out[444];
    assign layer2_out[197] = layer1_out[216] & ~layer1_out[217];
    assign layer2_out[198] = ~layer1_out[547];
    assign layer2_out[199] = layer1_out[503];
    assign layer2_out[200] = layer1_out[12] | layer1_out[13];
    assign layer2_out[201] = ~layer1_out[348];
    assign layer2_out[202] = ~layer1_out[302];
    assign layer2_out[203] = layer1_out[420];
    assign layer2_out[204] = ~(layer1_out[49] & layer1_out[50]);
    assign layer2_out[205] = layer1_out[336];
    assign layer2_out[206] = layer1_out[34] ^ layer1_out[35];
    assign layer2_out[207] = ~layer1_out[123];
    assign layer2_out[208] = layer1_out[329] & ~layer1_out[330];
    assign layer2_out[209] = ~layer1_out[182];
    assign layer2_out[210] = layer1_out[178] ^ layer1_out[179];
    assign layer2_out[211] = layer1_out[246] | layer1_out[247];
    assign layer2_out[212] = ~layer1_out[180];
    assign layer2_out[213] = layer1_out[117] | layer1_out[118];
    assign layer2_out[214] = layer1_out[35] & ~layer1_out[36];
    assign layer2_out[215] = layer1_out[422] & layer1_out[423];
    assign layer2_out[216] = ~(layer1_out[412] | layer1_out[413]);
    assign layer2_out[217] = 1'b1;
    assign layer2_out[218] = ~layer1_out[453];
    assign layer2_out[219] = layer1_out[479] & layer1_out[480];
    assign layer2_out[220] = layer1_out[4] ^ layer1_out[5];
    assign layer2_out[221] = layer1_out[305] | layer1_out[306];
    assign layer2_out[222] = layer1_out[148] ^ layer1_out[149];
    assign layer2_out[223] = ~(layer1_out[129] | layer1_out[130]);
    assign layer2_out[224] = layer1_out[121];
    assign layer2_out[225] = layer1_out[543] & layer1_out[544];
    assign layer2_out[226] = 1'b1;
    assign layer2_out[227] = ~layer1_out[455] | layer1_out[456];
    assign layer2_out[228] = layer1_out[150] | layer1_out[151];
    assign layer2_out[229] = ~layer1_out[312];
    assign layer2_out[230] = layer1_out[62];
    assign layer2_out[231] = ~(layer1_out[1] | layer1_out[2]);
    assign layer2_out[232] = 1'b0;
    assign layer2_out[233] = ~layer1_out[414];
    assign layer2_out[234] = layer1_out[527] | layer1_out[528];
    assign layer2_out[235] = 1'b1;
    assign layer2_out[236] = layer1_out[10] & layer1_out[11];
    assign layer2_out[237] = ~layer1_out[272];
    assign layer2_out[238] = ~(layer1_out[203] & layer1_out[204]);
    assign layer2_out[239] = layer1_out[524] & ~layer1_out[525];
    assign layer2_out[240] = layer1_out[446];
    assign layer2_out[241] = ~(layer1_out[547] | layer1_out[548]);
    assign layer2_out[242] = layer1_out[301];
    assign layer2_out[243] = layer1_out[110];
    assign layer2_out[244] = layer1_out[530];
    assign layer2_out[245] = ~layer1_out[258];
    assign layer2_out[246] = layer1_out[53] & ~layer1_out[52];
    assign layer2_out[247] = ~layer1_out[7];
    assign layer2_out[248] = ~(layer1_out[389] & layer1_out[390]);
    assign layer2_out[249] = 1'b0;
    assign layer2_out[250] = layer1_out[221];
    assign layer2_out[251] = layer1_out[153];
    assign layer2_out[252] = ~layer1_out[225];
    assign layer2_out[253] = layer1_out[363];
    assign layer2_out[254] = ~(layer1_out[257] | layer1_out[258]);
    assign layer2_out[255] = ~(layer1_out[36] | layer1_out[37]);
    assign layer2_out[256] = ~(layer1_out[105] | layer1_out[106]);
    assign layer2_out[257] = layer1_out[89] & layer1_out[90];
    assign layer2_out[258] = layer1_out[149] & ~layer1_out[150];
    assign layer2_out[259] = ~layer1_out[309] | layer1_out[308];
    assign layer2_out[260] = ~(layer1_out[21] | layer1_out[22]);
    assign layer2_out[261] = layer1_out[267] & ~layer1_out[266];
    assign layer2_out[262] = 1'b1;
    assign layer2_out[263] = 1'b1;
    assign layer2_out[264] = layer1_out[382] & layer1_out[383];
    assign layer2_out[265] = ~layer1_out[200];
    assign layer2_out[266] = layer1_out[63] & ~layer1_out[64];
    assign layer2_out[267] = layer1_out[40] | layer1_out[41];
    assign layer2_out[268] = 1'b0;
    assign layer2_out[269] = layer1_out[73] & ~layer1_out[72];
    assign layer2_out[270] = ~layer1_out[194];
    assign layer2_out[271] = ~layer1_out[437];
    assign layer2_out[272] = ~layer1_out[471];
    assign layer2_out[273] = layer1_out[154];
    assign layer2_out[274] = ~(layer1_out[201] & layer1_out[202]);
    assign layer2_out[275] = layer1_out[478];
    assign layer2_out[276] = 1'b0;
    assign layer2_out[277] = ~(layer1_out[261] & layer1_out[262]);
    assign layer2_out[278] = layer1_out[473] & ~layer1_out[472];
    assign layer2_out[279] = 1'b1;
    assign layer2_out[280] = layer1_out[199] & layer1_out[200];
    assign layer2_out[281] = ~layer1_out[522] | layer1_out[523];
    assign layer2_out[282] = ~layer1_out[240];
    assign layer2_out[283] = layer1_out[438] | layer1_out[439];
    assign layer2_out[284] = layer1_out[449] & ~layer1_out[448];
    assign layer2_out[285] = layer1_out[14];
    assign layer2_out[286] = layer1_out[517] & ~layer1_out[516];
    assign layer2_out[287] = ~(layer1_out[73] | layer1_out[74]);
    assign layer2_out[288] = ~layer1_out[298] | layer1_out[297];
    assign layer2_out[289] = ~layer1_out[156] | layer1_out[155];
    assign layer2_out[290] = ~layer1_out[443];
    assign layer2_out[291] = layer1_out[512];
    assign layer2_out[292] = layer1_out[28];
    assign layer2_out[293] = ~layer1_out[349] | layer1_out[348];
    assign layer2_out[294] = ~layer1_out[454] | layer1_out[455];
    assign layer2_out[295] = layer1_out[482] | layer1_out[483];
    assign layer2_out[296] = ~layer1_out[368];
    assign layer2_out[297] = layer1_out[304];
    assign layer2_out[298] = layer1_out[210] & ~layer1_out[211];
    assign layer2_out[299] = ~layer1_out[167] | layer1_out[168];
    assign layer2_out[300] = ~layer1_out[45];
    assign layer2_out[301] = layer1_out[406];
    assign layer2_out[302] = 1'b0;
    assign layer2_out[303] = ~(layer1_out[230] | layer1_out[231]);
    assign layer2_out[304] = layer1_out[287];
    assign layer2_out[305] = ~layer1_out[79];
    assign layer2_out[306] = layer1_out[415];
    assign layer2_out[307] = layer1_out[276];
    assign layer2_out[308] = ~(layer1_out[50] | layer1_out[51]);
    assign layer2_out[309] = ~layer1_out[477];
    assign layer2_out[310] = ~layer1_out[1];
    assign layer2_out[311] = ~(layer1_out[396] & layer1_out[397]);
    assign layer2_out[312] = ~layer1_out[8] | layer1_out[7];
    assign layer2_out[313] = layer1_out[263] & layer1_out[264];
    assign layer2_out[314] = layer1_out[102] & ~layer1_out[103];
    assign layer2_out[315] = layer1_out[186];
    assign layer2_out[316] = ~(layer1_out[379] | layer1_out[380]);
    assign layer2_out[317] = ~(layer1_out[354] | layer1_out[355]);
    assign layer2_out[318] = ~layer1_out[454] | layer1_out[453];
    assign layer2_out[319] = ~(layer1_out[23] | layer1_out[24]);
    assign layer2_out[320] = ~layer1_out[278];
    assign layer2_out[321] = ~layer1_out[142];
    assign layer2_out[322] = ~(layer1_out[177] | layer1_out[178]);
    assign layer2_out[323] = 1'b1;
    assign layer2_out[324] = ~(layer1_out[372] | layer1_out[373]);
    assign layer2_out[325] = ~layer1_out[338];
    assign layer2_out[326] = layer1_out[274] & ~layer1_out[273];
    assign layer2_out[327] = ~layer1_out[520];
    assign layer2_out[328] = ~layer1_out[192];
    assign layer2_out[329] = layer1_out[75] | layer1_out[76];
    assign layer2_out[330] = ~layer1_out[70];
    assign layer2_out[331] = layer1_out[54] & ~layer1_out[53];
    assign layer2_out[332] = 1'b0;
    assign layer2_out[333] = ~(layer1_out[274] & layer1_out[275]);
    assign layer2_out[334] = 1'b0;
    assign layer2_out[335] = layer1_out[256] & layer1_out[257];
    assign layer2_out[336] = ~layer1_out[483];
    assign layer2_out[337] = ~layer1_out[132] | layer1_out[133];
    assign layer2_out[338] = layer1_out[161];
    assign layer2_out[339] = layer1_out[413];
    assign layer2_out[340] = ~layer1_out[152] | layer1_out[151];
    assign layer2_out[341] = ~layer1_out[526];
    assign layer2_out[342] = 1'b1;
    assign layer2_out[343] = layer1_out[298];
    assign layer2_out[344] = ~layer1_out[94];
    assign layer2_out[345] = layer1_out[22] ^ layer1_out[23];
    assign layer2_out[346] = layer1_out[183] | layer1_out[184];
    assign layer2_out[347] = ~layer1_out[357] | layer1_out[358];
    assign layer2_out[348] = layer1_out[163] & ~layer1_out[162];
    assign layer2_out[349] = ~layer1_out[299] | layer1_out[300];
    assign layer2_out[350] = ~(layer1_out[168] | layer1_out[169]);
    assign layer2_out[351] = ~layer1_out[161];
    assign layer2_out[352] = 1'b1;
    assign layer2_out[353] = 1'b1;
    assign layer2_out[354] = layer1_out[94];
    assign layer2_out[355] = layer1_out[128];
    assign layer2_out[356] = ~(layer1_out[5] | layer1_out[6]);
    assign layer2_out[357] = ~(layer1_out[56] | layer1_out[57]);
    assign layer2_out[358] = ~layer1_out[66] | layer1_out[67];
    assign layer2_out[359] = layer1_out[341] & ~layer1_out[340];
    assign layer2_out[360] = ~layer1_out[281];
    assign layer2_out[361] = layer1_out[496];
    assign layer2_out[362] = 1'b1;
    assign layer2_out[363] = layer1_out[324];
    assign layer2_out[364] = 1'b1;
    assign layer2_out[365] = ~layer1_out[385];
    assign layer2_out[366] = ~layer1_out[457];
    assign layer2_out[367] = ~(layer1_out[231] & layer1_out[232]);
    assign layer2_out[368] = 1'b1;
    assign layer2_out[369] = layer1_out[296] | layer1_out[297];
    assign layer2_out[370] = layer1_out[255] & layer1_out[256];
    assign layer2_out[371] = ~layer1_out[450] | layer1_out[449];
    assign layer2_out[372] = ~layer1_out[42] | layer1_out[43];
    assign layer2_out[373] = layer1_out[403];
    assign layer2_out[374] = ~layer1_out[401];
    assign layer2_out[375] = ~layer1_out[363] | layer1_out[362];
    assign layer2_out[376] = ~layer1_out[109] | layer1_out[108];
    assign layer2_out[377] = layer1_out[288] | layer1_out[289];
    assign layer2_out[378] = layer1_out[494];
    assign layer2_out[379] = layer1_out[523] | layer1_out[524];
    assign layer2_out[380] = ~layer1_out[131] | layer1_out[130];
    assign layer2_out[381] = layer1_out[15] | layer1_out[16];
    assign layer2_out[382] = layer1_out[250];
    assign layer2_out[383] = layer1_out[52];
    assign layer2_out[384] = layer1_out[211] & layer1_out[212];
    assign layer2_out[385] = layer1_out[499] & ~layer1_out[500];
    assign layer2_out[386] = ~(layer1_out[38] & layer1_out[39]);
    assign layer2_out[387] = layer1_out[364] & layer1_out[365];
    assign layer2_out[388] = layer1_out[188] & ~layer1_out[189];
    assign layer2_out[389] = ~(layer1_out[529] & layer1_out[530]);
    assign layer2_out[390] = ~layer1_out[440];
    assign layer2_out[391] = layer1_out[387];
    assign layer2_out[392] = layer1_out[114] & ~layer1_out[115];
    assign layer2_out[393] = layer1_out[496];
    assign layer2_out[394] = ~(layer1_out[219] | layer1_out[220]);
    assign layer2_out[395] = layer1_out[251];
    assign layer2_out[396] = ~layer1_out[247];
    assign layer2_out[397] = ~layer1_out[508] | layer1_out[507];
    assign layer2_out[398] = layer1_out[33] | layer1_out[34];
    assign layer2_out[399] = ~layer1_out[372] | layer1_out[371];
    assign layer2_out[400] = ~layer1_out[66] | layer1_out[65];
    assign layer2_out[401] = ~layer1_out[209];
    assign layer2_out[402] = 1'b0;
    assign layer2_out[403] = layer1_out[99] & ~layer1_out[100];
    assign layer2_out[404] = layer1_out[338];
    assign layer2_out[405] = ~(layer1_out[163] | layer1_out[164]);
    assign layer2_out[406] = ~layer1_out[79] | layer1_out[78];
    assign layer2_out[407] = 1'b0;
    assign layer2_out[408] = layer1_out[433];
    assign layer2_out[409] = layer1_out[212];
    assign layer2_out[410] = layer1_out[491];
    assign layer2_out[411] = ~layer1_out[271] | layer1_out[270];
    assign layer2_out[412] = layer1_out[69];
    assign layer2_out[413] = ~layer1_out[236];
    assign layer2_out[414] = ~layer1_out[392];
    assign layer2_out[415] = layer1_out[265];
    assign layer2_out[416] = ~layer1_out[333];
    assign layer2_out[417] = ~layer1_out[315] | layer1_out[316];
    assign layer2_out[418] = ~layer1_out[233];
    assign layer2_out[419] = layer1_out[490] | layer1_out[491];
    assign layer2_out[420] = ~layer1_out[48];
    assign layer2_out[421] = ~(layer1_out[277] & layer1_out[278]);
    assign layer2_out[422] = ~layer1_out[502];
    assign layer2_out[423] = layer1_out[430] & ~layer1_out[429];
    assign layer2_out[424] = ~layer1_out[261];
    assign layer2_out[425] = layer1_out[406];
    assign layer2_out[426] = ~layer1_out[485] | layer1_out[484];
    assign layer2_out[427] = ~layer1_out[379];
    assign layer2_out[428] = ~layer1_out[520];
    assign layer2_out[429] = layer1_out[303] & ~layer1_out[304];
    assign layer2_out[430] = ~layer1_out[374];
    assign layer2_out[431] = ~layer1_out[301];
    assign layer2_out[432] = ~(layer1_out[316] | layer1_out[317]);
    assign layer2_out[433] = ~(layer1_out[381] & layer1_out[382]);
    assign layer2_out[434] = ~layer1_out[541];
    assign layer2_out[435] = layer1_out[548] & layer1_out[549];
    assign layer2_out[436] = layer1_out[47] & ~layer1_out[46];
    assign layer2_out[437] = ~(layer1_out[3] ^ layer1_out[4]);
    assign layer2_out[438] = ~layer1_out[433];
    assign layer2_out[439] = ~layer1_out[428];
    assign layer2_out[440] = ~(layer1_out[465] | layer1_out[466]);
    assign layer2_out[441] = layer1_out[475];
    assign layer2_out[442] = ~(layer1_out[375] | layer1_out[376]);
    assign layer2_out[443] = layer1_out[313];
    assign layer2_out[444] = layer1_out[242];
    assign layer2_out[445] = 1'b1;
    assign layer2_out[446] = layer1_out[432] & ~layer1_out[431];
    assign layer2_out[447] = ~layer1_out[476] | layer1_out[477];
    assign layer2_out[448] = ~layer1_out[159];
    assign layer2_out[449] = ~layer1_out[81];
    assign layer2_out[450] = ~layer1_out[245];
    assign layer2_out[451] = ~layer1_out[31];
    assign layer2_out[452] = ~layer1_out[228] | layer1_out[227];
    assign layer2_out[453] = ~(layer1_out[521] | layer1_out[522]);
    assign layer2_out[454] = ~layer1_out[136];
    assign layer2_out[455] = layer1_out[90] & ~layer1_out[91];
    assign layer2_out[456] = layer1_out[243];
    assign layer2_out[457] = ~(layer1_out[106] | layer1_out[107]);
    assign layer2_out[458] = layer1_out[380] | layer1_out[381];
    assign layer2_out[459] = layer1_out[84];
    assign layer2_out[460] = layer1_out[125];
    assign layer2_out[461] = layer1_out[265] & ~layer1_out[266];
    assign layer2_out[462] = layer1_out[408];
    assign layer2_out[463] = layer1_out[428];
    assign layer2_out[464] = 1'b1;
    assign layer2_out[465] = layer1_out[269] & ~layer1_out[270];
    assign layer2_out[466] = ~layer1_out[55] | layer1_out[56];
    assign layer2_out[467] = ~layer1_out[331];
    assign layer2_out[468] = ~layer1_out[470];
    assign layer2_out[469] = ~layer1_out[288];
    assign layer2_out[470] = ~(layer1_out[404] | layer1_out[405]);
    assign layer2_out[471] = layer1_out[80];
    assign layer2_out[472] = layer1_out[328];
    assign layer2_out[473] = ~(layer1_out[121] | layer1_out[122]);
    assign layer2_out[474] = layer1_out[388] & ~layer1_out[389];
    assign layer2_out[475] = ~layer1_out[481];
    assign layer2_out[476] = layer1_out[458] & layer1_out[459];
    assign layer2_out[477] = ~layer1_out[424];
    assign layer2_out[478] = layer1_out[166] | layer1_out[167];
    assign layer2_out[479] = 1'b0;
    assign layer2_out[480] = ~layer1_out[244] | layer1_out[243];
    assign layer2_out[481] = layer1_out[511] & ~layer1_out[510];
    assign layer2_out[482] = layer1_out[356] & ~layer1_out[357];
    assign layer2_out[483] = ~(layer1_out[374] | layer1_out[375]);
    assign layer2_out[484] = 1'b0;
    assign layer2_out[485] = layer1_out[346];
    assign layer2_out[486] = ~layer1_out[222];
    assign layer2_out[487] = layer1_out[292];
    assign layer2_out[488] = ~layer1_out[169] | layer1_out[170];
    assign layer2_out[489] = ~layer1_out[252];
    assign layer2_out[490] = ~layer1_out[335];
    assign layer2_out[491] = ~(layer1_out[317] & layer1_out[318]);
    assign layer2_out[492] = ~layer1_out[143];
    assign layer2_out[493] = layer1_out[41] & ~layer1_out[42];
    assign layer2_out[494] = layer1_out[105];
    assign layer2_out[495] = ~layer1_out[481];
    assign layer2_out[496] = layer1_out[487];
    assign layer2_out[497] = ~(layer1_out[474] & layer1_out[475]);
    assign layer2_out[498] = layer1_out[369];
    assign layer2_out[499] = ~layer1_out[474] | layer1_out[473];
    assign layer2_out[500] = layer1_out[176];
    assign layer2_out[501] = layer1_out[116];
    assign layer2_out[502] = layer1_out[417];
    assign layer2_out[503] = layer1_out[513] & ~layer1_out[514];
    assign layer2_out[504] = layer1_out[531] & layer1_out[532];
    assign layer2_out[505] = ~(layer1_out[192] & layer1_out[193]);
    assign layer2_out[506] = layer1_out[133] | layer1_out[134];
    assign layer2_out[507] = 1'b0;
    assign layer2_out[508] = layer1_out[320] & ~layer1_out[321];
    assign layer2_out[509] = ~(layer1_out[259] & layer1_out[260]);
    assign layer2_out[510] = 1'b1;
    assign layer2_out[511] = layer1_out[2];
    assign layer2_out[512] = layer1_out[123] | layer1_out[124];
    assign layer2_out[513] = ~layer1_out[515];
    assign layer2_out[514] = 1'b1;
    assign layer2_out[515] = ~layer1_out[445] | layer1_out[446];
    assign layer2_out[516] = ~layer1_out[253];
    assign layer2_out[517] = ~layer1_out[176];
    assign layer2_out[518] = layer1_out[466];
    assign layer2_out[519] = layer1_out[538];
    assign layer2_out[520] = ~(layer1_out[498] & layer1_out[499]);
    assign layer2_out[521] = layer1_out[360] & ~layer1_out[359];
    assign layer2_out[522] = ~layer1_out[456];
    assign layer2_out[523] = layer1_out[262] & layer1_out[263];
    assign layer2_out[524] = layer1_out[64] & ~layer1_out[65];
    assign layer2_out[525] = layer1_out[325] & ~layer1_out[326];
    assign layer2_out[526] = layer1_out[226];
    assign layer2_out[527] = layer1_out[98] & ~layer1_out[97];
    assign layer2_out[528] = layer1_out[425] & layer1_out[426];
    assign layer2_out[529] = ~(layer1_out[281] | layer1_out[282]);
    assign layer2_out[530] = layer1_out[156] ^ layer1_out[157];
    assign layer2_out[531] = layer1_out[59] ^ layer1_out[60];
    assign layer2_out[532] = layer1_out[377];
    assign layer2_out[533] = layer1_out[390] | layer1_out[391];
    assign layer2_out[534] = layer1_out[112];
    assign layer2_out[535] = ~layer1_out[218] | layer1_out[219];
    assign layer2_out[536] = layer1_out[537] & ~layer1_out[536];
    assign layer2_out[537] = layer1_out[224];
    assign layer2_out[538] = ~layer1_out[435];
    assign layer2_out[539] = layer1_out[198] & ~layer1_out[199];
    assign layer2_out[540] = ~(layer1_out[16] | layer1_out[17]);
    assign layer2_out[541] = ~layer1_out[538];
    assign layer2_out[542] = 1'b1;
    assign layer2_out[543] = layer1_out[166];
    assign layer2_out[544] = ~layer1_out[164];
    assign layer2_out[545] = ~(layer1_out[137] & layer1_out[138]);
    assign layer2_out[546] = ~(layer1_out[365] | layer1_out[366]);
    assign layer2_out[547] = ~layer1_out[0] | layer1_out[2];
    assign layer2_out[548] = layer1_out[328];
    assign layer2_out[549] = ~layer1_out[462];
    assign layer3_out[0] = layer2_out[446];
    assign layer3_out[1] = ~layer2_out[138] | layer2_out[139];
    assign layer3_out[2] = layer2_out[378] & ~layer2_out[379];
    assign layer3_out[3] = ~layer2_out[157] | layer2_out[156];
    assign layer3_out[4] = layer2_out[89] & ~layer2_out[88];
    assign layer3_out[5] = ~layer2_out[212];
    assign layer3_out[6] = layer2_out[425] & layer2_out[426];
    assign layer3_out[7] = layer2_out[317];
    assign layer3_out[8] = layer2_out[375] & layer2_out[376];
    assign layer3_out[9] = ~layer2_out[372];
    assign layer3_out[10] = layer2_out[444] & ~layer2_out[445];
    assign layer3_out[11] = ~layer2_out[341];
    assign layer3_out[12] = layer2_out[368] ^ layer2_out[369];
    assign layer3_out[13] = ~layer2_out[172];
    assign layer3_out[14] = ~(layer2_out[46] ^ layer2_out[47]);
    assign layer3_out[15] = ~layer2_out[536];
    assign layer3_out[16] = layer2_out[94];
    assign layer3_out[17] = layer2_out[332];
    assign layer3_out[18] = layer2_out[71] & ~layer2_out[72];
    assign layer3_out[19] = ~(layer2_out[189] & layer2_out[190]);
    assign layer3_out[20] = ~layer2_out[149];
    assign layer3_out[21] = layer2_out[545] | layer2_out[546];
    assign layer3_out[22] = ~layer2_out[348];
    assign layer3_out[23] = layer2_out[529] & layer2_out[530];
    assign layer3_out[24] = layer2_out[236] | layer2_out[237];
    assign layer3_out[25] = layer2_out[408];
    assign layer3_out[26] = ~layer2_out[462] | layer2_out[463];
    assign layer3_out[27] = 1'b0;
    assign layer3_out[28] = ~(layer2_out[192] | layer2_out[193]);
    assign layer3_out[29] = layer2_out[13];
    assign layer3_out[30] = layer2_out[413];
    assign layer3_out[31] = ~layer2_out[515];
    assign layer3_out[32] = ~layer2_out[287] | layer2_out[288];
    assign layer3_out[33] = ~layer2_out[4];
    assign layer3_out[34] = ~layer2_out[18] | layer2_out[17];
    assign layer3_out[35] = ~layer2_out[343];
    assign layer3_out[36] = layer2_out[521] & layer2_out[522];
    assign layer3_out[37] = ~(layer2_out[515] & layer2_out[516]);
    assign layer3_out[38] = ~layer2_out[141] | layer2_out[140];
    assign layer3_out[39] = layer2_out[241];
    assign layer3_out[40] = ~layer2_out[253];
    assign layer3_out[41] = layer2_out[382];
    assign layer3_out[42] = ~(layer2_out[533] | layer2_out[534]);
    assign layer3_out[43] = ~(layer2_out[260] ^ layer2_out[261]);
    assign layer3_out[44] = ~(layer2_out[415] & layer2_out[416]);
    assign layer3_out[45] = ~layer2_out[527];
    assign layer3_out[46] = ~layer2_out[466] | layer2_out[467];
    assign layer3_out[47] = layer2_out[106];
    assign layer3_out[48] = layer2_out[533];
    assign layer3_out[49] = ~layer2_out[365];
    assign layer3_out[50] = ~layer2_out[96];
    assign layer3_out[51] = ~(layer2_out[383] | layer2_out[384]);
    assign layer3_out[52] = layer2_out[236];
    assign layer3_out[53] = ~(layer2_out[128] & layer2_out[129]);
    assign layer3_out[54] = 1'b0;
    assign layer3_out[55] = 1'b0;
    assign layer3_out[56] = layer2_out[217];
    assign layer3_out[57] = ~layer2_out[263];
    assign layer3_out[58] = ~(layer2_out[430] & layer2_out[431]);
    assign layer3_out[59] = layer2_out[483];
    assign layer3_out[60] = ~(layer2_out[337] | layer2_out[338]);
    assign layer3_out[61] = layer2_out[321];
    assign layer3_out[62] = layer2_out[0];
    assign layer3_out[63] = layer2_out[220] & layer2_out[221];
    assign layer3_out[64] = layer2_out[341];
    assign layer3_out[65] = ~(layer2_out[534] | layer2_out[535]);
    assign layer3_out[66] = layer2_out[177] & layer2_out[178];
    assign layer3_out[67] = layer2_out[20] & layer2_out[21];
    assign layer3_out[68] = layer2_out[108];
    assign layer3_out[69] = layer2_out[200] & ~layer2_out[199];
    assign layer3_out[70] = ~layer2_out[526] | layer2_out[527];
    assign layer3_out[71] = ~(layer2_out[110] | layer2_out[111]);
    assign layer3_out[72] = ~layer2_out[477];
    assign layer3_out[73] = 1'b1;
    assign layer3_out[74] = layer2_out[377] & layer2_out[378];
    assign layer3_out[75] = layer2_out[496] & layer2_out[497];
    assign layer3_out[76] = layer2_out[384] | layer2_out[385];
    assign layer3_out[77] = layer2_out[274];
    assign layer3_out[78] = ~layer2_out[213] | layer2_out[214];
    assign layer3_out[79] = ~layer2_out[202];
    assign layer3_out[80] = ~layer2_out[275];
    assign layer3_out[81] = layer2_out[277] ^ layer2_out[278];
    assign layer3_out[82] = ~(layer2_out[525] | layer2_out[526]);
    assign layer3_out[83] = layer2_out[82] & layer2_out[83];
    assign layer3_out[84] = layer2_out[544];
    assign layer3_out[85] = layer2_out[264] & ~layer2_out[265];
    assign layer3_out[86] = layer2_out[441];
    assign layer3_out[87] = layer2_out[53];
    assign layer3_out[88] = layer2_out[66] & ~layer2_out[65];
    assign layer3_out[89] = layer2_out[73] | layer2_out[74];
    assign layer3_out[90] = ~layer2_out[206];
    assign layer3_out[91] = ~(layer2_out[271] & layer2_out[272]);
    assign layer3_out[92] = ~(layer2_out[539] | layer2_out[540]);
    assign layer3_out[93] = ~layer2_out[277];
    assign layer3_out[94] = ~layer2_out[216];
    assign layer3_out[95] = layer2_out[26] & ~layer2_out[27];
    assign layer3_out[96] = layer2_out[127];
    assign layer3_out[97] = ~layer2_out[485];
    assign layer3_out[98] = ~(layer2_out[7] | layer2_out[8]);
    assign layer3_out[99] = ~layer2_out[319];
    assign layer3_out[100] = 1'b1;
    assign layer3_out[101] = layer2_out[60] & ~layer2_out[61];
    assign layer3_out[102] = ~(layer2_out[142] & layer2_out[143]);
    assign layer3_out[103] = ~(layer2_out[315] | layer2_out[316]);
    assign layer3_out[104] = ~layer2_out[126] | layer2_out[125];
    assign layer3_out[105] = ~layer2_out[223];
    assign layer3_out[106] = layer2_out[406];
    assign layer3_out[107] = layer2_out[43] & ~layer2_out[44];
    assign layer3_out[108] = ~layer2_out[25];
    assign layer3_out[109] = ~layer2_out[325] | layer2_out[326];
    assign layer3_out[110] = ~layer2_out[362] | layer2_out[363];
    assign layer3_out[111] = layer2_out[87] & layer2_out[88];
    assign layer3_out[112] = layer2_out[508] & ~layer2_out[509];
    assign layer3_out[113] = ~(layer2_out[122] & layer2_out[123]);
    assign layer3_out[114] = layer2_out[405];
    assign layer3_out[115] = ~layer2_out[198];
    assign layer3_out[116] = 1'b0;
    assign layer3_out[117] = ~layer2_out[439];
    assign layer3_out[118] = layer2_out[41] & layer2_out[42];
    assign layer3_out[119] = ~layer2_out[438];
    assign layer3_out[120] = ~layer2_out[475];
    assign layer3_out[121] = ~layer2_out[66] | layer2_out[67];
    assign layer3_out[122] = ~layer2_out[447];
    assign layer3_out[123] = ~(layer2_out[442] ^ layer2_out[443]);
    assign layer3_out[124] = ~layer2_out[75];
    assign layer3_out[125] = ~layer2_out[91];
    assign layer3_out[126] = 1'b0;
    assign layer3_out[127] = layer2_out[311];
    assign layer3_out[128] = ~layer2_out[336];
    assign layer3_out[129] = ~layer2_out[7];
    assign layer3_out[130] = ~layer2_out[461] | layer2_out[462];
    assign layer3_out[131] = layer2_out[272] | layer2_out[273];
    assign layer3_out[132] = layer2_out[186];
    assign layer3_out[133] = layer2_out[547] & layer2_out[548];
    assign layer3_out[134] = ~layer2_out[501];
    assign layer3_out[135] = ~layer2_out[233] | layer2_out[234];
    assign layer3_out[136] = ~(layer2_out[360] | layer2_out[361]);
    assign layer3_out[137] = layer2_out[180];
    assign layer3_out[138] = layer2_out[240];
    assign layer3_out[139] = ~layer2_out[419];
    assign layer3_out[140] = ~layer2_out[29];
    assign layer3_out[141] = ~layer2_out[215];
    assign layer3_out[142] = layer2_out[464] & layer2_out[465];
    assign layer3_out[143] = 1'b0;
    assign layer3_out[144] = layer2_out[5] | layer2_out[6];
    assign layer3_out[145] = layer2_out[513] & layer2_out[514];
    assign layer3_out[146] = ~(layer2_out[279] | layer2_out[280]);
    assign layer3_out[147] = layer2_out[3];
    assign layer3_out[148] = ~layer2_out[2] | layer2_out[3];
    assign layer3_out[149] = ~layer2_out[266] | layer2_out[267];
    assign layer3_out[150] = ~layer2_out[247];
    assign layer3_out[151] = layer2_out[70] & layer2_out[71];
    assign layer3_out[152] = layer2_out[356] & layer2_out[357];
    assign layer3_out[153] = ~layer2_out[469] | layer2_out[470];
    assign layer3_out[154] = layer2_out[38];
    assign layer3_out[155] = ~(layer2_out[1] & layer2_out[2]);
    assign layer3_out[156] = ~(layer2_out[159] ^ layer2_out[160]);
    assign layer3_out[157] = ~layer2_out[518];
    assign layer3_out[158] = layer2_out[338];
    assign layer3_out[159] = ~layer2_out[218] | layer2_out[219];
    assign layer3_out[160] = layer2_out[156] & ~layer2_out[155];
    assign layer3_out[161] = ~layer2_out[175];
    assign layer3_out[162] = layer2_out[25];
    assign layer3_out[163] = layer2_out[122] & ~layer2_out[121];
    assign layer3_out[164] = layer2_out[154] & ~layer2_out[155];
    assign layer3_out[165] = ~layer2_out[374] | layer2_out[375];
    assign layer3_out[166] = ~layer2_out[263];
    assign layer3_out[167] = layer2_out[460];
    assign layer3_out[168] = layer2_out[490] & layer2_out[491];
    assign layer3_out[169] = layer2_out[229] ^ layer2_out[230];
    assign layer3_out[170] = ~layer2_out[285] | layer2_out[286];
    assign layer3_out[171] = ~(layer2_out[12] | layer2_out[13]);
    assign layer3_out[172] = layer2_out[169];
    assign layer3_out[173] = layer2_out[425] & ~layer2_out[424];
    assign layer3_out[174] = ~(layer2_out[173] | layer2_out[174]);
    assign layer3_out[175] = ~layer2_out[491] | layer2_out[492];
    assign layer3_out[176] = layer2_out[428];
    assign layer3_out[177] = ~layer2_out[454] | layer2_out[453];
    assign layer3_out[178] = layer2_out[439] & layer2_out[440];
    assign layer3_out[179] = ~layer2_out[240] | layer2_out[239];
    assign layer3_out[180] = layer2_out[59];
    assign layer3_out[181] = layer2_out[306];
    assign layer3_out[182] = ~layer2_out[311];
    assign layer3_out[183] = layer2_out[313];
    assign layer3_out[184] = layer2_out[499] & layer2_out[500];
    assign layer3_out[185] = layer2_out[90];
    assign layer3_out[186] = ~(layer2_out[296] | layer2_out[297]);
    assign layer3_out[187] = ~layer2_out[248];
    assign layer3_out[188] = layer2_out[80];
    assign layer3_out[189] = layer2_out[256] & ~layer2_out[255];
    assign layer3_out[190] = ~layer2_out[511];
    assign layer3_out[191] = ~(layer2_out[398] & layer2_out[399]);
    assign layer3_out[192] = ~layer2_out[117];
    assign layer3_out[193] = ~layer2_out[83] | layer2_out[84];
    assign layer3_out[194] = layer2_out[97] & layer2_out[98];
    assign layer3_out[195] = ~layer2_out[280];
    assign layer3_out[196] = ~layer2_out[400] | layer2_out[399];
    assign layer3_out[197] = layer2_out[393] & layer2_out[394];
    assign layer3_out[198] = layer2_out[126] & layer2_out[127];
    assign layer3_out[199] = ~(layer2_out[144] | layer2_out[145]);
    assign layer3_out[200] = ~(layer2_out[30] & layer2_out[31]);
    assign layer3_out[201] = 1'b1;
    assign layer3_out[202] = ~(layer2_out[143] | layer2_out[144]);
    assign layer3_out[203] = ~(layer2_out[157] | layer2_out[158]);
    assign layer3_out[204] = ~layer2_out[113];
    assign layer3_out[205] = ~layer2_out[58] | layer2_out[59];
    assign layer3_out[206] = ~layer2_out[209] | layer2_out[210];
    assign layer3_out[207] = layer2_out[134];
    assign layer3_out[208] = layer2_out[392] | layer2_out[393];
    assign layer3_out[209] = layer2_out[299];
    assign layer3_out[210] = layer2_out[543];
    assign layer3_out[211] = 1'b1;
    assign layer3_out[212] = layer2_out[470] | layer2_out[471];
    assign layer3_out[213] = ~(layer2_out[74] ^ layer2_out[75]);
    assign layer3_out[214] = ~layer2_out[141];
    assign layer3_out[215] = layer2_out[195] | layer2_out[196];
    assign layer3_out[216] = ~layer2_out[361];
    assign layer3_out[217] = ~(layer2_out[8] ^ layer2_out[9]);
    assign layer3_out[218] = ~layer2_out[254] | layer2_out[255];
    assign layer3_out[219] = ~layer2_out[92];
    assign layer3_out[220] = layer2_out[226];
    assign layer3_out[221] = ~layer2_out[108];
    assign layer3_out[222] = ~layer2_out[390];
    assign layer3_out[223] = ~layer2_out[50] | layer2_out[49];
    assign layer3_out[224] = ~layer2_out[256] | layer2_out[257];
    assign layer3_out[225] = ~layer2_out[279];
    assign layer3_out[226] = layer2_out[531];
    assign layer3_out[227] = ~layer2_out[180];
    assign layer3_out[228] = layer2_out[190];
    assign layer3_out[229] = layer2_out[19] ^ layer2_out[20];
    assign layer3_out[230] = ~layer2_out[145];
    assign layer3_out[231] = ~layer2_out[309] | layer2_out[308];
    assign layer3_out[232] = layer2_out[63];
    assign layer3_out[233] = layer2_out[293] & layer2_out[294];
    assign layer3_out[234] = layer2_out[163];
    assign layer3_out[235] = ~layer2_out[165] | layer2_out[164];
    assign layer3_out[236] = ~layer2_out[51];
    assign layer3_out[237] = ~layer2_out[208] | layer2_out[209];
    assign layer3_out[238] = ~layer2_out[115];
    assign layer3_out[239] = layer2_out[251];
    assign layer3_out[240] = layer2_out[45];
    assign layer3_out[241] = ~(layer2_out[302] & layer2_out[303]);
    assign layer3_out[242] = ~layer2_out[390];
    assign layer3_out[243] = ~layer2_out[284] | layer2_out[285];
    assign layer3_out[244] = ~(layer2_out[36] & layer2_out[37]);
    assign layer3_out[245] = layer2_out[250];
    assign layer3_out[246] = layer2_out[321];
    assign layer3_out[247] = ~(layer2_out[345] & layer2_out[346]);
    assign layer3_out[248] = ~(layer2_out[15] ^ layer2_out[16]);
    assign layer3_out[249] = ~(layer2_out[152] & layer2_out[153]);
    assign layer3_out[250] = 1'b1;
    assign layer3_out[251] = layer2_out[505] & ~layer2_out[504];
    assign layer3_out[252] = ~(layer2_out[147] ^ layer2_out[148]);
    assign layer3_out[253] = layer2_out[414];
    assign layer3_out[254] = layer2_out[15] & ~layer2_out[14];
    assign layer3_out[255] = layer2_out[168] & ~layer2_out[167];
    assign layer3_out[256] = ~layer2_out[472];
    assign layer3_out[257] = 1'b0;
    assign layer3_out[258] = ~layer2_out[420];
    assign layer3_out[259] = ~layer2_out[21];
    assign layer3_out[260] = ~(layer2_out[406] & layer2_out[407]);
    assign layer3_out[261] = ~(layer2_out[224] ^ layer2_out[225]);
    assign layer3_out[262] = ~layer2_out[290];
    assign layer3_out[263] = layer2_out[178] | layer2_out[179];
    assign layer3_out[264] = layer2_out[220] & ~layer2_out[219];
    assign layer3_out[265] = ~layer2_out[455] | layer2_out[456];
    assign layer3_out[266] = ~(layer2_out[149] & layer2_out[150]);
    assign layer3_out[267] = layer2_out[174] & layer2_out[175];
    assign layer3_out[268] = ~layer2_out[161];
    assign layer3_out[269] = ~(layer2_out[450] & layer2_out[451]);
    assign layer3_out[270] = ~(layer2_out[170] | layer2_out[171]);
    assign layer3_out[271] = layer2_out[476];
    assign layer3_out[272] = ~layer2_out[200] | layer2_out[201];
    assign layer3_out[273] = layer2_out[186];
    assign layer3_out[274] = ~layer2_out[41] | layer2_out[40];
    assign layer3_out[275] = layer2_out[261] & ~layer2_out[262];
    assign layer3_out[276] = ~(layer2_out[536] | layer2_out[537]);
    assign layer3_out[277] = layer2_out[47];
    assign layer3_out[278] = layer2_out[282];
    assign layer3_out[279] = ~(layer2_out[463] ^ layer2_out[464]);
    assign layer3_out[280] = layer2_out[486];
    assign layer3_out[281] = ~layer2_out[303];
    assign layer3_out[282] = ~(layer2_out[131] | layer2_out[132]);
    assign layer3_out[283] = ~(layer2_out[117] | layer2_out[118]);
    assign layer3_out[284] = layer2_out[227] | layer2_out[228];
    assign layer3_out[285] = ~layer2_out[129];
    assign layer3_out[286] = ~layer2_out[367];
    assign layer3_out[287] = layer2_out[351] & ~layer2_out[350];
    assign layer3_out[288] = layer2_out[188] ^ layer2_out[189];
    assign layer3_out[289] = ~layer2_out[442];
    assign layer3_out[290] = ~layer2_out[115];
    assign layer3_out[291] = ~layer2_out[513];
    assign layer3_out[292] = ~layer2_out[28];
    assign layer3_out[293] = layer2_out[548] | layer2_out[549];
    assign layer3_out[294] = ~(layer2_out[234] | layer2_out[235]);
    assign layer3_out[295] = layer2_out[238];
    assign layer3_out[296] = 1'b0;
    assign layer3_out[297] = ~layer2_out[58];
    assign layer3_out[298] = layer2_out[520];
    assign layer3_out[299] = layer2_out[169] & ~layer2_out[168];
    assign layer3_out[300] = ~(layer2_out[98] & layer2_out[99]);
    assign layer3_out[301] = ~layer2_out[337];
    assign layer3_out[302] = ~layer2_out[195] | layer2_out[194];
    assign layer3_out[303] = layer2_out[114] & ~layer2_out[113];
    assign layer3_out[304] = ~layer2_out[487] | layer2_out[488];
    assign layer3_out[305] = ~layer2_out[364] | layer2_out[363];
    assign layer3_out[306] = ~layer2_out[103];
    assign layer3_out[307] = ~layer2_out[35];
    assign layer3_out[308] = layer2_out[537] & ~layer2_out[538];
    assign layer3_out[309] = layer2_out[489] & ~layer2_out[488];
    assign layer3_out[310] = ~layer2_out[302] | layer2_out[301];
    assign layer3_out[311] = layer2_out[251];
    assign layer3_out[312] = layer2_out[475] & ~layer2_out[476];
    assign layer3_out[313] = layer2_out[305] & ~layer2_out[304];
    assign layer3_out[314] = layer2_out[135] | layer2_out[136];
    assign layer3_out[315] = ~layer2_out[301];
    assign layer3_out[316] = layer2_out[328] & layer2_out[329];
    assign layer3_out[317] = layer2_out[33];
    assign layer3_out[318] = layer2_out[182];
    assign layer3_out[319] = ~layer2_out[82];
    assign layer3_out[320] = ~layer2_out[70];
    assign layer3_out[321] = ~(layer2_out[423] & layer2_out[424]);
    assign layer3_out[322] = layer2_out[468] | layer2_out[469];
    assign layer3_out[323] = layer2_out[457];
    assign layer3_out[324] = layer2_out[54];
    assign layer3_out[325] = layer2_out[331] & ~layer2_out[330];
    assign layer3_out[326] = ~layer2_out[391];
    assign layer3_out[327] = ~layer2_out[400] | layer2_out[401];
    assign layer3_out[328] = ~layer2_out[237];
    assign layer3_out[329] = ~(layer2_out[61] | layer2_out[62]);
    assign layer3_out[330] = 1'b0;
    assign layer3_out[331] = layer2_out[258] | layer2_out[259];
    assign layer3_out[332] = layer2_out[481];
    assign layer3_out[333] = layer2_out[139] & ~layer2_out[140];
    assign layer3_out[334] = layer2_out[199];
    assign layer3_out[335] = layer2_out[467];
    assign layer3_out[336] = layer2_out[455];
    assign layer3_out[337] = ~layer2_out[52] | layer2_out[53];
    assign layer3_out[338] = ~layer2_out[495] | layer2_out[496];
    assign layer3_out[339] = layer2_out[101] & ~layer2_out[102];
    assign layer3_out[340] = layer2_out[473] & layer2_out[474];
    assign layer3_out[341] = ~layer2_out[67];
    assign layer3_out[342] = 1'b1;
    assign layer3_out[343] = layer2_out[221];
    assign layer3_out[344] = ~layer2_out[416] | layer2_out[417];
    assign layer3_out[345] = layer2_out[434] & ~layer2_out[435];
    assign layer3_out[346] = layer2_out[247] & ~layer2_out[248];
    assign layer3_out[347] = layer2_out[494];
    assign layer3_out[348] = layer2_out[335];
    assign layer3_out[349] = layer2_out[161] & ~layer2_out[162];
    assign layer3_out[350] = layer2_out[540];
    assign layer3_out[351] = ~layer2_out[51];
    assign layer3_out[352] = layer2_out[296];
    assign layer3_out[353] = layer2_out[203];
    assign layer3_out[354] = layer2_out[478];
    assign layer3_out[355] = layer2_out[31] & ~layer2_out[32];
    assign layer3_out[356] = layer2_out[328] & ~layer2_out[327];
    assign layer3_out[357] = ~(layer2_out[84] & layer2_out[85]);
    assign layer3_out[358] = layer2_out[520];
    assign layer3_out[359] = ~layer2_out[358] | layer2_out[357];
    assign layer3_out[360] = layer2_out[485];
    assign layer3_out[361] = ~layer2_out[81];
    assign layer3_out[362] = ~layer2_out[292] | layer2_out[291];
    assign layer3_out[363] = ~layer2_out[11];
    assign layer3_out[364] = layer2_out[267] | layer2_out[268];
    assign layer3_out[365] = ~layer2_out[105];
    assign layer3_out[366] = ~layer2_out[218];
    assign layer3_out[367] = layer2_out[365] & layer2_out[366];
    assign layer3_out[368] = ~layer2_out[204] | layer2_out[205];
    assign layer3_out[369] = layer2_out[77];
    assign layer3_out[370] = layer2_out[542];
    assign layer3_out[371] = ~(layer2_out[427] ^ layer2_out[428]);
    assign layer3_out[372] = 1'b1;
    assign layer3_out[373] = layer2_out[359];
    assign layer3_out[374] = 1'b1;
    assign layer3_out[375] = ~layer2_out[306];
    assign layer3_out[376] = layer2_out[377];
    assign layer3_out[377] = ~layer2_out[224];
    assign layer3_out[378] = layer2_out[62] | layer2_out[63];
    assign layer3_out[379] = ~(layer2_out[395] | layer2_out[396]);
    assign layer3_out[380] = ~layer2_out[231];
    assign layer3_out[381] = layer2_out[380];
    assign layer3_out[382] = layer2_out[397] ^ layer2_out[398];
    assign layer3_out[383] = layer2_out[245] & layer2_out[246];
    assign layer3_out[384] = ~layer2_out[530] | layer2_out[531];
    assign layer3_out[385] = layer2_out[245];
    assign layer3_out[386] = layer2_out[493];
    assign layer3_out[387] = layer2_out[353];
    assign layer3_out[388] = ~layer2_out[437];
    assign layer3_out[389] = ~layer2_out[187];
    assign layer3_out[390] = ~layer2_out[177];
    assign layer3_out[391] = layer2_out[494] & ~layer2_out[493];
    assign layer3_out[392] = ~layer2_out[433] | layer2_out[434];
    assign layer3_out[393] = ~(layer2_out[387] | layer2_out[388]);
    assign layer3_out[394] = ~layer2_out[346] | layer2_out[347];
    assign layer3_out[395] = ~layer2_out[146];
    assign layer3_out[396] = layer2_out[451] | layer2_out[452];
    assign layer3_out[397] = ~layer2_out[191] | layer2_out[192];
    assign layer3_out[398] = layer2_out[481] & ~layer2_out[480];
    assign layer3_out[399] = layer2_out[449];
    assign layer3_out[400] = ~(layer2_out[386] | layer2_out[387]);
    assign layer3_out[401] = ~layer2_out[329] | layer2_out[330];
    assign layer3_out[402] = ~(layer2_out[242] | layer2_out[243]);
    assign layer3_out[403] = 1'b1;
    assign layer3_out[404] = ~layer2_out[347];
    assign layer3_out[405] = layer2_out[432];
    assign layer3_out[406] = ~layer2_out[324];
    assign layer3_out[407] = layer2_out[354];
    assign layer3_out[408] = layer2_out[286] ^ layer2_out[287];
    assign layer3_out[409] = layer2_out[396];
    assign layer3_out[410] = ~(layer2_out[93] | layer2_out[94]);
    assign layer3_out[411] = layer2_out[422] & layer2_out[423];
    assign layer3_out[412] = ~(layer2_out[426] & layer2_out[427]);
    assign layer3_out[413] = ~(layer2_out[403] & layer2_out[404]);
    assign layer3_out[414] = layer2_out[203] & ~layer2_out[204];
    assign layer3_out[415] = layer2_out[368] & ~layer2_out[367];
    assign layer3_out[416] = layer2_out[162] & layer2_out[163];
    assign layer3_out[417] = layer2_out[411];
    assign layer3_out[418] = layer2_out[48];
    assign layer3_out[419] = layer2_out[503] & ~layer2_out[504];
    assign layer3_out[420] = ~(layer2_out[471] | layer2_out[472]);
    assign layer3_out[421] = ~(layer2_out[516] & layer2_out[517]);
    assign layer3_out[422] = layer2_out[332];
    assign layer3_out[423] = ~layer2_out[517] | layer2_out[518];
    assign layer3_out[424] = layer2_out[77] & ~layer2_out[76];
    assign layer3_out[425] = ~layer2_out[119] | layer2_out[118];
    assign layer3_out[426] = ~(layer2_out[385] & layer2_out[386]);
    assign layer3_out[427] = layer2_out[523] | layer2_out[524];
    assign layer3_out[428] = ~(layer2_out[373] & layer2_out[374]);
    assign layer3_out[429] = layer2_out[228] | layer2_out[229];
    assign layer3_out[430] = layer2_out[408] & ~layer2_out[409];
    assign layer3_out[431] = ~(layer2_out[133] & layer2_out[134]);
    assign layer3_out[432] = layer2_out[307];
    assign layer3_out[433] = 1'b0;
    assign layer3_out[434] = layer2_out[153] & layer2_out[154];
    assign layer3_out[435] = ~layer2_out[283];
    assign layer3_out[436] = layer2_out[324] & ~layer2_out[325];
    assign layer3_out[437] = ~layer2_out[33];
    assign layer3_out[438] = ~layer2_out[260];
    assign layer3_out[439] = layer2_out[421];
    assign layer3_out[440] = ~layer2_out[45] | layer2_out[44];
    assign layer3_out[441] = ~layer2_out[258];
    assign layer3_out[442] = ~layer2_out[183];
    assign layer3_out[443] = layer2_out[85] & ~layer2_out[86];
    assign layer3_out[444] = 1'b0;
    assign layer3_out[445] = ~(layer2_out[290] ^ layer2_out[291]);
    assign layer3_out[446] = layer2_out[294];
    assign layer3_out[447] = ~layer2_out[410];
    assign layer3_out[448] = layer2_out[502] & layer2_out[503];
    assign layer3_out[449] = layer2_out[420] & ~layer2_out[419];
    assign layer3_out[450] = layer2_out[166];
    assign layer3_out[451] = layer2_out[42] & layer2_out[43];
    assign layer3_out[452] = layer2_out[270] & ~layer2_out[269];
    assign layer3_out[453] = ~(layer2_out[196] & layer2_out[197]);
    assign layer3_out[454] = layer2_out[345] & ~layer2_out[344];
    assign layer3_out[455] = layer2_out[432];
    assign layer3_out[456] = layer2_out[289];
    assign layer3_out[457] = ~layer2_out[351];
    assign layer3_out[458] = layer2_out[56];
    assign layer3_out[459] = ~(layer2_out[124] & layer2_out[125]);
    assign layer3_out[460] = ~(layer2_out[369] | layer2_out[370]);
    assign layer3_out[461] = layer2_out[68] ^ layer2_out[69];
    assign layer3_out[462] = layer2_out[505] & ~layer2_out[506];
    assign layer3_out[463] = layer2_out[546] & layer2_out[547];
    assign layer3_out[464] = layer2_out[226] ^ layer2_out[227];
    assign layer3_out[465] = layer2_out[266];
    assign layer3_out[466] = layer2_out[158];
    assign layer3_out[467] = ~layer2_out[166] | layer2_out[165];
    assign layer3_out[468] = layer2_out[95];
    assign layer3_out[469] = ~(layer2_out[193] | layer2_out[194]);
    assign layer3_out[470] = ~layer2_out[212] | layer2_out[211];
    assign layer3_out[471] = layer2_out[78] & layer2_out[79];
    assign layer3_out[472] = ~(layer2_out[123] & layer2_out[124]);
    assign layer3_out[473] = ~layer2_out[208];
    assign layer3_out[474] = layer2_out[449];
    assign layer3_out[475] = layer2_out[22] | layer2_out[23];
    assign layer3_out[476] = layer2_out[352] | layer2_out[353];
    assign layer3_out[477] = ~layer2_out[410];
    assign layer3_out[478] = 1'b0;
    assign layer3_out[479] = ~layer2_out[506];
    assign layer3_out[480] = layer2_out[500] & layer2_out[501];
    assign layer3_out[481] = layer2_out[152] & ~layer2_out[151];
    assign layer3_out[482] = ~layer2_out[207] | layer2_out[206];
    assign layer3_out[483] = layer2_out[34];
    assign layer3_out[484] = layer2_out[489] | layer2_out[490];
    assign layer3_out[485] = layer2_out[418];
    assign layer3_out[486] = ~layer2_out[479] | layer2_out[480];
    assign layer3_out[487] = ~(layer2_out[38] & layer2_out[39]);
    assign layer3_out[488] = layer2_out[243];
    assign layer3_out[489] = layer2_out[508];
    assign layer3_out[490] = ~(layer2_out[498] & layer2_out[499]);
    assign layer3_out[491] = layer2_out[275];
    assign layer3_out[492] = ~layer2_out[452];
    assign layer3_out[493] = layer2_out[90];
    assign layer3_out[494] = ~layer2_out[457];
    assign layer3_out[495] = ~layer2_out[511];
    assign layer3_out[496] = layer2_out[150] | layer2_out[151];
    assign layer3_out[497] = ~layer2_out[310] | layer2_out[309];
    assign layer3_out[498] = layer2_out[382] & ~layer2_out[383];
    assign layer3_out[499] = layer2_out[326];
    assign layer3_out[500] = ~(layer2_out[318] | layer2_out[319]);
    assign layer3_out[501] = ~layer2_out[371] | layer2_out[370];
    assign layer3_out[502] = ~layer2_out[282] | layer2_out[283];
    assign layer3_out[503] = ~(layer2_out[528] & layer2_out[529]);
    assign layer3_out[504] = layer2_out[360];
    assign layer3_out[505] = ~(layer2_out[55] ^ layer2_out[56]);
    assign layer3_out[506] = ~(layer2_out[268] | layer2_out[269]);
    assign layer3_out[507] = ~layer2_out[18];
    assign layer3_out[508] = layer2_out[312] & ~layer2_out[313];
    assign layer3_out[509] = ~(layer2_out[509] | layer2_out[510]);
    assign layer3_out[510] = layer2_out[403];
    assign layer3_out[511] = ~layer2_out[394];
    assign layer3_out[512] = ~(layer2_out[184] & layer2_out[185]);
    assign layer3_out[513] = layer2_out[65];
    assign layer3_out[514] = ~layer2_out[136];
    assign layer3_out[515] = ~layer2_out[299] | layer2_out[300];
    assign layer3_out[516] = layer2_out[0] & ~layer2_out[2];
    assign layer3_out[517] = ~(layer2_out[23] ^ layer2_out[24]);
    assign layer3_out[518] = ~layer2_out[210];
    assign layer3_out[519] = 1'b1;
    assign layer3_out[520] = ~(layer2_out[443] | layer2_out[444]);
    assign layer3_out[521] = layer2_out[446];
    assign layer3_out[522] = layer2_out[86] & layer2_out[87];
    assign layer3_out[523] = ~layer2_out[270] | layer2_out[271];
    assign layer3_out[524] = ~(layer2_out[230] & layer2_out[231]);
    assign layer3_out[525] = layer2_out[109] & ~layer2_out[110];
    assign layer3_out[526] = layer2_out[232];
    assign layer3_out[527] = layer2_out[525];
    assign layer3_out[528] = ~layer2_out[104];
    assign layer3_out[529] = 1'b1;
    assign layer3_out[530] = layer2_out[388];
    assign layer3_out[531] = ~layer2_out[137];
    assign layer3_out[532] = layer2_out[111] & ~layer2_out[112];
    assign layer3_out[533] = layer2_out[182] & ~layer2_out[181];
    assign layer3_out[534] = 1'b0;
    assign layer3_out[535] = ~layer2_out[322];
    assign layer3_out[536] = layer2_out[30];
    assign layer3_out[537] = layer2_out[356];
    assign layer3_out[538] = ~(layer2_out[458] & layer2_out[459]);
    assign layer3_out[539] = ~(layer2_out[9] & layer2_out[10]);
    assign layer3_out[540] = ~layer2_out[73];
    assign layer3_out[541] = layer2_out[465];
    assign layer3_out[542] = ~layer2_out[339];
    assign layer3_out[543] = ~(layer2_out[171] & layer2_out[172]);
    assign layer3_out[544] = ~layer2_out[380] | layer2_out[381];
    assign layer3_out[545] = ~layer2_out[372];
    assign layer3_out[546] = layer2_out[484];
    assign layer3_out[547] = layer2_out[10] & layer2_out[11];
    assign layer3_out[548] = layer2_out[314] & ~layer2_out[315];
    assign layer3_out[549] = layer2_out[39] & ~layer2_out[40];
    assign layer4_out[0] = ~(layer3_out[248] & layer3_out[249]);
    assign layer4_out[1] = layer3_out[493] & ~layer3_out[492];
    assign layer4_out[2] = layer3_out[405] | layer3_out[406];
    assign layer4_out[3] = ~layer3_out[523] | layer3_out[524];
    assign layer4_out[4] = ~layer3_out[290];
    assign layer4_out[5] = layer3_out[406] | layer3_out[407];
    assign layer4_out[6] = layer3_out[336] ^ layer3_out[337];
    assign layer4_out[7] = ~(layer3_out[384] & layer3_out[385]);
    assign layer4_out[8] = layer3_out[105] & layer3_out[106];
    assign layer4_out[9] = layer3_out[313];
    assign layer4_out[10] = layer3_out[463];
    assign layer4_out[11] = ~layer3_out[277];
    assign layer4_out[12] = layer3_out[316] & ~layer3_out[317];
    assign layer4_out[13] = ~layer3_out[129];
    assign layer4_out[14] = ~(layer3_out[418] & layer3_out[419]);
    assign layer4_out[15] = ~layer3_out[487];
    assign layer4_out[16] = layer3_out[531];
    assign layer4_out[17] = layer3_out[128];
    assign layer4_out[18] = ~layer3_out[494] | layer3_out[493];
    assign layer4_out[19] = ~(layer3_out[314] & layer3_out[315]);
    assign layer4_out[20] = ~layer3_out[0] | layer3_out[2];
    assign layer4_out[21] = 1'b0;
    assign layer4_out[22] = ~layer3_out[518];
    assign layer4_out[23] = layer3_out[78];
    assign layer4_out[24] = ~layer3_out[473] | layer3_out[472];
    assign layer4_out[25] = ~layer3_out[527];
    assign layer4_out[26] = layer3_out[294];
    assign layer4_out[27] = ~layer3_out[349];
    assign layer4_out[28] = ~layer3_out[81] | layer3_out[80];
    assign layer4_out[29] = layer3_out[4] & ~layer3_out[5];
    assign layer4_out[30] = ~layer3_out[273];
    assign layer4_out[31] = ~layer3_out[70];
    assign layer4_out[32] = ~layer3_out[219];
    assign layer4_out[33] = layer3_out[399] & ~layer3_out[400];
    assign layer4_out[34] = ~layer3_out[535];
    assign layer4_out[35] = layer3_out[114];
    assign layer4_out[36] = layer3_out[408] & ~layer3_out[409];
    assign layer4_out[37] = ~layer3_out[296] | layer3_out[295];
    assign layer4_out[38] = ~layer3_out[530];
    assign layer4_out[39] = ~layer3_out[300] | layer3_out[299];
    assign layer4_out[40] = layer3_out[355];
    assign layer4_out[41] = layer3_out[291];
    assign layer4_out[42] = layer3_out[97];
    assign layer4_out[43] = layer3_out[535];
    assign layer4_out[44] = layer3_out[429] & layer3_out[430];
    assign layer4_out[45] = layer3_out[537] & layer3_out[538];
    assign layer4_out[46] = layer3_out[246] & ~layer3_out[247];
    assign layer4_out[47] = layer3_out[356] & ~layer3_out[357];
    assign layer4_out[48] = ~layer3_out[113];
    assign layer4_out[49] = layer3_out[232];
    assign layer4_out[50] = layer3_out[66];
    assign layer4_out[51] = layer3_out[20] | layer3_out[21];
    assign layer4_out[52] = layer3_out[190];
    assign layer4_out[53] = layer3_out[280] & ~layer3_out[279];
    assign layer4_out[54] = ~layer3_out[428];
    assign layer4_out[55] = ~layer3_out[202];
    assign layer4_out[56] = layer3_out[88] & layer3_out[89];
    assign layer4_out[57] = layer3_out[140] & layer3_out[141];
    assign layer4_out[58] = layer3_out[358] & ~layer3_out[359];
    assign layer4_out[59] = ~layer3_out[86];
    assign layer4_out[60] = layer3_out[540];
    assign layer4_out[61] = layer3_out[290];
    assign layer4_out[62] = layer3_out[342] & ~layer3_out[341];
    assign layer4_out[63] = ~(layer3_out[445] & layer3_out[446]);
    assign layer4_out[64] = 1'b1;
    assign layer4_out[65] = ~layer3_out[273];
    assign layer4_out[66] = ~(layer3_out[16] ^ layer3_out[17]);
    assign layer4_out[67] = layer3_out[240] & ~layer3_out[239];
    assign layer4_out[68] = layer3_out[9];
    assign layer4_out[69] = layer3_out[480] | layer3_out[481];
    assign layer4_out[70] = layer3_out[147] & layer3_out[148];
    assign layer4_out[71] = ~layer3_out[540];
    assign layer4_out[72] = layer3_out[541];
    assign layer4_out[73] = ~layer3_out[238] | layer3_out[239];
    assign layer4_out[74] = ~(layer3_out[275] ^ layer3_out[276]);
    assign layer4_out[75] = layer3_out[119];
    assign layer4_out[76] = ~layer3_out[545];
    assign layer4_out[77] = ~layer3_out[200];
    assign layer4_out[78] = layer3_out[498] & ~layer3_out[497];
    assign layer4_out[79] = layer3_out[417] | layer3_out[418];
    assign layer4_out[80] = layer3_out[214];
    assign layer4_out[81] = ~(layer3_out[412] & layer3_out[413]);
    assign layer4_out[82] = ~layer3_out[345];
    assign layer4_out[83] = layer3_out[173] & ~layer3_out[174];
    assign layer4_out[84] = ~layer3_out[182];
    assign layer4_out[85] = layer3_out[467] & ~layer3_out[468];
    assign layer4_out[86] = ~layer3_out[30] | layer3_out[31];
    assign layer4_out[87] = ~layer3_out[423];
    assign layer4_out[88] = layer3_out[192] & ~layer3_out[191];
    assign layer4_out[89] = ~layer3_out[437];
    assign layer4_out[90] = layer3_out[50] & ~layer3_out[49];
    assign layer4_out[91] = ~layer3_out[195];
    assign layer4_out[92] = layer3_out[83] & layer3_out[84];
    assign layer4_out[93] = ~layer3_out[466] | layer3_out[465];
    assign layer4_out[94] = ~layer3_out[48];
    assign layer4_out[95] = layer3_out[58];
    assign layer4_out[96] = ~layer3_out[172];
    assign layer4_out[97] = ~layer3_out[391];
    assign layer4_out[98] = layer3_out[218];
    assign layer4_out[99] = ~layer3_out[12];
    assign layer4_out[100] = ~(layer3_out[298] | layer3_out[299]);
    assign layer4_out[101] = ~(layer3_out[249] ^ layer3_out[250]);
    assign layer4_out[102] = ~layer3_out[165];
    assign layer4_out[103] = layer3_out[267] | layer3_out[268];
    assign layer4_out[104] = layer3_out[402] | layer3_out[403];
    assign layer4_out[105] = layer3_out[369];
    assign layer4_out[106] = layer3_out[415] | layer3_out[416];
    assign layer4_out[107] = 1'b1;
    assign layer4_out[108] = ~layer3_out[402];
    assign layer4_out[109] = layer3_out[310] & ~layer3_out[309];
    assign layer4_out[110] = ~layer3_out[226] | layer3_out[227];
    assign layer4_out[111] = layer3_out[43] ^ layer3_out[44];
    assign layer4_out[112] = layer3_out[504] & ~layer3_out[505];
    assign layer4_out[113] = layer3_out[334];
    assign layer4_out[114] = ~(layer3_out[447] & layer3_out[448]);
    assign layer4_out[115] = ~(layer3_out[61] | layer3_out[62]);
    assign layer4_out[116] = ~(layer3_out[84] ^ layer3_out[85]);
    assign layer4_out[117] = layer3_out[519] & layer3_out[520];
    assign layer4_out[118] = layer3_out[38] & ~layer3_out[37];
    assign layer4_out[119] = layer3_out[46];
    assign layer4_out[120] = ~(layer3_out[548] & layer3_out[549]);
    assign layer4_out[121] = ~layer3_out[547];
    assign layer4_out[122] = layer3_out[148] ^ layer3_out[149];
    assign layer4_out[123] = layer3_out[327] & layer3_out[328];
    assign layer4_out[124] = ~layer3_out[253];
    assign layer4_out[125] = layer3_out[90] & ~layer3_out[91];
    assign layer4_out[126] = layer3_out[141] & layer3_out[142];
    assign layer4_out[127] = layer3_out[527];
    assign layer4_out[128] = ~layer3_out[347];
    assign layer4_out[129] = layer3_out[388];
    assign layer4_out[130] = ~layer3_out[469];
    assign layer4_out[131] = ~layer3_out[436] | layer3_out[435];
    assign layer4_out[132] = layer3_out[455] | layer3_out[456];
    assign layer4_out[133] = ~layer3_out[380];
    assign layer4_out[134] = layer3_out[263] & ~layer3_out[264];
    assign layer4_out[135] = ~layer3_out[64];
    assign layer4_out[136] = 1'b1;
    assign layer4_out[137] = ~layer3_out[152] | layer3_out[153];
    assign layer4_out[138] = ~(layer3_out[542] & layer3_out[543]);
    assign layer4_out[139] = layer3_out[475] ^ layer3_out[476];
    assign layer4_out[140] = layer3_out[57];
    assign layer4_out[141] = ~layer3_out[256];
    assign layer4_out[142] = ~layer3_out[14] | layer3_out[13];
    assign layer4_out[143] = layer3_out[15] & ~layer3_out[16];
    assign layer4_out[144] = ~layer3_out[96] | layer3_out[95];
    assign layer4_out[145] = ~(layer3_out[301] ^ layer3_out[302]);
    assign layer4_out[146] = ~(layer3_out[27] | layer3_out[28]);
    assign layer4_out[147] = ~(layer3_out[306] | layer3_out[307]);
    assign layer4_out[148] = layer3_out[494] & layer3_out[495];
    assign layer4_out[149] = ~layer3_out[58];
    assign layer4_out[150] = ~(layer3_out[416] ^ layer3_out[417]);
    assign layer4_out[151] = layer3_out[98] & layer3_out[99];
    assign layer4_out[152] = ~(layer3_out[188] | layer3_out[189]);
    assign layer4_out[153] = ~(layer3_out[502] ^ layer3_out[503]);
    assign layer4_out[154] = ~layer3_out[66];
    assign layer4_out[155] = ~layer3_out[363] | layer3_out[364];
    assign layer4_out[156] = layer3_out[241] & ~layer3_out[242];
    assign layer4_out[157] = layer3_out[147];
    assign layer4_out[158] = 1'b1;
    assign layer4_out[159] = ~(layer3_out[305] ^ layer3_out[306]);
    assign layer4_out[160] = layer3_out[79] & layer3_out[80];
    assign layer4_out[161] = layer3_out[145];
    assign layer4_out[162] = ~layer3_out[265];
    assign layer4_out[163] = ~(layer3_out[367] ^ layer3_out[368]);
    assign layer4_out[164] = ~(layer3_out[261] & layer3_out[262]);
    assign layer4_out[165] = layer3_out[138] | layer3_out[139];
    assign layer4_out[166] = ~layer3_out[36];
    assign layer4_out[167] = layer3_out[153];
    assign layer4_out[168] = layer3_out[287] & ~layer3_out[286];
    assign layer4_out[169] = ~layer3_out[369];
    assign layer4_out[170] = layer3_out[51] | layer3_out[52];
    assign layer4_out[171] = layer3_out[29];
    assign layer4_out[172] = 1'b0;
    assign layer4_out[173] = ~(layer3_out[143] | layer3_out[144]);
    assign layer4_out[174] = ~layer3_out[489];
    assign layer4_out[175] = layer3_out[434];
    assign layer4_out[176] = ~layer3_out[85];
    assign layer4_out[177] = layer3_out[331];
    assign layer4_out[178] = 1'b0;
    assign layer4_out[179] = ~layer3_out[251];
    assign layer4_out[180] = layer3_out[319] & layer3_out[320];
    assign layer4_out[181] = ~layer3_out[362];
    assign layer4_out[182] = ~layer3_out[97];
    assign layer4_out[183] = layer3_out[54] ^ layer3_out[55];
    assign layer4_out[184] = layer3_out[61];
    assign layer4_out[185] = layer3_out[25] | layer3_out[26];
    assign layer4_out[186] = layer3_out[107] | layer3_out[108];
    assign layer4_out[187] = layer3_out[21];
    assign layer4_out[188] = ~(layer3_out[292] ^ layer3_out[293]);
    assign layer4_out[189] = layer3_out[448] & ~layer3_out[449];
    assign layer4_out[190] = ~layer3_out[530];
    assign layer4_out[191] = ~layer3_out[271];
    assign layer4_out[192] = ~layer3_out[349];
    assign layer4_out[193] = layer3_out[501] | layer3_out[502];
    assign layer4_out[194] = ~layer3_out[197];
    assign layer4_out[195] = ~layer3_out[404] | layer3_out[405];
    assign layer4_out[196] = ~layer3_out[366] | layer3_out[365];
    assign layer4_out[197] = layer3_out[377];
    assign layer4_out[198] = layer3_out[324] | layer3_out[325];
    assign layer4_out[199] = ~layer3_out[303] | layer3_out[304];
    assign layer4_out[200] = ~(layer3_out[205] & layer3_out[206]);
    assign layer4_out[201] = ~layer3_out[221];
    assign layer4_out[202] = ~layer3_out[142] | layer3_out[143];
    assign layer4_out[203] = ~(layer3_out[491] & layer3_out[492]);
    assign layer4_out[204] = layer3_out[167] & ~layer3_out[168];
    assign layer4_out[205] = ~(layer3_out[476] ^ layer3_out[477]);
    assign layer4_out[206] = layer3_out[93] & ~layer3_out[92];
    assign layer4_out[207] = ~layer3_out[77];
    assign layer4_out[208] = ~(layer3_out[70] & layer3_out[71]);
    assign layer4_out[209] = layer3_out[456] & layer3_out[457];
    assign layer4_out[210] = ~layer3_out[154];
    assign layer4_out[211] = layer3_out[244];
    assign layer4_out[212] = layer3_out[484] & ~layer3_out[485];
    assign layer4_out[213] = ~layer3_out[385] | layer3_out[386];
    assign layer4_out[214] = ~layer3_out[174] | layer3_out[175];
    assign layer4_out[215] = layer3_out[121] & layer3_out[122];
    assign layer4_out[216] = ~layer3_out[161] | layer3_out[160];
    assign layer4_out[217] = ~layer3_out[41];
    assign layer4_out[218] = ~layer3_out[521] | layer3_out[522];
    assign layer4_out[219] = layer3_out[428];
    assign layer4_out[220] = ~(layer3_out[179] & layer3_out[180]);
    assign layer4_out[221] = ~(layer3_out[460] & layer3_out[461]);
    assign layer4_out[222] = ~layer3_out[127];
    assign layer4_out[223] = ~layer3_out[7] | layer3_out[6];
    assign layer4_out[224] = layer3_out[498] & ~layer3_out[499];
    assign layer4_out[225] = layer3_out[217] | layer3_out[218];
    assign layer4_out[226] = ~(layer3_out[318] & layer3_out[319]);
    assign layer4_out[227] = ~layer3_out[40] | layer3_out[39];
    assign layer4_out[228] = 1'b1;
    assign layer4_out[229] = layer3_out[254] & ~layer3_out[255];
    assign layer4_out[230] = ~layer3_out[228];
    assign layer4_out[231] = ~layer3_out[103];
    assign layer4_out[232] = layer3_out[339];
    assign layer4_out[233] = layer3_out[244];
    assign layer4_out[234] = ~layer3_out[286];
    assign layer4_out[235] = layer3_out[149] & layer3_out[150];
    assign layer4_out[236] = layer3_out[471];
    assign layer4_out[237] = ~(layer3_out[517] & layer3_out[518]);
    assign layer4_out[238] = ~layer3_out[322];
    assign layer4_out[239] = ~layer3_out[352];
    assign layer4_out[240] = layer3_out[110];
    assign layer4_out[241] = ~layer3_out[22] | layer3_out[23];
    assign layer4_out[242] = layer3_out[374] ^ layer3_out[375];
    assign layer4_out[243] = ~layer3_out[443];
    assign layer4_out[244] = layer3_out[282] | layer3_out[283];
    assign layer4_out[245] = ~(layer3_out[481] | layer3_out[482]);
    assign layer4_out[246] = ~(layer3_out[512] ^ layer3_out[513]);
    assign layer4_out[247] = layer3_out[302];
    assign layer4_out[248] = ~layer3_out[166] | layer3_out[167];
    assign layer4_out[249] = ~layer3_out[23] | layer3_out[24];
    assign layer4_out[250] = layer3_out[252];
    assign layer4_out[251] = layer3_out[18];
    assign layer4_out[252] = ~layer3_out[19];
    assign layer4_out[253] = ~(layer3_out[362] & layer3_out[363]);
    assign layer4_out[254] = ~(layer3_out[48] & layer3_out[49]);
    assign layer4_out[255] = ~layer3_out[62] | layer3_out[63];
    assign layer4_out[256] = layer3_out[501];
    assign layer4_out[257] = layer3_out[52];
    assign layer4_out[258] = layer3_out[14] & ~layer3_out[15];
    assign layer4_out[259] = ~(layer3_out[287] & layer3_out[288]);
    assign layer4_out[260] = ~layer3_out[1];
    assign layer4_out[261] = ~layer3_out[507] | layer3_out[508];
    assign layer4_out[262] = 1'b1;
    assign layer4_out[263] = ~(layer3_out[18] ^ layer3_out[19]);
    assign layer4_out[264] = layer3_out[255] | layer3_out[256];
    assign layer4_out[265] = ~layer3_out[434];
    assign layer4_out[266] = ~layer3_out[231];
    assign layer4_out[267] = layer3_out[54] & ~layer3_out[53];
    assign layer4_out[268] = ~layer3_out[415];
    assign layer4_out[269] = layer3_out[189] & layer3_out[190];
    assign layer4_out[270] = ~layer3_out[157];
    assign layer4_out[271] = ~(layer3_out[464] | layer3_out[465]);
    assign layer4_out[272] = layer3_out[298] & ~layer3_out[297];
    assign layer4_out[273] = ~(layer3_out[209] & layer3_out[210]);
    assign layer4_out[274] = layer3_out[162];
    assign layer4_out[275] = layer3_out[72] & layer3_out[73];
    assign layer4_out[276] = layer3_out[30];
    assign layer4_out[277] = ~layer3_out[305];
    assign layer4_out[278] = layer3_out[111];
    assign layer4_out[279] = layer3_out[262] & ~layer3_out[263];
    assign layer4_out[280] = layer3_out[295];
    assign layer4_out[281] = ~layer3_out[373];
    assign layer4_out[282] = ~layer3_out[187];
    assign layer4_out[283] = ~(layer3_out[419] | layer3_out[420]);
    assign layer4_out[284] = ~layer3_out[424];
    assign layer4_out[285] = ~(layer3_out[236] & layer3_out[237]);
    assign layer4_out[286] = ~layer3_out[452] | layer3_out[453];
    assign layer4_out[287] = ~layer3_out[216];
    assign layer4_out[288] = layer3_out[74] & ~layer3_out[75];
    assign layer4_out[289] = ~layer3_out[60];
    assign layer4_out[290] = ~layer3_out[392];
    assign layer4_out[291] = layer3_out[42];
    assign layer4_out[292] = layer3_out[335];
    assign layer4_out[293] = layer3_out[24] | layer3_out[25];
    assign layer4_out[294] = layer3_out[225] & ~layer3_out[226];
    assign layer4_out[295] = layer3_out[371];
    assign layer4_out[296] = layer3_out[185] & ~layer3_out[184];
    assign layer4_out[297] = 1'b0;
    assign layer4_out[298] = ~layer3_out[69];
    assign layer4_out[299] = ~layer3_out[373];
    assign layer4_out[300] = layer3_out[343];
    assign layer4_out[301] = layer3_out[137] & ~layer3_out[136];
    assign layer4_out[302] = layer3_out[268];
    assign layer4_out[303] = layer3_out[412] & ~layer3_out[411];
    assign layer4_out[304] = layer3_out[528] | layer3_out[529];
    assign layer4_out[305] = layer3_out[176] | layer3_out[177];
    assign layer4_out[306] = ~layer3_out[393] | layer3_out[394];
    assign layer4_out[307] = ~layer3_out[437] | layer3_out[436];
    assign layer4_out[308] = layer3_out[35] & ~layer3_out[36];
    assign layer4_out[309] = ~layer3_out[6];
    assign layer4_out[310] = layer3_out[258] | layer3_out[259];
    assign layer4_out[311] = ~layer3_out[152] | layer3_out[151];
    assign layer4_out[312] = ~layer3_out[539];
    assign layer4_out[313] = ~layer3_out[526] | layer3_out[525];
    assign layer4_out[314] = layer3_out[479] | layer3_out[480];
    assign layer4_out[315] = layer3_out[516];
    assign layer4_out[316] = layer3_out[203] & ~layer3_out[202];
    assign layer4_out[317] = layer3_out[3];
    assign layer4_out[318] = layer3_out[522] & layer3_out[523];
    assign layer4_out[319] = ~layer3_out[3] | layer3_out[2];
    assign layer4_out[320] = ~(layer3_out[344] ^ layer3_out[345]);
    assign layer4_out[321] = layer3_out[459];
    assign layer4_out[322] = ~(layer3_out[134] & layer3_out[135]);
    assign layer4_out[323] = ~layer3_out[50];
    assign layer4_out[324] = ~layer3_out[169] | layer3_out[168];
    assign layer4_out[325] = layer3_out[384] & ~layer3_out[383];
    assign layer4_out[326] = ~layer3_out[457];
    assign layer4_out[327] = ~layer3_out[128];
    assign layer4_out[328] = layer3_out[477];
    assign layer4_out[329] = layer3_out[247];
    assign layer4_out[330] = ~(layer3_out[320] & layer3_out[321]);
    assign layer4_out[331] = layer3_out[350];
    assign layer4_out[332] = ~layer3_out[468] | layer3_out[469];
    assign layer4_out[333] = layer3_out[104] & layer3_out[105];
    assign layer4_out[334] = 1'b0;
    assign layer4_out[335] = ~layer3_out[124] | layer3_out[123];
    assign layer4_out[336] = layer3_out[197];
    assign layer4_out[337] = layer3_out[259];
    assign layer4_out[338] = ~layer3_out[459];
    assign layer4_out[339] = layer3_out[139];
    assign layer4_out[340] = ~layer3_out[325];
    assign layer4_out[341] = ~layer3_out[157];
    assign layer4_out[342] = ~layer3_out[266] | layer3_out[267];
    assign layer4_out[343] = layer3_out[81] | layer3_out[82];
    assign layer4_out[344] = layer3_out[378] & layer3_out[379];
    assign layer4_out[345] = layer3_out[401];
    assign layer4_out[346] = layer3_out[160];
    assign layer4_out[347] = layer3_out[311] & layer3_out[312];
    assign layer4_out[348] = ~(layer3_out[499] ^ layer3_out[500]);
    assign layer4_out[349] = ~layer3_out[68];
    assign layer4_out[350] = layer3_out[338];
    assign layer4_out[351] = layer3_out[317] & layer3_out[318];
    assign layer4_out[352] = ~layer3_out[120];
    assign layer4_out[353] = ~(layer3_out[177] | layer3_out[178]);
    assign layer4_out[354] = layer3_out[272];
    assign layer4_out[355] = layer3_out[495];
    assign layer4_out[356] = ~layer3_out[94] | layer3_out[95];
    assign layer4_out[357] = ~layer3_out[163] | layer3_out[164];
    assign layer4_out[358] = ~(layer3_out[124] | layer3_out[125]);
    assign layer4_out[359] = layer3_out[536] & ~layer3_out[537];
    assign layer4_out[360] = layer3_out[314];
    assign layer4_out[361] = ~layer3_out[212];
    assign layer4_out[362] = ~(layer3_out[351] & layer3_out[352]);
    assign layer4_out[363] = layer3_out[183];
    assign layer4_out[364] = layer3_out[33];
    assign layer4_out[365] = ~layer3_out[145] | layer3_out[144];
    assign layer4_out[366] = layer3_out[138];
    assign layer4_out[367] = layer3_out[130] | layer3_out[131];
    assign layer4_out[368] = layer3_out[442] & ~layer3_out[441];
    assign layer4_out[369] = ~layer3_out[389];
    assign layer4_out[370] = layer3_out[347] & ~layer3_out[346];
    assign layer4_out[371] = ~(layer3_out[296] & layer3_out[297]);
    assign layer4_out[372] = ~layer3_out[170];
    assign layer4_out[373] = ~layer3_out[516];
    assign layer4_out[374] = ~layer3_out[170] | layer3_out[169];
    assign layer4_out[375] = layer3_out[103] & layer3_out[104];
    assign layer4_out[376] = ~layer3_out[510];
    assign layer4_out[377] = layer3_out[322];
    assign layer4_out[378] = ~layer3_out[300];
    assign layer4_out[379] = layer3_out[207] & layer3_out[208];
    assign layer4_out[380] = layer3_out[450];
    assign layer4_out[381] = layer3_out[278] | layer3_out[279];
    assign layer4_out[382] = layer3_out[235] | layer3_out[236];
    assign layer4_out[383] = layer3_out[432];
    assign layer4_out[384] = 1'b0;
    assign layer4_out[385] = ~layer3_out[354] | layer3_out[355];
    assign layer4_out[386] = ~(layer3_out[110] ^ layer3_out[111]);
    assign layer4_out[387] = layer3_out[311];
    assign layer4_out[388] = ~layer3_out[224] | layer3_out[223];
    assign layer4_out[389] = ~layer3_out[472] | layer3_out[471];
    assign layer4_out[390] = ~(layer3_out[442] | layer3_out[443]);
    assign layer4_out[391] = layer3_out[399];
    assign layer4_out[392] = ~(layer3_out[264] | layer3_out[265]);
    assign layer4_out[393] = 1'b1;
    assign layer4_out[394] = layer3_out[397] & layer3_out[398];
    assign layer4_out[395] = layer3_out[155] | layer3_out[156];
    assign layer4_out[396] = layer3_out[210] & layer3_out[211];
    assign layer4_out[397] = ~layer3_out[224];
    assign layer4_out[398] = ~layer3_out[533];
    assign layer4_out[399] = ~layer3_out[396];
    assign layer4_out[400] = ~layer3_out[394] | layer3_out[395];
    assign layer4_out[401] = ~layer3_out[440];
    assign layer4_out[402] = ~layer3_out[454];
    assign layer4_out[403] = ~layer3_out[232];
    assign layer4_out[404] = ~layer3_out[192] | layer3_out[193];
    assign layer4_out[405] = ~layer3_out[172] | layer3_out[171];
    assign layer4_out[406] = layer3_out[440] & ~layer3_out[441];
    assign layer4_out[407] = layer3_out[431];
    assign layer4_out[408] = ~layer3_out[422];
    assign layer4_out[409] = layer3_out[445];
    assign layer4_out[410] = layer3_out[109] & ~layer3_out[108];
    assign layer4_out[411] = layer3_out[200];
    assign layer4_out[412] = layer3_out[371];
    assign layer4_out[413] = ~layer3_out[113];
    assign layer4_out[414] = layer3_out[315];
    assign layer4_out[415] = layer3_out[7] & layer3_out[8];
    assign layer4_out[416] = layer3_out[181];
    assign layer4_out[417] = ~layer3_out[425] | layer3_out[426];
    assign layer4_out[418] = layer3_out[382];
    assign layer4_out[419] = ~layer3_out[353];
    assign layer4_out[420] = layer3_out[508] ^ layer3_out[509];
    assign layer4_out[421] = ~(layer3_out[473] & layer3_out[474]);
    assign layer4_out[422] = ~layer3_out[451];
    assign layer4_out[423] = ~layer3_out[341];
    assign layer4_out[424] = ~layer3_out[193];
    assign layer4_out[425] = ~layer3_out[490];
    assign layer4_out[426] = ~layer3_out[430];
    assign layer4_out[427] = ~layer3_out[222];
    assign layer4_out[428] = layer3_out[34];
    assign layer4_out[429] = layer3_out[389];
    assign layer4_out[430] = layer3_out[77];
    assign layer4_out[431] = ~layer3_out[76] | layer3_out[75];
    assign layer4_out[432] = ~layer3_out[246];
    assign layer4_out[433] = ~layer3_out[475];
    assign layer4_out[434] = layer3_out[308];
    assign layer4_out[435] = ~layer3_out[31];
    assign layer4_out[436] = ~layer3_out[366] | layer3_out[367];
    assign layer4_out[437] = layer3_out[175] ^ layer3_out[176];
    assign layer4_out[438] = layer3_out[276] ^ layer3_out[277];
    assign layer4_out[439] = layer3_out[309];
    assign layer4_out[440] = layer3_out[233];
    assign layer4_out[441] = layer3_out[284] & ~layer3_out[283];
    assign layer4_out[442] = ~layer3_out[339];
    assign layer4_out[443] = ~layer3_out[510];
    assign layer4_out[444] = ~(layer3_out[446] & layer3_out[447]);
    assign layer4_out[445] = ~(layer3_out[520] | layer3_out[521]);
    assign layer4_out[446] = ~layer3_out[125];
    assign layer4_out[447] = ~layer3_out[333];
    assign layer4_out[448] = layer3_out[91] ^ layer3_out[92];
    assign layer4_out[449] = layer3_out[74];
    assign layer4_out[450] = 1'b1;
    assign layer4_out[451] = layer3_out[196] & ~layer3_out[195];
    assign layer4_out[452] = ~layer3_out[165] | layer3_out[164];
    assign layer4_out[453] = layer3_out[258] & ~layer3_out[257];
    assign layer4_out[454] = ~(layer3_out[132] | layer3_out[133]);
    assign layer4_out[455] = layer3_out[63] | layer3_out[64];
    assign layer4_out[456] = ~(layer3_out[332] | layer3_out[333]);
    assign layer4_out[457] = ~layer3_out[214] | layer3_out[215];
    assign layer4_out[458] = layer3_out[133] ^ layer3_out[134];
    assign layer4_out[459] = ~(layer3_out[288] & layer3_out[289]);
    assign layer4_out[460] = layer3_out[122] & ~layer3_out[123];
    assign layer4_out[461] = ~layer3_out[454];
    assign layer4_out[462] = ~layer3_out[490];
    assign layer4_out[463] = ~layer3_out[281];
    assign layer4_out[464] = layer3_out[485];
    assign layer4_out[465] = layer3_out[120] | layer3_out[121];
    assign layer4_out[466] = layer3_out[242];
    assign layer4_out[467] = layer3_out[484];
    assign layer4_out[468] = layer3_out[217];
    assign layer4_out[469] = ~layer3_out[503];
    assign layer4_out[470] = layer3_out[227] & layer3_out[228];
    assign layer4_out[471] = layer3_out[420];
    assign layer4_out[472] = ~(layer3_out[284] & layer3_out[285]);
    assign layer4_out[473] = layer3_out[377] & layer3_out[378];
    assign layer4_out[474] = ~(layer3_out[87] | layer3_out[88]);
    assign layer4_out[475] = ~(layer3_out[451] | layer3_out[452]);
    assign layer4_out[476] = ~(layer3_out[375] ^ layer3_out[376]);
    assign layer4_out[477] = ~layer3_out[182];
    assign layer4_out[478] = layer3_out[116] & ~layer3_out[117];
    assign layer4_out[479] = ~(layer3_out[131] & layer3_out[132]);
    assign layer4_out[480] = layer3_out[229] & ~layer3_out[230];
    assign layer4_out[481] = layer3_out[260] & ~layer3_out[261];
    assign layer4_out[482] = ~(layer3_out[466] & layer3_out[467]);
    assign layer4_out[483] = layer3_out[396] & ~layer3_out[397];
    assign layer4_out[484] = layer3_out[89] & ~layer3_out[90];
    assign layer4_out[485] = layer3_out[100];
    assign layer4_out[486] = layer3_out[328] & ~layer3_out[329];
    assign layer4_out[487] = ~layer3_out[33];
    assign layer4_out[488] = layer3_out[45];
    assign layer4_out[489] = ~layer3_out[101] | layer3_out[102];
    assign layer4_out[490] = layer3_out[360];
    assign layer4_out[491] = layer3_out[487] & ~layer3_out[488];
    assign layer4_out[492] = layer3_out[329];
    assign layer4_out[493] = ~layer3_out[274] | layer3_out[275];
    assign layer4_out[494] = layer3_out[26];
    assign layer4_out[495] = ~layer3_out[327];
    assign layer4_out[496] = ~layer3_out[545];
    assign layer4_out[497] = ~layer3_out[404];
    assign layer4_out[498] = layer3_out[511];
    assign layer4_out[499] = 1'b0;
    assign layer4_out[500] = ~layer3_out[0];
    assign layer4_out[501] = ~layer3_out[212];
    assign layer4_out[502] = layer3_out[118] & ~layer3_out[117];
    assign layer4_out[503] = layer3_out[135] ^ layer3_out[136];
    assign layer4_out[504] = layer3_out[410] ^ layer3_out[411];
    assign layer4_out[505] = ~layer3_out[496];
    assign layer4_out[506] = ~(layer3_out[115] ^ layer3_out[116]);
    assign layer4_out[507] = ~layer3_out[281];
    assign layer4_out[508] = layer3_out[199];
    assign layer4_out[509] = layer3_out[463] | layer3_out[464];
    assign layer4_out[510] = ~layer3_out[72] | layer3_out[71];
    assign layer4_out[511] = layer3_out[525];
    assign layer4_out[512] = layer3_out[222] | layer3_out[223];
    assign layer4_out[513] = layer3_out[240];
    assign layer4_out[514] = ~layer3_out[101];
    assign layer4_out[515] = ~layer3_out[514] | layer3_out[515];
    assign layer4_out[516] = ~layer3_out[413];
    assign layer4_out[517] = ~layer3_out[483];
    assign layer4_out[518] = layer3_out[187] | layer3_out[188];
    assign layer4_out[519] = layer3_out[514];
    assign layer4_out[520] = 1'b0;
    assign layer4_out[521] = ~layer3_out[506];
    assign layer4_out[522] = ~layer3_out[479];
    assign layer4_out[523] = ~layer3_out[38] | layer3_out[39];
    assign layer4_out[524] = layer3_out[461] ^ layer3_out[462];
    assign layer4_out[525] = ~layer3_out[178];
    assign layer4_out[526] = ~layer3_out[408];
    assign layer4_out[527] = layer3_out[386];
    assign layer4_out[528] = layer3_out[505] | layer3_out[506];
    assign layer4_out[529] = ~layer3_out[364] | layer3_out[365];
    assign layer4_out[530] = layer3_out[11];
    assign layer4_out[531] = layer3_out[207] & ~layer3_out[206];
    assign layer4_out[532] = ~layer3_out[158];
    assign layer4_out[533] = layer3_out[546] & layer3_out[547];
    assign layer4_out[534] = ~layer3_out[8] | layer3_out[9];
    assign layer4_out[535] = layer3_out[393];
    assign layer4_out[536] = ~(layer3_out[93] & layer3_out[94]);
    assign layer4_out[537] = layer3_out[357] & ~layer3_out[358];
    assign layer4_out[538] = layer3_out[380] | layer3_out[381];
    assign layer4_out[539] = ~layer3_out[237] | layer3_out[238];
    assign layer4_out[540] = layer3_out[150] & ~layer3_out[151];
    assign layer4_out[541] = ~layer3_out[543];
    assign layer4_out[542] = layer3_out[204];
    assign layer4_out[543] = layer3_out[234] & ~layer3_out[235];
    assign layer4_out[544] = ~layer3_out[383] | layer3_out[382];
    assign layer4_out[545] = layer3_out[532] & layer3_out[533];
    assign layer4_out[546] = ~layer3_out[323];
    assign layer4_out[547] = layer3_out[360] ^ layer3_out[361];
    assign layer4_out[548] = ~layer3_out[269];
    assign layer4_out[549] = layer3_out[55] & ~layer3_out[56];
    assign layer5_out[0] = ~layer4_out[116];
    assign layer5_out[1] = ~(layer4_out[338] | layer4_out[339]);
    assign layer5_out[2] = layer4_out[318];
    assign layer5_out[3] = layer4_out[44];
    assign layer5_out[4] = ~layer4_out[197];
    assign layer5_out[5] = layer4_out[540];
    assign layer5_out[6] = layer4_out[283];
    assign layer5_out[7] = ~(layer4_out[533] ^ layer4_out[534]);
    assign layer5_out[8] = ~layer4_out[52];
    assign layer5_out[9] = ~(layer4_out[253] & layer4_out[254]);
    assign layer5_out[10] = ~layer4_out[410];
    assign layer5_out[11] = layer4_out[452] & ~layer4_out[453];
    assign layer5_out[12] = ~layer4_out[532];
    assign layer5_out[13] = ~(layer4_out[486] | layer4_out[487]);
    assign layer5_out[14] = ~(layer4_out[425] | layer4_out[426]);
    assign layer5_out[15] = ~(layer4_out[487] | layer4_out[488]);
    assign layer5_out[16] = ~layer4_out[332];
    assign layer5_out[17] = layer4_out[159];
    assign layer5_out[18] = ~layer4_out[18];
    assign layer5_out[19] = layer4_out[528] & ~layer4_out[529];
    assign layer5_out[20] = ~layer4_out[394];
    assign layer5_out[21] = ~(layer4_out[531] | layer4_out[532]);
    assign layer5_out[22] = layer4_out[447];
    assign layer5_out[23] = layer4_out[417] & layer4_out[418];
    assign layer5_out[24] = ~layer4_out[355];
    assign layer5_out[25] = ~layer4_out[510];
    assign layer5_out[26] = layer4_out[340] & ~layer4_out[339];
    assign layer5_out[27] = ~layer4_out[326];
    assign layer5_out[28] = ~(layer4_out[123] | layer4_out[124]);
    assign layer5_out[29] = layer4_out[474];
    assign layer5_out[30] = ~(layer4_out[60] | layer4_out[61]);
    assign layer5_out[31] = layer4_out[364] & layer4_out[365];
    assign layer5_out[32] = ~layer4_out[9];
    assign layer5_out[33] = layer4_out[243] & ~layer4_out[244];
    assign layer5_out[34] = ~(layer4_out[101] | layer4_out[102]);
    assign layer5_out[35] = layer4_out[32] & ~layer4_out[33];
    assign layer5_out[36] = ~layer4_out[224];
    assign layer5_out[37] = ~(layer4_out[133] | layer4_out[134]);
    assign layer5_out[38] = layer4_out[239];
    assign layer5_out[39] = layer4_out[65] & ~layer4_out[66];
    assign layer5_out[40] = layer4_out[278];
    assign layer5_out[41] = ~(layer4_out[53] | layer4_out[54]);
    assign layer5_out[42] = ~layer4_out[521] | layer4_out[520];
    assign layer5_out[43] = layer4_out[461] & ~layer4_out[462];
    assign layer5_out[44] = layer4_out[459];
    assign layer5_out[45] = ~(layer4_out[94] ^ layer4_out[95]);
    assign layer5_out[46] = layer4_out[75] & layer4_out[76];
    assign layer5_out[47] = layer4_out[514] ^ layer4_out[515];
    assign layer5_out[48] = layer4_out[235];
    assign layer5_out[49] = ~layer4_out[276] | layer4_out[275];
    assign layer5_out[50] = layer4_out[144];
    assign layer5_out[51] = layer4_out[431] & ~layer4_out[430];
    assign layer5_out[52] = layer4_out[259] & layer4_out[260];
    assign layer5_out[53] = ~(layer4_out[265] | layer4_out[266]);
    assign layer5_out[54] = layer4_out[356] & layer4_out[357];
    assign layer5_out[55] = ~layer4_out[20];
    assign layer5_out[56] = ~layer4_out[395] | layer4_out[394];
    assign layer5_out[57] = layer4_out[200];
    assign layer5_out[58] = ~(layer4_out[464] | layer4_out[465]);
    assign layer5_out[59] = layer4_out[222] & ~layer4_out[223];
    assign layer5_out[60] = ~(layer4_out[114] | layer4_out[115]);
    assign layer5_out[61] = layer4_out[414] & layer4_out[415];
    assign layer5_out[62] = ~layer4_out[357];
    assign layer5_out[63] = layer4_out[473];
    assign layer5_out[64] = ~layer4_out[441];
    assign layer5_out[65] = ~layer4_out[176];
    assign layer5_out[66] = layer4_out[530] & layer4_out[531];
    assign layer5_out[67] = ~(layer4_out[248] & layer4_out[249]);
    assign layer5_out[68] = ~layer4_out[477];
    assign layer5_out[69] = layer4_out[100];
    assign layer5_out[70] = layer4_out[206];
    assign layer5_out[71] = layer4_out[158] ^ layer4_out[159];
    assign layer5_out[72] = layer4_out[23] & ~layer4_out[24];
    assign layer5_out[73] = ~(layer4_out[527] | layer4_out[528]);
    assign layer5_out[74] = layer4_out[247] ^ layer4_out[248];
    assign layer5_out[75] = layer4_out[548];
    assign layer5_out[76] = layer4_out[212] & ~layer4_out[213];
    assign layer5_out[77] = ~layer4_out[383];
    assign layer5_out[78] = ~layer4_out[544];
    assign layer5_out[79] = ~(layer4_out[371] ^ layer4_out[372]);
    assign layer5_out[80] = layer4_out[125];
    assign layer5_out[81] = ~(layer4_out[305] | layer4_out[306]);
    assign layer5_out[82] = layer4_out[8] ^ layer4_out[9];
    assign layer5_out[83] = layer4_out[45];
    assign layer5_out[84] = ~(layer4_out[195] | layer4_out[196]);
    assign layer5_out[85] = layer4_out[331];
    assign layer5_out[86] = layer4_out[60] & ~layer4_out[59];
    assign layer5_out[87] = layer4_out[233] & ~layer4_out[234];
    assign layer5_out[88] = ~layer4_out[544];
    assign layer5_out[89] = ~layer4_out[381];
    assign layer5_out[90] = layer4_out[480] & ~layer4_out[481];
    assign layer5_out[91] = ~(layer4_out[284] | layer4_out[285]);
    assign layer5_out[92] = layer4_out[473] & ~layer4_out[474];
    assign layer5_out[93] = ~layer4_out[74];
    assign layer5_out[94] = layer4_out[47];
    assign layer5_out[95] = ~layer4_out[335];
    assign layer5_out[96] = ~layer4_out[213];
    assign layer5_out[97] = layer4_out[392];
    assign layer5_out[98] = ~(layer4_out[217] | layer4_out[218]);
    assign layer5_out[99] = layer4_out[23] & ~layer4_out[22];
    assign layer5_out[100] = ~layer4_out[76];
    assign layer5_out[101] = layer4_out[13] & ~layer4_out[14];
    assign layer5_out[102] = ~layer4_out[371] | layer4_out[370];
    assign layer5_out[103] = ~(layer4_out[108] | layer4_out[109]);
    assign layer5_out[104] = layer4_out[493] & ~layer4_out[494];
    assign layer5_out[105] = ~(layer4_out[120] & layer4_out[121]);
    assign layer5_out[106] = ~layer4_out[311];
    assign layer5_out[107] = layer4_out[129] & ~layer4_out[130];
    assign layer5_out[108] = layer4_out[135];
    assign layer5_out[109] = ~layer4_out[137];
    assign layer5_out[110] = ~layer4_out[19];
    assign layer5_out[111] = layer4_out[475] & layer4_out[476];
    assign layer5_out[112] = layer4_out[41];
    assign layer5_out[113] = layer4_out[134] & layer4_out[135];
    assign layer5_out[114] = layer4_out[268] & ~layer4_out[269];
    assign layer5_out[115] = layer4_out[36];
    assign layer5_out[116] = ~layer4_out[103] | layer4_out[102];
    assign layer5_out[117] = layer4_out[448];
    assign layer5_out[118] = layer4_out[57] & ~layer4_out[58];
    assign layer5_out[119] = layer4_out[165] & layer4_out[166];
    assign layer5_out[120] = ~(layer4_out[274] | layer4_out[275]);
    assign layer5_out[121] = ~layer4_out[6];
    assign layer5_out[122] = layer4_out[447];
    assign layer5_out[123] = layer4_out[194];
    assign layer5_out[124] = layer4_out[7];
    assign layer5_out[125] = layer4_out[50] & ~layer4_out[49];
    assign layer5_out[126] = layer4_out[105] & ~layer4_out[106];
    assign layer5_out[127] = layer4_out[481] ^ layer4_out[482];
    assign layer5_out[128] = layer4_out[332] & ~layer4_out[333];
    assign layer5_out[129] = ~layer4_out[198];
    assign layer5_out[130] = ~(layer4_out[395] & layer4_out[396]);
    assign layer5_out[131] = layer4_out[296];
    assign layer5_out[132] = ~(layer4_out[206] | layer4_out[207]);
    assign layer5_out[133] = ~(layer4_out[317] | layer4_out[318]);
    assign layer5_out[134] = layer4_out[345] & ~layer4_out[346];
    assign layer5_out[135] = ~(layer4_out[420] & layer4_out[421]);
    assign layer5_out[136] = ~layer4_out[242];
    assign layer5_out[137] = ~(layer4_out[302] | layer4_out[303]);
    assign layer5_out[138] = ~layer4_out[86];
    assign layer5_out[139] = layer4_out[246];
    assign layer5_out[140] = layer4_out[403];
    assign layer5_out[141] = layer4_out[205];
    assign layer5_out[142] = layer4_out[514];
    assign layer5_out[143] = ~(layer4_out[526] | layer4_out[527]);
    assign layer5_out[144] = layer4_out[490] & layer4_out[491];
    assign layer5_out[145] = ~layer4_out[228] | layer4_out[229];
    assign layer5_out[146] = ~layer4_out[114];
    assign layer5_out[147] = ~layer4_out[518];
    assign layer5_out[148] = layer4_out[256];
    assign layer5_out[149] = layer4_out[16] & ~layer4_out[15];
    assign layer5_out[150] = layer4_out[365] & layer4_out[366];
    assign layer5_out[151] = layer4_out[389];
    assign layer5_out[152] = ~(layer4_out[112] | layer4_out[113]);
    assign layer5_out[153] = layer4_out[236];
    assign layer5_out[154] = ~(layer4_out[280] & layer4_out[281]);
    assign layer5_out[155] = layer4_out[362];
    assign layer5_out[156] = ~layer4_out[112];
    assign layer5_out[157] = ~layer4_out[27];
    assign layer5_out[158] = ~layer4_out[192];
    assign layer5_out[159] = ~layer4_out[382];
    assign layer5_out[160] = ~layer4_out[342] | layer4_out[341];
    assign layer5_out[161] = layer4_out[98];
    assign layer5_out[162] = layer4_out[390] | layer4_out[391];
    assign layer5_out[163] = layer4_out[152] & layer4_out[153];
    assign layer5_out[164] = ~(layer4_out[478] ^ layer4_out[479]);
    assign layer5_out[165] = layer4_out[491] & layer4_out[492];
    assign layer5_out[166] = layer4_out[379];
    assign layer5_out[167] = layer4_out[40] & ~layer4_out[41];
    assign layer5_out[168] = layer4_out[372];
    assign layer5_out[169] = layer4_out[149] | layer4_out[150];
    assign layer5_out[170] = layer4_out[28] & ~layer4_out[27];
    assign layer5_out[171] = layer4_out[257] & ~layer4_out[256];
    assign layer5_out[172] = ~layer4_out[155];
    assign layer5_out[173] = layer4_out[179];
    assign layer5_out[174] = ~layer4_out[326] | layer4_out[327];
    assign layer5_out[175] = layer4_out[519];
    assign layer5_out[176] = layer4_out[67];
    assign layer5_out[177] = ~layer4_out[397];
    assign layer5_out[178] = layer4_out[307] & ~layer4_out[308];
    assign layer5_out[179] = layer4_out[145] & ~layer4_out[146];
    assign layer5_out[180] = layer4_out[359];
    assign layer5_out[181] = layer4_out[401];
    assign layer5_out[182] = layer4_out[495] ^ layer4_out[496];
    assign layer5_out[183] = layer4_out[72];
    assign layer5_out[184] = layer4_out[303];
    assign layer5_out[185] = ~layer4_out[35];
    assign layer5_out[186] = layer4_out[142] & ~layer4_out[141];
    assign layer5_out[187] = layer4_out[379] & ~layer4_out[380];
    assign layer5_out[188] = ~layer4_out[212];
    assign layer5_out[189] = ~layer4_out[71];
    assign layer5_out[190] = ~layer4_out[273];
    assign layer5_out[191] = layer4_out[489] & layer4_out[490];
    assign layer5_out[192] = layer4_out[126];
    assign layer5_out[193] = layer4_out[84] & layer4_out[85];
    assign layer5_out[194] = ~layer4_out[404];
    assign layer5_out[195] = ~layer4_out[38];
    assign layer5_out[196] = ~layer4_out[97];
    assign layer5_out[197] = layer4_out[343] & layer4_out[344];
    assign layer5_out[198] = layer4_out[169] & layer4_out[170];
    assign layer5_out[199] = ~layer4_out[535];
    assign layer5_out[200] = layer4_out[431] & layer4_out[432];
    assign layer5_out[201] = ~layer4_out[190];
    assign layer5_out[202] = ~(layer4_out[538] & layer4_out[539]);
    assign layer5_out[203] = ~layer4_out[83];
    assign layer5_out[204] = layer4_out[80] & ~layer4_out[79];
    assign layer5_out[205] = layer4_out[160] & layer4_out[161];
    assign layer5_out[206] = layer4_out[548];
    assign layer5_out[207] = ~(layer4_out[174] | layer4_out[175]);
    assign layer5_out[208] = layer4_out[454];
    assign layer5_out[209] = ~layer4_out[35];
    assign layer5_out[210] = layer4_out[63] & ~layer4_out[62];
    assign layer5_out[211] = ~layer4_out[521];
    assign layer5_out[212] = layer4_out[540] & ~layer4_out[541];
    assign layer5_out[213] = ~layer4_out[32];
    assign layer5_out[214] = layer4_out[413];
    assign layer5_out[215] = ~layer4_out[456];
    assign layer5_out[216] = ~(layer4_out[61] | layer4_out[62]);
    assign layer5_out[217] = layer4_out[151] & layer4_out[152];
    assign layer5_out[218] = layer4_out[536];
    assign layer5_out[219] = ~layer4_out[138];
    assign layer5_out[220] = ~layer4_out[428];
    assign layer5_out[221] = layer4_out[317];
    assign layer5_out[222] = layer4_out[203] & ~layer4_out[204];
    assign layer5_out[223] = ~layer4_out[177];
    assign layer5_out[224] = layer4_out[516];
    assign layer5_out[225] = layer4_out[128];
    assign layer5_out[226] = layer4_out[42] & layer4_out[43];
    assign layer5_out[227] = ~layer4_out[305];
    assign layer5_out[228] = ~layer4_out[122];
    assign layer5_out[229] = layer4_out[484];
    assign layer5_out[230] = ~layer4_out[498];
    assign layer5_out[231] = layer4_out[300] & ~layer4_out[301];
    assign layer5_out[232] = ~layer4_out[310];
    assign layer5_out[233] = layer4_out[358];
    assign layer5_out[234] = ~layer4_out[402];
    assign layer5_out[235] = ~layer4_out[461];
    assign layer5_out[236] = layer4_out[15];
    assign layer5_out[237] = ~(layer4_out[210] | layer4_out[211]);
    assign layer5_out[238] = layer4_out[323];
    assign layer5_out[239] = ~layer4_out[422] | layer4_out[423];
    assign layer5_out[240] = layer4_out[171] & ~layer4_out[172];
    assign layer5_out[241] = layer4_out[108];
    assign layer5_out[242] = layer4_out[208] & ~layer4_out[207];
    assign layer5_out[243] = ~layer4_out[472];
    assign layer5_out[244] = ~(layer4_out[386] | layer4_out[387]);
    assign layer5_out[245] = layer4_out[346];
    assign layer5_out[246] = layer4_out[74] & ~layer4_out[75];
    assign layer5_out[247] = layer4_out[12];
    assign layer5_out[248] = ~(layer4_out[477] ^ layer4_out[478]);
    assign layer5_out[249] = ~layer4_out[376];
    assign layer5_out[250] = ~layer4_out[187];
    assign layer5_out[251] = layer4_out[6] & ~layer4_out[7];
    assign layer5_out[252] = layer4_out[458] & layer4_out[459];
    assign layer5_out[253] = ~layer4_out[376];
    assign layer5_out[254] = ~layer4_out[292];
    assign layer5_out[255] = ~layer4_out[220];
    assign layer5_out[256] = ~layer4_out[292];
    assign layer5_out[257] = ~(layer4_out[157] ^ layer4_out[158]);
    assign layer5_out[258] = layer4_out[523];
    assign layer5_out[259] = layer4_out[263];
    assign layer5_out[260] = layer4_out[186] & ~layer4_out[185];
    assign layer5_out[261] = layer4_out[470];
    assign layer5_out[262] = ~layer4_out[546];
    assign layer5_out[263] = layer4_out[56];
    assign layer5_out[264] = ~layer4_out[230];
    assign layer5_out[265] = ~layer4_out[4];
    assign layer5_out[266] = layer4_out[488] & ~layer4_out[489];
    assign layer5_out[267] = ~layer4_out[500];
    assign layer5_out[268] = ~layer4_out[278] | layer4_out[277];
    assign layer5_out[269] = layer4_out[467] & layer4_out[468];
    assign layer5_out[270] = layer4_out[449];
    assign layer5_out[271] = ~layer4_out[200];
    assign layer5_out[272] = layer4_out[258] | layer4_out[259];
    assign layer5_out[273] = layer4_out[288] & layer4_out[289];
    assign layer5_out[274] = layer4_out[220] ^ layer4_out[221];
    assign layer5_out[275] = ~layer4_out[255];
    assign layer5_out[276] = layer4_out[181];
    assign layer5_out[277] = ~layer4_out[458];
    assign layer5_out[278] = ~layer4_out[309];
    assign layer5_out[279] = ~layer4_out[39];
    assign layer5_out[280] = layer4_out[83] & layer4_out[84];
    assign layer5_out[281] = layer4_out[133];
    assign layer5_out[282] = ~layer4_out[354];
    assign layer5_out[283] = layer4_out[89];
    assign layer5_out[284] = layer4_out[406];
    assign layer5_out[285] = layer4_out[494];
    assign layer5_out[286] = layer4_out[409];
    assign layer5_out[287] = layer4_out[503] & ~layer4_out[504];
    assign layer5_out[288] = layer4_out[119] & ~layer4_out[118];
    assign layer5_out[289] = ~layer4_out[110];
    assign layer5_out[290] = layer4_out[250] ^ layer4_out[251];
    assign layer5_out[291] = ~layer4_out[335];
    assign layer5_out[292] = layer4_out[89];
    assign layer5_out[293] = ~layer4_out[512];
    assign layer5_out[294] = ~(layer4_out[229] | layer4_out[230]);
    assign layer5_out[295] = ~(layer4_out[28] ^ layer4_out[29]);
    assign layer5_out[296] = ~layer4_out[173];
    assign layer5_out[297] = layer4_out[368] & ~layer4_out[369];
    assign layer5_out[298] = ~layer4_out[110];
    assign layer5_out[299] = layer4_out[537];
    assign layer5_out[300] = layer4_out[223] & layer4_out[224];
    assign layer5_out[301] = ~(layer4_out[388] | layer4_out[389]);
    assign layer5_out[302] = layer4_out[315] | layer4_out[316];
    assign layer5_out[303] = ~(layer4_out[289] & layer4_out[290]);
    assign layer5_out[304] = ~layer4_out[412];
    assign layer5_out[305] = layer4_out[419] | layer4_out[420];
    assign layer5_out[306] = ~layer4_out[428];
    assign layer5_out[307] = layer4_out[100];
    assign layer5_out[308] = layer4_out[320];
    assign layer5_out[309] = ~layer4_out[105];
    assign layer5_out[310] = ~(layer4_out[21] ^ layer4_out[22]);
    assign layer5_out[311] = ~(layer4_out[276] | layer4_out[277]);
    assign layer5_out[312] = layer4_out[500] | layer4_out[501];
    assign layer5_out[313] = ~layer4_out[378];
    assign layer5_out[314] = ~(layer4_out[294] ^ layer4_out[295]);
    assign layer5_out[315] = ~(layer4_out[143] | layer4_out[144]);
    assign layer5_out[316] = layer4_out[168];
    assign layer5_out[317] = ~(layer4_out[445] ^ layer4_out[446]);
    assign layer5_out[318] = layer4_out[202] & layer4_out[203];
    assign layer5_out[319] = ~layer4_out[244] | layer4_out[245];
    assign layer5_out[320] = layer4_out[424];
    assign layer5_out[321] = layer4_out[547];
    assign layer5_out[322] = layer4_out[131] ^ layer4_out[132];
    assign layer5_out[323] = ~layer4_out[219];
    assign layer5_out[324] = layer4_out[347];
    assign layer5_out[325] = ~layer4_out[3];
    assign layer5_out[326] = layer4_out[34] & ~layer4_out[33];
    assign layer5_out[327] = layer4_out[352] & ~layer4_out[353];
    assign layer5_out[328] = layer4_out[264] & ~layer4_out[265];
    assign layer5_out[329] = ~layer4_out[392];
    assign layer5_out[330] = ~(layer4_out[208] | layer4_out[209]);
    assign layer5_out[331] = layer4_out[407];
    assign layer5_out[332] = layer4_out[68];
    assign layer5_out[333] = ~layer4_out[169];
    assign layer5_out[334] = layer4_out[429] & layer4_out[430];
    assign layer5_out[335] = ~layer4_out[63];
    assign layer5_out[336] = layer4_out[151];
    assign layer5_out[337] = layer4_out[399];
    assign layer5_out[338] = layer4_out[78];
    assign layer5_out[339] = layer4_out[93];
    assign layer5_out[340] = layer4_out[139];
    assign layer5_out[341] = layer4_out[497] & ~layer4_out[496];
    assign layer5_out[342] = ~layer4_out[287];
    assign layer5_out[343] = layer4_out[443] & ~layer4_out[444];
    assign layer5_out[344] = layer4_out[328] & layer4_out[329];
    assign layer5_out[345] = ~(layer4_out[367] ^ layer4_out[368]);
    assign layer5_out[346] = ~(layer4_out[37] ^ layer4_out[38]);
    assign layer5_out[347] = layer4_out[243] & ~layer4_out[242];
    assign layer5_out[348] = layer4_out[397];
    assign layer5_out[349] = layer4_out[351] ^ layer4_out[352];
    assign layer5_out[350] = layer4_out[269] | layer4_out[270];
    assign layer5_out[351] = layer4_out[181] & layer4_out[182];
    assign layer5_out[352] = ~layer4_out[166];
    assign layer5_out[353] = ~(layer4_out[156] | layer4_out[157]);
    assign layer5_out[354] = layer4_out[141];
    assign layer5_out[355] = ~layer4_out[225];
    assign layer5_out[356] = layer4_out[95] & ~layer4_out[96];
    assign layer5_out[357] = layer4_out[462] & ~layer4_out[463];
    assign layer5_out[358] = ~layer4_out[247];
    assign layer5_out[359] = layer4_out[312] & layer4_out[313];
    assign layer5_out[360] = layer4_out[343] & ~layer4_out[342];
    assign layer5_out[361] = ~(layer4_out[161] | layer4_out[162]);
    assign layer5_out[362] = layer4_out[511] & layer4_out[512];
    assign layer5_out[363] = ~layer4_out[325];
    assign layer5_out[364] = layer4_out[10];
    assign layer5_out[365] = layer4_out[423] ^ layer4_out[424];
    assign layer5_out[366] = layer4_out[399];
    assign layer5_out[367] = layer4_out[466] & layer4_out[467];
    assign layer5_out[368] = ~layer4_out[350];
    assign layer5_out[369] = ~(layer4_out[216] | layer4_out[217]);
    assign layer5_out[370] = ~layer4_out[307];
    assign layer5_out[371] = ~(layer4_out[122] ^ layer4_out[123]);
    assign layer5_out[372] = ~layer4_out[82];
    assign layer5_out[373] = ~(layer4_out[369] | layer4_out[370]);
    assign layer5_out[374] = ~(layer4_out[410] | layer4_out[411]);
    assign layer5_out[375] = layer4_out[257] | layer4_out[258];
    assign layer5_out[376] = ~layer4_out[237];
    assign layer5_out[377] = layer4_out[440];
    assign layer5_out[378] = ~(layer4_out[363] | layer4_out[364]);
    assign layer5_out[379] = layer4_out[542];
    assign layer5_out[380] = layer4_out[509] & layer4_out[510];
    assign layer5_out[381] = layer4_out[65];
    assign layer5_out[382] = ~(layer4_out[146] ^ layer4_out[147]);
    assign layer5_out[383] = layer4_out[227];
    assign layer5_out[384] = ~layer4_out[436];
    assign layer5_out[385] = layer4_out[66];
    assign layer5_out[386] = ~layer4_out[455];
    assign layer5_out[387] = ~layer4_out[518] | layer4_out[519];
    assign layer5_out[388] = ~(layer4_out[50] ^ layer4_out[51]);
    assign layer5_out[389] = ~layer4_out[216];
    assign layer5_out[390] = ~layer4_out[443];
    assign layer5_out[391] = layer4_out[266] ^ layer4_out[267];
    assign layer5_out[392] = layer4_out[330] & ~layer4_out[329];
    assign layer5_out[393] = layer4_out[190] & ~layer4_out[191];
    assign layer5_out[394] = layer4_out[1] & ~layer4_out[2];
    assign layer5_out[395] = layer4_out[301];
    assign layer5_out[396] = layer4_out[70] & ~layer4_out[69];
    assign layer5_out[397] = layer4_out[501] & layer4_out[502];
    assign layer5_out[398] = layer4_out[327];
    assign layer5_out[399] = ~(layer4_out[194] | layer4_out[195]);
    assign layer5_out[400] = ~layer4_out[107] | layer4_out[106];
    assign layer5_out[401] = layer4_out[43] & ~layer4_out[44];
    assign layer5_out[402] = ~layer4_out[103];
    assign layer5_out[403] = layer4_out[290];
    assign layer5_out[404] = ~layer4_out[482];
    assign layer5_out[405] = layer4_out[456] & ~layer4_out[457];
    assign layer5_out[406] = ~layer4_out[17];
    assign layer5_out[407] = ~(layer4_out[298] & layer4_out[299]);
    assign layer5_out[408] = ~layer4_out[525];
    assign layer5_out[409] = layer4_out[1];
    assign layer5_out[410] = layer4_out[143];
    assign layer5_out[411] = ~layer4_out[407];
    assign layer5_out[412] = layer4_out[87] & layer4_out[88];
    assign layer5_out[413] = ~(layer4_out[524] | layer4_out[525]);
    assign layer5_out[414] = layer4_out[272];
    assign layer5_out[415] = ~(layer4_out[497] | layer4_out[498]);
    assign layer5_out[416] = layer4_out[118];
    assign layer5_out[417] = ~(layer4_out[506] | layer4_out[507]);
    assign layer5_out[418] = layer4_out[58] | layer4_out[59];
    assign layer5_out[419] = layer4_out[48];
    assign layer5_out[420] = ~(layer4_out[505] | layer4_out[506]);
    assign layer5_out[421] = layer4_out[52] & layer4_out[53];
    assign layer5_out[422] = layer4_out[416] & layer4_out[417];
    assign layer5_out[423] = ~layer4_out[542];
    assign layer5_out[424] = ~layer4_out[466];
    assign layer5_out[425] = layer4_out[87] & ~layer4_out[86];
    assign layer5_out[426] = ~(layer4_out[385] | layer4_out[386]);
    assign layer5_out[427] = layer4_out[155] & ~layer4_out[154];
    assign layer5_out[428] = layer4_out[418] | layer4_out[419];
    assign layer5_out[429] = ~(layer4_out[313] & layer4_out[314]);
    assign layer5_out[430] = layer4_out[436] & layer4_out[437];
    assign layer5_out[431] = layer4_out[438] & ~layer4_out[439];
    assign layer5_out[432] = layer4_out[300];
    assign layer5_out[433] = ~layer4_out[452];
    assign layer5_out[434] = layer4_out[361];
    assign layer5_out[435] = layer4_out[416] & ~layer4_out[415];
    assign layer5_out[436] = ~layer4_out[170];
    assign layer5_out[437] = ~layer4_out[30];
    assign layer5_out[438] = layer4_out[322] & ~layer4_out[321];
    assign layer5_out[439] = layer4_out[148];
    assign layer5_out[440] = ~(layer4_out[319] | layer4_out[320]);
    assign layer5_out[441] = layer4_out[282] | layer4_out[283];
    assign layer5_out[442] = layer4_out[385];
    assign layer5_out[443] = layer4_out[197] & layer4_out[198];
    assign layer5_out[444] = ~layer4_out[253];
    assign layer5_out[445] = ~layer4_out[17];
    assign layer5_out[446] = layer4_out[80] & ~layer4_out[81];
    assign layer5_out[447] = ~(layer4_out[535] | layer4_out[536]);
    assign layer5_out[448] = layer4_out[97];
    assign layer5_out[449] = ~(layer4_out[433] | layer4_out[434]);
    assign layer5_out[450] = ~layer4_out[387];
    assign layer5_out[451] = layer4_out[240] & ~layer4_out[239];
    assign layer5_out[452] = layer4_out[363];
    assign layer5_out[453] = layer4_out[445];
    assign layer5_out[454] = ~layer4_out[261];
    assign layer5_out[455] = layer4_out[174];
    assign layer5_out[456] = ~(layer4_out[434] | layer4_out[435]);
    assign layer5_out[457] = ~layer4_out[348];
    assign layer5_out[458] = layer4_out[92];
    assign layer5_out[459] = layer4_out[492] & ~layer4_out[493];
    assign layer5_out[460] = ~(layer4_out[260] | layer4_out[261]);
    assign layer5_out[461] = layer4_out[13];
    assign layer5_out[462] = layer4_out[438] & ~layer4_out[437];
    assign layer5_out[463] = layer4_out[137] & layer4_out[138];
    assign layer5_out[464] = layer4_out[179] & ~layer4_out[180];
    assign layer5_out[465] = layer4_out[426] & ~layer4_out[427];
    assign layer5_out[466] = layer4_out[147];
    assign layer5_out[467] = layer4_out[350];
    assign layer5_out[468] = ~layer4_out[274];
    assign layer5_out[469] = ~layer4_out[309] | layer4_out[308];
    assign layer5_out[470] = layer4_out[282];
    assign layer5_out[471] = ~(layer4_out[336] ^ layer4_out[337]);
    assign layer5_out[472] = layer4_out[119] & layer4_out[120];
    assign layer5_out[473] = ~(layer4_out[164] | layer4_out[165]);
    assign layer5_out[474] = layer4_out[432] & ~layer4_out[433];
    assign layer5_out[475] = ~layer4_out[471];
    assign layer5_out[476] = ~layer4_out[464];
    assign layer5_out[477] = ~layer4_out[184];
    assign layer5_out[478] = ~layer4_out[231];
    assign layer5_out[479] = layer4_out[279] & layer4_out[280];
    assign layer5_out[480] = layer4_out[267] ^ layer4_out[268];
    assign layer5_out[481] = ~layer4_out[184];
    assign layer5_out[482] = layer4_out[366] ^ layer4_out[367];
    assign layer5_out[483] = layer4_out[382] & ~layer4_out[383];
    assign layer5_out[484] = ~layer4_out[414];
    assign layer5_out[485] = layer4_out[507] | layer4_out[508];
    assign layer5_out[486] = layer4_out[402] & ~layer4_out[401];
    assign layer5_out[487] = layer4_out[505];
    assign layer5_out[488] = layer4_out[240] & ~layer4_out[241];
    assign layer5_out[489] = layer4_out[129];
    assign layer5_out[490] = ~layer4_out[49];
    assign layer5_out[491] = layer4_out[189] & ~layer4_out[188];
    assign layer5_out[492] = layer4_out[72];
    assign layer5_out[493] = layer4_out[77] & ~layer4_out[78];
    assign layer5_out[494] = ~layer4_out[479];
    assign layer5_out[495] = layer4_out[56] & ~layer4_out[55];
    assign layer5_out[496] = layer4_out[127];
    assign layer5_out[497] = layer4_out[338];
    assign layer5_out[498] = layer4_out[340] & ~layer4_out[341];
    assign layer5_out[499] = layer4_out[468] & layer4_out[469];
    assign layer5_out[500] = ~(layer4_out[450] ^ layer4_out[451]);
    assign layer5_out[501] = layer4_out[374] & layer4_out[375];
    assign layer5_out[502] = ~layer4_out[202];
    assign layer5_out[503] = layer4_out[163] & ~layer4_out[164];
    assign layer5_out[504] = layer4_out[441] & layer4_out[442];
    assign layer5_out[505] = ~layer4_out[153];
    assign layer5_out[506] = layer4_out[188] & ~layer4_out[187];
    assign layer5_out[507] = layer4_out[314] & ~layer4_out[315];
    assign layer5_out[508] = layer4_out[486];
    assign layer5_out[509] = layer4_out[333];
    assign layer5_out[510] = layer4_out[115];
    assign layer5_out[511] = ~layer4_out[25];
    assign layer5_out[512] = layer4_out[373] & layer4_out[374];
    assign layer5_out[513] = layer4_out[90];
    assign layer5_out[514] = ~(layer4_out[508] | layer4_out[509]);
    assign layer5_out[515] = layer4_out[295] & ~layer4_out[296];
    assign layer5_out[516] = ~(layer4_out[293] ^ layer4_out[294]);
    assign layer5_out[517] = layer4_out[355];
    assign layer5_out[518] = ~layer4_out[55];
    assign layer5_out[519] = ~layer4_out[182];
    assign layer5_out[520] = ~(layer4_out[232] ^ layer4_out[233]);
    assign layer5_out[521] = layer4_out[235] & ~layer4_out[234];
    assign layer5_out[522] = layer4_out[271] & ~layer4_out[270];
    assign layer5_out[523] = ~layer4_out[30] | layer4_out[31];
    assign layer5_out[524] = layer4_out[250];
    assign layer5_out[525] = ~layer4_out[529];
    assign layer5_out[526] = layer4_out[502] & layer4_out[503];
    assign layer5_out[527] = ~layer4_out[5];
    assign layer5_out[528] = ~layer4_out[422];
    assign layer5_out[529] = ~layer4_out[285];
    assign layer5_out[530] = ~layer4_out[210];
    assign layer5_out[531] = layer4_out[24] & ~layer4_out[25];
    assign layer5_out[532] = ~(layer4_out[0] | layer4_out[2]);
    assign layer5_out[533] = layer4_out[163] & ~layer4_out[162];
    assign layer5_out[534] = layer4_out[516];
    assign layer5_out[535] = layer4_out[287] & ~layer4_out[288];
    assign layer5_out[536] = ~(layer4_out[323] & layer4_out[324]);
    assign layer5_out[537] = layer4_out[130] & ~layer4_out[131];
    assign layer5_out[538] = layer4_out[215];
    assign layer5_out[539] = layer4_out[483] | layer4_out[484];
    assign layer5_out[540] = ~(layer4_out[93] | layer4_out[94]);
    assign layer5_out[541] = layer4_out[192] & ~layer4_out[191];
    assign layer5_out[542] = layer4_out[344];
    assign layer5_out[543] = ~(layer4_out[221] ^ layer4_out[222]);
    assign layer5_out[544] = layer4_out[263];
    assign layer5_out[545] = ~layer4_out[176];
    assign layer5_out[546] = ~(layer4_out[522] | layer4_out[523]);
    assign layer5_out[547] = layer4_out[227] ^ layer4_out[228];
    assign layer5_out[548] = layer4_out[298];
    assign layer5_out[549] = layer4_out[251] ^ layer4_out[252];
      wire [549:0] last_layer_output;
      assign last_layer_output = layer5_out;
      wire [5:0] result [9:0];

      assign result[0] = last_layer_output[0] + last_layer_output[1] + last_layer_output[2] + last_layer_output[3] + last_layer_output[4] + last_layer_output[5] + last_layer_output[6] + last_layer_output[7] + last_layer_output[8] + last_layer_output[9] + last_layer_output[10] + last_layer_output[11] + last_layer_output[12] + last_layer_output[13] + last_layer_output[14] + last_layer_output[15] + last_layer_output[16] + last_layer_output[17] + last_layer_output[18] + last_layer_output[19] + last_layer_output[20] + last_layer_output[21] + last_layer_output[22] + last_layer_output[23] + last_layer_output[24] + last_layer_output[25] + last_layer_output[26] + last_layer_output[27] + last_layer_output[28] + last_layer_output[29] + last_layer_output[30] + last_layer_output[31] + last_layer_output[32] + last_layer_output[33] + last_layer_output[34] + last_layer_output[35] + last_layer_output[36] + last_layer_output[37] + last_layer_output[38] + last_layer_output[39] + last_layer_output[40] + last_layer_output[41] + last_layer_output[42] + last_layer_output[43] + last_layer_output[44] + last_layer_output[45] + last_layer_output[46] + last_layer_output[47] + last_layer_output[48] + last_layer_output[49] + last_layer_output[50] + last_layer_output[51] + last_layer_output[52] + last_layer_output[53] + last_layer_output[54];
      assign result[1] = last_layer_output[55] + last_layer_output[56] + last_layer_output[57] + last_layer_output[58] + last_layer_output[59] + last_layer_output[60] + last_layer_output[61] + last_layer_output[62] + last_layer_output[63] + last_layer_output[64] + last_layer_output[65] + last_layer_output[66] + last_layer_output[67] + last_layer_output[68] + last_layer_output[69] + last_layer_output[70] + last_layer_output[71] + last_layer_output[72] + last_layer_output[73] + last_layer_output[74] + last_layer_output[75] + last_layer_output[76] + last_layer_output[77] + last_layer_output[78] + last_layer_output[79] + last_layer_output[80] + last_layer_output[81] + last_layer_output[82] + last_layer_output[83] + last_layer_output[84] + last_layer_output[85] + last_layer_output[86] + last_layer_output[87] + last_layer_output[88] + last_layer_output[89] + last_layer_output[90] + last_layer_output[91] + last_layer_output[92] + last_layer_output[93] + last_layer_output[94] + last_layer_output[95] + last_layer_output[96] + last_layer_output[97] + last_layer_output[98] + last_layer_output[99] + last_layer_output[100] + last_layer_output[101] + last_layer_output[102] + last_layer_output[103] + last_layer_output[104] + last_layer_output[105] + last_layer_output[106] + last_layer_output[107] + last_layer_output[108] + last_layer_output[109];
      assign result[2] = last_layer_output[110] + last_layer_output[111] + last_layer_output[112] + last_layer_output[113] + last_layer_output[114] + last_layer_output[115] + last_layer_output[116] + last_layer_output[117] + last_layer_output[118] + last_layer_output[119] + last_layer_output[120] + last_layer_output[121] + last_layer_output[122] + last_layer_output[123] + last_layer_output[124] + last_layer_output[125] + last_layer_output[126] + last_layer_output[127] + last_layer_output[128] + last_layer_output[129] + last_layer_output[130] + last_layer_output[131] + last_layer_output[132] + last_layer_output[133] + last_layer_output[134] + last_layer_output[135] + last_layer_output[136] + last_layer_output[137] + last_layer_output[138] + last_layer_output[139] + last_layer_output[140] + last_layer_output[141] + last_layer_output[142] + last_layer_output[143] + last_layer_output[144] + last_layer_output[145] + last_layer_output[146] + last_layer_output[147] + last_layer_output[148] + last_layer_output[149] + last_layer_output[150] + last_layer_output[151] + last_layer_output[152] + last_layer_output[153] + last_layer_output[154] + last_layer_output[155] + last_layer_output[156] + last_layer_output[157] + last_layer_output[158] + last_layer_output[159] + last_layer_output[160] + last_layer_output[161] + last_layer_output[162] + last_layer_output[163] + last_layer_output[164];
      assign result[3] = last_layer_output[165] + last_layer_output[166] + last_layer_output[167] + last_layer_output[168] + last_layer_output[169] + last_layer_output[170] + last_layer_output[171] + last_layer_output[172] + last_layer_output[173] + last_layer_output[174] + last_layer_output[175] + last_layer_output[176] + last_layer_output[177] + last_layer_output[178] + last_layer_output[179] + last_layer_output[180] + last_layer_output[181] + last_layer_output[182] + last_layer_output[183] + last_layer_output[184] + last_layer_output[185] + last_layer_output[186] + last_layer_output[187] + last_layer_output[188] + last_layer_output[189] + last_layer_output[190] + last_layer_output[191] + last_layer_output[192] + last_layer_output[193] + last_layer_output[194] + last_layer_output[195] + last_layer_output[196] + last_layer_output[197] + last_layer_output[198] + last_layer_output[199] + last_layer_output[200] + last_layer_output[201] + last_layer_output[202] + last_layer_output[203] + last_layer_output[204] + last_layer_output[205] + last_layer_output[206] + last_layer_output[207] + last_layer_output[208] + last_layer_output[209] + last_layer_output[210] + last_layer_output[211] + last_layer_output[212] + last_layer_output[213] + last_layer_output[214] + last_layer_output[215] + last_layer_output[216] + last_layer_output[217] + last_layer_output[218] + last_layer_output[219];
      assign result[4] = last_layer_output[220] + last_layer_output[221] + last_layer_output[222] + last_layer_output[223] + last_layer_output[224] + last_layer_output[225] + last_layer_output[226] + last_layer_output[227] + last_layer_output[228] + last_layer_output[229] + last_layer_output[230] + last_layer_output[231] + last_layer_output[232] + last_layer_output[233] + last_layer_output[234] + last_layer_output[235] + last_layer_output[236] + last_layer_output[237] + last_layer_output[238] + last_layer_output[239] + last_layer_output[240] + last_layer_output[241] + last_layer_output[242] + last_layer_output[243] + last_layer_output[244] + last_layer_output[245] + last_layer_output[246] + last_layer_output[247] + last_layer_output[248] + last_layer_output[249] + last_layer_output[250] + last_layer_output[251] + last_layer_output[252] + last_layer_output[253] + last_layer_output[254] + last_layer_output[255] + last_layer_output[256] + last_layer_output[257] + last_layer_output[258] + last_layer_output[259] + last_layer_output[260] + last_layer_output[261] + last_layer_output[262] + last_layer_output[263] + last_layer_output[264] + last_layer_output[265] + last_layer_output[266] + last_layer_output[267] + last_layer_output[268] + last_layer_output[269] + last_layer_output[270] + last_layer_output[271] + last_layer_output[272] + last_layer_output[273] + last_layer_output[274];
      assign result[5] = last_layer_output[275] + last_layer_output[276] + last_layer_output[277] + last_layer_output[278] + last_layer_output[279] + last_layer_output[280] + last_layer_output[281] + last_layer_output[282] + last_layer_output[283] + last_layer_output[284] + last_layer_output[285] + last_layer_output[286] + last_layer_output[287] + last_layer_output[288] + last_layer_output[289] + last_layer_output[290] + last_layer_output[291] + last_layer_output[292] + last_layer_output[293] + last_layer_output[294] + last_layer_output[295] + last_layer_output[296] + last_layer_output[297] + last_layer_output[298] + last_layer_output[299] + last_layer_output[300] + last_layer_output[301] + last_layer_output[302] + last_layer_output[303] + last_layer_output[304] + last_layer_output[305] + last_layer_output[306] + last_layer_output[307] + last_layer_output[308] + last_layer_output[309] + last_layer_output[310] + last_layer_output[311] + last_layer_output[312] + last_layer_output[313] + last_layer_output[314] + last_layer_output[315] + last_layer_output[316] + last_layer_output[317] + last_layer_output[318] + last_layer_output[319] + last_layer_output[320] + last_layer_output[321] + last_layer_output[322] + last_layer_output[323] + last_layer_output[324] + last_layer_output[325] + last_layer_output[326] + last_layer_output[327] + last_layer_output[328] + last_layer_output[329];
      assign result[6] = last_layer_output[330] + last_layer_output[331] + last_layer_output[332] + last_layer_output[333] + last_layer_output[334] + last_layer_output[335] + last_layer_output[336] + last_layer_output[337] + last_layer_output[338] + last_layer_output[339] + last_layer_output[340] + last_layer_output[341] + last_layer_output[342] + last_layer_output[343] + last_layer_output[344] + last_layer_output[345] + last_layer_output[346] + last_layer_output[347] + last_layer_output[348] + last_layer_output[349] + last_layer_output[350] + last_layer_output[351] + last_layer_output[352] + last_layer_output[353] + last_layer_output[354] + last_layer_output[355] + last_layer_output[356] + last_layer_output[357] + last_layer_output[358] + last_layer_output[359] + last_layer_output[360] + last_layer_output[361] + last_layer_output[362] + last_layer_output[363] + last_layer_output[364] + last_layer_output[365] + last_layer_output[366] + last_layer_output[367] + last_layer_output[368] + last_layer_output[369] + last_layer_output[370] + last_layer_output[371] + last_layer_output[372] + last_layer_output[373] + last_layer_output[374] + last_layer_output[375] + last_layer_output[376] + last_layer_output[377] + last_layer_output[378] + last_layer_output[379] + last_layer_output[380] + last_layer_output[381] + last_layer_output[382] + last_layer_output[383] + last_layer_output[384];
      assign result[7] = last_layer_output[385] + last_layer_output[386] + last_layer_output[387] + last_layer_output[388] + last_layer_output[389] + last_layer_output[390] + last_layer_output[391] + last_layer_output[392] + last_layer_output[393] + last_layer_output[394] + last_layer_output[395] + last_layer_output[396] + last_layer_output[397] + last_layer_output[398] + last_layer_output[399] + last_layer_output[400] + last_layer_output[401] + last_layer_output[402] + last_layer_output[403] + last_layer_output[404] + last_layer_output[405] + last_layer_output[406] + last_layer_output[407] + last_layer_output[408] + last_layer_output[409] + last_layer_output[410] + last_layer_output[411] + last_layer_output[412] + last_layer_output[413] + last_layer_output[414] + last_layer_output[415] + last_layer_output[416] + last_layer_output[417] + last_layer_output[418] + last_layer_output[419] + last_layer_output[420] + last_layer_output[421] + last_layer_output[422] + last_layer_output[423] + last_layer_output[424] + last_layer_output[425] + last_layer_output[426] + last_layer_output[427] + last_layer_output[428] + last_layer_output[429] + last_layer_output[430] + last_layer_output[431] + last_layer_output[432] + last_layer_output[433] + last_layer_output[434] + last_layer_output[435] + last_layer_output[436] + last_layer_output[437] + last_layer_output[438] + last_layer_output[439];
      assign result[8] = last_layer_output[440] + last_layer_output[441] + last_layer_output[442] + last_layer_output[443] + last_layer_output[444] + last_layer_output[445] + last_layer_output[446] + last_layer_output[447] + last_layer_output[448] + last_layer_output[449] + last_layer_output[450] + last_layer_output[451] + last_layer_output[452] + last_layer_output[453] + last_layer_output[454] + last_layer_output[455] + last_layer_output[456] + last_layer_output[457] + last_layer_output[458] + last_layer_output[459] + last_layer_output[460] + last_layer_output[461] + last_layer_output[462] + last_layer_output[463] + last_layer_output[464] + last_layer_output[465] + last_layer_output[466] + last_layer_output[467] + last_layer_output[468] + last_layer_output[469] + last_layer_output[470] + last_layer_output[471] + last_layer_output[472] + last_layer_output[473] + last_layer_output[474] + last_layer_output[475] + last_layer_output[476] + last_layer_output[477] + last_layer_output[478] + last_layer_output[479] + last_layer_output[480] + last_layer_output[481] + last_layer_output[482] + last_layer_output[483] + last_layer_output[484] + last_layer_output[485] + last_layer_output[486] + last_layer_output[487] + last_layer_output[488] + last_layer_output[489] + last_layer_output[490] + last_layer_output[491] + last_layer_output[492] + last_layer_output[493] + last_layer_output[494];
      assign result[9] = last_layer_output[495] + last_layer_output[496] + last_layer_output[497] + last_layer_output[498] + last_layer_output[499] + last_layer_output[500] + last_layer_output[501] + last_layer_output[502] + last_layer_output[503] + last_layer_output[504] + last_layer_output[505] + last_layer_output[506] + last_layer_output[507] + last_layer_output[508] + last_layer_output[509] + last_layer_output[510] + last_layer_output[511] + last_layer_output[512] + last_layer_output[513] + last_layer_output[514] + last_layer_output[515] + last_layer_output[516] + last_layer_output[517] + last_layer_output[518] + last_layer_output[519] + last_layer_output[520] + last_layer_output[521] + last_layer_output[522] + last_layer_output[523] + last_layer_output[524] + last_layer_output[525] + last_layer_output[526] + last_layer_output[527] + last_layer_output[528] + last_layer_output[529] + last_layer_output[530] + last_layer_output[531] + last_layer_output[532] + last_layer_output[533] + last_layer_output[534] + last_layer_output[535] + last_layer_output[536] + last_layer_output[537] + last_layer_output[538] + last_layer_output[539] + last_layer_output[540] + last_layer_output[541] + last_layer_output[542] + last_layer_output[543] + last_layer_output[544] + last_layer_output[545] + last_layer_output[546] + last_layer_output[547] + last_layer_output[548] + last_layer_output[549];
      assign y[59:55]=result[0];
      assign y[54:50]=result[1];
      assign y[49:45]=result[2];
      assign y[44:40]=result[3];
      assign y[39:35]=result[4];
      assign y[34:30]=result[5];
      assign y[29:25]=result[6];
      assign y[24:20]=result[7];
      assign y[19:15]=result[8];
      assign y[14:10]=result[9];
      assign y[9:5]=result[10];
      assign y[4:0]=result[11];
endmodule