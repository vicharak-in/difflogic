module logic_network (    input clk,
    input wire [399:0] x,
    output wire [79:0] y
);
      reg [1499:0] layer0_out = 0;
      reg [1499:0] layer1_out = 0;
      reg [1499:0] layer2_out = 0;
      reg [1499:0] layer3_out = 0;
      reg [1499:0] layer4_out = 0;
      reg [1499:0] layer5_out = 0;
      reg [1499:0] layer6_out = 0;
      reg [1499:0] layer7_out = 0;
      reg [1499:0] last_layer_output = 0;
      reg [7:0] result [9:0];
      always @(posedge clk) begin
     layer0_out[0] <= ~(x[156] | x[159]);
     layer0_out[1] <= ~(x[149] & x[151]);
     layer0_out[2] <= x[24] | x[26];
     layer0_out[3] <= ~x[22] | x[18];
     layer0_out[4] <= ~x[207];
     layer0_out[5] <= ~x[51] | x[50];
     layer0_out[6] <= x[189] | x[190];
     layer0_out[7] <= 1'b0;
     layer0_out[8] <= 1'b1;
     layer0_out[9] <= 1'b0;
     layer0_out[10] <= 1'b0;
     layer0_out[11] <= x[89] & x[91];
     layer0_out[12] <= ~x[348] | x[345];
     layer0_out[13] <= ~(x[303] | x[305]);
     layer0_out[14] <= x[317] & ~x[316];
     layer0_out[15] <= ~(x[223] | x[225]);
     layer0_out[16] <= x[388] & x[391];
     layer0_out[17] <= ~(x[78] ^ x[82]);
     layer0_out[18] <= 1'b0;
     layer0_out[19] <= ~x[322] | x[323];
     layer0_out[20] <= 1'b0;
     layer0_out[21] <= 1'b0;
     layer0_out[22] <= ~(x[329] | x[330]);
     layer0_out[23] <= x[155] | x[158];
     layer0_out[24] <= 1'b0;
     layer0_out[25] <= x[86] & x[90];
     layer0_out[26] <= x[218] & ~x[214];
     layer0_out[27] <= ~(x[164] | x[167]);
     layer0_out[28] <= ~x[363] | x[365];
     layer0_out[29] <= 1'b0;
     layer0_out[30] <= x[393] & ~x[391];
     layer0_out[31] <= ~(x[85] | x[86]);
     layer0_out[32] <= x[224] ^ x[228];
     layer0_out[33] <= 1'b0;
     layer0_out[34] <= x[392];
     layer0_out[35] <= x[348] | x[350];
     layer0_out[36] <= 1'b1;
     layer0_out[37] <= ~(x[38] | x[41]);
     layer0_out[38] <= ~(x[66] & x[70]);
     layer0_out[39] <= ~(x[265] | x[269]);
     layer0_out[40] <= ~x[234] | x[238];
     layer0_out[41] <= x[14] | x[16];
     layer0_out[42] <= x[94] ^ x[97];
     layer0_out[43] <= x[302] & ~x[299];
     layer0_out[44] <= x[128];
     layer0_out[45] <= 1'b0;
     layer0_out[46] <= 1'b1;
     layer0_out[47] <= x[84] & ~x[88];
     layer0_out[48] <= ~(x[261] ^ x[262]);
     layer0_out[49] <= x[295] | x[296];
     layer0_out[50] <= ~x[249];
     layer0_out[51] <= x[172] & ~x[171];
     layer0_out[52] <= x[159] & x[160];
     layer0_out[53] <= 1'b0;
     layer0_out[54] <= ~(x[340] & x[343]);
     layer0_out[55] <= ~(x[156] | x[158]);
     layer0_out[56] <= x[197] | x[200];
     layer0_out[57] <= x[276] & x[278];
     layer0_out[58] <= 1'b0;
     layer0_out[59] <= x[220] & ~x[222];
     layer0_out[60] <= x[36] & ~x[40];
     layer0_out[61] <= ~(x[298] | x[299]);
     layer0_out[62] <= x[215] | x[219];
     layer0_out[63] <= x[153] & ~x[152];
     layer0_out[64] <= x[248] | x[249];
     layer0_out[65] <= ~x[127] | x[123];
     layer0_out[66] <= x[175] | x[176];
     layer0_out[67] <= x[122] | x[123];
     layer0_out[68] <= 1'b0;
     layer0_out[69] <= x[92] & x[96];
     layer0_out[70] <= x[204] & ~x[205];
     layer0_out[71] <= x[0] ^ x[4];
     layer0_out[72] <= 1'b1;
     layer0_out[73] <= 1'b1;
     layer0_out[74] <= x[110] | x[112];
     layer0_out[75] <= ~(x[235] | x[237]);
     layer0_out[76] <= ~x[250];
     layer0_out[77] <= ~(x[340] | x[342]);
     layer0_out[78] <= ~(x[10] & x[13]);
     layer0_out[79] <= 1'b0;
     layer0_out[80] <= 1'b1;
     layer0_out[81] <= ~(x[250] | x[251]);
     layer0_out[82] <= x[227] & ~x[228];
     layer0_out[83] <= x[310] & x[312];
     layer0_out[84] <= x[180] & x[182];
     layer0_out[85] <= ~(x[367] | x[368]);
     layer0_out[86] <= ~x[95] | x[92];
     layer0_out[87] <= x[218] & ~x[215];
     layer0_out[88] <= ~(x[12] & x[16]);
     layer0_out[89] <= ~(x[193] | x[194]);
     layer0_out[90] <= x[26] & x[28];
     layer0_out[91] <= ~(x[203] | x[205]);
     layer0_out[92] <= 1'b1;
     layer0_out[93] <= ~x[299];
     layer0_out[94] <= x[307] & ~x[306];
     layer0_out[95] <= 1'b0;
     layer0_out[96] <= ~(x[104] | x[106]);
     layer0_out[97] <= 1'b1;
     layer0_out[98] <= ~x[39] | x[38];
     layer0_out[99] <= 1'b0;
     layer0_out[100] <= ~x[196] | x[192];
     layer0_out[101] <= ~x[181] | x[182];
     layer0_out[102] <= 1'b0;
     layer0_out[103] <= ~x[142];
     layer0_out[104] <= x[360] | x[362];
     layer0_out[105] <= ~x[289] | x[292];
     layer0_out[106] <= x[103] & ~x[105];
     layer0_out[107] <= 1'b1;
     layer0_out[108] <= ~x[336] | x[337];
     layer0_out[109] <= 1'b1;
     layer0_out[110] <= 1'b1;
     layer0_out[111] <= x[87] & x[88];
     layer0_out[112] <= ~(x[327] ^ x[329]);
     layer0_out[113] <= x[308] | x[311];
     layer0_out[114] <= 1'b0;
     layer0_out[115] <= x[138] | x[139];
     layer0_out[116] <= ~x[160];
     layer0_out[117] <= ~x[360];
     layer0_out[118] <= x[248];
     layer0_out[119] <= 1'b0;
     layer0_out[120] <= 1'b0;
     layer0_out[121] <= ~x[41] | x[43];
     layer0_out[122] <= 1'b0;
     layer0_out[123] <= 1'b0;
     layer0_out[124] <= 1'b0;
     layer0_out[125] <= ~(x[233] & x[236]);
     layer0_out[126] <= ~(x[94] | x[96]);
     layer0_out[127] <= 1'b1;
     layer0_out[128] <= 1'b0;
     layer0_out[129] <= x[217];
     layer0_out[130] <= x[232];
     layer0_out[131] <= ~(x[19] & x[21]);
     layer0_out[132] <= x[72];
     layer0_out[133] <= ~(x[26] | x[27]);
     layer0_out[134] <= ~x[170];
     layer0_out[135] <= ~(x[174] | x[176]);
     layer0_out[136] <= x[99] & ~x[98];
     layer0_out[137] <= ~x[252];
     layer0_out[138] <= ~x[262];
     layer0_out[139] <= 1'b0;
     layer0_out[140] <= x[290] ^ x[293];
     layer0_out[141] <= ~(x[214] | x[217]);
     layer0_out[142] <= 1'b0;
     layer0_out[143] <= ~(x[249] | x[250]);
     layer0_out[144] <= x[377] | x[380];
     layer0_out[145] <= ~x[333];
     layer0_out[146] <= ~(x[144] | x[148]);
     layer0_out[147] <= x[199] | x[202];
     layer0_out[148] <= ~(x[292] & x[294]);
     layer0_out[149] <= ~x[181] | x[178];
     layer0_out[150] <= 1'b1;
     layer0_out[151] <= ~x[173];
     layer0_out[152] <= 1'b0;
     layer0_out[153] <= x[277] & x[279];
     layer0_out[154] <= 1'b1;
     layer0_out[155] <= ~(x[267] | x[269]);
     layer0_out[156] <= 1'b1;
     layer0_out[157] <= x[283] | x[285];
     layer0_out[158] <= x[188] & x[191];
     layer0_out[159] <= 1'b1;
     layer0_out[160] <= 1'b0;
     layer0_out[161] <= ~(x[72] & x[75]);
     layer0_out[162] <= x[263] ^ x[264];
     layer0_out[163] <= ~(x[36] | x[39]);
     layer0_out[164] <= ~(x[335] | x[337]);
     layer0_out[165] <= ~x[91];
     layer0_out[166] <= x[371] & ~x[372];
     layer0_out[167] <= 1'b0;
     layer0_out[168] <= x[351] | x[352];
     layer0_out[169] <= x[354];
     layer0_out[170] <= x[138] | x[141];
     layer0_out[171] <= x[224] & ~x[221];
     layer0_out[172] <= ~(x[267] | x[268]);
     layer0_out[173] <= 1'b1;
     layer0_out[174] <= ~(x[132] & x[133]);
     layer0_out[175] <= 1'b1;
     layer0_out[176] <= x[63];
     layer0_out[177] <= ~x[200];
     layer0_out[178] <= 1'b1;
     layer0_out[179] <= ~x[216] | x[213];
     layer0_out[180] <= x[314] | x[315];
     layer0_out[181] <= 1'b1;
     layer0_out[182] <= ~(x[161] & x[164]);
     layer0_out[183] <= 1'b1;
     layer0_out[184] <= ~(x[1] | x[5]);
     layer0_out[185] <= x[120] & ~x[124];
     layer0_out[186] <= 1'b1;
     layer0_out[187] <= x[320] | x[322];
     layer0_out[188] <= ~(x[238] & x[240]);
     layer0_out[189] <= 1'b0;
     layer0_out[190] <= x[4] | x[5];
     layer0_out[191] <= ~x[109];
     layer0_out[192] <= x[322] | x[324];
     layer0_out[193] <= 1'b0;
     layer0_out[194] <= 1'b1;
     layer0_out[195] <= x[225];
     layer0_out[196] <= ~(x[17] & x[21]);
     layer0_out[197] <= 1'b1;
     layer0_out[198] <= x[300] | x[302];
     layer0_out[199] <= x[264] | x[266];
     layer0_out[200] <= x[117] & x[121];
     layer0_out[201] <= 1'b0;
     layer0_out[202] <= ~x[151] | x[152];
     layer0_out[203] <= x[83] & ~x[84];
     layer0_out[204] <= ~(x[273] | x[274]);
     layer0_out[205] <= ~(x[185] ^ x[188]);
     layer0_out[206] <= x[165] ^ x[166];
     layer0_out[207] <= x[276] & ~x[273];
     layer0_out[208] <= x[124] | x[126];
     layer0_out[209] <= x[109] & x[113];
     layer0_out[210] <= ~(x[119] & x[120]);
     layer0_out[211] <= x[197];
     layer0_out[212] <= ~(x[273] | x[275]);
     layer0_out[213] <= x[302] | x[303];
     layer0_out[214] <= ~(x[292] & x[296]);
     layer0_out[215] <= ~(x[17] | x[20]);
     layer0_out[216] <= ~(x[165] | x[167]);
     layer0_out[217] <= x[128];
     layer0_out[218] <= ~(x[345] | x[347]);
     layer0_out[219] <= ~(x[125] & x[127]);
     layer0_out[220] <= x[380] | x[383];
     layer0_out[221] <= ~x[372];
     layer0_out[222] <= x[190];
     layer0_out[223] <= x[98];
     layer0_out[224] <= ~x[152] | x[156];
     layer0_out[225] <= ~x[50];
     layer0_out[226] <= ~(x[379] & x[381]);
     layer0_out[227] <= 1'b0;
     layer0_out[228] <= ~(x[381] | x[382]);
     layer0_out[229] <= x[225] & ~x[221];
     layer0_out[230] <= x[57] | x[59];
     layer0_out[231] <= 1'b1;
     layer0_out[232] <= x[84] | x[85];
     layer0_out[233] <= x[391] & x[394];
     layer0_out[234] <= x[318] | x[321];
     layer0_out[235] <= 1'b1;
     layer0_out[236] <= 1'b1;
     layer0_out[237] <= x[243] ^ x[246];
     layer0_out[238] <= ~x[207] | x[210];
     layer0_out[239] <= ~x[129];
     layer0_out[240] <= x[148];
     layer0_out[241] <= 1'b0;
     layer0_out[242] <= x[76] | x[78];
     layer0_out[243] <= ~(x[81] | x[83]);
     layer0_out[244] <= x[386] & x[389];
     layer0_out[245] <= ~(x[364] | x[367]);
     layer0_out[246] <= x[60] | x[64];
     layer0_out[247] <= ~(x[8] | x[10]);
     layer0_out[248] <= x[69];
     layer0_out[249] <= ~x[79] | x[76];
     layer0_out[250] <= 1'b1;
     layer0_out[251] <= 1'b0;
     layer0_out[252] <= x[395] & ~x[397];
     layer0_out[253] <= ~x[259];
     layer0_out[254] <= ~(x[380] | x[381]);
     layer0_out[255] <= x[118] & x[119];
     layer0_out[256] <= 1'b1;
     layer0_out[257] <= x[196] | x[198];
     layer0_out[258] <= x[142] | x[144];
     layer0_out[259] <= x[181] | x[184];
     layer0_out[260] <= ~x[238];
     layer0_out[261] <= x[205] ^ x[209];
     layer0_out[262] <= ~(x[177] | x[179]);
     layer0_out[263] <= x[13] & ~x[17];
     layer0_out[264] <= ~(x[103] | x[107]);
     layer0_out[265] <= 1'b0;
     layer0_out[266] <= x[50];
     layer0_out[267] <= ~x[196];
     layer0_out[268] <= ~x[222];
     layer0_out[269] <= ~(x[195] | x[197]);
     layer0_out[270] <= ~(x[128] & x[131]);
     layer0_out[271] <= x[113] & x[116];
     layer0_out[272] <= x[266] | x[270];
     layer0_out[273] <= 1'b0;
     layer0_out[274] <= ~x[353] | x[350];
     layer0_out[275] <= 1'b0;
     layer0_out[276] <= x[376] & ~x[378];
     layer0_out[277] <= x[397] | x[399];
     layer0_out[278] <= ~(x[155] | x[156]);
     layer0_out[279] <= x[343] | x[344];
     layer0_out[280] <= 1'b0;
     layer0_out[281] <= 1'b0;
     layer0_out[282] <= x[372];
     layer0_out[283] <= 1'b0;
     layer0_out[284] <= x[375] | x[378];
     layer0_out[285] <= 1'b1;
     layer0_out[286] <= 1'b1;
     layer0_out[287] <= ~x[219];
     layer0_out[288] <= 1'b1;
     layer0_out[289] <= x[161];
     layer0_out[290] <= x[299] | x[300];
     layer0_out[291] <= x[243] & x[245];
     layer0_out[292] <= x[92] & ~x[94];
     layer0_out[293] <= x[72] | x[76];
     layer0_out[294] <= ~(x[343] | x[345]);
     layer0_out[295] <= x[34] | x[37];
     layer0_out[296] <= 1'b0;
     layer0_out[297] <= x[120] & ~x[118];
     layer0_out[298] <= 1'b0;
     layer0_out[299] <= 1'b0;
     layer0_out[300] <= 1'b0;
     layer0_out[301] <= ~(x[275] ^ x[278]);
     layer0_out[302] <= x[219] & ~x[217];
     layer0_out[303] <= x[181] | x[183];
     layer0_out[304] <= x[330] | x[333];
     layer0_out[305] <= x[29] & x[33];
     layer0_out[306] <= x[35] & ~x[33];
     layer0_out[307] <= x[349] & ~x[351];
     layer0_out[308] <= 1'b0;
     layer0_out[309] <= x[351] | x[354];
     layer0_out[310] <= x[171];
     layer0_out[311] <= 1'b1;
     layer0_out[312] <= ~(x[185] | x[186]);
     layer0_out[313] <= x[47] & x[51];
     layer0_out[314] <= 1'b1;
     layer0_out[315] <= 1'b1;
     layer0_out[316] <= x[366] & ~x[368];
     layer0_out[317] <= ~x[146] | x[142];
     layer0_out[318] <= ~(x[129] | x[132]);
     layer0_out[319] <= ~x[112];
     layer0_out[320] <= ~x[142];
     layer0_out[321] <= ~(x[226] | x[227]);
     layer0_out[322] <= x[222] | x[225];
     layer0_out[323] <= ~(x[153] | x[155]);
     layer0_out[324] <= ~(x[337] & x[340]);
     layer0_out[325] <= 1'b1;
     layer0_out[326] <= ~x[161];
     layer0_out[327] <= ~(x[247] | x[249]);
     layer0_out[328] <= x[40];
     layer0_out[329] <= ~(x[321] | x[324]);
     layer0_out[330] <= x[259];
     layer0_out[331] <= x[261] & x[265];
     layer0_out[332] <= 1'b1;
     layer0_out[333] <= x[154];
     layer0_out[334] <= ~(x[20] | x[22]);
     layer0_out[335] <= ~(x[75] & x[77]);
     layer0_out[336] <= ~x[190];
     layer0_out[337] <= x[54] & ~x[52];
     layer0_out[338] <= x[238] | x[242];
     layer0_out[339] <= x[341];
     layer0_out[340] <= x[378] | x[381];
     layer0_out[341] <= ~x[285] | x[282];
     layer0_out[342] <= x[30] | x[32];
     layer0_out[343] <= x[345] | x[346];
     layer0_out[344] <= 1'b0;
     layer0_out[345] <= x[80];
     layer0_out[346] <= x[288] & ~x[290];
     layer0_out[347] <= x[67] & x[71];
     layer0_out[348] <= x[80];
     layer0_out[349] <= 1'b0;
     layer0_out[350] <= 1'b1;
     layer0_out[351] <= x[71];
     layer0_out[352] <= ~x[191] | x[187];
     layer0_out[353] <= x[271] ^ x[275];
     layer0_out[354] <= ~x[150] | x[151];
     layer0_out[355] <= x[86] & ~x[82];
     layer0_out[356] <= 1'b0;
     layer0_out[357] <= ~(x[262] | x[263]);
     layer0_out[358] <= 1'b1;
     layer0_out[359] <= x[45] | x[47];
     layer0_out[360] <= x[100] | x[102];
     layer0_out[361] <= ~(x[394] ^ x[397]);
     layer0_out[362] <= ~(x[259] | x[262]);
     layer0_out[363] <= x[301];
     layer0_out[364] <= x[99];
     layer0_out[365] <= ~x[5] | x[9];
     layer0_out[366] <= ~x[227];
     layer0_out[367] <= 1'b1;
     layer0_out[368] <= ~(x[303] | x[304]);
     layer0_out[369] <= x[246] | x[249];
     layer0_out[370] <= x[372] & x[375];
     layer0_out[371] <= ~(x[169] & x[173]);
     layer0_out[372] <= ~(x[158] | x[162]);
     layer0_out[373] <= ~x[301];
     layer0_out[374] <= x[271];
     layer0_out[375] <= 1'b1;
     layer0_out[376] <= 1'b0;
     layer0_out[377] <= 1'b1;
     layer0_out[378] <= 1'b1;
     layer0_out[379] <= x[133] & ~x[135];
     layer0_out[380] <= ~(x[369] | x[370]);
     layer0_out[381] <= ~(x[103] | x[106]);
     layer0_out[382] <= x[212];
     layer0_out[383] <= ~x[240] | x[241];
     layer0_out[384] <= ~x[242] | x[241];
     layer0_out[385] <= x[319];
     layer0_out[386] <= 1'b1;
     layer0_out[387] <= x[272] ^ x[276];
     layer0_out[388] <= 1'b0;
     layer0_out[389] <= 1'b0;
     layer0_out[390] <= x[81] & ~x[82];
     layer0_out[391] <= x[233] | x[237];
     layer0_out[392] <= x[360] & ~x[357];
     layer0_out[393] <= 1'b0;
     layer0_out[394] <= 1'b1;
     layer0_out[395] <= x[287] | x[291];
     layer0_out[396] <= ~(x[142] | x[145]);
     layer0_out[397] <= ~x[263] | x[267];
     layer0_out[398] <= x[338] | x[341];
     layer0_out[399] <= x[63] | x[64];
     layer0_out[400] <= ~x[232] | x[231];
     layer0_out[401] <= ~x[254];
     layer0_out[402] <= x[248];
     layer0_out[403] <= x[189];
     layer0_out[404] <= ~(x[235] | x[239]);
     layer0_out[405] <= x[325] & ~x[326];
     layer0_out[406] <= ~x[59];
     layer0_out[407] <= x[172] | x[174];
     layer0_out[408] <= 1'b0;
     layer0_out[409] <= 1'b1;
     layer0_out[410] <= ~(x[150] & x[154]);
     layer0_out[411] <= ~(x[7] & x[8]);
     layer0_out[412] <= ~(x[91] & x[95]);
     layer0_out[413] <= x[34] | x[38];
     layer0_out[414] <= x[45] | x[49];
     layer0_out[415] <= ~(x[297] | x[300]);
     layer0_out[416] <= x[334] | x[335];
     layer0_out[417] <= 1'b0;
     layer0_out[418] <= ~(x[31] & x[33]);
     layer0_out[419] <= x[119];
     layer0_out[420] <= ~x[3];
     layer0_out[421] <= x[182] | x[186];
     layer0_out[422] <= 1'b1;
     layer0_out[423] <= x[275];
     layer0_out[424] <= x[120] | x[123];
     layer0_out[425] <= ~(x[374] | x[376]);
     layer0_out[426] <= 1'b1;
     layer0_out[427] <= x[2] | x[4];
     layer0_out[428] <= 1'b1;
     layer0_out[429] <= 1'b0;
     layer0_out[430] <= x[305];
     layer0_out[431] <= ~x[48];
     layer0_out[432] <= x[308];
     layer0_out[433] <= 1'b1;
     layer0_out[434] <= x[231] & ~x[229];
     layer0_out[435] <= 1'b1;
     layer0_out[436] <= ~(x[61] & x[64]);
     layer0_out[437] <= ~(x[149] & x[153]);
     layer0_out[438] <= ~x[295];
     layer0_out[439] <= x[124] | x[125];
     layer0_out[440] <= ~x[287] | x[288];
     layer0_out[441] <= x[157] & ~x[160];
     layer0_out[442] <= x[122] ^ x[125];
     layer0_out[443] <= 1'b1;
     layer0_out[444] <= ~x[159] | x[163];
     layer0_out[445] <= x[316];
     layer0_out[446] <= x[159] & x[162];
     layer0_out[447] <= x[219] | x[222];
     layer0_out[448] <= x[51] ^ x[53];
     layer0_out[449] <= x[235] & ~x[233];
     layer0_out[450] <= ~(x[229] ^ x[230]);
     layer0_out[451] <= 1'b1;
     layer0_out[452] <= ~(x[178] | x[179]);
     layer0_out[453] <= ~x[187];
     layer0_out[454] <= x[299] | x[301];
     layer0_out[455] <= 1'b1;
     layer0_out[456] <= 1'b1;
     layer0_out[457] <= ~(x[136] ^ x[137]);
     layer0_out[458] <= x[90] & x[93];
     layer0_out[459] <= x[18];
     layer0_out[460] <= ~x[58];
     layer0_out[461] <= x[53];
     layer0_out[462] <= ~x[180] | x[183];
     layer0_out[463] <= 1'b0;
     layer0_out[464] <= x[18] | x[21];
     layer0_out[465] <= ~x[95];
     layer0_out[466] <= x[163] | x[164];
     layer0_out[467] <= x[206] & ~x[207];
     layer0_out[468] <= ~x[241];
     layer0_out[469] <= x[180] & ~x[177];
     layer0_out[470] <= ~(x[236] | x[238]);
     layer0_out[471] <= x[309];
     layer0_out[472] <= 1'b1;
     layer0_out[473] <= ~(x[194] & x[197]);
     layer0_out[474] <= ~(x[371] ^ x[373]);
     layer0_out[475] <= ~x[314] | x[316];
     layer0_out[476] <= 1'b1;
     layer0_out[477] <= x[310] & x[313];
     layer0_out[478] <= 1'b0;
     layer0_out[479] <= ~x[53] | x[50];
     layer0_out[480] <= ~(x[20] & x[23]);
     layer0_out[481] <= ~x[244];
     layer0_out[482] <= x[67];
     layer0_out[483] <= ~x[384];
     layer0_out[484] <= x[153] | x[157];
     layer0_out[485] <= x[396] | x[397];
     layer0_out[486] <= ~x[311] | x[310];
     layer0_out[487] <= x[274] | x[276];
     layer0_out[488] <= ~(x[63] & x[66]);
     layer0_out[489] <= ~(x[392] | x[394]);
     layer0_out[490] <= x[26];
     layer0_out[491] <= ~x[1] | x[4];
     layer0_out[492] <= ~(x[243] ^ x[247]);
     layer0_out[493] <= x[216] | x[219];
     layer0_out[494] <= ~x[63];
     layer0_out[495] <= x[8] & x[11];
     layer0_out[496] <= 1'b1;
     layer0_out[497] <= ~x[59];
     layer0_out[498] <= ~x[93];
     layer0_out[499] <= 1'b0;
     layer0_out[500] <= x[314] & x[317];
     layer0_out[501] <= ~(x[217] | x[221]);
     layer0_out[502] <= x[325] | x[327];
     layer0_out[503] <= x[326] & ~x[324];
     layer0_out[504] <= ~(x[215] | x[216]);
     layer0_out[505] <= ~x[147];
     layer0_out[506] <= 1'b0;
     layer0_out[507] <= ~x[80];
     layer0_out[508] <= x[33] | x[37];
     layer0_out[509] <= ~(x[46] | x[48]);
     layer0_out[510] <= x[121] | x[124];
     layer0_out[511] <= x[88];
     layer0_out[512] <= x[78] & ~x[81];
     layer0_out[513] <= ~(x[194] | x[196]);
     layer0_out[514] <= x[283] ^ x[284];
     layer0_out[515] <= ~(x[200] | x[201]);
     layer0_out[516] <= 1'b0;
     layer0_out[517] <= ~(x[123] | x[125]);
     layer0_out[518] <= x[28];
     layer0_out[519] <= x[341] | x[342];
     layer0_out[520] <= ~x[370];
     layer0_out[521] <= ~(x[211] ^ x[215]);
     layer0_out[522] <= 1'b0;
     layer0_out[523] <= ~x[277] | x[273];
     layer0_out[524] <= x[136] & ~x[135];
     layer0_out[525] <= x[105] | x[106];
     layer0_out[526] <= ~x[157] | x[155];
     layer0_out[527] <= ~(x[327] ^ x[328]);
     layer0_out[528] <= ~(x[350] ^ x[352]);
     layer0_out[529] <= ~x[115] | x[111];
     layer0_out[530] <= 1'b0;
     layer0_out[531] <= ~(x[165] & x[169]);
     layer0_out[532] <= 1'b1;
     layer0_out[533] <= x[343] & x[346];
     layer0_out[534] <= x[384];
     layer0_out[535] <= ~x[173];
     layer0_out[536] <= x[381] & x[383];
     layer0_out[537] <= ~x[210];
     layer0_out[538] <= x[254] & x[257];
     layer0_out[539] <= 1'b0;
     layer0_out[540] <= x[139] ^ x[140];
     layer0_out[541] <= 1'b1;
     layer0_out[542] <= 1'b0;
     layer0_out[543] <= 1'b1;
     layer0_out[544] <= x[398];
     layer0_out[545] <= ~(x[208] | x[209]);
     layer0_out[546] <= x[111] | x[113];
     layer0_out[547] <= ~x[323];
     layer0_out[548] <= x[368] | x[370];
     layer0_out[549] <= x[223] & ~x[224];
     layer0_out[550] <= ~(x[263] | x[266]);
     layer0_out[551] <= 1'b1;
     layer0_out[552] <= 1'b1;
     layer0_out[553] <= 1'b0;
     layer0_out[554] <= 1'b1;
     layer0_out[555] <= x[17];
     layer0_out[556] <= x[44] | x[47];
     layer0_out[557] <= ~(x[120] | x[122]);
     layer0_out[558] <= x[234] | x[235];
     layer0_out[559] <= 1'b1;
     layer0_out[560] <= x[40] & ~x[38];
     layer0_out[561] <= x[118] & ~x[115];
     layer0_out[562] <= x[286] | x[289];
     layer0_out[563] <= x[191] | x[195];
     layer0_out[564] <= x[200] & ~x[204];
     layer0_out[565] <= x[272];
     layer0_out[566] <= ~x[39];
     layer0_out[567] <= x[334] & ~x[332];
     layer0_out[568] <= x[134] ^ x[138];
     layer0_out[569] <= 1'b0;
     layer0_out[570] <= x[307] & x[309];
     layer0_out[571] <= x[114] & x[116];
     layer0_out[572] <= 1'b1;
     layer0_out[573] <= x[259];
     layer0_out[574] <= x[231];
     layer0_out[575] <= x[243] & ~x[244];
     layer0_out[576] <= x[2] & x[6];
     layer0_out[577] <= x[182] | x[184];
     layer0_out[578] <= 1'b0;
     layer0_out[579] <= ~(x[148] | x[150]);
     layer0_out[580] <= 1'b1;
     layer0_out[581] <= ~(x[270] ^ x[271]);
     layer0_out[582] <= ~(x[289] & x[293]);
     layer0_out[583] <= 1'b1;
     layer0_out[584] <= ~x[212];
     layer0_out[585] <= ~(x[358] | x[361]);
     layer0_out[586] <= x[71] ^ x[74];
     layer0_out[587] <= x[66] | x[68];
     layer0_out[588] <= ~(x[147] ^ x[151]);
     layer0_out[589] <= ~(x[201] | x[203]);
     layer0_out[590] <= 1'b1;
     layer0_out[591] <= ~x[344] | x[342];
     layer0_out[592] <= ~x[233];
     layer0_out[593] <= 1'b0;
     layer0_out[594] <= 1'b1;
     layer0_out[595] <= 1'b0;
     layer0_out[596] <= x[315] ^ x[317];
     layer0_out[597] <= x[11] & ~x[12];
     layer0_out[598] <= ~(x[326] & x[328]);
     layer0_out[599] <= x[251] | x[253];
     layer0_out[600] <= ~x[173];
     layer0_out[601] <= 1'b0;
     layer0_out[602] <= x[182] | x[185];
     layer0_out[603] <= ~x[321];
     layer0_out[604] <= x[77] & x[80];
     layer0_out[605] <= x[247] | x[248];
     layer0_out[606] <= ~(x[177] | x[178]);
     layer0_out[607] <= 1'b1;
     layer0_out[608] <= x[112] | x[116];
     layer0_out[609] <= x[101] | x[104];
     layer0_out[610] <= 1'b0;
     layer0_out[611] <= 1'b1;
     layer0_out[612] <= x[34] | x[36];
     layer0_out[613] <= x[353] | x[355];
     layer0_out[614] <= x[132] | x[134];
     layer0_out[615] <= ~x[205];
     layer0_out[616] <= ~(x[303] | x[306]);
     layer0_out[617] <= ~(x[373] | x[375]);
     layer0_out[618] <= ~x[366];
     layer0_out[619] <= x[241] & x[245];
     layer0_out[620] <= x[21] & ~x[24];
     layer0_out[621] <= x[292] & ~x[293];
     layer0_out[622] <= x[342] & ~x[343];
     layer0_out[623] <= x[162] & x[166];
     layer0_out[624] <= x[280] & x[281];
     layer0_out[625] <= ~(x[370] | x[372]);
     layer0_out[626] <= 1'b1;
     layer0_out[627] <= ~x[258];
     layer0_out[628] <= ~(x[74] & x[76]);
     layer0_out[629] <= ~(x[30] | x[31]);
     layer0_out[630] <= 1'b1;
     layer0_out[631] <= ~(x[125] ^ x[128]);
     layer0_out[632] <= ~(x[239] & x[243]);
     layer0_out[633] <= ~x[301] | x[302];
     layer0_out[634] <= ~x[377];
     layer0_out[635] <= 1'b0;
     layer0_out[636] <= ~x[176] | x[179];
     layer0_out[637] <= ~(x[278] | x[281]);
     layer0_out[638] <= ~x[208];
     layer0_out[639] <= x[167] & ~x[163];
     layer0_out[640] <= x[20] & ~x[16];
     layer0_out[641] <= x[244];
     layer0_out[642] <= 1'b1;
     layer0_out[643] <= 1'b0;
     layer0_out[644] <= x[221] & x[223];
     layer0_out[645] <= x[254] ^ x[256];
     layer0_out[646] <= 1'b1;
     layer0_out[647] <= 1'b0;
     layer0_out[648] <= 1'b0;
     layer0_out[649] <= ~(x[64] & x[67]);
     layer0_out[650] <= x[73] | x[76];
     layer0_out[651] <= ~(x[44] & x[48]);
     layer0_out[652] <= x[320] | x[323];
     layer0_out[653] <= x[146] & ~x[144];
     layer0_out[654] <= x[395];
     layer0_out[655] <= x[228] | x[230];
     layer0_out[656] <= 1'b0;
     layer0_out[657] <= 1'b0;
     layer0_out[658] <= x[336];
     layer0_out[659] <= 1'b1;
     layer0_out[660] <= x[255] | x[257];
     layer0_out[661] <= ~x[227];
     layer0_out[662] <= x[38] & x[42];
     layer0_out[663] <= x[234] & ~x[231];
     layer0_out[664] <= ~x[240] | x[242];
     layer0_out[665] <= ~x[344] | x[347];
     layer0_out[666] <= ~(x[283] ^ x[286]);
     layer0_out[667] <= x[111] & ~x[114];
     layer0_out[668] <= 1'b1;
     layer0_out[669] <= ~x[124];
     layer0_out[670] <= x[34];
     layer0_out[671] <= ~(x[141] | x[143]);
     layer0_out[672] <= ~(x[104] | x[107]);
     layer0_out[673] <= x[112] ^ x[115];
     layer0_out[674] <= 1'b1;
     layer0_out[675] <= ~(x[383] & x[385]);
     layer0_out[676] <= x[80] ^ x[84];
     layer0_out[677] <= ~x[291];
     layer0_out[678] <= 1'b0;
     layer0_out[679] <= x[273] & ~x[269];
     layer0_out[680] <= x[240];
     layer0_out[681] <= ~x[379];
     layer0_out[682] <= x[202] | x[203];
     layer0_out[683] <= x[231] | x[233];
     layer0_out[684] <= 1'b0;
     layer0_out[685] <= 1'b1;
     layer0_out[686] <= ~x[260];
     layer0_out[687] <= x[288] & x[292];
     layer0_out[688] <= ~(x[225] | x[227]);
     layer0_out[689] <= ~(x[263] | x[265]);
     layer0_out[690] <= x[197] & ~x[196];
     layer0_out[691] <= ~x[265];
     layer0_out[692] <= x[384];
     layer0_out[693] <= ~x[308];
     layer0_out[694] <= ~(x[116] ^ x[120]);
     layer0_out[695] <= x[160] & ~x[164];
     layer0_out[696] <= x[61] & ~x[65];
     layer0_out[697] <= x[103] ^ x[104];
     layer0_out[698] <= x[143] | x[144];
     layer0_out[699] <= x[190] | x[192];
     layer0_out[700] <= x[186] | x[189];
     layer0_out[701] <= ~x[43];
     layer0_out[702] <= x[2] | x[3];
     layer0_out[703] <= ~x[391] | x[389];
     layer0_out[704] <= ~(x[120] | x[121]);
     layer0_out[705] <= 1'b0;
     layer0_out[706] <= x[220] & ~x[224];
     layer0_out[707] <= 1'b1;
     layer0_out[708] <= 1'b0;
     layer0_out[709] <= x[368] | x[371];
     layer0_out[710] <= x[227];
     layer0_out[711] <= x[204] ^ x[206];
     layer0_out[712] <= 1'b0;
     layer0_out[713] <= x[116] | x[118];
     layer0_out[714] <= x[378] | x[380];
     layer0_out[715] <= x[55] & x[58];
     layer0_out[716] <= ~(x[224] | x[226]);
     layer0_out[717] <= x[136] & ~x[134];
     layer0_out[718] <= x[73] | x[75];
     layer0_out[719] <= x[137] & ~x[134];
     layer0_out[720] <= x[271];
     layer0_out[721] <= x[282];
     layer0_out[722] <= 1'b0;
     layer0_out[723] <= x[15] & x[18];
     layer0_out[724] <= ~x[44] | x[45];
     layer0_out[725] <= x[386] & ~x[388];
     layer0_out[726] <= ~(x[294] | x[296]);
     layer0_out[727] <= ~(x[72] ^ x[74]);
     layer0_out[728] <= 1'b1;
     layer0_out[729] <= 1'b0;
     layer0_out[730] <= 1'b0;
     layer0_out[731] <= x[347] | x[348];
     layer0_out[732] <= 1'b0;
     layer0_out[733] <= 1'b1;
     layer0_out[734] <= x[57] & ~x[53];
     layer0_out[735] <= 1'b0;
     layer0_out[736] <= 1'b0;
     layer0_out[737] <= ~x[57] | x[56];
     layer0_out[738] <= ~(x[162] | x[163]);
     layer0_out[739] <= x[168] & ~x[170];
     layer0_out[740] <= 1'b0;
     layer0_out[741] <= x[172] | x[173];
     layer0_out[742] <= ~(x[56] | x[59]);
     layer0_out[743] <= ~(x[32] | x[34]);
     layer0_out[744] <= x[44];
     layer0_out[745] <= ~(x[223] | x[226]);
     layer0_out[746] <= ~x[282];
     layer0_out[747] <= ~(x[195] ^ x[198]);
     layer0_out[748] <= 1'b1;
     layer0_out[749] <= ~x[3];
     layer0_out[750] <= ~(x[109] & x[112]);
     layer0_out[751] <= ~(x[269] | x[270]);
     layer0_out[752] <= x[82] | x[84];
     layer0_out[753] <= 1'b0;
     layer0_out[754] <= ~x[331];
     layer0_out[755] <= ~x[378];
     layer0_out[756] <= ~(x[31] | x[32]);
     layer0_out[757] <= x[15] ^ x[19];
     layer0_out[758] <= x[77] | x[79];
     layer0_out[759] <= x[366] | x[369];
     layer0_out[760] <= ~x[140];
     layer0_out[761] <= x[79] & ~x[78];
     layer0_out[762] <= ~x[10] | x[11];
     layer0_out[763] <= 1'b0;
     layer0_out[764] <= 1'b1;
     layer0_out[765] <= ~x[123] | x[126];
     layer0_out[766] <= ~(x[324] | x[327]);
     layer0_out[767] <= x[119] | x[122];
     layer0_out[768] <= ~x[166] | x[164];
     layer0_out[769] <= x[261] & x[264];
     layer0_out[770] <= x[22] | x[25];
     layer0_out[771] <= 1'b0;
     layer0_out[772] <= ~(x[247] & x[250]);
     layer0_out[773] <= ~(x[127] & x[130]);
     layer0_out[774] <= 1'b1;
     layer0_out[775] <= x[6];
     layer0_out[776] <= ~(x[379] | x[380]);
     layer0_out[777] <= 1'b1;
     layer0_out[778] <= ~x[236];
     layer0_out[779] <= ~x[1] | x[0];
     layer0_out[780] <= 1'b1;
     layer0_out[781] <= x[352] | x[355];
     layer0_out[782] <= 1'b1;
     layer0_out[783] <= x[32] & x[35];
     layer0_out[784] <= 1'b1;
     layer0_out[785] <= ~(x[70] & x[73]);
     layer0_out[786] <= x[87];
     layer0_out[787] <= x[305] & x[308];
     layer0_out[788] <= 1'b1;
     layer0_out[789] <= x[385] | x[388];
     layer0_out[790] <= ~(x[356] | x[358]);
     layer0_out[791] <= 1'b1;
     layer0_out[792] <= x[342] | x[345];
     layer0_out[793] <= x[107] | x[108];
     layer0_out[794] <= x[318] | x[320];
     layer0_out[795] <= x[114] | x[115];
     layer0_out[796] <= ~(x[285] | x[286]);
     layer0_out[797] <= ~x[229] | x[226];
     layer0_out[798] <= 1'b1;
     layer0_out[799] <= ~x[174];
     layer0_out[800] <= ~(x[245] | x[246]);
     layer0_out[801] <= ~(x[229] & x[232]);
     layer0_out[802] <= x[301] | x[303];
     layer0_out[803] <= ~x[357];
     layer0_out[804] <= x[385] & ~x[387];
     layer0_out[805] <= 1'b1;
     layer0_out[806] <= x[330] & ~x[327];
     layer0_out[807] <= ~(x[161] | x[163]);
     layer0_out[808] <= x[180] | x[184];
     layer0_out[809] <= ~x[28];
     layer0_out[810] <= x[64] | x[66];
     layer0_out[811] <= ~(x[130] | x[131]);
     layer0_out[812] <= x[58] | x[62];
     layer0_out[813] <= ~(x[104] ^ x[108]);
     layer0_out[814] <= 1'b0;
     layer0_out[815] <= x[36] | x[37];
     layer0_out[816] <= 1'b1;
     layer0_out[817] <= ~(x[121] | x[123]);
     layer0_out[818] <= 1'b0;
     layer0_out[819] <= x[192];
     layer0_out[820] <= ~x[319];
     layer0_out[821] <= 1'b1;
     layer0_out[822] <= 1'b0;
     layer0_out[823] <= x[310];
     layer0_out[824] <= ~(x[54] & x[57]);
     layer0_out[825] <= 1'b0;
     layer0_out[826] <= 1'b0;
     layer0_out[827] <= x[374] ^ x[377];
     layer0_out[828] <= x[205] | x[207];
     layer0_out[829] <= 1'b1;
     layer0_out[830] <= ~(x[107] & x[111]);
     layer0_out[831] <= 1'b1;
     layer0_out[832] <= 1'b1;
     layer0_out[833] <= x[180];
     layer0_out[834] <= x[162];
     layer0_out[835] <= x[256] & x[260];
     layer0_out[836] <= 1'b1;
     layer0_out[837] <= x[129];
     layer0_out[838] <= ~(x[207] | x[209]);
     layer0_out[839] <= x[300] | x[303];
     layer0_out[840] <= x[395];
     layer0_out[841] <= ~(x[265] & x[267]);
     layer0_out[842] <= x[141] | x[144];
     layer0_out[843] <= 1'b0;
     layer0_out[844] <= 1'b1;
     layer0_out[845] <= x[202];
     layer0_out[846] <= ~(x[360] | x[361]);
     layer0_out[847] <= 1'b0;
     layer0_out[848] <= x[254];
     layer0_out[849] <= ~x[213];
     layer0_out[850] <= x[201] | x[202];
     layer0_out[851] <= x[90] & x[91];
     layer0_out[852] <= ~(x[136] & x[140]);
     layer0_out[853] <= x[29];
     layer0_out[854] <= x[9];
     layer0_out[855] <= ~(x[211] | x[212]);
     layer0_out[856] <= ~x[309];
     layer0_out[857] <= 1'b1;
     layer0_out[858] <= x[139] & ~x[143];
     layer0_out[859] <= x[236] | x[237];
     layer0_out[860] <= x[146] | x[148];
     layer0_out[861] <= ~x[61];
     layer0_out[862] <= ~x[291] | x[295];
     layer0_out[863] <= x[6] & ~x[8];
     layer0_out[864] <= x[188];
     layer0_out[865] <= 1'b1;
     layer0_out[866] <= ~(x[260] | x[262]);
     layer0_out[867] <= 1'b1;
     layer0_out[868] <= x[179] | x[182];
     layer0_out[869] <= 1'b0;
     layer0_out[870] <= x[363] & ~x[361];
     layer0_out[871] <= ~x[87] | x[86];
     layer0_out[872] <= 1'b0;
     layer0_out[873] <= x[7] & x[10];
     layer0_out[874] <= ~x[101] | x[97];
     layer0_out[875] <= 1'b1;
     layer0_out[876] <= ~(x[353] | x[354]);
     layer0_out[877] <= x[35] | x[37];
     layer0_out[878] <= 1'b1;
     layer0_out[879] <= 1'b1;
     layer0_out[880] <= 1'b0;
     layer0_out[881] <= x[313] & ~x[315];
     layer0_out[882] <= 1'b1;
     layer0_out[883] <= x[131] | x[133];
     layer0_out[884] <= ~(x[284] | x[288]);
     layer0_out[885] <= 1'b1;
     layer0_out[886] <= ~(x[332] | x[333]);
     layer0_out[887] <= x[171];
     layer0_out[888] <= x[281] & x[284];
     layer0_out[889] <= ~x[225] | x[229];
     layer0_out[890] <= x[232] | x[234];
     layer0_out[891] <= 1'b0;
     layer0_out[892] <= 1'b0;
     layer0_out[893] <= ~x[171];
     layer0_out[894] <= 1'b0;
     layer0_out[895] <= x[57];
     layer0_out[896] <= x[167] & ~x[168];
     layer0_out[897] <= ~x[56];
     layer0_out[898] <= 1'b0;
     layer0_out[899] <= 1'b0;
     layer0_out[900] <= ~x[297] | x[295];
     layer0_out[901] <= ~x[11];
     layer0_out[902] <= ~x[172];
     layer0_out[903] <= ~(x[323] | x[325]);
     layer0_out[904] <= x[268] | x[270];
     layer0_out[905] <= ~(x[274] | x[278]);
     layer0_out[906] <= ~(x[166] | x[168]);
     layer0_out[907] <= x[226] & ~x[230];
     layer0_out[908] <= x[108];
     layer0_out[909] <= ~x[371];
     layer0_out[910] <= x[81] & ~x[84];
     layer0_out[911] <= 1'b1;
     layer0_out[912] <= ~(x[244] | x[246]);
     layer0_out[913] <= x[163] & ~x[165];
     layer0_out[914] <= ~(x[170] | x[174]);
     layer0_out[915] <= 1'b0;
     layer0_out[916] <= x[332] & x[335];
     layer0_out[917] <= x[276] | x[277];
     layer0_out[918] <= x[361] | x[364];
     layer0_out[919] <= ~(x[344] | x[346]);
     layer0_out[920] <= x[279] & ~x[276];
     layer0_out[921] <= x[175] & x[177];
     layer0_out[922] <= ~(x[213] & x[215]);
     layer0_out[923] <= x[280] | x[283];
     layer0_out[924] <= x[257] & ~x[258];
     layer0_out[925] <= x[109] | x[110];
     layer0_out[926] <= x[30];
     layer0_out[927] <= x[301] & x[304];
     layer0_out[928] <= x[100] & ~x[97];
     layer0_out[929] <= ~(x[193] | x[195]);
     layer0_out[930] <= 1'b1;
     layer0_out[931] <= x[40] & ~x[44];
     layer0_out[932] <= x[279] & ~x[278];
     layer0_out[933] <= ~(x[154] & x[158]);
     layer0_out[934] <= ~x[356] | x[354];
     layer0_out[935] <= x[74] ^ x[75];
     layer0_out[936] <= x[135] | x[137];
     layer0_out[937] <= x[152] & x[154];
     layer0_out[938] <= ~(x[237] | x[238]);
     layer0_out[939] <= 1'b1;
     layer0_out[940] <= x[313] & ~x[311];
     layer0_out[941] <= 1'b1;
     layer0_out[942] <= ~(x[134] | x[135]);
     layer0_out[943] <= ~(x[341] | x[344]);
     layer0_out[944] <= 1'b0;
     layer0_out[945] <= 1'b1;
     layer0_out[946] <= 1'b1;
     layer0_out[947] <= 1'b0;
     layer0_out[948] <= ~x[73] | x[71];
     layer0_out[949] <= ~(x[285] | x[287]);
     layer0_out[950] <= ~(x[66] & x[69]);
     layer0_out[951] <= x[24] | x[25];
     layer0_out[952] <= ~(x[147] | x[149]);
     layer0_out[953] <= 1'b1;
     layer0_out[954] <= ~(x[230] | x[232]);
     layer0_out[955] <= 1'b1;
     layer0_out[956] <= ~x[21] | x[22];
     layer0_out[957] <= x[143] & x[145];
     layer0_out[958] <= x[302] | x[304];
     layer0_out[959] <= 1'b1;
     layer0_out[960] <= x[227] | x[231];
     layer0_out[961] <= ~x[267];
     layer0_out[962] <= x[278];
     layer0_out[963] <= 1'b1;
     layer0_out[964] <= 1'b0;
     layer0_out[965] <= ~x[87] | x[89];
     layer0_out[966] <= x[76] & x[77];
     layer0_out[967] <= ~x[96];
     layer0_out[968] <= x[119] | x[121];
     layer0_out[969] <= x[294] | x[295];
     layer0_out[970] <= ~(x[31] | x[35]);
     layer0_out[971] <= 1'b0;
     layer0_out[972] <= ~x[226];
     layer0_out[973] <= x[192] & x[194];
     layer0_out[974] <= ~x[279] | x[282];
     layer0_out[975] <= x[68] & x[72];
     layer0_out[976] <= x[110];
     layer0_out[977] <= ~(x[368] ^ x[369]);
     layer0_out[978] <= 1'b0;
     layer0_out[979] <= ~x[150];
     layer0_out[980] <= ~(x[224] | x[225]);
     layer0_out[981] <= ~x[339];
     layer0_out[982] <= ~x[177] | x[173];
     layer0_out[983] <= x[54] & x[56];
     layer0_out[984] <= 1'b1;
     layer0_out[985] <= x[113];
     layer0_out[986] <= ~x[149] | x[152];
     layer0_out[987] <= 1'b1;
     layer0_out[988] <= x[115] | x[116];
     layer0_out[989] <= x[238] & ~x[241];
     layer0_out[990] <= x[264];
     layer0_out[991] <= ~x[242];
     layer0_out[992] <= ~(x[383] & x[384]);
     layer0_out[993] <= x[162];
     layer0_out[994] <= ~x[151] | x[148];
     layer0_out[995] <= ~(x[21] & x[23]);
     layer0_out[996] <= ~x[362];
     layer0_out[997] <= 1'b0;
     layer0_out[998] <= ~(x[91] & x[93]);
     layer0_out[999] <= 1'b1;
     layer0_out[1000] <= ~x[118] | x[122];
     layer0_out[1001] <= ~(x[313] | x[314]);
     layer0_out[1002] <= x[296] | x[300];
     layer0_out[1003] <= ~(x[57] | x[61]);
     layer0_out[1004] <= x[374];
     layer0_out[1005] <= ~(x[284] | x[287]);
     layer0_out[1006] <= x[215] & ~x[217];
     layer0_out[1007] <= x[255] | x[258];
     layer0_out[1008] <= x[160];
     layer0_out[1009] <= x[192];
     layer0_out[1010] <= ~x[367];
     layer0_out[1011] <= x[127] | x[131];
     layer0_out[1012] <= 1'b1;
     layer0_out[1013] <= x[11];
     layer0_out[1014] <= 1'b1;
     layer0_out[1015] <= x[172] ^ x[175];
     layer0_out[1016] <= x[95] | x[98];
     layer0_out[1017] <= x[98];
     layer0_out[1018] <= x[198] & x[199];
     layer0_out[1019] <= 1'b0;
     layer0_out[1020] <= ~x[185];
     layer0_out[1021] <= x[214] & x[215];
     layer0_out[1022] <= x[104];
     layer0_out[1023] <= 1'b1;
     layer0_out[1024] <= ~(x[20] | x[21]);
     layer0_out[1025] <= x[296] | x[298];
     layer0_out[1026] <= 1'b0;
     layer0_out[1027] <= ~x[300] | x[298];
     layer0_out[1028] <= x[218];
     layer0_out[1029] <= 1'b0;
     layer0_out[1030] <= x[259];
     layer0_out[1031] <= ~x[13] | x[16];
     layer0_out[1032] <= x[184] | x[188];
     layer0_out[1033] <= ~x[161];
     layer0_out[1034] <= 1'b1;
     layer0_out[1035] <= x[377] | x[379];
     layer0_out[1036] <= 1'b0;
     layer0_out[1037] <= 1'b1;
     layer0_out[1038] <= x[364];
     layer0_out[1039] <= ~(x[217] | x[218]);
     layer0_out[1040] <= ~(x[85] & x[88]);
     layer0_out[1041] <= 1'b1;
     layer0_out[1042] <= x[92] & ~x[89];
     layer0_out[1043] <= ~(x[18] | x[20]);
     layer0_out[1044] <= x[167];
     layer0_out[1045] <= x[222] & ~x[223];
     layer0_out[1046] <= x[157] | x[158];
     layer0_out[1047] <= ~x[259];
     layer0_out[1048] <= x[15] ^ x[16];
     layer0_out[1049] <= ~(x[238] ^ x[239]);
     layer0_out[1050] <= x[43] & ~x[46];
     layer0_out[1051] <= x[367] | x[370];
     layer0_out[1052] <= 1'b0;
     layer0_out[1053] <= 1'b1;
     layer0_out[1054] <= x[46] & ~x[47];
     layer0_out[1055] <= 1'b0;
     layer0_out[1056] <= ~(x[49] & x[52]);
     layer0_out[1057] <= 1'b1;
     layer0_out[1058] <= ~x[208] | x[204];
     layer0_out[1059] <= ~x[30] | x[34];
     layer0_out[1060] <= x[85];
     layer0_out[1061] <= x[279] | x[283];
     layer0_out[1062] <= ~(x[98] | x[101]);
     layer0_out[1063] <= 1'b0;
     layer0_out[1064] <= ~x[239];
     layer0_out[1065] <= ~(x[135] | x[139]);
     layer0_out[1066] <= x[277] & ~x[275];
     layer0_out[1067] <= x[117] & ~x[119];
     layer0_out[1068] <= x[137] | x[140];
     layer0_out[1069] <= ~(x[267] & x[270]);
     layer0_out[1070] <= ~x[12];
     layer0_out[1071] <= ~(x[232] | x[235]);
     layer0_out[1072] <= x[142] | x[143];
     layer0_out[1073] <= ~x[268] | x[272];
     layer0_out[1074] <= ~(x[136] ^ x[139]);
     layer0_out[1075] <= x[62];
     layer0_out[1076] <= ~(x[268] ^ x[271]);
     layer0_out[1077] <= 1'b0;
     layer0_out[1078] <= 1'b1;
     layer0_out[1079] <= ~(x[241] | x[244]);
     layer0_out[1080] <= x[64] | x[65];
     layer0_out[1081] <= ~x[257] | x[260];
     layer0_out[1082] <= ~x[78] | x[74];
     layer0_out[1083] <= 1'b1;
     layer0_out[1084] <= x[60];
     layer0_out[1085] <= 1'b0;
     layer0_out[1086] <= 1'b0;
     layer0_out[1087] <= 1'b0;
     layer0_out[1088] <= x[326];
     layer0_out[1089] <= x[31] & x[34];
     layer0_out[1090] <= x[81] | x[85];
     layer0_out[1091] <= x[99];
     layer0_out[1092] <= ~(x[2] | x[5]);
     layer0_out[1093] <= ~(x[97] & x[99]);
     layer0_out[1094] <= x[96] & x[100];
     layer0_out[1095] <= x[98] | x[100];
     layer0_out[1096] <= ~(x[185] & x[189]);
     layer0_out[1097] <= 1'b0;
     layer0_out[1098] <= ~x[4] | x[7];
     layer0_out[1099] <= ~(x[360] | x[363]);
     layer0_out[1100] <= 1'b1;
     layer0_out[1101] <= ~x[293] | x[296];
     layer0_out[1102] <= x[55] | x[56];
     layer0_out[1103] <= x[49];
     layer0_out[1104] <= x[147] | x[148];
     layer0_out[1105] <= 1'b0;
     layer0_out[1106] <= ~(x[264] | x[265]);
     layer0_out[1107] <= x[171] | x[175];
     layer0_out[1108] <= ~(x[241] | x[243]);
     layer0_out[1109] <= x[286] | x[288];
     layer0_out[1110] <= x[185] & x[187];
     layer0_out[1111] <= 1'b0;
     layer0_out[1112] <= x[19];
     layer0_out[1113] <= ~(x[206] | x[210]);
     layer0_out[1114] <= x[130] ^ x[134];
     layer0_out[1115] <= 1'b1;
     layer0_out[1116] <= ~(x[253] & x[257]);
     layer0_out[1117] <= ~x[140];
     layer0_out[1118] <= x[88] & ~x[86];
     layer0_out[1119] <= ~x[149];
     layer0_out[1120] <= 1'b0;
     layer0_out[1121] <= 1'b0;
     layer0_out[1122] <= ~(x[75] & x[79]);
     layer0_out[1123] <= ~(x[24] | x[27]);
     layer0_out[1124] <= ~(x[305] | x[306]);
     layer0_out[1125] <= 1'b1;
     layer0_out[1126] <= 1'b1;
     layer0_out[1127] <= x[207];
     layer0_out[1128] <= x[117];
     layer0_out[1129] <= ~(x[106] & x[107]);
     layer0_out[1130] <= x[374] | x[375];
     layer0_out[1131] <= ~(x[108] | x[109]);
     layer0_out[1132] <= ~x[119];
     layer0_out[1133] <= x[284] & ~x[286];
     layer0_out[1134] <= 1'b0;
     layer0_out[1135] <= 1'b0;
     layer0_out[1136] <= x[309] & x[310];
     layer0_out[1137] <= x[348] & x[351];
     layer0_out[1138] <= x[287] | x[290];
     layer0_out[1139] <= ~x[117];
     layer0_out[1140] <= ~(x[349] | x[352]);
     layer0_out[1141] <= ~x[258];
     layer0_out[1142] <= x[176] | x[178];
     layer0_out[1143] <= x[306];
     layer0_out[1144] <= 1'b1;
     layer0_out[1145] <= x[62];
     layer0_out[1146] <= x[6] & ~x[5];
     layer0_out[1147] <= ~(x[245] | x[248]);
     layer0_out[1148] <= ~(x[388] | x[390]);
     layer0_out[1149] <= 1'b0;
     layer0_out[1150] <= ~(x[295] | x[299]);
     layer0_out[1151] <= ~x[68] | x[71];
     layer0_out[1152] <= ~(x[291] | x[292]);
     layer0_out[1153] <= ~x[358];
     layer0_out[1154] <= 1'b1;
     layer0_out[1155] <= ~(x[281] | x[283]);
     layer0_out[1156] <= 1'b1;
     layer0_out[1157] <= ~(x[149] | x[150]);
     layer0_out[1158] <= x[233] & ~x[234];
     layer0_out[1159] <= x[131] | x[134];
     layer0_out[1160] <= ~(x[346] | x[348]);
     layer0_out[1161] <= x[183] | x[184];
     layer0_out[1162] <= ~x[358];
     layer0_out[1163] <= ~(x[282] | x[283]);
     layer0_out[1164] <= ~(x[40] | x[43]);
     layer0_out[1165] <= x[143] ^ x[146];
     layer0_out[1166] <= 1'b0;
     layer0_out[1167] <= 1'b0;
     layer0_out[1168] <= 1'b0;
     layer0_out[1169] <= 1'b1;
     layer0_out[1170] <= 1'b1;
     layer0_out[1171] <= x[212];
     layer0_out[1172] <= x[249] & ~x[251];
     layer0_out[1173] <= 1'b0;
     layer0_out[1174] <= x[90];
     layer0_out[1175] <= ~(x[140] | x[142]);
     layer0_out[1176] <= x[1] | x[2];
     layer0_out[1177] <= 1'b1;
     layer0_out[1178] <= ~x[190] | x[187];
     layer0_out[1179] <= x[0] ^ x[3];
     layer0_out[1180] <= x[359];
     layer0_out[1181] <= ~x[155] | x[154];
     layer0_out[1182] <= ~(x[138] & x[140]);
     layer0_out[1183] <= ~x[298] | x[295];
     layer0_out[1184] <= 1'b0;
     layer0_out[1185] <= 1'b1;
     layer0_out[1186] <= 1'b0;
     layer0_out[1187] <= ~(x[244] & x[247]);
     layer0_out[1188] <= ~x[176] | x[180];
     layer0_out[1189] <= ~x[194];
     layer0_out[1190] <= ~x[303];
     layer0_out[1191] <= x[319] | x[320];
     layer0_out[1192] <= ~(x[177] | x[181]);
     layer0_out[1193] <= ~(x[210] & x[213]);
     layer0_out[1194] <= ~x[13];
     layer0_out[1195] <= x[132] ^ x[136];
     layer0_out[1196] <= 1'b1;
     layer0_out[1197] <= ~x[166] | x[167];
     layer0_out[1198] <= ~(x[166] & x[169]);
     layer0_out[1199] <= ~(x[373] & x[376]);
     layer0_out[1200] <= ~(x[84] | x[86]);
     layer0_out[1201] <= x[394] | x[396];
     layer0_out[1202] <= ~x[102] | x[106];
     layer0_out[1203] <= 1'b1;
     layer0_out[1204] <= ~x[211];
     layer0_out[1205] <= ~(x[338] | x[340]);
     layer0_out[1206] <= x[0] | x[2];
     layer0_out[1207] <= ~x[226];
     layer0_out[1208] <= 1'b0;
     layer0_out[1209] <= ~(x[166] | x[170]);
     layer0_out[1210] <= ~(x[363] | x[364]);
     layer0_out[1211] <= 1'b1;
     layer0_out[1212] <= 1'b1;
     layer0_out[1213] <= x[65] & ~x[66];
     layer0_out[1214] <= ~x[79];
     layer0_out[1215] <= 1'b0;
     layer0_out[1216] <= x[52];
     layer0_out[1217] <= 1'b0;
     layer0_out[1218] <= 1'b0;
     layer0_out[1219] <= x[243];
     layer0_out[1220] <= ~x[213];
     layer0_out[1221] <= x[186] & ~x[183];
     layer0_out[1222] <= x[256] | x[258];
     layer0_out[1223] <= ~x[248] | x[246];
     layer0_out[1224] <= ~x[230];
     layer0_out[1225] <= 1'b0;
     layer0_out[1226] <= x[38];
     layer0_out[1227] <= x[261] & ~x[258];
     layer0_out[1228] <= ~x[156];
     layer0_out[1229] <= x[179] & ~x[175];
     layer0_out[1230] <= x[35] & ~x[34];
     layer0_out[1231] <= 1'b0;
     layer0_out[1232] <= x[137] | x[138];
     layer0_out[1233] <= ~(x[181] & x[185]);
     layer0_out[1234] <= ~(x[188] | x[190]);
     layer0_out[1235] <= x[317] | x[318];
     layer0_out[1236] <= ~(x[384] | x[385]);
     layer0_out[1237] <= 1'b0;
     layer0_out[1238] <= 1'b1;
     layer0_out[1239] <= ~(x[312] | x[315]);
     layer0_out[1240] <= x[188] | x[192];
     layer0_out[1241] <= x[198];
     layer0_out[1242] <= x[16] | x[18];
     layer0_out[1243] <= ~(x[266] | x[268]);
     layer0_out[1244] <= ~(x[190] | x[191]);
     layer0_out[1245] <= ~(x[127] | x[128]);
     layer0_out[1246] <= ~(x[152] | x[155]);
     layer0_out[1247] <= x[140] | x[141];
     layer0_out[1248] <= 1'b0;
     layer0_out[1249] <= ~x[172];
     layer0_out[1250] <= x[319] & x[321];
     layer0_out[1251] <= 1'b1;
     layer0_out[1252] <= 1'b1;
     layer0_out[1253] <= 1'b0;
     layer0_out[1254] <= x[70] | x[72];
     layer0_out[1255] <= ~x[189];
     layer0_out[1256] <= ~(x[264] | x[268]);
     layer0_out[1257] <= x[41] | x[44];
     layer0_out[1258] <= x[55] | x[57];
     layer0_out[1259] <= ~x[206];
     layer0_out[1260] <= ~(x[296] | x[299]);
     layer0_out[1261] <= ~x[225] | x[226];
     layer0_out[1262] <= x[336] & x[339];
     layer0_out[1263] <= ~x[130] | x[126];
     layer0_out[1264] <= 1'b0;
     layer0_out[1265] <= x[161] | x[165];
     layer0_out[1266] <= 1'b0;
     layer0_out[1267] <= x[305] & ~x[302];
     layer0_out[1268] <= x[298] ^ x[302];
     layer0_out[1269] <= ~x[119];
     layer0_out[1270] <= ~x[314];
     layer0_out[1271] <= ~(x[359] | x[362]);
     layer0_out[1272] <= ~(x[55] | x[59]);
     layer0_out[1273] <= x[269] & x[272];
     layer0_out[1274] <= x[201] | x[205];
     layer0_out[1275] <= ~(x[220] | x[223]);
     layer0_out[1276] <= x[164] & x[165];
     layer0_out[1277] <= x[281] | x[285];
     layer0_out[1278] <= x[289] | x[291];
     layer0_out[1279] <= 1'b1;
     layer0_out[1280] <= x[358] | x[359];
     layer0_out[1281] <= ~x[168];
     layer0_out[1282] <= 1'b0;
     layer0_out[1283] <= 1'b0;
     layer0_out[1284] <= ~(x[280] & x[284]);
     layer0_out[1285] <= ~(x[330] | x[331]);
     layer0_out[1286] <= ~(x[250] | x[253]);
     layer0_out[1287] <= ~(x[258] | x[259]);
     layer0_out[1288] <= ~(x[101] & x[105]);
     layer0_out[1289] <= ~(x[183] ^ x[185]);
     layer0_out[1290] <= ~x[45];
     layer0_out[1291] <= x[42] & ~x[44];
     layer0_out[1292] <= 1'b0;
     layer0_out[1293] <= 1'b0;
     layer0_out[1294] <= x[170] & ~x[171];
     layer0_out[1295] <= 1'b1;
     layer0_out[1296] <= ~(x[70] & x[71]);
     layer0_out[1297] <= ~x[346];
     layer0_out[1298] <= ~(x[304] | x[305]);
     layer0_out[1299] <= 1'b1;
     layer0_out[1300] <= x[122] ^ x[126];
     layer0_out[1301] <= ~x[150] | x[146];
     layer0_out[1302] <= 1'b1;
     layer0_out[1303] <= x[317] | x[320];
     layer0_out[1304] <= ~(x[130] | x[133]);
     layer0_out[1305] <= x[104];
     layer0_out[1306] <= x[106] | x[109];
     layer0_out[1307] <= x[150];
     layer0_out[1308] <= x[189];
     layer0_out[1309] <= 1'b0;
     layer0_out[1310] <= ~(x[352] ^ x[353]);
     layer0_out[1311] <= ~x[146];
     layer0_out[1312] <= x[131];
     layer0_out[1313] <= ~(x[209] | x[211]);
     layer0_out[1314] <= x[106] | x[110];
     layer0_out[1315] <= 1'b1;
     layer0_out[1316] <= ~x[266];
     layer0_out[1317] <= ~(x[137] | x[139]);
     layer0_out[1318] <= x[202] & ~x[206];
     layer0_out[1319] <= x[85];
     layer0_out[1320] <= ~(x[191] ^ x[194]);
     layer0_out[1321] <= x[206] & ~x[208];
     layer0_out[1322] <= ~(x[339] | x[342]);
     layer0_out[1323] <= x[29] | x[30];
     layer0_out[1324] <= 1'b1;
     layer0_out[1325] <= x[82] & ~x[83];
     layer0_out[1326] <= ~(x[148] | x[149]);
     layer0_out[1327] <= ~(x[40] | x[41]);
     layer0_out[1328] <= ~(x[17] | x[18]);
     layer0_out[1329] <= ~(x[96] | x[98]);
     layer0_out[1330] <= ~x[210];
     layer0_out[1331] <= ~(x[252] | x[253]);
     layer0_out[1332] <= 1'b1;
     layer0_out[1333] <= 1'b1;
     layer0_out[1334] <= ~(x[74] | x[77]);
     layer0_out[1335] <= 1'b1;
     layer0_out[1336] <= 1'b0;
     layer0_out[1337] <= x[93] & x[97];
     layer0_out[1338] <= 1'b0;
     layer0_out[1339] <= 1'b1;
     layer0_out[1340] <= 1'b0;
     layer0_out[1341] <= ~x[249] | x[253];
     layer0_out[1342] <= x[386] | x[387];
     layer0_out[1343] <= ~(x[387] | x[388]);
     layer0_out[1344] <= ~(x[144] | x[145]);
     layer0_out[1345] <= x[51] & x[54];
     layer0_out[1346] <= ~(x[390] | x[393]);
     layer0_out[1347] <= 1'b0;
     layer0_out[1348] <= x[62] & x[64];
     layer0_out[1349] <= x[317] | x[319];
     layer0_out[1350] <= x[286] & x[287];
     layer0_out[1351] <= 1'b0;
     layer0_out[1352] <= x[158] & x[161];
     layer0_out[1353] <= 1'b0;
     layer0_out[1354] <= x[387];
     layer0_out[1355] <= 1'b1;
     layer0_out[1356] <= 1'b1;
     layer0_out[1357] <= ~x[255] | x[254];
     layer0_out[1358] <= ~(x[132] & x[135]);
     layer0_out[1359] <= 1'b1;
     layer0_out[1360] <= ~(x[382] & x[385]);
     layer0_out[1361] <= ~x[72] | x[73];
     layer0_out[1362] <= x[48] & x[51];
     layer0_out[1363] <= 1'b1;
     layer0_out[1364] <= 1'b0;
     layer0_out[1365] <= x[280] & ~x[276];
     layer0_out[1366] <= ~x[22] | x[23];
     layer0_out[1367] <= ~(x[315] | x[318]);
     layer0_out[1368] <= ~(x[157] | x[159]);
     layer0_out[1369] <= x[397] | x[398];
     layer0_out[1370] <= ~(x[242] | x[243]);
     layer0_out[1371] <= ~x[141] | x[139];
     layer0_out[1372] <= 1'b0;
     layer0_out[1373] <= 1'b0;
     layer0_out[1374] <= ~x[370] | x[373];
     layer0_out[1375] <= x[156];
     layer0_out[1376] <= 1'b1;
     layer0_out[1377] <= ~(x[355] | x[356]);
     layer0_out[1378] <= 1'b0;
     layer0_out[1379] <= 1'b0;
     layer0_out[1380] <= ~(x[396] & x[399]);
     layer0_out[1381] <= 1'b1;
     layer0_out[1382] <= ~(x[65] ^ x[68]);
     layer0_out[1383] <= x[339] & ~x[341];
     layer0_out[1384] <= ~x[168];
     layer0_out[1385] <= x[368];
     layer0_out[1386] <= ~(x[200] | x[202]);
     layer0_out[1387] <= ~(x[60] | x[63]);
     layer0_out[1388] <= ~x[147];
     layer0_out[1389] <= x[312] | x[313];
     layer0_out[1390] <= x[200] | x[203];
     layer0_out[1391] <= 1'b1;
     layer0_out[1392] <= x[48] & x[52];
     layer0_out[1393] <= 1'b1;
     layer0_out[1394] <= x[304] & ~x[307];
     layer0_out[1395] <= ~(x[59] | x[63]);
     layer0_out[1396] <= 1'b0;
     layer0_out[1397] <= x[128] & x[130];
     layer0_out[1398] <= x[363] | x[366];
     layer0_out[1399] <= ~(x[293] | x[297]);
     layer0_out[1400] <= ~(x[89] & x[90]);
     layer0_out[1401] <= x[369] & x[371];
     layer0_out[1402] <= ~x[49] | x[48];
     layer0_out[1403] <= ~(x[265] | x[266]);
     layer0_out[1404] <= 1'b0;
     layer0_out[1405] <= x[60];
     layer0_out[1406] <= x[252] | x[256];
     layer0_out[1407] <= 1'b1;
     layer0_out[1408] <= ~(x[197] ^ x[201]);
     layer0_out[1409] <= x[40] | x[42];
     layer0_out[1410] <= ~x[219] | x[221];
     layer0_out[1411] <= 1'b1;
     layer0_out[1412] <= x[357] & x[359];
     layer0_out[1413] <= x[181];
     layer0_out[1414] <= 1'b1;
     layer0_out[1415] <= ~(x[394] | x[395]);
     layer0_out[1416] <= x[221];
     layer0_out[1417] <= x[234] | x[236];
     layer0_out[1418] <= x[295];
     layer0_out[1419] <= ~(x[321] | x[322]);
     layer0_out[1420] <= ~(x[339] | x[340]);
     layer0_out[1421] <= x[197];
     layer0_out[1422] <= ~(x[70] | x[74]);
     layer0_out[1423] <= ~(x[101] | x[102]);
     layer0_out[1424] <= ~x[319];
     layer0_out[1425] <= x[19] & ~x[18];
     layer0_out[1426] <= x[47];
     layer0_out[1427] <= ~x[338];
     layer0_out[1428] <= 1'b0;
     layer0_out[1429] <= 1'b0;
     layer0_out[1430] <= x[294] | x[297];
     layer0_out[1431] <= ~(x[100] ^ x[104]);
     layer0_out[1432] <= x[282] | x[284];
     layer0_out[1433] <= x[5] & ~x[8];
     layer0_out[1434] <= x[58] | x[59];
     layer0_out[1435] <= ~x[83] | x[86];
     layer0_out[1436] <= x[22] | x[24];
     layer0_out[1437] <= 1'b0;
     layer0_out[1438] <= ~x[27];
     layer0_out[1439] <= ~x[222];
     layer0_out[1440] <= ~x[359];
     layer0_out[1441] <= x[135] | x[138];
     layer0_out[1442] <= 1'b1;
     layer0_out[1443] <= x[26] & x[29];
     layer0_out[1444] <= x[336] | x[338];
     layer0_out[1445] <= x[127];
     layer0_out[1446] <= x[179] | x[180];
     layer0_out[1447] <= x[297] | x[298];
     layer0_out[1448] <= x[218] | x[219];
     layer0_out[1449] <= x[312] | x[314];
     layer0_out[1450] <= ~x[15];
     layer0_out[1451] <= x[94];
     layer0_out[1452] <= 1'b1;
     layer0_out[1453] <= x[220] & ~x[216];
     layer0_out[1454] <= 1'b1;
     layer0_out[1455] <= x[208] | x[210];
     layer0_out[1456] <= ~(x[316] | x[318]);
     layer0_out[1457] <= x[112] | x[114];
     layer0_out[1458] <= 1'b0;
     layer0_out[1459] <= ~(x[354] & x[357]);
     layer0_out[1460] <= x[340] | x[341];
     layer0_out[1461] <= x[179];
     layer0_out[1462] <= x[240];
     layer0_out[1463] <= x[184] | x[187];
     layer0_out[1464] <= 1'b0;
     layer0_out[1465] <= ~x[78];
     layer0_out[1466] <= 1'b0;
     layer0_out[1467] <= ~(x[376] | x[379]);
     layer0_out[1468] <= ~x[364];
     layer0_out[1469] <= ~(x[234] | x[237]);
     layer0_out[1470] <= ~x[64] | x[68];
     layer0_out[1471] <= x[143] & ~x[147];
     layer0_out[1472] <= 1'b1;
     layer0_out[1473] <= x[280] | x[282];
     layer0_out[1474] <= x[379];
     layer0_out[1475] <= ~x[200];
     layer0_out[1476] <= x[176];
     layer0_out[1477] <= 1'b1;
     layer0_out[1478] <= x[41] | x[42];
     layer0_out[1479] <= x[62] | x[63];
     layer0_out[1480] <= x[42] & x[46];
     layer0_out[1481] <= x[101] & ~x[103];
     layer0_out[1482] <= 1'b1;
     layer0_out[1483] <= x[327];
     layer0_out[1484] <= x[281];
     layer0_out[1485] <= 1'b1;
     layer0_out[1486] <= 1'b1;
     layer0_out[1487] <= 1'b1;
     layer0_out[1488] <= ~(x[355] & x[357]);
     layer0_out[1489] <= ~(x[76] & x[80]);
     layer0_out[1490] <= ~(x[29] | x[31]);
     layer0_out[1491] <= ~(x[216] | x[218]);
     layer0_out[1492] <= x[153] | x[154];
     layer0_out[1493] <= 1'b1;
     layer0_out[1494] <= 1'b1;
     layer0_out[1495] <= x[8] & ~x[9];
     layer0_out[1496] <= x[81] & ~x[77];
     layer0_out[1497] <= ~(x[197] | x[198]);
     layer0_out[1498] <= ~x[36];
     layer0_out[1499] <= ~x[82];
     layer1_out[0] <= layer0_out[1195] & ~layer0_out[1194];
     layer1_out[1] <= ~layer0_out[550];
     layer1_out[2] <= layer0_out[74] & ~layer0_out[75];
     layer1_out[3] <= layer0_out[418];
     layer1_out[4] <= layer0_out[90];
     layer1_out[5] <= ~(layer0_out[662] & layer0_out[663]);
     layer1_out[6] <= ~layer0_out[356];
     layer1_out[7] <= ~layer0_out[99] | layer0_out[98];
     layer1_out[8] <= 1'b1;
     layer1_out[9] <= layer0_out[895] ^ layer0_out[896];
     layer1_out[10] <= layer0_out[199] & ~layer0_out[198];
     layer1_out[11] <= 1'b0;
     layer1_out[12] <= ~layer0_out[411] | layer0_out[410];
     layer1_out[13] <= ~(layer0_out[1013] | layer0_out[1014]);
     layer1_out[14] <= ~(layer0_out[179] & layer0_out[180]);
     layer1_out[15] <= 1'b0;
     layer1_out[16] <= layer0_out[104] | layer0_out[105];
     layer1_out[17] <= ~layer0_out[1278] | layer0_out[1279];
     layer1_out[18] <= layer0_out[1254];
     layer1_out[19] <= layer0_out[1377];
     layer1_out[20] <= ~layer0_out[589];
     layer1_out[21] <= layer0_out[337] & layer0_out[338];
     layer1_out[22] <= 1'b1;
     layer1_out[23] <= ~layer0_out[509] | layer0_out[510];
     layer1_out[24] <= 1'b1;
     layer1_out[25] <= ~layer0_out[25];
     layer1_out[26] <= layer0_out[709] ^ layer0_out[710];
     layer1_out[27] <= 1'b0;
     layer1_out[28] <= layer0_out[50];
     layer1_out[29] <= ~layer0_out[1142];
     layer1_out[30] <= 1'b1;
     layer1_out[31] <= ~layer0_out[1330];
     layer1_out[32] <= 1'b0;
     layer1_out[33] <= ~(layer0_out[529] & layer0_out[530]);
     layer1_out[34] <= ~layer0_out[720] | layer0_out[719];
     layer1_out[35] <= layer0_out[1345] | layer0_out[1346];
     layer1_out[36] <= layer0_out[277];
     layer1_out[37] <= ~(layer0_out[823] & layer0_out[824]);
     layer1_out[38] <= ~(layer0_out[692] & layer0_out[693]);
     layer1_out[39] <= ~layer0_out[1232] | layer0_out[1233];
     layer1_out[40] <= layer0_out[993] & ~layer0_out[994];
     layer1_out[41] <= ~layer0_out[94];
     layer1_out[42] <= ~layer0_out[1221] | layer0_out[1220];
     layer1_out[43] <= ~(layer0_out[425] | layer0_out[426]);
     layer1_out[44] <= ~layer0_out[630] | layer0_out[629];
     layer1_out[45] <= ~layer0_out[357];
     layer1_out[46] <= layer0_out[693] | layer0_out[694];
     layer1_out[47] <= 1'b0;
     layer1_out[48] <= 1'b1;
     layer1_out[49] <= 1'b1;
     layer1_out[50] <= layer0_out[445] & layer0_out[446];
     layer1_out[51] <= ~(layer0_out[1275] & layer0_out[1276]);
     layer1_out[52] <= ~(layer0_out[1426] | layer0_out[1427]);
     layer1_out[53] <= ~(layer0_out[1072] & layer0_out[1073]);
     layer1_out[54] <= 1'b1;
     layer1_out[55] <= ~(layer0_out[269] | layer0_out[270]);
     layer1_out[56] <= ~(layer0_out[1266] & layer0_out[1267]);
     layer1_out[57] <= layer0_out[187] & layer0_out[188];
     layer1_out[58] <= layer0_out[674] | layer0_out[675];
     layer1_out[59] <= layer0_out[912] | layer0_out[913];
     layer1_out[60] <= 1'b1;
     layer1_out[61] <= ~(layer0_out[714] ^ layer0_out[715]);
     layer1_out[62] <= layer0_out[472] & ~layer0_out[471];
     layer1_out[63] <= ~layer0_out[1210];
     layer1_out[64] <= 1'b0;
     layer1_out[65] <= ~(layer0_out[1356] | layer0_out[1357]);
     layer1_out[66] <= ~(layer0_out[1062] | layer0_out[1063]);
     layer1_out[67] <= layer0_out[957] & ~layer0_out[958];
     layer1_out[68] <= layer0_out[468];
     layer1_out[69] <= layer0_out[56] & ~layer0_out[55];
     layer1_out[70] <= ~layer0_out[1431] | layer0_out[1432];
     layer1_out[71] <= ~(layer0_out[554] & layer0_out[555]);
     layer1_out[72] <= ~layer0_out[1398] | layer0_out[1399];
     layer1_out[73] <= layer0_out[629];
     layer1_out[74] <= 1'b1;
     layer1_out[75] <= 1'b1;
     layer1_out[76] <= ~(layer0_out[514] | layer0_out[515]);
     layer1_out[77] <= 1'b0;
     layer1_out[78] <= layer0_out[207];
     layer1_out[79] <= layer0_out[859];
     layer1_out[80] <= ~(layer0_out[138] | layer0_out[139]);
     layer1_out[81] <= ~layer0_out[1109];
     layer1_out[82] <= layer0_out[570] & ~layer0_out[569];
     layer1_out[83] <= layer0_out[688] & ~layer0_out[687];
     layer1_out[84] <= ~layer0_out[1344] | layer0_out[1345];
     layer1_out[85] <= layer0_out[450] | layer0_out[451];
     layer1_out[86] <= 1'b1;
     layer1_out[87] <= ~layer0_out[309];
     layer1_out[88] <= 1'b0;
     layer1_out[89] <= 1'b0;
     layer1_out[90] <= layer0_out[1388] & ~layer0_out[1389];
     layer1_out[91] <= ~layer0_out[1395];
     layer1_out[92] <= layer0_out[1047] | layer0_out[1048];
     layer1_out[93] <= ~layer0_out[359];
     layer1_out[94] <= 1'b0;
     layer1_out[95] <= layer0_out[1086] & layer0_out[1087];
     layer1_out[96] <= ~layer0_out[665];
     layer1_out[97] <= layer0_out[624] & layer0_out[625];
     layer1_out[98] <= ~layer0_out[51] | layer0_out[50];
     layer1_out[99] <= layer0_out[670] & ~layer0_out[671];
     layer1_out[100] <= layer0_out[369];
     layer1_out[101] <= layer0_out[42];
     layer1_out[102] <= layer0_out[1240];
     layer1_out[103] <= ~layer0_out[1228] | layer0_out[1227];
     layer1_out[104] <= layer0_out[575] & layer0_out[576];
     layer1_out[105] <= layer0_out[293] | layer0_out[294];
     layer1_out[106] <= layer0_out[290] & ~layer0_out[291];
     layer1_out[107] <= layer0_out[731];
     layer1_out[108] <= layer0_out[43] | layer0_out[44];
     layer1_out[109] <= ~layer0_out[66];
     layer1_out[110] <= layer0_out[1174];
     layer1_out[111] <= layer0_out[1201] & layer0_out[1202];
     layer1_out[112] <= layer0_out[1409];
     layer1_out[113] <= 1'b0;
     layer1_out[114] <= layer0_out[512];
     layer1_out[115] <= ~(layer0_out[1150] & layer0_out[1151]);
     layer1_out[116] <= 1'b1;
     layer1_out[117] <= 1'b0;
     layer1_out[118] <= layer0_out[1212] | layer0_out[1213];
     layer1_out[119] <= ~layer0_out[648] | layer0_out[649];
     layer1_out[120] <= ~layer0_out[316] | layer0_out[315];
     layer1_out[121] <= layer0_out[1214];
     layer1_out[122] <= layer0_out[1390] & layer0_out[1391];
     layer1_out[123] <= ~(layer0_out[442] & layer0_out[443]);
     layer1_out[124] <= 1'b0;
     layer1_out[125] <= layer0_out[328] | layer0_out[329];
     layer1_out[126] <= ~(layer0_out[1071] & layer0_out[1072]);
     layer1_out[127] <= ~layer0_out[480];
     layer1_out[128] <= layer0_out[953] | layer0_out[954];
     layer1_out[129] <= ~layer0_out[35] | layer0_out[36];
     layer1_out[130] <= layer0_out[92];
     layer1_out[131] <= ~(layer0_out[617] ^ layer0_out[618]);
     layer1_out[132] <= 1'b1;
     layer1_out[133] <= layer0_out[330] & layer0_out[331];
     layer1_out[134] <= ~layer0_out[1405];
     layer1_out[135] <= layer0_out[1324];
     layer1_out[136] <= ~layer0_out[1013];
     layer1_out[137] <= layer0_out[515] | layer0_out[516];
     layer1_out[138] <= ~(layer0_out[484] & layer0_out[485]);
     layer1_out[139] <= ~(layer0_out[720] & layer0_out[721]);
     layer1_out[140] <= ~layer0_out[222] | layer0_out[221];
     layer1_out[141] <= layer0_out[59];
     layer1_out[142] <= ~layer0_out[332] | layer0_out[331];
     layer1_out[143] <= ~layer0_out[1245];
     layer1_out[144] <= ~layer0_out[1319] | layer0_out[1318];
     layer1_out[145] <= layer0_out[965];
     layer1_out[146] <= ~(layer0_out[1229] | layer0_out[1230]);
     layer1_out[147] <= layer0_out[631] & layer0_out[632];
     layer1_out[148] <= ~(layer0_out[682] & layer0_out[683]);
     layer1_out[149] <= ~layer0_out[1137];
     layer1_out[150] <= ~layer0_out[1327] | layer0_out[1326];
     layer1_out[151] <= ~layer0_out[424] | layer0_out[423];
     layer1_out[152] <= layer0_out[362];
     layer1_out[153] <= 1'b1;
     layer1_out[154] <= layer0_out[1495] & layer0_out[1496];
     layer1_out[155] <= layer0_out[1147] | layer0_out[1148];
     layer1_out[156] <= layer0_out[321] & ~layer0_out[322];
     layer1_out[157] <= layer0_out[830] | layer0_out[831];
     layer1_out[158] <= layer0_out[976] & ~layer0_out[977];
     layer1_out[159] <= 1'b1;
     layer1_out[160] <= layer0_out[177];
     layer1_out[161] <= ~layer0_out[882] | layer0_out[883];
     layer1_out[162] <= ~layer0_out[212] | layer0_out[211];
     layer1_out[163] <= layer0_out[1295] & layer0_out[1296];
     layer1_out[164] <= layer0_out[595] & ~layer0_out[594];
     layer1_out[165] <= ~(layer0_out[947] & layer0_out[948]);
     layer1_out[166] <= ~(layer0_out[840] ^ layer0_out[841]);
     layer1_out[167] <= layer0_out[27] & ~layer0_out[26];
     layer1_out[168] <= ~(layer0_out[1169] | layer0_out[1170]);
     layer1_out[169] <= layer0_out[806] & ~layer0_out[807];
     layer1_out[170] <= layer0_out[181] ^ layer0_out[182];
     layer1_out[171] <= layer0_out[324] & ~layer0_out[323];
     layer1_out[172] <= ~layer0_out[1446];
     layer1_out[173] <= ~layer0_out[165];
     layer1_out[174] <= 1'b1;
     layer1_out[175] <= 1'b0;
     layer1_out[176] <= ~(layer0_out[952] & layer0_out[953]);
     layer1_out[177] <= ~(layer0_out[1466] | layer0_out[1467]);
     layer1_out[178] <= 1'b0;
     layer1_out[179] <= layer0_out[145] & ~layer0_out[146];
     layer1_out[180] <= layer0_out[272];
     layer1_out[181] <= 1'b1;
     layer1_out[182] <= layer0_out[354] & layer0_out[355];
     layer1_out[183] <= layer0_out[1264] | layer0_out[1265];
     layer1_out[184] <= ~(layer0_out[503] | layer0_out[504]);
     layer1_out[185] <= layer0_out[247] & layer0_out[248];
     layer1_out[186] <= ~layer0_out[809];
     layer1_out[187] <= layer0_out[1284] & ~layer0_out[1285];
     layer1_out[188] <= ~layer0_out[1005] | layer0_out[1004];
     layer1_out[189] <= ~layer0_out[170] | layer0_out[171];
     layer1_out[190] <= ~(layer0_out[139] & layer0_out[140]);
     layer1_out[191] <= layer0_out[961];
     layer1_out[192] <= ~(layer0_out[1396] & layer0_out[1397]);
     layer1_out[193] <= ~layer0_out[362] | layer0_out[363];
     layer1_out[194] <= ~(layer0_out[252] | layer0_out[253]);
     layer1_out[195] <= ~layer0_out[540];
     layer1_out[196] <= layer0_out[1440] ^ layer0_out[1441];
     layer1_out[197] <= 1'b0;
     layer1_out[198] <= ~(layer0_out[653] & layer0_out[654]);
     layer1_out[199] <= ~(layer0_out[350] | layer0_out[351]);
     layer1_out[200] <= ~(layer0_out[386] | layer0_out[387]);
     layer1_out[201] <= layer0_out[193] & ~layer0_out[194];
     layer1_out[202] <= ~layer0_out[191];
     layer1_out[203] <= layer0_out[682];
     layer1_out[204] <= ~layer0_out[1058];
     layer1_out[205] <= ~layer0_out[550] | layer0_out[549];
     layer1_out[206] <= layer0_out[1];
     layer1_out[207] <= layer0_out[289] & layer0_out[290];
     layer1_out[208] <= layer0_out[300];
     layer1_out[209] <= layer0_out[1280];
     layer1_out[210] <= layer0_out[190] | layer0_out[191];
     layer1_out[211] <= 1'b1;
     layer1_out[212] <= 1'b0;
     layer1_out[213] <= 1'b0;
     layer1_out[214] <= ~layer0_out[548];
     layer1_out[215] <= ~(layer0_out[982] & layer0_out[983]);
     layer1_out[216] <= ~layer0_out[914] | layer0_out[915];
     layer1_out[217] <= layer0_out[544] | layer0_out[545];
     layer1_out[218] <= ~layer0_out[380];
     layer1_out[219] <= ~layer0_out[985] | layer0_out[984];
     layer1_out[220] <= ~(layer0_out[1330] & layer0_out[1331]);
     layer1_out[221] <= layer0_out[61];
     layer1_out[222] <= 1'b0;
     layer1_out[223] <= 1'b0;
     layer1_out[224] <= layer0_out[189] & ~layer0_out[188];
     layer1_out[225] <= layer0_out[1039] | layer0_out[1040];
     layer1_out[226] <= layer0_out[1378] & layer0_out[1379];
     layer1_out[227] <= ~layer0_out[224] | layer0_out[225];
     layer1_out[228] <= ~layer0_out[980] | layer0_out[981];
     layer1_out[229] <= ~(layer0_out[805] & layer0_out[806]);
     layer1_out[230] <= layer0_out[1479] & ~layer0_out[1480];
     layer1_out[231] <= ~layer0_out[1416] | layer0_out[1417];
     layer1_out[232] <= layer0_out[172];
     layer1_out[233] <= ~(layer0_out[769] & layer0_out[770]);
     layer1_out[234] <= layer0_out[1341] & layer0_out[1342];
     layer1_out[235] <= ~layer0_out[268] | layer0_out[269];
     layer1_out[236] <= layer0_out[716];
     layer1_out[237] <= 1'b0;
     layer1_out[238] <= ~layer0_out[1219] | layer0_out[1218];
     layer1_out[239] <= ~(layer0_out[1498] & layer0_out[1499]);
     layer1_out[240] <= ~layer0_out[106] | layer0_out[105];
     layer1_out[241] <= layer0_out[367] & ~layer0_out[368];
     layer1_out[242] <= ~layer0_out[1460] | layer0_out[1461];
     layer1_out[243] <= ~layer0_out[1200];
     layer1_out[244] <= ~(layer0_out[505] | layer0_out[506]);
     layer1_out[245] <= layer0_out[1301];
     layer1_out[246] <= layer0_out[756] & layer0_out[757];
     layer1_out[247] <= layer0_out[873] | layer0_out[874];
     layer1_out[248] <= ~(layer0_out[578] | layer0_out[579]);
     layer1_out[249] <= ~(layer0_out[851] & layer0_out[852]);
     layer1_out[250] <= ~(layer0_out[1310] & layer0_out[1311]);
     layer1_out[251] <= layer0_out[1298];
     layer1_out[252] <= ~(layer0_out[203] | layer0_out[204]);
     layer1_out[253] <= layer0_out[532] & ~layer0_out[531];
     layer1_out[254] <= 1'b1;
     layer1_out[255] <= layer0_out[866] | layer0_out[867];
     layer1_out[256] <= 1'b1;
     layer1_out[257] <= ~layer0_out[148];
     layer1_out[258] <= ~layer0_out[571] | layer0_out[572];
     layer1_out[259] <= 1'b0;
     layer1_out[260] <= layer0_out[270] & ~layer0_out[271];
     layer1_out[261] <= layer0_out[1008] & ~layer0_out[1009];
     layer1_out[262] <= layer0_out[1462];
     layer1_out[263] <= layer0_out[84] | layer0_out[85];
     layer1_out[264] <= layer0_out[3] & ~layer0_out[2];
     layer1_out[265] <= 1'b0;
     layer1_out[266] <= layer0_out[20];
     layer1_out[267] <= 1'b0;
     layer1_out[268] <= layer0_out[1242] | layer0_out[1243];
     layer1_out[269] <= layer0_out[97] | layer0_out[98];
     layer1_out[270] <= ~layer0_out[614];
     layer1_out[271] <= layer0_out[1382] | layer0_out[1383];
     layer1_out[272] <= ~layer0_out[245];
     layer1_out[273] <= layer0_out[747] & ~layer0_out[746];
     layer1_out[274] <= ~(layer0_out[742] | layer0_out[743]);
     layer1_out[275] <= ~(layer0_out[233] | layer0_out[234]);
     layer1_out[276] <= 1'b1;
     layer1_out[277] <= ~layer0_out[1082] | layer0_out[1083];
     layer1_out[278] <= ~(layer0_out[831] | layer0_out[832]);
     layer1_out[279] <= 1'b0;
     layer1_out[280] <= layer0_out[225];
     layer1_out[281] <= layer0_out[1269] & ~layer0_out[1268];
     layer1_out[282] <= ~(layer0_out[1074] | layer0_out[1075]);
     layer1_out[283] <= layer0_out[1120] & layer0_out[1121];
     layer1_out[284] <= ~(layer0_out[110] | layer0_out[111]);
     layer1_out[285] <= layer0_out[1178] & ~layer0_out[1177];
     layer1_out[286] <= layer0_out[611];
     layer1_out[287] <= layer0_out[739];
     layer1_out[288] <= layer0_out[638] ^ layer0_out[639];
     layer1_out[289] <= ~layer0_out[853];
     layer1_out[290] <= ~layer0_out[418] | layer0_out[419];
     layer1_out[291] <= ~(layer0_out[1444] | layer0_out[1445]);
     layer1_out[292] <= layer0_out[229] & ~layer0_out[228];
     layer1_out[293] <= layer0_out[1467] | layer0_out[1468];
     layer1_out[294] <= 1'b1;
     layer1_out[295] <= 1'b0;
     layer1_out[296] <= ~layer0_out[1133];
     layer1_out[297] <= ~layer0_out[1392];
     layer1_out[298] <= ~layer0_out[79];
     layer1_out[299] <= ~layer0_out[256] | layer0_out[255];
     layer1_out[300] <= ~(layer0_out[125] & layer0_out[126]);
     layer1_out[301] <= ~layer0_out[1176];
     layer1_out[302] <= layer0_out[971] & ~layer0_out[970];
     layer1_out[303] <= layer0_out[655] & ~layer0_out[654];
     layer1_out[304] <= ~(layer0_out[340] & layer0_out[341]);
     layer1_out[305] <= 1'b1;
     layer1_out[306] <= ~layer0_out[404];
     layer1_out[307] <= layer0_out[602];
     layer1_out[308] <= ~layer0_out[454];
     layer1_out[309] <= ~layer0_out[195] | layer0_out[194];
     layer1_out[310] <= layer0_out[481];
     layer1_out[311] <= layer0_out[881];
     layer1_out[312] <= 1'b0;
     layer1_out[313] <= ~layer0_out[923] | layer0_out[924];
     layer1_out[314] <= layer0_out[310] & ~layer0_out[309];
     layer1_out[315] <= ~(layer0_out[16] | layer0_out[17]);
     layer1_out[316] <= ~layer0_out[1219] | layer0_out[1220];
     layer1_out[317] <= ~(layer0_out[604] | layer0_out[605]);
     layer1_out[318] <= layer0_out[151] | layer0_out[152];
     layer1_out[319] <= ~layer0_out[955];
     layer1_out[320] <= layer0_out[672] & ~layer0_out[671];
     layer1_out[321] <= ~layer0_out[660];
     layer1_out[322] <= 1'b1;
     layer1_out[323] <= ~layer0_out[493] | layer0_out[492];
     layer1_out[324] <= layer0_out[382];
     layer1_out[325] <= ~layer0_out[489] | layer0_out[490];
     layer1_out[326] <= 1'b0;
     layer1_out[327] <= layer0_out[253] | layer0_out[254];
     layer1_out[328] <= 1'b1;
     layer1_out[329] <= 1'b1;
     layer1_out[330] <= ~layer0_out[336];
     layer1_out[331] <= 1'b1;
     layer1_out[332] <= ~layer0_out[1021] | layer0_out[1020];
     layer1_out[333] <= ~(layer0_out[1476] | layer0_out[1477]);
     layer1_out[334] <= layer0_out[1241] | layer0_out[1242];
     layer1_out[335] <= layer0_out[1473] & ~layer0_out[1474];
     layer1_out[336] <= 1'b1;
     layer1_out[337] <= layer0_out[729] & layer0_out[730];
     layer1_out[338] <= layer0_out[298] & layer0_out[299];
     layer1_out[339] <= layer0_out[22] & ~layer0_out[21];
     layer1_out[340] <= layer0_out[352] & ~layer0_out[351];
     layer1_out[341] <= ~(layer0_out[88] ^ layer0_out[89]);
     layer1_out[342] <= ~layer0_out[120] | layer0_out[121];
     layer1_out[343] <= layer0_out[1385];
     layer1_out[344] <= layer0_out[972] & layer0_out[973];
     layer1_out[345] <= ~layer0_out[65];
     layer1_out[346] <= ~layer0_out[460] | layer0_out[459];
     layer1_out[347] <= ~layer0_out[583] | layer0_out[582];
     layer1_out[348] <= 1'b0;
     layer1_out[349] <= 1'b1;
     layer1_out[350] <= ~(layer0_out[768] & layer0_out[769]);
     layer1_out[351] <= ~layer0_out[408];
     layer1_out[352] <= 1'b1;
     layer1_out[353] <= 1'b0;
     layer1_out[354] <= 1'b1;
     layer1_out[355] <= ~layer0_out[1239];
     layer1_out[356] <= ~layer0_out[489];
     layer1_out[357] <= 1'b1;
     layer1_out[358] <= 1'b0;
     layer1_out[359] <= ~(layer0_out[992] ^ layer0_out[993]);
     layer1_out[360] <= layer0_out[1411] & ~layer0_out[1410];
     layer1_out[361] <= 1'b0;
     layer1_out[362] <= layer0_out[1443] & layer0_out[1444];
     layer1_out[363] <= 1'b0;
     layer1_out[364] <= layer0_out[1235];
     layer1_out[365] <= ~(layer0_out[998] | layer0_out[999]);
     layer1_out[366] <= 1'b0;
     layer1_out[367] <= 1'b1;
     layer1_out[368] <= 1'b0;
     layer1_out[369] <= 1'b0;
     layer1_out[370] <= 1'b0;
     layer1_out[371] <= ~(layer0_out[523] | layer0_out[524]);
     layer1_out[372] <= ~layer0_out[497];
     layer1_out[373] <= layer0_out[374];
     layer1_out[374] <= layer0_out[118] & layer0_out[119];
     layer1_out[375] <= ~layer0_out[214] | layer0_out[215];
     layer1_out[376] <= layer0_out[591] | layer0_out[592];
     layer1_out[377] <= 1'b0;
     layer1_out[378] <= ~layer0_out[520] | layer0_out[519];
     layer1_out[379] <= ~layer0_out[375];
     layer1_out[380] <= layer0_out[1025] & ~layer0_out[1026];
     layer1_out[381] <= layer0_out[279] & layer0_out[280];
     layer1_out[382] <= layer0_out[785];
     layer1_out[383] <= 1'b0;
     layer1_out[384] <= 1'b1;
     layer1_out[385] <= layer0_out[1453] & ~layer0_out[1452];
     layer1_out[386] <= layer0_out[281] & ~layer0_out[280];
     layer1_out[387] <= layer0_out[564];
     layer1_out[388] <= layer0_out[1227];
     layer1_out[389] <= layer0_out[709];
     layer1_out[390] <= layer0_out[938];
     layer1_out[391] <= ~layer0_out[262] | layer0_out[261];
     layer1_out[392] <= layer0_out[1449];
     layer1_out[393] <= ~layer0_out[780] | layer0_out[779];
     layer1_out[394] <= ~layer0_out[123] | layer0_out[124];
     layer1_out[395] <= layer0_out[91];
     layer1_out[396] <= 1'b0;
     layer1_out[397] <= ~layer0_out[943];
     layer1_out[398] <= ~layer0_out[741];
     layer1_out[399] <= layer0_out[1360];
     layer1_out[400] <= 1'b1;
     layer1_out[401] <= 1'b0;
     layer1_out[402] <= ~layer0_out[1147] | layer0_out[1146];
     layer1_out[403] <= layer0_out[568];
     layer1_out[404] <= ~layer0_out[1278] | layer0_out[1277];
     layer1_out[405] <= ~layer0_out[277];
     layer1_out[406] <= ~layer0_out[1032];
     layer1_out[407] <= layer0_out[1070] & ~layer0_out[1069];
     layer1_out[408] <= 1'b1;
     layer1_out[409] <= layer0_out[849];
     layer1_out[410] <= ~layer0_out[1132];
     layer1_out[411] <= ~(layer0_out[590] ^ layer0_out[591]);
     layer1_out[412] <= ~(layer0_out[1021] & layer0_out[1022]);
     layer1_out[413] <= layer0_out[1287];
     layer1_out[414] <= layer0_out[1175] & layer0_out[1176];
     layer1_out[415] <= ~(layer0_out[466] & layer0_out[467]);
     layer1_out[416] <= ~layer0_out[1134];
     layer1_out[417] <= layer0_out[726] & ~layer0_out[727];
     layer1_out[418] <= ~(layer0_out[140] & layer0_out[141]);
     layer1_out[419] <= layer0_out[339] | layer0_out[340];
     layer1_out[420] <= layer0_out[755] & ~layer0_out[754];
     layer1_out[421] <= layer0_out[773];
     layer1_out[422] <= ~(layer0_out[790] & layer0_out[791]);
     layer1_out[423] <= ~(layer0_out[1455] & layer0_out[1456]);
     layer1_out[424] <= 1'b0;
     layer1_out[425] <= layer0_out[1195];
     layer1_out[426] <= ~(layer0_out[152] & layer0_out[153]);
     layer1_out[427] <= layer0_out[304] & ~layer0_out[305];
     layer1_out[428] <= layer0_out[1201];
     layer1_out[429] <= layer0_out[14] ^ layer0_out[15];
     layer1_out[430] <= ~layer0_out[1437] | layer0_out[1438];
     layer1_out[431] <= 1'b1;
     layer1_out[432] <= layer0_out[792];
     layer1_out[433] <= ~(layer0_out[1123] | layer0_out[1124]);
     layer1_out[434] <= 1'b1;
     layer1_out[435] <= ~layer0_out[922] | layer0_out[921];
     layer1_out[436] <= ~layer0_out[904] | layer0_out[905];
     layer1_out[437] <= 1'b1;
     layer1_out[438] <= ~(layer0_out[1029] | layer0_out[1030]);
     layer1_out[439] <= ~layer0_out[127] | layer0_out[126];
     layer1_out[440] <= layer0_out[808] | layer0_out[809];
     layer1_out[441] <= layer0_out[1151] | layer0_out[1152];
     layer1_out[442] <= ~(layer0_out[1406] & layer0_out[1407]);
     layer1_out[443] <= 1'b1;
     layer1_out[444] <= 1'b0;
     layer1_out[445] <= layer0_out[160];
     layer1_out[446] <= ~layer0_out[645] | layer0_out[646];
     layer1_out[447] <= layer0_out[1362];
     layer1_out[448] <= 1'b0;
     layer1_out[449] <= ~(layer0_out[204] | layer0_out[205]);
     layer1_out[450] <= ~(layer0_out[1114] | layer0_out[1115]);
     layer1_out[451] <= layer0_out[1386];
     layer1_out[452] <= layer0_out[1368] & ~layer0_out[1369];
     layer1_out[453] <= layer0_out[910] & ~layer0_out[911];
     layer1_out[454] <= layer0_out[1081] | layer0_out[1082];
     layer1_out[455] <= layer0_out[1054] & ~layer0_out[1053];
     layer1_out[456] <= ~layer0_out[68] | layer0_out[69];
     layer1_out[457] <= ~layer0_out[284] | layer0_out[285];
     layer1_out[458] <= 1'b1;
     layer1_out[459] <= 1'b1;
     layer1_out[460] <= ~layer0_out[1293];
     layer1_out[461] <= layer0_out[318];
     layer1_out[462] <= layer0_out[502];
     layer1_out[463] <= layer0_out[1033];
     layer1_out[464] <= layer0_out[1350] & layer0_out[1351];
     layer1_out[465] <= layer0_out[743] & ~layer0_out[744];
     layer1_out[466] <= 1'b0;
     layer1_out[467] <= ~layer0_out[218];
     layer1_out[468] <= 1'b0;
     layer1_out[469] <= layer0_out[1475] | layer0_out[1476];
     layer1_out[470] <= ~(layer0_out[345] | layer0_out[346]);
     layer1_out[471] <= layer0_out[1491] ^ layer0_out[1492];
     layer1_out[472] <= layer0_out[275] & ~layer0_out[274];
     layer1_out[473] <= ~layer0_out[484];
     layer1_out[474] <= ~layer0_out[673];
     layer1_out[475] <= 1'b1;
     layer1_out[476] <= ~layer0_out[1038] | layer0_out[1039];
     layer1_out[477] <= 1'b1;
     layer1_out[478] <= 1'b1;
     layer1_out[479] <= ~layer0_out[664];
     layer1_out[480] <= layer0_out[607] & layer0_out[608];
     layer1_out[481] <= ~layer0_out[838];
     layer1_out[482] <= layer0_out[981] | layer0_out[982];
     layer1_out[483] <= layer0_out[788] & ~layer0_out[789];
     layer1_out[484] <= ~layer0_out[1421];
     layer1_out[485] <= layer0_out[420] & layer0_out[421];
     layer1_out[486] <= layer0_out[1256];
     layer1_out[487] <= ~(layer0_out[1009] | layer0_out[1010]);
     layer1_out[488] <= layer0_out[612] & layer0_out[613];
     layer1_out[489] <= ~layer0_out[976] | layer0_out[975];
     layer1_out[490] <= ~layer0_out[1209];
     layer1_out[491] <= layer0_out[82] ^ layer0_out[83];
     layer1_out[492] <= 1'b1;
     layer1_out[493] <= ~layer0_out[495];
     layer1_out[494] <= ~(layer0_out[537] | layer0_out[538]);
     layer1_out[495] <= layer0_out[856];
     layer1_out[496] <= 1'b1;
     layer1_out[497] <= layer0_out[1370] & ~layer0_out[1371];
     layer1_out[498] <= 1'b1;
     layer1_out[499] <= 1'b1;
     layer1_out[500] <= layer0_out[686];
     layer1_out[501] <= ~(layer0_out[482] | layer0_out[483]);
     layer1_out[502] <= layer0_out[1334];
     layer1_out[503] <= ~layer0_out[477];
     layer1_out[504] <= ~(layer0_out[1113] | layer0_out[1114]);
     layer1_out[505] <= layer0_out[1311] | layer0_out[1312];
     layer1_out[506] <= ~layer0_out[994] | layer0_out[995];
     layer1_out[507] <= 1'b0;
     layer1_out[508] <= layer0_out[228];
     layer1_out[509] <= 1'b1;
     layer1_out[510] <= 1'b0;
     layer1_out[511] <= layer0_out[1312] & ~layer0_out[1313];
     layer1_out[512] <= layer0_out[1349];
     layer1_out[513] <= layer0_out[1416];
     layer1_out[514] <= layer0_out[639] | layer0_out[640];
     layer1_out[515] <= ~(layer0_out[909] & layer0_out[910]);
     layer1_out[516] <= ~layer0_out[1490];
     layer1_out[517] <= layer0_out[440] & ~layer0_out[439];
     layer1_out[518] <= ~layer0_out[1300];
     layer1_out[519] <= ~layer0_out[669] | layer0_out[670];
     layer1_out[520] <= ~layer0_out[1434];
     layer1_out[521] <= layer0_out[407];
     layer1_out[522] <= layer0_out[281] & ~layer0_out[282];
     layer1_out[523] <= layer0_out[329] & layer0_out[330];
     layer1_out[524] <= layer0_out[1246];
     layer1_out[525] <= layer0_out[819] | layer0_out[820];
     layer1_out[526] <= layer0_out[437];
     layer1_out[527] <= layer0_out[1125] & ~layer0_out[1124];
     layer1_out[528] <= ~layer0_out[615];
     layer1_out[529] <= 1'b0;
     layer1_out[530] <= 1'b1;
     layer1_out[531] <= 1'b0;
     layer1_out[532] <= ~(layer0_out[757] & layer0_out[758]);
     layer1_out[533] <= layer0_out[1472];
     layer1_out[534] <= layer0_out[619] & layer0_out[620];
     layer1_out[535] <= 1'b1;
     layer1_out[536] <= layer0_out[1318];
     layer1_out[537] <= 1'b0;
     layer1_out[538] <= ~(layer0_out[1383] | layer0_out[1384]);
     layer1_out[539] <= layer0_out[15];
     layer1_out[540] <= 1'b0;
     layer1_out[541] <= layer0_out[1211] | layer0_out[1212];
     layer1_out[542] <= 1'b1;
     layer1_out[543] <= ~(layer0_out[102] | layer0_out[103]);
     layer1_out[544] <= layer0_out[373] & ~layer0_out[374];
     layer1_out[545] <= layer0_out[1158] & ~layer0_out[1157];
     layer1_out[546] <= 1'b1;
     layer1_out[547] <= layer0_out[584];
     layer1_out[548] <= ~layer0_out[795] | layer0_out[794];
     layer1_out[549] <= ~(layer0_out[254] | layer0_out[255]);
     layer1_out[550] <= layer0_out[1349];
     layer1_out[551] <= ~layer0_out[861] | layer0_out[860];
     layer1_out[552] <= 1'b0;
     layer1_out[553] <= layer0_out[906] | layer0_out[907];
     layer1_out[554] <= ~(layer0_out[173] & layer0_out[174]);
     layer1_out[555] <= ~(layer0_out[333] | layer0_out[334]);
     layer1_out[556] <= layer0_out[1260] & ~layer0_out[1259];
     layer1_out[557] <= layer0_out[558];
     layer1_out[558] <= layer0_out[567] & ~layer0_out[566];
     layer1_out[559] <= layer0_out[867];
     layer1_out[560] <= layer0_out[570];
     layer1_out[561] <= ~layer0_out[549] | layer0_out[548];
     layer1_out[562] <= 1'b1;
     layer1_out[563] <= layer0_out[272] & ~layer0_out[271];
     layer1_out[564] <= ~layer0_out[950];
     layer1_out[565] <= ~layer0_out[137];
     layer1_out[566] <= 1'b0;
     layer1_out[567] <= layer0_out[1389] | layer0_out[1390];
     layer1_out[568] <= ~layer0_out[1043];
     layer1_out[569] <= layer0_out[546] & layer0_out[547];
     layer1_out[570] <= ~layer0_out[607] | layer0_out[606];
     layer1_out[571] <= ~(layer0_out[900] & layer0_out[901]);
     layer1_out[572] <= layer0_out[958] & layer0_out[959];
     layer1_out[573] <= ~layer0_out[397] | layer0_out[396];
     layer1_out[574] <= ~(layer0_out[244] | layer0_out[245]);
     layer1_out[575] <= layer0_out[1471];
     layer1_out[576] <= ~(layer0_out[415] | layer0_out[416]);
     layer1_out[577] <= layer0_out[1204];
     layer1_out[578] <= 1'b1;
     layer1_out[579] <= ~layer0_out[162] | layer0_out[163];
     layer1_out[580] <= ~(layer0_out[1019] & layer0_out[1020]);
     layer1_out[581] <= 1'b1;
     layer1_out[582] <= ~layer0_out[1275] | layer0_out[1274];
     layer1_out[583] <= layer0_out[839] & ~layer0_out[840];
     layer1_out[584] <= ~layer0_out[616];
     layer1_out[585] <= ~layer0_out[686];
     layer1_out[586] <= layer0_out[1289] & layer0_out[1290];
     layer1_out[587] <= ~layer0_out[1488] | layer0_out[1487];
     layer1_out[588] <= 1'b0;
     layer1_out[589] <= ~layer0_out[1294] | layer0_out[1295];
     layer1_out[590] <= ~layer0_out[647];
     layer1_out[591] <= ~(layer0_out[1091] ^ layer0_out[1092]);
     layer1_out[592] <= ~layer0_out[979];
     layer1_out[593] <= 1'b1;
     layer1_out[594] <= ~(layer0_out[96] | layer0_out[97]);
     layer1_out[595] <= 1'b0;
     layer1_out[596] <= ~layer0_out[70] | layer0_out[71];
     layer1_out[597] <= ~layer0_out[116] | layer0_out[117];
     layer1_out[598] <= 1'b1;
     layer1_out[599] <= ~(layer0_out[861] ^ layer0_out[862]);
     layer1_out[600] <= ~layer0_out[1092];
     layer1_out[601] <= layer0_out[1138] & layer0_out[1139];
     layer1_out[602] <= 1'b1;
     layer1_out[603] <= layer0_out[893] | layer0_out[894];
     layer1_out[604] <= ~layer0_out[668] | layer0_out[669];
     layer1_out[605] <= 1'b0;
     layer1_out[606] <= layer0_out[766] & ~layer0_out[765];
     layer1_out[607] <= 1'b1;
     layer1_out[608] <= ~(layer0_out[195] & layer0_out[196]);
     layer1_out[609] <= ~(layer0_out[133] | layer0_out[134]);
     layer1_out[610] <= 1'b0;
     layer1_out[611] <= ~layer0_out[49] | layer0_out[48];
     layer1_out[612] <= 1'b0;
     layer1_out[613] <= 1'b1;
     layer1_out[614] <= ~(layer0_out[1462] ^ layer0_out[1463]);
     layer1_out[615] <= 1'b0;
     layer1_out[616] <= layer0_out[533] & layer0_out[534];
     layer1_out[617] <= ~(layer0_out[395] & layer0_out[396]);
     layer1_out[618] <= layer0_out[531];
     layer1_out[619] <= layer0_out[1367];
     layer1_out[620] <= 1'b0;
     layer1_out[621] <= layer0_out[209] & ~layer0_out[210];
     layer1_out[622] <= 1'b0;
     layer1_out[623] <= 1'b0;
     layer1_out[624] <= 1'b0;
     layer1_out[625] <= 1'b1;
     layer1_out[626] <= ~(layer0_out[475] | layer0_out[476]);
     layer1_out[627] <= layer0_out[858] & ~layer0_out[857];
     layer1_out[628] <= ~layer0_out[286] | layer0_out[287];
     layer1_out[629] <= layer0_out[23];
     layer1_out[630] <= layer0_out[1430] | layer0_out[1431];
     layer1_out[631] <= layer0_out[795] | layer0_out[796];
     layer1_out[632] <= ~layer0_out[176];
     layer1_out[633] <= layer0_out[1071] & ~layer0_out[1070];
     layer1_out[634] <= layer0_out[753] & ~layer0_out[754];
     layer1_out[635] <= layer0_out[1117] & ~layer0_out[1118];
     layer1_out[636] <= 1'b1;
     layer1_out[637] <= layer0_out[574];
     layer1_out[638] <= ~(layer0_out[143] | layer0_out[144]);
     layer1_out[639] <= 1'b0;
     layer1_out[640] <= ~(layer0_out[858] | layer0_out[859]);
     layer1_out[641] <= layer0_out[763] & ~layer0_out[764];
     layer1_out[642] <= ~layer0_out[577];
     layer1_out[643] <= ~(layer0_out[12] | layer0_out[13]);
     layer1_out[644] <= ~(layer0_out[651] & layer0_out[652]);
     layer1_out[645] <= layer0_out[302] | layer0_out[303];
     layer1_out[646] <= layer0_out[284];
     layer1_out[647] <= ~layer0_out[1035];
     layer1_out[648] <= layer0_out[1247];
     layer1_out[649] <= layer0_out[969] & ~layer0_out[970];
     layer1_out[650] <= ~layer0_out[103];
     layer1_out[651] <= ~(layer0_out[815] & layer0_out[816]);
     layer1_out[652] <= ~layer0_out[1365];
     layer1_out[653] <= layer0_out[1456] & layer0_out[1457];
     layer1_out[654] <= layer0_out[1414] & ~layer0_out[1415];
     layer1_out[655] <= layer0_out[1380] | layer0_out[1381];
     layer1_out[656] <= 1'b0;
     layer1_out[657] <= layer0_out[979] & ~layer0_out[980];
     layer1_out[658] <= layer0_out[1433] & layer0_out[1434];
     layer1_out[659] <= layer0_out[698] & ~layer0_out[697];
     layer1_out[660] <= layer0_out[85];
     layer1_out[661] <= layer0_out[223];
     layer1_out[662] <= ~(layer0_out[883] & layer0_out[884]);
     layer1_out[663] <= 1'b1;
     layer1_out[664] <= ~layer0_out[727];
     layer1_out[665] <= ~layer0_out[34];
     layer1_out[666] <= layer0_out[1418] | layer0_out[1419];
     layer1_out[667] <= ~layer0_out[70] | layer0_out[69];
     layer1_out[668] <= ~layer0_out[273] | layer0_out[274];
     layer1_out[669] <= layer0_out[527] & layer0_out[528];
     layer1_out[670] <= 1'b1;
     layer1_out[671] <= ~(layer0_out[130] & layer0_out[131]);
     layer1_out[672] <= 1'b1;
     layer1_out[673] <= layer0_out[916] & ~layer0_out[915];
     layer1_out[674] <= layer0_out[249];
     layer1_out[675] <= layer0_out[897] & ~layer0_out[896];
     layer1_out[676] <= layer0_out[987] & ~layer0_out[986];
     layer1_out[677] <= layer0_out[1066] & layer0_out[1067];
     layer1_out[678] <= layer0_out[1174] & layer0_out[1175];
     layer1_out[679] <= ~layer0_out[1128] | layer0_out[1129];
     layer1_out[680] <= 1'b0;
     layer1_out[681] <= ~layer0_out[634];
     layer1_out[682] <= ~layer0_out[425] | layer0_out[424];
     layer1_out[683] <= ~layer0_out[403];
     layer1_out[684] <= layer0_out[1481];
     layer1_out[685] <= ~layer0_out[1024];
     layer1_out[686] <= 1'b1;
     layer1_out[687] <= layer0_out[295];
     layer1_out[688] <= layer0_out[320] ^ layer0_out[321];
     layer1_out[689] <= ~(layer0_out[608] | layer0_out[609]);
     layer1_out[690] <= layer0_out[1408] & ~layer0_out[1407];
     layer1_out[691] <= ~layer0_out[436];
     layer1_out[692] <= layer0_out[143];
     layer1_out[693] <= ~(layer0_out[1435] & layer0_out[1436]);
     layer1_out[694] <= ~layer0_out[1104];
     layer1_out[695] <= layer0_out[465] & ~layer0_out[466];
     layer1_out[696] <= layer0_out[609];
     layer1_out[697] <= layer0_out[385] & ~layer0_out[386];
     layer1_out[698] <= layer0_out[837];
     layer1_out[699] <= layer0_out[902] & ~layer0_out[903];
     layer1_out[700] <= ~layer0_out[1309];
     layer1_out[701] <= 1'b0;
     layer1_out[702] <= 1'b1;
     layer1_out[703] <= ~layer0_out[1379] | layer0_out[1380];
     layer1_out[704] <= 1'b1;
     layer1_out[705] <= layer0_out[27];
     layer1_out[706] <= layer0_out[199];
     layer1_out[707] <= layer0_out[1392];
     layer1_out[708] <= 1'b1;
     layer1_out[709] <= layer0_out[170] & ~layer0_out[169];
     layer1_out[710] <= layer0_out[1207] & ~layer0_out[1206];
     layer1_out[711] <= layer0_out[412];
     layer1_out[712] <= layer0_out[862];
     layer1_out[713] <= 1'b1;
     layer1_out[714] <= ~layer0_out[888] | layer0_out[887];
     layer1_out[715] <= 1'b0;
     layer1_out[716] <= layer0_out[853] | layer0_out[854];
     layer1_out[717] <= 1'b1;
     layer1_out[718] <= ~(layer0_out[77] & layer0_out[78]);
     layer1_out[719] <= layer0_out[1007] & layer0_out[1008];
     layer1_out[720] <= ~layer0_out[978];
     layer1_out[721] <= layer0_out[1028] & layer0_out[1029];
     layer1_out[722] <= layer0_out[684];
     layer1_out[723] <= ~layer0_out[147];
     layer1_out[724] <= layer0_out[436];
     layer1_out[725] <= ~(layer0_out[1179] ^ layer0_out[1180]);
     layer1_out[726] <= layer0_out[486] & ~layer0_out[487];
     layer1_out[727] <= ~layer0_out[215] | layer0_out[216];
     layer1_out[728] <= layer0_out[735] | layer0_out[736];
     layer1_out[729] <= 1'b0;
     layer1_out[730] <= layer0_out[1064];
     layer1_out[731] <= layer0_out[1216];
     layer1_out[732] <= layer0_out[1068] | layer0_out[1069];
     layer1_out[733] <= layer0_out[917] & layer0_out[918];
     layer1_out[734] <= ~(layer0_out[175] & layer0_out[176]);
     layer1_out[735] <= ~(layer0_out[713] | layer0_out[714]);
     layer1_out[736] <= 1'b1;
     layer1_out[737] <= 1'b1;
     layer1_out[738] <= ~(layer0_out[584] | layer0_out[585]);
     layer1_out[739] <= layer0_out[1058];
     layer1_out[740] <= ~(layer0_out[1006] & layer0_out[1007]);
     layer1_out[741] <= ~(layer0_out[1002] | layer0_out[1003]);
     layer1_out[742] <= ~(layer0_out[1167] & layer0_out[1168]);
     layer1_out[743] <= ~layer0_out[1303] | layer0_out[1304];
     layer1_out[744] <= layer0_out[427];
     layer1_out[745] <= layer0_out[602];
     layer1_out[746] <= layer0_out[312];
     layer1_out[747] <= layer0_out[1109];
     layer1_out[748] <= ~(layer0_out[25] | layer0_out[26]);
     layer1_out[749] <= ~(layer0_out[855] & layer0_out[856]);
     layer1_out[750] <= ~layer0_out[38];
     layer1_out[751] <= ~layer0_out[546];
     layer1_out[752] <= ~layer0_out[1102] | layer0_out[1103];
     layer1_out[753] <= layer0_out[723] & ~layer0_out[724];
     layer1_out[754] <= 1'b1;
     layer1_out[755] <= ~(layer0_out[1484] ^ layer0_out[1485]);
     layer1_out[756] <= layer0_out[620] & ~layer0_out[621];
     layer1_out[757] <= layer0_out[88];
     layer1_out[758] <= layer0_out[776] & ~layer0_out[775];
     layer1_out[759] <= layer0_out[1068] & ~layer0_out[1067];
     layer1_out[760] <= layer0_out[348];
     layer1_out[761] <= layer0_out[1251] | layer0_out[1252];
     layer1_out[762] <= ~(layer0_out[937] ^ layer0_out[938]);
     layer1_out[763] <= ~(layer0_out[1253] ^ layer0_out[1254]);
     layer1_out[764] <= ~layer0_out[1190] | layer0_out[1191];
     layer1_out[765] <= layer0_out[238] & layer0_out[239];
     layer1_out[766] <= ~layer0_out[1044] | layer0_out[1045];
     layer1_out[767] <= layer0_out[945] | layer0_out[946];
     layer1_out[768] <= layer0_out[134] & ~layer0_out[135];
     layer1_out[769] <= 1'b0;
     layer1_out[770] <= layer0_out[348];
     layer1_out[771] <= 1'b1;
     layer1_out[772] <= 1'b0;
     layer1_out[773] <= 1'b1;
     layer1_out[774] <= ~(layer0_out[5] | layer0_out[6]);
     layer1_out[775] <= layer0_out[213] & ~layer0_out[212];
     layer1_out[776] <= ~layer0_out[301] | layer0_out[302];
     layer1_out[777] <= layer0_out[1222];
     layer1_out[778] <= layer0_out[1447] ^ layer0_out[1448];
     layer1_out[779] <= layer0_out[1382];
     layer1_out[780] <= layer0_out[1270] & layer0_out[1271];
     layer1_out[781] <= 1'b0;
     layer1_out[782] <= ~layer0_out[165];
     layer1_out[783] <= 1'b0;
     layer1_out[784] <= 1'b0;
     layer1_out[785] <= layer0_out[636] | layer0_out[637];
     layer1_out[786] <= ~layer0_out[1141] | layer0_out[1142];
     layer1_out[787] <= layer0_out[1183] ^ layer0_out[1184];
     layer1_out[788] <= 1'b1;
     layer1_out[789] <= 1'b0;
     layer1_out[790] <= ~layer0_out[389];
     layer1_out[791] <= layer0_out[297];
     layer1_out[792] <= ~(layer0_out[778] | layer0_out[779]);
     layer1_out[793] <= 1'b0;
     layer1_out[794] <= layer0_out[845];
     layer1_out[795] <= ~layer0_out[1388] | layer0_out[1387];
     layer1_out[796] <= layer0_out[114] | layer0_out[115];
     layer1_out[797] <= 1'b1;
     layer1_out[798] <= layer0_out[960] & ~layer0_out[961];
     layer1_out[799] <= layer0_out[77] & ~layer0_out[76];
     layer1_out[800] <= 1'b1;
     layer1_out[801] <= layer0_out[1261] ^ layer0_out[1262];
     layer1_out[802] <= ~(layer0_out[874] | layer0_out[875]);
     layer1_out[803] <= ~(layer0_out[342] | layer0_out[343]);
     layer1_out[804] <= ~(layer0_out[1196] | layer0_out[1197]);
     layer1_out[805] <= 1'b1;
     layer1_out[806] <= layer0_out[1453];
     layer1_out[807] <= ~(layer0_out[407] & layer0_out[408]);
     layer1_out[808] <= ~layer0_out[3];
     layer1_out[809] <= ~(layer0_out[817] | layer0_out[818]);
     layer1_out[810] <= ~layer0_out[702] | layer0_out[703];
     layer1_out[811] <= ~(layer0_out[1486] | layer0_out[1487]);
     layer1_out[812] <= ~(layer0_out[1307] | layer0_out[1308]);
     layer1_out[813] <= ~layer0_out[1376];
     layer1_out[814] <= ~layer0_out[1108] | layer0_out[1107];
     layer1_out[815] <= ~layer0_out[1459];
     layer1_out[816] <= ~layer0_out[323];
     layer1_out[817] <= 1'b0;
     layer1_out[818] <= layer0_out[759] & ~layer0_out[758];
     layer1_out[819] <= 1'b1;
     layer1_out[820] <= ~layer0_out[1131] | layer0_out[1130];
     layer1_out[821] <= layer0_out[991] & ~layer0_out[990];
     layer1_out[822] <= layer0_out[1289] & ~layer0_out[1288];
     layer1_out[823] <= layer0_out[875] | layer0_out[876];
     layer1_out[824] <= layer0_out[398];
     layer1_out[825] <= layer0_out[414] & ~layer0_out[413];
     layer1_out[826] <= 1'b0;
     layer1_out[827] <= 1'b1;
     layer1_out[828] <= 1'b0;
     layer1_out[829] <= ~layer0_out[264];
     layer1_out[830] <= ~layer0_out[1044] | layer0_out[1043];
     layer1_out[831] <= 1'b1;
     layer1_out[832] <= ~(layer0_out[1279] & layer0_out[1280]);
     layer1_out[833] <= 1'b0;
     layer1_out[834] <= 1'b0;
     layer1_out[835] <= layer0_out[150];
     layer1_out[836] <= layer0_out[1094] & layer0_out[1095];
     layer1_out[837] <= layer0_out[8];
     layer1_out[838] <= layer0_out[1477] & layer0_out[1478];
     layer1_out[839] <= 1'b1;
     layer1_out[840] <= 1'b1;
     layer1_out[841] <= ~layer0_out[1413];
     layer1_out[842] <= ~layer0_out[1100] | layer0_out[1099];
     layer1_out[843] <= layer0_out[448];
     layer1_out[844] <= layer0_out[1119];
     layer1_out[845] <= ~layer0_out[421];
     layer1_out[846] <= layer0_out[559] | layer0_out[560];
     layer1_out[847] <= ~(layer0_out[251] & layer0_out[252]);
     layer1_out[848] <= ~(layer0_out[1272] | layer0_out[1273]);
     layer1_out[849] <= ~(layer0_out[1419] & layer0_out[1420]);
     layer1_out[850] <= layer0_out[755] & layer0_out[756];
     layer1_out[851] <= ~layer0_out[558] | layer0_out[557];
     layer1_out[852] <= 1'b1;
     layer1_out[853] <= 1'b0;
     layer1_out[854] <= ~layer0_out[371] | layer0_out[370];
     layer1_out[855] <= ~layer0_out[266];
     layer1_out[856] <= ~layer0_out[934] | layer0_out[933];
     layer1_out[857] <= layer0_out[460] | layer0_out[461];
     layer1_out[858] <= 1'b0;
     layer1_out[859] <= layer0_out[232] & ~layer0_out[233];
     layer1_out[860] <= ~layer0_out[1475];
     layer1_out[861] <= ~(layer0_out[208] | layer0_out[209]);
     layer1_out[862] <= ~layer0_out[1079] | layer0_out[1080];
     layer1_out[863] <= 1'b1;
     layer1_out[864] <= layer0_out[172];
     layer1_out[865] <= layer0_out[1165];
     layer1_out[866] <= layer0_out[1243] & layer0_out[1244];
     layer1_out[867] <= ~layer0_out[783];
     layer1_out[868] <= layer0_out[868] & ~layer0_out[869];
     layer1_out[869] <= ~(layer0_out[1320] & layer0_out[1321]);
     layer1_out[870] <= ~layer0_out[409] | layer0_out[410];
     layer1_out[871] <= ~(layer0_out[1397] ^ layer0_out[1398]);
     layer1_out[872] <= 1'b0;
     layer1_out[873] <= layer0_out[834] & layer0_out[835];
     layer1_out[874] <= ~(layer0_out[86] & layer0_out[87]);
     layer1_out[875] <= ~layer0_out[1065];
     layer1_out[876] <= ~layer0_out[420] | layer0_out[419];
     layer1_out[877] <= layer0_out[477];
     layer1_out[878] <= layer0_out[276];
     layer1_out[879] <= ~layer0_out[649] | layer0_out[650];
     layer1_out[880] <= 1'b1;
     layer1_out[881] <= 1'b1;
     layer1_out[882] <= ~layer0_out[651] | layer0_out[650];
     layer1_out[883] <= layer0_out[1160];
     layer1_out[884] <= ~(layer0_out[1286] | layer0_out[1287]);
     layer1_out[885] <= 1'b0;
     layer1_out[886] <= layer0_out[332] | layer0_out[333];
     layer1_out[887] <= 1'b0;
     layer1_out[888] <= layer0_out[1189] & ~layer0_out[1190];
     layer1_out[889] <= layer0_out[919] & ~layer0_out[918];
     layer1_out[890] <= ~(layer0_out[634] & layer0_out[635]);
     layer1_out[891] <= layer0_out[744];
     layer1_out[892] <= ~layer0_out[1417];
     layer1_out[893] <= layer0_out[363] | layer0_out[364];
     layer1_out[894] <= layer0_out[353];
     layer1_out[895] <= ~(layer0_out[643] & layer0_out[644]);
     layer1_out[896] <= ~layer0_out[645] | layer0_out[644];
     layer1_out[897] <= layer0_out[402];
     layer1_out[898] <= layer0_out[573];
     layer1_out[899] <= layer0_out[487] & layer0_out[488];
     layer1_out[900] <= layer0_out[1439] & ~layer0_out[1438];
     layer1_out[901] <= 1'b0;
     layer1_out[902] <= layer0_out[1015] | layer0_out[1016];
     layer1_out[903] <= ~(layer0_out[1159] | layer0_out[1160]);
     layer1_out[904] <= layer0_out[793] & ~layer0_out[794];
     layer1_out[905] <= 1'b0;
     layer1_out[906] <= 1'b1;
     layer1_out[907] <= ~(layer0_out[598] & layer0_out[599]);
     layer1_out[908] <= 1'b0;
     layer1_out[909] <= layer0_out[1178] | layer0_out[1179];
     layer1_out[910] <= ~layer0_out[462];
     layer1_out[911] <= layer0_out[991];
     layer1_out[912] <= layer0_out[214];
     layer1_out[913] <= layer0_out[632];
     layer1_out[914] <= layer0_out[1153];
     layer1_out[915] <= ~layer0_out[1150];
     layer1_out[916] <= 1'b0;
     layer1_out[917] <= layer0_out[712] & ~layer0_out[711];
     layer1_out[918] <= 1'b1;
     layer1_out[919] <= layer0_out[920] & ~layer0_out[919];
     layer1_out[920] <= ~layer0_out[1457];
     layer1_out[921] <= 1'b0;
     layer1_out[922] <= 1'b1;
     layer1_out[923] <= 1'b0;
     layer1_out[924] <= ~layer0_out[464];
     layer1_out[925] <= layer0_out[201];
     layer1_out[926] <= layer0_out[560] & ~layer0_out[561];
     layer1_out[927] <= ~layer0_out[353] | layer0_out[354];
     layer1_out[928] <= ~layer0_out[556];
     layer1_out[929] <= layer0_out[163] & ~layer0_out[164];
     layer1_out[930] <= 1'b1;
     layer1_out[931] <= ~layer0_out[951];
     layer1_out[932] <= ~(layer0_out[955] | layer0_out[956]);
     layer1_out[933] <= layer0_out[998];
     layer1_out[934] <= layer0_out[904];
     layer1_out[935] <= ~layer0_out[1494] | layer0_out[1493];
     layer1_out[936] <= 1'b1;
     layer1_out[937] <= layer0_out[265] & layer0_out[266];
     layer1_out[938] <= 1'b0;
     layer1_out[939] <= ~layer0_out[1411];
     layer1_out[940] <= ~(layer0_out[1285] & layer0_out[1286]);
     layer1_out[941] <= layer0_out[1450] | layer0_out[1451];
     layer1_out[942] <= ~layer0_out[1088] | layer0_out[1087];
     layer1_out[943] <= ~layer0_out[1003];
     layer1_out[944] <= ~(layer0_out[524] | layer0_out[525]);
     layer1_out[945] <= ~layer0_out[523];
     layer1_out[946] <= layer0_out[849] & ~layer0_out[848];
     layer1_out[947] <= ~layer0_out[400] | layer0_out[401];
     layer1_out[948] <= 1'b1;
     layer1_out[949] <= ~(layer0_out[816] | layer0_out[817]);
     layer1_out[950] <= 1'b0;
     layer1_out[951] <= ~(layer0_out[683] & layer0_out[684]);
     layer1_out[952] <= 1'b0;
     layer1_out[953] <= ~(layer0_out[1432] | layer0_out[1433]);
     layer1_out[954] <= layer0_out[33] & layer0_out[34];
     layer1_out[955] <= ~(layer0_out[1257] & layer0_out[1258]);
     layer1_out[956] <= ~layer0_out[987] | layer0_out[988];
     layer1_out[957] <= ~(layer0_out[532] & layer0_out[533]);
     layer1_out[958] <= ~(layer0_out[1420] | layer0_out[1421]);
     layer1_out[959] <= 1'b0;
     layer1_out[960] <= ~layer0_out[843] | layer0_out[844];
     layer1_out[961] <= ~layer0_out[1161];
     layer1_out[962] <= ~layer0_out[1022] | layer0_out[1023];
     layer1_out[963] <= layer0_out[1230] | layer0_out[1231];
     layer1_out[964] <= layer0_out[799];
     layer1_out[965] <= 1'b0;
     layer1_out[966] <= ~(layer0_out[38] | layer0_out[39]);
     layer1_out[967] <= ~(layer0_out[1248] | layer0_out[1249]);
     layer1_out[968] <= 1'b0;
     layer1_out[969] <= layer0_out[1273] & ~layer0_out[1274];
     layer1_out[970] <= layer0_out[556] ^ layer0_out[557];
     layer1_out[971] <= ~(layer0_out[587] | layer0_out[588]);
     layer1_out[972] <= 1'b0;
     layer1_out[973] <= layer0_out[846] | layer0_out[847];
     layer1_out[974] <= ~layer0_out[807];
     layer1_out[975] <= ~(layer0_out[905] & layer0_out[906]);
     layer1_out[976] <= 1'b0;
     layer1_out[977] <= 1'b1;
     layer1_out[978] <= layer0_out[236] | layer0_out[237];
     layer1_out[979] <= ~layer0_out[1112];
     layer1_out[980] <= ~(layer0_out[493] | layer0_out[494]);
     layer1_out[981] <= ~(layer0_out[597] | layer0_out[598]);
     layer1_out[982] <= ~layer0_out[387];
     layer1_out[983] <= layer0_out[925] ^ layer0_out[926];
     layer1_out[984] <= ~layer0_out[431] | layer0_out[430];
     layer1_out[985] <= ~(layer0_out[577] | layer0_out[578]);
     layer1_out[986] <= layer0_out[952];
     layer1_out[987] <= ~layer0_out[13] | layer0_out[14];
     layer1_out[988] <= 1'b1;
     layer1_out[989] <= 1'b1;
     layer1_out[990] <= ~(layer0_out[1252] & layer0_out[1253]);
     layer1_out[991] <= layer0_out[217];
     layer1_out[992] <= layer0_out[946] ^ layer0_out[947];
     layer1_out[993] <= layer0_out[20] & layer0_out[21];
     layer1_out[994] <= layer0_out[1047] & ~layer0_out[1046];
     layer1_out[995] <= layer0_out[1187] | layer0_out[1188];
     layer1_out[996] <= 1'b0;
     layer1_out[997] <= 1'b1;
     layer1_out[998] <= 1'b1;
     layer1_out[999] <= ~layer0_out[748] | layer0_out[747];
     layer1_out[1000] <= ~(layer0_out[1100] | layer0_out[1101]);
     layer1_out[1001] <= ~(layer0_out[392] & layer0_out[393]);
     layer1_out[1002] <= layer0_out[510] & ~layer0_out[511];
     layer1_out[1003] <= 1'b1;
     layer1_out[1004] <= layer0_out[248] & layer0_out[249];
     layer1_out[1005] <= ~layer0_out[137];
     layer1_out[1006] <= 1'b1;
     layer1_out[1007] <= ~(layer0_out[789] & layer0_out[790]);
     layer1_out[1008] <= layer0_out[316] & ~layer0_out[317];
     layer1_out[1009] <= ~layer0_out[1268] | layer0_out[1267];
     layer1_out[1010] <= layer0_out[469] & layer0_out[470];
     layer1_out[1011] <= ~layer0_out[452] | layer0_out[453];
     layer1_out[1012] <= layer0_out[185];
     layer1_out[1013] <= ~layer0_out[585];
     layer1_out[1014] <= 1'b1;
     layer1_out[1015] <= ~(layer0_out[928] & layer0_out[929]);
     layer1_out[1016] <= 1'b0;
     layer1_out[1017] <= 1'b0;
     layer1_out[1018] <= layer0_out[1308] & ~layer0_out[1309];
     layer1_out[1019] <= layer0_out[1159];
     layer1_out[1020] <= layer0_out[589] | layer0_out[590];
     layer1_out[1021] <= ~layer0_out[251] | layer0_out[250];
     layer1_out[1022] <= 1'b1;
     layer1_out[1023] <= layer0_out[1325];
     layer1_out[1024] <= ~layer0_out[706] | layer0_out[707];
     layer1_out[1025] <= 1'b0;
     layer1_out[1026] <= layer0_out[931] & ~layer0_out[930];
     layer1_out[1027] <= ~(layer0_out[491] | layer0_out[492]);
     layer1_out[1028] <= ~layer0_out[144] | layer0_out[145];
     layer1_out[1029] <= layer0_out[812] | layer0_out[813];
     layer1_out[1030] <= ~layer0_out[1465];
     layer1_out[1031] <= layer0_out[1478] | layer0_out[1479];
     layer1_out[1032] <= layer0_out[1208] & ~layer0_out[1207];
     layer1_out[1033] <= layer0_out[520];
     layer1_out[1034] <= layer0_out[282];
     layer1_out[1035] <= layer0_out[1277];
     layer1_out[1036] <= 1'b1;
     layer1_out[1037] <= 1'b0;
     layer1_out[1038] <= 1'b0;
     layer1_out[1039] <= ~layer0_out[923] | layer0_out[922];
     layer1_out[1040] <= layer0_out[1098] | layer0_out[1099];
     layer1_out[1041] <= ~layer0_out[1332] | layer0_out[1331];
     layer1_out[1042] <= ~(layer0_out[1182] | layer0_out[1183]);
     layer1_out[1043] <= ~layer0_out[1346];
     layer1_out[1044] <= layer0_out[1344] & ~layer0_out[1343];
     layer1_out[1045] <= layer0_out[1262] | layer0_out[1263];
     layer1_out[1046] <= 1'b1;
     layer1_out[1047] <= layer0_out[378] & ~layer0_out[379];
     layer1_out[1048] <= layer0_out[942];
     layer1_out[1049] <= ~layer0_out[1441];
     layer1_out[1050] <= 1'b1;
     layer1_out[1051] <= 1'b0;
     layer1_out[1052] <= ~(layer0_out[1171] | layer0_out[1172]);
     layer1_out[1053] <= layer0_out[368];
     layer1_out[1054] <= 1'b0;
     layer1_out[1055] <= layer0_out[216] ^ layer0_out[217];
     layer1_out[1056] <= layer0_out[168] | layer0_out[169];
     layer1_out[1057] <= ~layer0_out[1321];
     layer1_out[1058] <= ~layer0_out[380];
     layer1_out[1059] <= 1'b1;
     layer1_out[1060] <= layer0_out[95] | layer0_out[96];
     layer1_out[1061] <= layer0_out[1001] & ~layer0_out[1002];
     layer1_out[1062] <= ~(layer0_out[398] & layer0_out[399]);
     layer1_out[1063] <= layer0_out[700] & layer0_out[701];
     layer1_out[1064] <= layer0_out[1197] | layer0_out[1198];
     layer1_out[1065] <= 1'b1;
     layer1_out[1066] <= layer0_out[625] | layer0_out[626];
     layer1_out[1067] <= layer0_out[220] | layer0_out[221];
     layer1_out[1068] <= layer0_out[186] & layer0_out[187];
     layer1_out[1069] <= 1'b0;
     layer1_out[1070] <= ~layer0_out[372] | layer0_out[371];
     layer1_out[1071] <= ~layer0_out[1422] | layer0_out[1423];
     layer1_out[1072] <= layer0_out[1400] & ~layer0_out[1401];
     layer1_out[1073] <= layer0_out[422] & ~layer0_out[423];
     layer1_out[1074] <= ~layer0_out[1140] | layer0_out[1141];
     layer1_out[1075] <= 1'b0;
     layer1_out[1076] <= layer0_out[911] & ~layer0_out[912];
     layer1_out[1077] <= 1'b0;
     layer1_out[1078] <= layer0_out[1052] & ~layer0_out[1051];
     layer1_out[1079] <= ~(layer0_out[234] & layer0_out[235]);
     layer1_out[1080] <= 1'b1;
     layer1_out[1081] <= 1'b1;
     layer1_out[1082] <= ~layer0_out[63] | layer0_out[62];
     layer1_out[1083] <= ~layer0_out[1358];
     layer1_out[1084] <= ~layer0_out[1374] | layer0_out[1375];
     layer1_out[1085] <= ~layer0_out[31] | layer0_out[30];
     layer1_out[1086] <= ~(layer0_out[1106] | layer0_out[1107]);
     layer1_out[1087] <= layer0_out[802];
     layer1_out[1088] <= layer0_out[935] | layer0_out[936];
     layer1_out[1089] <= 1'b1;
     layer1_out[1090] <= ~(layer0_out[66] & layer0_out[67]);
     layer1_out[1091] <= ~(layer0_out[36] | layer0_out[37]);
     layer1_out[1092] <= layer0_out[1156] & ~layer0_out[1155];
     layer1_out[1093] <= 1'b1;
     layer1_out[1094] <= 1'b0;
     layer1_out[1095] <= layer0_out[41] & ~layer0_out[42];
     layer1_out[1096] <= 1'b1;
     layer1_out[1097] <= layer0_out[908];
     layer1_out[1098] <= ~layer0_out[877] | layer0_out[876];
     layer1_out[1099] <= layer0_out[1480] | layer0_out[1481];
     layer1_out[1100] <= ~(layer0_out[891] & layer0_out[892]);
     layer1_out[1101] <= layer0_out[1425] & layer0_out[1426];
     layer1_out[1102] <= 1'b1;
     layer1_out[1103] <= layer0_out[825] & layer0_out[826];
     layer1_out[1104] <= 1'b1;
     layer1_out[1105] <= ~layer0_out[242] | layer0_out[241];
     layer1_out[1106] <= 1'b1;
     layer1_out[1107] <= ~layer0_out[125];
     layer1_out[1108] <= ~layer0_out[926] | layer0_out[927];
     layer1_out[1109] <= layer0_out[1497] & layer0_out[1498];
     layer1_out[1110] <= layer0_out[1137];
     layer1_out[1111] <= layer0_out[432];
     layer1_out[1112] <= ~layer0_out[802];
     layer1_out[1113] <= layer0_out[1323];
     layer1_out[1114] <= 1'b1;
     layer1_out[1115] <= ~layer0_out[760] | layer0_out[759];
     layer1_out[1116] <= layer0_out[1352] & layer0_out[1353];
     layer1_out[1117] <= 1'b1;
     layer1_out[1118] <= ~layer0_out[677] | layer0_out[676];
     layer1_out[1119] <= 1'b0;
     layer1_out[1120] <= layer0_out[344] & layer0_out[345];
     layer1_out[1121] <= layer0_out[72] | layer0_out[73];
     layer1_out[1122] <= ~(layer0_out[434] & layer0_out[435]);
     layer1_out[1123] <= layer0_out[395];
     layer1_out[1124] <= ~(layer0_out[962] & layer0_out[963]);
     layer1_out[1125] <= 1'b0;
     layer1_out[1126] <= ~(layer0_out[499] & layer0_out[500]);
     layer1_out[1127] <= layer0_out[722] & layer0_out[723];
     layer1_out[1128] <= 1'b0;
     layer1_out[1129] <= 1'b0;
     layer1_out[1130] <= ~(layer0_out[1061] & layer0_out[1062]);
     layer1_out[1131] <= layer0_out[63] & ~layer0_out[64];
     layer1_out[1132] <= layer0_out[734] & ~layer0_out[733];
     layer1_out[1133] <= ~layer0_out[1236];
     layer1_out[1134] <= layer0_out[198] & ~layer0_out[197];
     layer1_out[1135] <= 1'b1;
     layer1_out[1136] <= ~(layer0_out[974] & layer0_out[975]);
     layer1_out[1137] <= ~layer0_out[610] | layer0_out[611];
     layer1_out[1138] <= 1'b0;
     layer1_out[1139] <= 1'b0;
     layer1_out[1140] <= 1'b1;
     layer1_out[1141] <= layer0_out[262] ^ layer0_out[263];
     layer1_out[1142] <= ~(layer0_out[749] | layer0_out[750]);
     layer1_out[1143] <= ~layer0_out[1117];
     layer1_out[1144] <= ~(layer0_out[885] | layer0_out[886]);
     layer1_out[1145] <= ~(layer0_out[600] & layer0_out[601]);
     layer1_out[1146] <= 1'b0;
     layer1_out[1147] <= 1'b0;
     layer1_out[1148] <= layer0_out[286];
     layer1_out[1149] <= ~(layer0_out[1260] | layer0_out[1261]);
     layer1_out[1150] <= 1'b0;
     layer1_out[1151] <= ~layer0_out[878];
     layer1_out[1152] <= 1'b1;
     layer1_out[1153] <= ~layer0_out[382] | layer0_out[383];
     layer1_out[1154] <= 1'b0;
     layer1_out[1155] <= layer0_out[593] & ~layer0_out[594];
     layer1_out[1156] <= layer0_out[315] & ~layer0_out[314];
     layer1_out[1157] <= ~(layer0_out[844] ^ layer0_out[845]);
     layer1_out[1158] <= layer0_out[376] & ~layer0_out[377];
     layer1_out[1159] <= 1'b0;
     layer1_out[1160] <= 1'b1;
     layer1_out[1161] <= layer0_out[703] & ~layer0_out[704];
     layer1_out[1162] <= ~layer0_out[948] | layer0_out[949];
     layer1_out[1163] <= ~layer0_out[1409];
     layer1_out[1164] <= ~(layer0_out[107] | layer0_out[108]);
     layer1_out[1165] <= ~layer0_out[706];
     layer1_out[1166] <= ~layer0_out[881] | layer0_out[882];
     layer1_out[1167] <= ~(layer0_out[463] & layer0_out[464]);
     layer1_out[1168] <= 1'b1;
     layer1_out[1169] <= layer0_out[835];
     layer1_out[1170] <= ~(layer0_out[1205] | layer0_out[1206]);
     layer1_out[1171] <= 1'b0;
     layer1_out[1172] <= layer0_out[1463] | layer0_out[1464];
     layer1_out[1173] <= layer0_out[641] & layer0_out[642];
     layer1_out[1174] <= 1'b1;
     layer1_out[1175] <= 1'b0;
     layer1_out[1176] <= ~layer0_out[701] | layer0_out[702];
     layer1_out[1177] <= ~layer0_out[967] | layer0_out[968];
     layer1_out[1178] <= layer0_out[1327] & ~layer0_out[1328];
     layer1_out[1179] <= layer0_out[636];
     layer1_out[1180] <= layer0_out[1497];
     layer1_out[1181] <= 1'b0;
     layer1_out[1182] <= 1'b0;
     layer1_out[1183] <= layer0_out[448] & layer0_out[449];
     layer1_out[1184] <= ~layer0_out[1313];
     layer1_out[1185] <= layer0_out[1223] & layer0_out[1224];
     layer1_out[1186] <= ~(layer0_out[1413] | layer0_out[1414]);
     layer1_out[1187] <= layer0_out[1035] & ~layer0_out[1036];
     layer1_out[1188] <= layer0_out[787] & ~layer0_out[786];
     layer1_out[1189] <= ~layer0_out[325] | layer0_out[326];
     layer1_out[1190] <= 1'b0;
     layer1_out[1191] <= 1'b1;
     layer1_out[1192] <= ~(layer0_out[907] | layer0_out[908]);
     layer1_out[1193] <= ~(layer0_out[776] | layer0_out[777]);
     layer1_out[1194] <= ~(layer0_out[1163] | layer0_out[1164]);
     layer1_out[1195] <= layer0_out[359] | layer0_out[360];
     layer1_out[1196] <= ~layer0_out[814];
     layer1_out[1197] <= layer0_out[1298] & ~layer0_out[1297];
     layer1_out[1198] <= layer0_out[1059];
     layer1_out[1199] <= ~(layer0_out[561] & layer0_out[562]);
     layer1_out[1200] <= layer0_out[313] & layer0_out[314];
     layer1_out[1201] <= ~layer0_out[1052] | layer0_out[1053];
     layer1_out[1202] <= 1'b0;
     layer1_out[1203] <= ~layer0_out[890];
     layer1_out[1204] <= layer0_out[666] & ~layer0_out[667];
     layer1_out[1205] <= 1'b0;
     layer1_out[1206] <= layer0_out[501] & ~layer0_out[500];
     layer1_out[1207] <= ~layer0_out[748] | layer0_out[749];
     layer1_out[1208] <= ~layer0_out[372];
     layer1_out[1209] <= layer0_out[60] & ~layer0_out[61];
     layer1_out[1210] <= ~layer0_out[1403];
     layer1_out[1211] <= ~layer0_out[289];
     layer1_out[1212] <= 1'b0;
     layer1_out[1213] <= layer0_out[1140];
     layer1_out[1214] <= 1'b1;
     layer1_out[1215] <= 1'b1;
     layer1_out[1216] <= layer0_out[536] | layer0_out[537];
     layer1_out[1217] <= ~layer0_out[752] | layer0_out[751];
     layer1_out[1218] <= 1'b1;
     layer1_out[1219] <= layer0_out[837];
     layer1_out[1220] <= layer0_out[183] | layer0_out[184];
     layer1_out[1221] <= layer0_out[1228];
     layer1_out[1222] <= ~layer0_out[40] | layer0_out[39];
     layer1_out[1223] <= ~layer0_out[1046];
     layer1_out[1224] <= layer0_out[1127];
     layer1_out[1225] <= layer0_out[914] & ~layer0_out[913];
     layer1_out[1226] <= layer0_out[1180] | layer0_out[1181];
     layer1_out[1227] <= ~layer0_out[940] | layer0_out[939];
     layer1_out[1228] <= layer0_out[111] | layer0_out[112];
     layer1_out[1229] <= ~layer0_out[783];
     layer1_out[1230] <= ~layer0_out[1483] | layer0_out[1482];
     layer1_out[1231] <= 1'b0;
     layer1_out[1232] <= 1'b1;
     layer1_out[1233] <= 1'b0;
     layer1_out[1234] <= ~(layer0_out[341] | layer0_out[342]);
     layer1_out[1235] <= 1'b0;
     layer1_out[1236] <= ~layer0_out[336];
     layer1_out[1237] <= layer0_out[897] | layer0_out[898];
     layer1_out[1238] <= ~(layer0_out[1296] | layer0_out[1297]);
     layer1_out[1239] <= 1'b1;
     layer1_out[1240] <= layer0_out[490] & ~layer0_out[491];
     layer1_out[1241] <= ~layer0_out[1025] | layer0_out[1024];
     layer1_out[1242] <= 1'b0;
     layer1_out[1243] <= ~layer0_out[93];
     layer1_out[1244] <= layer0_out[1401];
     layer1_out[1245] <= ~layer0_out[944] | layer0_out[945];
     layer1_out[1246] <= layer0_out[660];
     layer1_out[1247] <= layer0_out[1329] & ~layer0_out[1328];
     layer1_out[1248] <= layer0_out[79] & ~layer0_out[78];
     layer1_out[1249] <= ~layer0_out[1265];
     layer1_out[1250] <= 1'b1;
     layer1_out[1251] <= layer0_out[574] & ~layer0_out[575];
     layer1_out[1252] <= 1'b1;
     layer1_out[1253] <= layer0_out[1145];
     layer1_out[1254] <= ~layer0_out[230];
     layer1_out[1255] <= ~layer0_out[691] | layer0_out[692];
     layer1_out[1256] <= ~(layer0_out[1271] ^ layer0_out[1272]);
     layer1_out[1257] <= 1'b0;
     layer1_out[1258] <= ~(layer0_out[259] | layer0_out[260]);
     layer1_out[1259] <= ~(layer0_out[675] & layer0_out[676]);
     layer1_out[1260] <= ~(layer0_out[603] | layer0_out[604]);
     layer1_out[1261] <= layer0_out[509] & ~layer0_out[508];
     layer1_out[1262] <= layer0_out[1466];
     layer1_out[1263] <= layer0_out[637];
     layer1_out[1264] <= 1'b0;
     layer1_out[1265] <= layer0_out[128] & ~layer0_out[127];
     layer1_out[1266] <= 1'b0;
     layer1_out[1267] <= 1'b0;
     layer1_out[1268] <= 1'b1;
     layer1_out[1269] <= 1'b0;
     layer1_out[1270] <= ~(layer0_out[1075] | layer0_out[1076]);
     layer1_out[1271] <= 1'b0;
     layer1_out[1272] <= ~layer0_out[393] | layer0_out[394];
     layer1_out[1273] <= layer0_out[48];
     layer1_out[1274] <= ~layer0_out[1354];
     layer1_out[1275] <= layer0_out[1488] | layer0_out[1489];
     layer1_out[1276] <= ~layer0_out[902];
     layer1_out[1277] <= ~(layer0_out[1439] & layer0_out[1440]);
     layer1_out[1278] <= ~layer0_out[1255] | layer0_out[1256];
     layer1_out[1279] <= layer0_out[1492];
     layer1_out[1280] <= layer0_out[129];
     layer1_out[1281] <= ~layer0_out[414];
     layer1_out[1282] <= ~layer0_out[694] | layer0_out[695];
     layer1_out[1283] <= layer0_out[17];
     layer1_out[1284] <= layer0_out[1060] & ~layer0_out[1061];
     layer1_out[1285] <= layer0_out[1027] | layer0_out[1028];
     layer1_out[1286] <= ~(layer0_out[307] & layer0_out[308]);
     layer1_out[1287] <= 1'b0;
     layer1_out[1288] <= ~(layer0_out[1014] | layer0_out[1015]);
     layer1_out[1289] <= 1'b1;
     layer1_out[1290] <= ~layer0_out[357];
     layer1_out[1291] <= 1'b0;
     layer1_out[1292] <= ~layer0_out[1122];
     layer1_out[1293] <= layer0_out[1199];
     layer1_out[1294] <= ~(layer0_out[764] | layer0_out[765]);
     layer1_out[1295] <= ~layer0_out[84] | layer0_out[83];
     layer1_out[1296] <= 1'b1;
     layer1_out[1297] <= layer0_out[842];
     layer1_out[1298] <= layer0_out[222];
     layer1_out[1299] <= ~layer0_out[1079];
     layer1_out[1300] <= layer0_out[367] & ~layer0_out[366];
     layer1_out[1301] <= ~layer0_out[622] | layer0_out[623];
     layer1_out[1302] <= layer0_out[504] & ~layer0_out[505];
     layer1_out[1303] <= ~(layer0_out[888] ^ layer0_out[889]);
     layer1_out[1304] <= 1'b1;
     layer1_out[1305] <= layer0_out[810] & ~layer0_out[811];
     layer1_out[1306] <= 1'b1;
     layer1_out[1307] <= layer0_out[884];
     layer1_out[1308] <= layer0_out[791] & ~layer0_out[792];
     layer1_out[1309] <= ~(layer0_out[1080] & layer0_out[1081]);
     layer1_out[1310] <= layer0_out[319] & ~layer0_out[320];
     layer1_out[1311] <= layer0_out[1051];
     layer1_out[1312] <= layer0_out[150] & ~layer0_out[151];
     layer1_out[1313] <= 1'b0;
     layer1_out[1314] <= layer0_out[1083] & layer0_out[1084];
     layer1_out[1315] <= layer0_out[722] & ~layer0_out[721];
     layer1_out[1316] <= 1'b0;
     layer1_out[1317] <= ~layer0_out[1470] | layer0_out[1469];
     layer1_out[1318] <= layer0_out[1234] & ~layer0_out[1233];
     layer1_out[1319] <= ~(layer0_out[497] | layer0_out[498]);
     layer1_out[1320] <= 1'b0;
     layer1_out[1321] <= layer0_out[1049];
     layer1_out[1322] <= 1'b1;
     layer1_out[1323] <= layer0_out[122] & layer0_out[123];
     layer1_out[1324] <= 1'b1;
     layer1_out[1325] <= 1'b0;
     layer1_out[1326] <= ~layer0_out[326];
     layer1_out[1327] <= 1'b1;
     layer1_out[1328] <= layer0_out[116];
     layer1_out[1329] <= layer0_out[535] & layer0_out[536];
     layer1_out[1330] <= layer0_out[983];
     layer1_out[1331] <= 1'b1;
     layer1_out[1332] <= layer0_out[1097] & ~layer0_out[1098];
     layer1_out[1333] <= 1'b0;
     layer1_out[1334] <= layer0_out[343] & layer0_out[344];
     layer1_out[1335] <= ~layer0_out[732];
     layer1_out[1336] <= ~(layer0_out[1304] | layer0_out[1305]);
     layer1_out[1337] <= 1'b0;
     layer1_out[1338] <= layer0_out[916] & layer0_out[917];
     layer1_out[1339] <= layer0_out[745] & layer0_out[746];
     layer1_out[1340] <= layer0_out[122] & ~layer0_out[121];
     layer1_out[1341] <= layer0_out[688] | layer0_out[689];
     layer1_out[1342] <= 1'b0;
     layer1_out[1343] <= layer0_out[564] & ~layer0_out[565];
     layer1_out[1344] <= layer0_out[630] | layer0_out[631];
     layer1_out[1345] <= ~layer0_out[652];
     layer1_out[1346] <= layer0_out[887];
     layer1_out[1347] <= ~(layer0_out[1357] | layer0_out[1358]);
     layer1_out[1348] <= ~layer0_out[517];
     layer1_out[1349] <= layer0_out[822] & ~layer0_out[821];
     layer1_out[1350] <= ~(layer0_out[196] | layer0_out[197]);
     layer1_out[1351] <= 1'b1;
     layer1_out[1352] <= 1'b0;
     layer1_out[1353] <= ~(layer0_out[932] ^ layer0_out[933]);
     layer1_out[1354] <= ~layer0_out[190];
     layer1_out[1355] <= layer0_out[246] & ~layer0_out[247];
     layer1_out[1356] <= layer0_out[11];
     layer1_out[1357] <= ~layer0_out[1443];
     layer1_out[1358] <= 1'b1;
     layer1_out[1359] <= ~layer0_out[1038];
     layer1_out[1360] <= layer0_out[9] & layer0_out[10];
     layer1_out[1361] <= ~layer0_out[579];
     layer1_out[1362] <= 1'b0;
     layer1_out[1363] <= 1'b1;
     layer1_out[1364] <= ~layer0_out[364] | layer0_out[365];
     layer1_out[1365] <= layer0_out[192] | layer0_out[193];
     layer1_out[1366] <= layer0_out[1323];
     layer1_out[1367] <= layer0_out[117];
     layer1_out[1368] <= layer0_out[1135] | layer0_out[1136];
     layer1_out[1369] <= 1'b0;
     layer1_out[1370] <= ~layer0_out[361] | layer0_out[360];
     layer1_out[1371] <= 1'b0;
     layer1_out[1372] <= layer0_out[481] | layer0_out[482];
     layer1_out[1373] <= ~layer0_out[527] | layer0_out[526];
     layer1_out[1374] <= 1'b1;
     layer1_out[1375] <= ~(layer0_out[1405] & layer0_out[1406]);
     layer1_out[1376] <= ~layer0_out[220] | layer0_out[219];
     layer1_out[1377] <= layer0_out[989] & ~layer0_out[988];
     layer1_out[1378] <= 1'b1;
     layer1_out[1379] <= 1'b0;
     layer1_out[1380] <= ~(layer0_out[1423] | layer0_out[1424]);
     layer1_out[1381] <= ~(layer0_out[210] ^ layer0_out[211]);
     layer1_out[1382] <= 1'b1;
     layer1_out[1383] <= layer0_out[447];
     layer1_out[1384] <= ~layer0_out[821];
     layer1_out[1385] <= layer0_out[892] | layer0_out[893];
     layer1_out[1386] <= ~layer0_out[785] | layer0_out[786];
     layer1_out[1387] <= layer0_out[402] | layer0_out[403];
     layer1_out[1388] <= 1'b0;
     layer1_out[1389] <= layer0_out[235] | layer0_out[236];
     layer1_out[1390] <= ~layer0_out[705] | layer0_out[704];
     layer1_out[1391] <= ~(layer0_out[455] | layer0_out[456]);
     layer1_out[1392] <= ~(layer0_out[787] & layer0_out[788]);
     layer1_out[1393] <= layer0_out[470] & layer0_out[471];
     layer1_out[1394] <= layer0_out[1249] | layer0_out[1250];
     layer1_out[1395] <= layer0_out[552] & ~layer0_out[551];
     layer1_out[1396] <= ~layer0_out[864];
     layer1_out[1397] <= ~(layer0_out[586] & layer0_out[587]);
     layer1_out[1398] <= layer0_out[1283] & ~layer0_out[1284];
     layer1_out[1399] <= ~(layer0_out[1055] ^ layer0_out[1056]);
     layer1_out[1400] <= ~(layer0_out[427] | layer0_out[428]);
     layer1_out[1401] <= ~(layer0_out[1143] & layer0_out[1144]);
     layer1_out[1402] <= layer0_out[313] & ~layer0_out[312];
     layer1_out[1403] <= layer0_out[1222];
     layer1_out[1404] <= layer0_out[441];
     layer1_out[1405] <= ~(layer0_out[780] & layer0_out[781]);
     layer1_out[1406] <= 1'b1;
     layer1_out[1407] <= 1'b1;
     layer1_out[1408] <= ~layer0_out[1040] | layer0_out[1041];
     layer1_out[1409] <= layer0_out[324] & ~layer0_out[325];
     layer1_out[1410] <= 1'b0;
     layer1_out[1411] <= ~(layer0_out[243] | layer0_out[244]);
     layer1_out[1412] <= 1'b1;
     layer1_out[1413] <= 1'b1;
     layer1_out[1414] <= layer0_out[256] & layer0_out[257];
     layer1_out[1415] <= ~layer0_out[800] | layer0_out[799];
     layer1_out[1416] <= layer0_out[829] & ~layer0_out[830];
     layer1_out[1417] <= layer0_out[259];
     layer1_out[1418] <= layer0_out[1011];
     layer1_out[1419] <= ~(layer0_out[1090] | layer0_out[1091]);
     layer1_out[1420] <= layer0_out[438];
     layer1_out[1421] <= layer0_out[157];
     layer1_out[1422] <= 1'b1;
     layer1_out[1423] <= 1'b0;
     layer1_out[1424] <= 1'b1;
     layer1_out[1425] <= ~layer0_out[31] | layer0_out[32];
     layer1_out[1426] <= 1'b0;
     layer1_out[1427] <= ~layer0_out[154] | layer0_out[155];
     layer1_out[1428] <= 1'b0;
     layer1_out[1429] <= layer0_out[1202] & ~layer0_out[1203];
     layer1_out[1430] <= 1'b0;
     layer1_out[1431] <= layer0_out[1240] & ~layer0_out[1241];
     layer1_out[1432] <= layer0_out[1449] & ~layer0_out[1448];
     layer1_out[1433] <= 1'b0;
     layer1_out[1434] <= layer0_out[1395];
     layer1_out[1435] <= 1'b0;
     layer1_out[1436] <= 1'b0;
     layer1_out[1437] <= ~layer0_out[0] | layer0_out[2];
     layer1_out[1438] <= ~(layer0_out[803] ^ layer0_out[804]);
     layer1_out[1439] <= 1'b0;
     layer1_out[1440] <= ~layer0_out[8] | layer0_out[7];
     layer1_out[1441] <= layer0_out[278] | layer0_out[279];
     layer1_out[1442] <= 1'b0;
     layer1_out[1443] <= 1'b0;
     layer1_out[1444] <= 1'b0;
     layer1_out[1445] <= 1'b0;
     layer1_out[1446] <= 1'b0;
     layer1_out[1447] <= ~layer0_out[828] | layer0_out[827];
     layer1_out[1448] <= ~layer0_out[132] | layer0_out[131];
     layer1_out[1449] <= layer0_out[543] | layer0_out[544];
     layer1_out[1450] <= ~layer0_out[1336] | layer0_out[1335];
     layer1_out[1451] <= 1'b0;
     layer1_out[1452] <= 1'b0;
     layer1_out[1453] <= ~layer0_out[258];
     layer1_out[1454] <= 1'b1;
     layer1_out[1455] <= ~layer0_out[606];
     layer1_out[1456] <= ~layer0_out[513];
     layer1_out[1457] <= ~(layer0_out[1316] ^ layer0_out[1317]);
     layer1_out[1458] <= layer0_out[1282] & layer0_out[1283];
     layer1_out[1459] <= 1'b1;
     layer1_out[1460] <= ~(layer0_out[1089] | layer0_out[1090]);
     layer1_out[1461] <= layer0_out[959] & ~layer0_out[960];
     layer1_out[1462] <= 1'b0;
     layer1_out[1463] <= layer0_out[110];
     layer1_out[1464] <= layer0_out[699] & ~layer0_out[698];
     layer1_out[1465] <= layer0_out[132] & ~layer0_out[133];
     layer1_out[1466] <= layer0_out[592] & ~layer0_out[593];
     layer1_out[1467] <= ~layer0_out[818];
     layer1_out[1468] <= 1'b1;
     layer1_out[1469] <= 1'b0;
     layer1_out[1470] <= ~layer0_out[850];
     layer1_out[1471] <= layer0_out[114] & ~layer0_out[113];
     layer1_out[1472] <= ~(layer0_out[334] & layer0_out[335]);
     layer1_out[1473] <= ~layer0_out[392] | layer0_out[391];
     layer1_out[1474] <= layer0_out[1115] | layer0_out[1116];
     layer1_out[1475] <= ~(layer0_out[1336] & layer0_out[1337]);
     layer1_out[1476] <= layer0_out[1232];
     layer1_out[1477] <= layer0_out[699];
     layer1_out[1478] <= layer0_out[327];
     layer1_out[1479] <= layer0_out[767] | layer0_out[768];
     layer1_out[1480] <= layer0_out[130];
     layer1_out[1481] <= 1'b1;
     layer1_out[1482] <= 1'b1;
     layer1_out[1483] <= layer0_out[1184] & ~layer0_out[1185];
     layer1_out[1484] <= layer0_out[718] & ~layer0_out[719];
     layer1_out[1485] <= layer0_out[184] | layer0_out[185];
     layer1_out[1486] <= ~(layer0_out[738] | layer0_out[739]);
     layer1_out[1487] <= ~(layer0_out[1483] | layer0_out[1484]);
     layer1_out[1488] <= layer0_out[1165] & ~layer0_out[1166];
     layer1_out[1489] <= layer0_out[1189] & ~layer0_out[1188];
     layer1_out[1490] <= ~(layer0_out[865] & layer0_out[866]);
     layer1_out[1491] <= ~(layer0_out[1095] | layer0_out[1096]);
     layer1_out[1492] <= ~layer0_out[1455] | layer0_out[1454];
     layer1_out[1493] <= 1'b1;
     layer1_out[1494] <= 1'b1;
     layer1_out[1495] <= ~(layer0_out[1305] ^ layer0_out[1306]);
     layer1_out[1496] <= ~layer0_out[1370] | layer0_out[1369];
     layer1_out[1497] <= ~layer0_out[1093];
     layer1_out[1498] <= ~(layer0_out[239] & layer0_out[240]);
     layer1_out[1499] <= 1'b0;
     layer2_out[0] <= ~(layer1_out[146] & layer1_out[147]);
     layer2_out[1] <= ~(layer1_out[1166] | layer1_out[1167]);
     layer2_out[2] <= layer1_out[733] & ~layer1_out[734];
     layer2_out[3] <= layer1_out[1223];
     layer2_out[4] <= ~layer1_out[768] | layer1_out[769];
     layer2_out[5] <= 1'b0;
     layer2_out[6] <= layer1_out[487] & layer1_out[488];
     layer2_out[7] <= ~layer1_out[839];
     layer2_out[8] <= layer1_out[375];
     layer2_out[9] <= ~layer1_out[738];
     layer2_out[10] <= layer1_out[954];
     layer2_out[11] <= 1'b1;
     layer2_out[12] <= layer1_out[1355] & layer1_out[1356];
     layer2_out[13] <= layer1_out[1121] | layer1_out[1122];
     layer2_out[14] <= layer1_out[525] | layer1_out[526];
     layer2_out[15] <= 1'b0;
     layer2_out[16] <= 1'b0;
     layer2_out[17] <= ~(layer1_out[562] & layer1_out[563]);
     layer2_out[18] <= layer1_out[1486] | layer1_out[1487];
     layer2_out[19] <= layer1_out[570] & layer1_out[571];
     layer2_out[20] <= layer1_out[544] | layer1_out[545];
     layer2_out[21] <= layer1_out[585] ^ layer1_out[586];
     layer2_out[22] <= layer1_out[1480];
     layer2_out[23] <= ~layer1_out[831] | layer1_out[830];
     layer2_out[24] <= layer1_out[1287] & layer1_out[1288];
     layer2_out[25] <= ~layer1_out[105];
     layer2_out[26] <= layer1_out[0] | layer1_out[2];
     layer2_out[27] <= ~layer1_out[1460];
     layer2_out[28] <= ~layer1_out[961];
     layer2_out[29] <= layer1_out[330];
     layer2_out[30] <= layer1_out[929] & ~layer1_out[930];
     layer2_out[31] <= ~layer1_out[1147];
     layer2_out[32] <= layer1_out[185] | layer1_out[186];
     layer2_out[33] <= ~layer1_out[938] | layer1_out[939];
     layer2_out[34] <= ~(layer1_out[988] | layer1_out[989]);
     layer2_out[35] <= ~(layer1_out[590] & layer1_out[591]);
     layer2_out[36] <= layer1_out[339];
     layer2_out[37] <= layer1_out[1221] & ~layer1_out[1222];
     layer2_out[38] <= 1'b0;
     layer2_out[39] <= ~layer1_out[1];
     layer2_out[40] <= layer1_out[314] | layer1_out[315];
     layer2_out[41] <= 1'b0;
     layer2_out[42] <= layer1_out[1200] & ~layer1_out[1201];
     layer2_out[43] <= ~layer1_out[126];
     layer2_out[44] <= ~layer1_out[599];
     layer2_out[45] <= ~layer1_out[147];
     layer2_out[46] <= ~(layer1_out[1258] | layer1_out[1259]);
     layer2_out[47] <= 1'b0;
     layer2_out[48] <= 1'b1;
     layer2_out[49] <= ~layer1_out[36] | layer1_out[37];
     layer2_out[50] <= 1'b1;
     layer2_out[51] <= ~layer1_out[497];
     layer2_out[52] <= ~layer1_out[1106] | layer1_out[1105];
     layer2_out[53] <= layer1_out[1052];
     layer2_out[54] <= 1'b1;
     layer2_out[55] <= layer1_out[1033];
     layer2_out[56] <= 1'b1;
     layer2_out[57] <= ~layer1_out[1184] | layer1_out[1183];
     layer2_out[58] <= layer1_out[397];
     layer2_out[59] <= layer1_out[465] & ~layer1_out[466];
     layer2_out[60] <= layer1_out[938];
     layer2_out[61] <= ~(layer1_out[955] | layer1_out[956]);
     layer2_out[62] <= ~layer1_out[1304];
     layer2_out[63] <= layer1_out[1422] & layer1_out[1423];
     layer2_out[64] <= ~(layer1_out[782] & layer1_out[783]);
     layer2_out[65] <= layer1_out[366] & ~layer1_out[367];
     layer2_out[66] <= ~layer1_out[730];
     layer2_out[67] <= layer1_out[877];
     layer2_out[68] <= layer1_out[980] & layer1_out[981];
     layer2_out[69] <= 1'b0;
     layer2_out[70] <= ~layer1_out[138];
     layer2_out[71] <= ~layer1_out[723] | layer1_out[722];
     layer2_out[72] <= 1'b1;
     layer2_out[73] <= layer1_out[179] & ~layer1_out[178];
     layer2_out[74] <= layer1_out[694] & ~layer1_out[693];
     layer2_out[75] <= layer1_out[1155] ^ layer1_out[1156];
     layer2_out[76] <= 1'b0;
     layer2_out[77] <= layer1_out[644];
     layer2_out[78] <= 1'b0;
     layer2_out[79] <= layer1_out[1417] & ~layer1_out[1418];
     layer2_out[80] <= 1'b1;
     layer2_out[81] <= layer1_out[173];
     layer2_out[82] <= layer1_out[956] | layer1_out[957];
     layer2_out[83] <= 1'b0;
     layer2_out[84] <= layer1_out[111] & layer1_out[112];
     layer2_out[85] <= layer1_out[1223] | layer1_out[1224];
     layer2_out[86] <= ~(layer1_out[1104] | layer1_out[1105]);
     layer2_out[87] <= ~layer1_out[1359] | layer1_out[1358];
     layer2_out[88] <= ~layer1_out[11];
     layer2_out[89] <= layer1_out[153] | layer1_out[154];
     layer2_out[90] <= ~layer1_out[558] | layer1_out[559];
     layer2_out[91] <= 1'b1;
     layer2_out[92] <= ~(layer1_out[1346] | layer1_out[1347]);
     layer2_out[93] <= layer1_out[382] & ~layer1_out[383];
     layer2_out[94] <= layer1_out[868] & ~layer1_out[869];
     layer2_out[95] <= ~layer1_out[900] | layer1_out[901];
     layer2_out[96] <= layer1_out[226] & ~layer1_out[227];
     layer2_out[97] <= ~layer1_out[407] | layer1_out[408];
     layer2_out[98] <= layer1_out[166];
     layer2_out[99] <= layer1_out[419];
     layer2_out[100] <= ~(layer1_out[1316] & layer1_out[1317]);
     layer2_out[101] <= ~layer1_out[1136];
     layer2_out[102] <= ~layer1_out[7] | layer1_out[6];
     layer2_out[103] <= layer1_out[351] | layer1_out[352];
     layer2_out[104] <= layer1_out[78];
     layer2_out[105] <= layer1_out[890] | layer1_out[891];
     layer2_out[106] <= layer1_out[758] | layer1_out[759];
     layer2_out[107] <= layer1_out[542] & layer1_out[543];
     layer2_out[108] <= layer1_out[310] & ~layer1_out[311];
     layer2_out[109] <= 1'b0;
     layer2_out[110] <= layer1_out[553];
     layer2_out[111] <= ~layer1_out[764];
     layer2_out[112] <= layer1_out[748] & ~layer1_out[747];
     layer2_out[113] <= ~layer1_out[1179] | layer1_out[1178];
     layer2_out[114] <= layer1_out[681] & layer1_out[682];
     layer2_out[115] <= layer1_out[296] & ~layer1_out[297];
     layer2_out[116] <= 1'b0;
     layer2_out[117] <= 1'b1;
     layer2_out[118] <= layer1_out[1088];
     layer2_out[119] <= ~layer1_out[28] | layer1_out[29];
     layer2_out[120] <= 1'b0;
     layer2_out[121] <= ~layer1_out[552] | layer1_out[551];
     layer2_out[122] <= layer1_out[1004] & layer1_out[1005];
     layer2_out[123] <= layer1_out[652];
     layer2_out[124] <= ~layer1_out[91] | layer1_out[90];
     layer2_out[125] <= ~(layer1_out[577] | layer1_out[578]);
     layer2_out[126] <= layer1_out[1323] & layer1_out[1324];
     layer2_out[127] <= ~layer1_out[772];
     layer2_out[128] <= 1'b0;
     layer2_out[129] <= layer1_out[894] & ~layer1_out[895];
     layer2_out[130] <= ~layer1_out[401] | layer1_out[400];
     layer2_out[131] <= layer1_out[1136] | layer1_out[1137];
     layer2_out[132] <= ~layer1_out[1072];
     layer2_out[133] <= layer1_out[1143] & layer1_out[1144];
     layer2_out[134] <= 1'b0;
     layer2_out[135] <= ~layer1_out[875] | layer1_out[876];
     layer2_out[136] <= layer1_out[787] & ~layer1_out[788];
     layer2_out[137] <= layer1_out[1206] & layer1_out[1207];
     layer2_out[138] <= 1'b0;
     layer2_out[139] <= layer1_out[666] & ~layer1_out[667];
     layer2_out[140] <= ~layer1_out[1307];
     layer2_out[141] <= 1'b0;
     layer2_out[142] <= ~layer1_out[249];
     layer2_out[143] <= layer1_out[163] & ~layer1_out[164];
     layer2_out[144] <= ~layer1_out[186] | layer1_out[187];
     layer2_out[145] <= ~(layer1_out[644] & layer1_out[645]);
     layer2_out[146] <= ~(layer1_out[1273] | layer1_out[1274]);
     layer2_out[147] <= layer1_out[1485];
     layer2_out[148] <= ~(layer1_out[1336] ^ layer1_out[1337]);
     layer2_out[149] <= ~(layer1_out[1463] & layer1_out[1464]);
     layer2_out[150] <= layer1_out[1271] & ~layer1_out[1272];
     layer2_out[151] <= layer1_out[439] & layer1_out[440];
     layer2_out[152] <= ~layer1_out[356];
     layer2_out[153] <= layer1_out[1230] & ~layer1_out[1229];
     layer2_out[154] <= 1'b0;
     layer2_out[155] <= layer1_out[182] | layer1_out[183];
     layer2_out[156] <= ~layer1_out[1124];
     layer2_out[157] <= layer1_out[745] & ~layer1_out[744];
     layer2_out[158] <= ~layer1_out[53];
     layer2_out[159] <= ~(layer1_out[891] & layer1_out[892]);
     layer2_out[160] <= ~layer1_out[45];
     layer2_out[161] <= ~layer1_out[171] | layer1_out[172];
     layer2_out[162] <= layer1_out[1356] | layer1_out[1357];
     layer2_out[163] <= ~layer1_out[1251];
     layer2_out[164] <= layer1_out[460] & ~layer1_out[459];
     layer2_out[165] <= ~layer1_out[701] | layer1_out[700];
     layer2_out[166] <= ~(layer1_out[701] | layer1_out[702]);
     layer2_out[167] <= layer1_out[128] | layer1_out[129];
     layer2_out[168] <= layer1_out[1252] & layer1_out[1253];
     layer2_out[169] <= ~(layer1_out[428] | layer1_out[429]);
     layer2_out[170] <= ~layer1_out[796];
     layer2_out[171] <= ~layer1_out[107];
     layer2_out[172] <= ~layer1_out[1184];
     layer2_out[173] <= 1'b1;
     layer2_out[174] <= 1'b1;
     layer2_out[175] <= 1'b0;
     layer2_out[176] <= ~layer1_out[1131];
     layer2_out[177] <= ~(layer1_out[7] | layer1_out[8]);
     layer2_out[178] <= layer1_out[450] & ~layer1_out[451];
     layer2_out[179] <= layer1_out[972] & ~layer1_out[971];
     layer2_out[180] <= layer1_out[1216];
     layer2_out[181] <= layer1_out[1039];
     layer2_out[182] <= layer1_out[1129] & layer1_out[1130];
     layer2_out[183] <= 1'b0;
     layer2_out[184] <= layer1_out[2] | layer1_out[3];
     layer2_out[185] <= ~(layer1_out[748] & layer1_out[749]);
     layer2_out[186] <= 1'b0;
     layer2_out[187] <= ~layer1_out[1414] | layer1_out[1413];
     layer2_out[188] <= 1'b0;
     layer2_out[189] <= layer1_out[399] & ~layer1_out[398];
     layer2_out[190] <= ~layer1_out[521];
     layer2_out[191] <= layer1_out[819] & ~layer1_out[818];
     layer2_out[192] <= ~(layer1_out[933] & layer1_out[934]);
     layer2_out[193] <= layer1_out[1245] | layer1_out[1246];
     layer2_out[194] <= 1'b1;
     layer2_out[195] <= layer1_out[231] ^ layer1_out[232];
     layer2_out[196] <= ~(layer1_out[1448] | layer1_out[1449]);
     layer2_out[197] <= ~(layer1_out[212] & layer1_out[213]);
     layer2_out[198] <= layer1_out[51] & ~layer1_out[52];
     layer2_out[199] <= ~layer1_out[671];
     layer2_out[200] <= layer1_out[930] | layer1_out[931];
     layer2_out[201] <= 1'b1;
     layer2_out[202] <= ~layer1_out[1221];
     layer2_out[203] <= layer1_out[31];
     layer2_out[204] <= ~layer1_out[403];
     layer2_out[205] <= ~layer1_out[866];
     layer2_out[206] <= ~(layer1_out[1438] | layer1_out[1439]);
     layer2_out[207] <= ~layer1_out[242];
     layer2_out[208] <= ~layer1_out[199] | layer1_out[198];
     layer2_out[209] <= layer1_out[627] ^ layer1_out[628];
     layer2_out[210] <= layer1_out[468] | layer1_out[469];
     layer2_out[211] <= ~layer1_out[746] | layer1_out[747];
     layer2_out[212] <= ~(layer1_out[106] | layer1_out[107]);
     layer2_out[213] <= layer1_out[289];
     layer2_out[214] <= layer1_out[1330];
     layer2_out[215] <= layer1_out[144] & layer1_out[145];
     layer2_out[216] <= ~(layer1_out[602] | layer1_out[603]);
     layer2_out[217] <= layer1_out[841] & ~layer1_out[842];
     layer2_out[218] <= ~layer1_out[869] | layer1_out[870];
     layer2_out[219] <= 1'b1;
     layer2_out[220] <= layer1_out[1365];
     layer2_out[221] <= ~layer1_out[188] | layer1_out[189];
     layer2_out[222] <= layer1_out[1477];
     layer2_out[223] <= ~layer1_out[889] | layer1_out[888];
     layer2_out[224] <= 1'b0;
     layer2_out[225] <= ~(layer1_out[292] | layer1_out[293]);
     layer2_out[226] <= ~(layer1_out[832] | layer1_out[833]);
     layer2_out[227] <= layer1_out[92];
     layer2_out[228] <= 1'b0;
     layer2_out[229] <= ~(layer1_out[713] | layer1_out[714]);
     layer2_out[230] <= layer1_out[705];
     layer2_out[231] <= ~layer1_out[968];
     layer2_out[232] <= layer1_out[17] & ~layer1_out[16];
     layer2_out[233] <= ~(layer1_out[1455] | layer1_out[1456]);
     layer2_out[234] <= 1'b0;
     layer2_out[235] <= layer1_out[244];
     layer2_out[236] <= layer1_out[844] & layer1_out[845];
     layer2_out[237] <= ~(layer1_out[1214] | layer1_out[1215]);
     layer2_out[238] <= layer1_out[282] & ~layer1_out[283];
     layer2_out[239] <= layer1_out[161] & ~layer1_out[162];
     layer2_out[240] <= 1'b0;
     layer2_out[241] <= ~layer1_out[371];
     layer2_out[242] <= ~layer1_out[1498];
     layer2_out[243] <= layer1_out[25] & layer1_out[26];
     layer2_out[244] <= layer1_out[967] & ~layer1_out[966];
     layer2_out[245] <= layer1_out[651] & layer1_out[652];
     layer2_out[246] <= 1'b1;
     layer2_out[247] <= 1'b1;
     layer2_out[248] <= layer1_out[409] | layer1_out[410];
     layer2_out[249] <= layer1_out[879];
     layer2_out[250] <= layer1_out[502];
     layer2_out[251] <= 1'b1;
     layer2_out[252] <= ~layer1_out[1495] | layer1_out[1496];
     layer2_out[253] <= layer1_out[827];
     layer2_out[254] <= layer1_out[1156] & layer1_out[1157];
     layer2_out[255] <= 1'b0;
     layer2_out[256] <= ~(layer1_out[945] ^ layer1_out[946]);
     layer2_out[257] <= 1'b1;
     layer2_out[258] <= ~layer1_out[848] | layer1_out[847];
     layer2_out[259] <= ~layer1_out[841];
     layer2_out[260] <= ~(layer1_out[1107] | layer1_out[1108]);
     layer2_out[261] <= ~layer1_out[114] | layer1_out[115];
     layer2_out[262] <= ~layer1_out[101];
     layer2_out[263] <= layer1_out[1018];
     layer2_out[264] <= layer1_out[596] & layer1_out[597];
     layer2_out[265] <= layer1_out[1003] & ~layer1_out[1004];
     layer2_out[266] <= layer1_out[1236] & ~layer1_out[1237];
     layer2_out[267] <= 1'b0;
     layer2_out[268] <= 1'b1;
     layer2_out[269] <= layer1_out[180] & ~layer1_out[179];
     layer2_out[270] <= ~layer1_out[1473];
     layer2_out[271] <= ~layer1_out[1425] | layer1_out[1424];
     layer2_out[272] <= layer1_out[1383];
     layer2_out[273] <= ~(layer1_out[1234] & layer1_out[1235]);
     layer2_out[274] <= ~layer1_out[60] | layer1_out[59];
     layer2_out[275] <= 1'b1;
     layer2_out[276] <= ~(layer1_out[1062] & layer1_out[1063]);
     layer2_out[277] <= ~(layer1_out[1123] | layer1_out[1124]);
     layer2_out[278] <= layer1_out[1112];
     layer2_out[279] <= ~(layer1_out[1067] & layer1_out[1068]);
     layer2_out[280] <= ~(layer1_out[690] | layer1_out[691]);
     layer2_out[281] <= ~layer1_out[512] | layer1_out[513];
     layer2_out[282] <= ~layer1_out[690];
     layer2_out[283] <= layer1_out[715] & ~layer1_out[716];
     layer2_out[284] <= 1'b0;
     layer2_out[285] <= 1'b0;
     layer2_out[286] <= ~layer1_out[464];
     layer2_out[287] <= ~layer1_out[556] | layer1_out[555];
     layer2_out[288] <= layer1_out[1029] & layer1_out[1030];
     layer2_out[289] <= ~layer1_out[1400];
     layer2_out[290] <= ~(layer1_out[1219] & layer1_out[1220]);
     layer2_out[291] <= ~(layer1_out[1406] | layer1_out[1407]);
     layer2_out[292] <= ~layer1_out[499];
     layer2_out[293] <= ~layer1_out[348] | layer1_out[347];
     layer2_out[294] <= ~layer1_out[1000] | layer1_out[1001];
     layer2_out[295] <= 1'b1;
     layer2_out[296] <= ~layer1_out[1181];
     layer2_out[297] <= 1'b1;
     layer2_out[298] <= ~(layer1_out[1378] & layer1_out[1379]);
     layer2_out[299] <= layer1_out[582] & ~layer1_out[583];
     layer2_out[300] <= ~layer1_out[1480];
     layer2_out[301] <= ~(layer1_out[1400] | layer1_out[1401]);
     layer2_out[302] <= layer1_out[664] & ~layer1_out[663];
     layer2_out[303] <= ~layer1_out[653] | layer1_out[654];
     layer2_out[304] <= layer1_out[1269];
     layer2_out[305] <= layer1_out[536];
     layer2_out[306] <= ~(layer1_out[1367] | layer1_out[1368]);
     layer2_out[307] <= 1'b0;
     layer2_out[308] <= ~(layer1_out[639] | layer1_out[640]);
     layer2_out[309] <= 1'b0;
     layer2_out[310] <= ~layer1_out[708] | layer1_out[707];
     layer2_out[311] <= ~(layer1_out[559] | layer1_out[560]);
     layer2_out[312] <= layer1_out[1375] | layer1_out[1376];
     layer2_out[313] <= layer1_out[1187];
     layer2_out[314] <= layer1_out[1377] & layer1_out[1378];
     layer2_out[315] <= layer1_out[633] & ~layer1_out[632];
     layer2_out[316] <= ~(layer1_out[442] | layer1_out[443]);
     layer2_out[317] <= ~layer1_out[977];
     layer2_out[318] <= layer1_out[139] | layer1_out[140];
     layer2_out[319] <= ~layer1_out[358] | layer1_out[359];
     layer2_out[320] <= ~layer1_out[1370] | layer1_out[1369];
     layer2_out[321] <= 1'b0;
     layer2_out[322] <= layer1_out[1420] & ~layer1_out[1421];
     layer2_out[323] <= layer1_out[1472] | layer1_out[1473];
     layer2_out[324] <= ~layer1_out[1192];
     layer2_out[325] <= layer1_out[569] & ~layer1_out[570];
     layer2_out[326] <= layer1_out[656] & ~layer1_out[655];
     layer2_out[327] <= layer1_out[609] & layer1_out[610];
     layer2_out[328] <= ~layer1_out[236];
     layer2_out[329] <= ~(layer1_out[683] & layer1_out[684]);
     layer2_out[330] <= ~layer1_out[785] | layer1_out[784];
     layer2_out[331] <= layer1_out[313];
     layer2_out[332] <= ~(layer1_out[757] ^ layer1_out[758]);
     layer2_out[333] <= ~layer1_out[368] | layer1_out[367];
     layer2_out[334] <= layer1_out[979];
     layer2_out[335] <= layer1_out[238];
     layer2_out[336] <= ~layer1_out[565];
     layer2_out[337] <= ~layer1_out[727] | layer1_out[728];
     layer2_out[338] <= layer1_out[516];
     layer2_out[339] <= 1'b0;
     layer2_out[340] <= ~(layer1_out[50] | layer1_out[51]);
     layer2_out[341] <= ~(layer1_out[823] & layer1_out[824]);
     layer2_out[342] <= layer1_out[908] & ~layer1_out[909];
     layer2_out[343] <= layer1_out[120] & ~layer1_out[121];
     layer2_out[344] <= ~layer1_out[1493];
     layer2_out[345] <= ~layer1_out[43];
     layer2_out[346] <= layer1_out[1329] & layer1_out[1330];
     layer2_out[347] <= ~layer1_out[850];
     layer2_out[348] <= ~layer1_out[1317];
     layer2_out[349] <= ~layer1_out[1447] | layer1_out[1448];
     layer2_out[350] <= ~(layer1_out[984] | layer1_out[985]);
     layer2_out[351] <= ~layer1_out[243] | layer1_out[242];
     layer2_out[352] <= ~layer1_out[849];
     layer2_out[353] <= ~(layer1_out[692] & layer1_out[693]);
     layer2_out[354] <= layer1_out[860];
     layer2_out[355] <= layer1_out[497];
     layer2_out[356] <= ~(layer1_out[1497] | layer1_out[1498]);
     layer2_out[357] <= ~layer1_out[218];
     layer2_out[358] <= ~(layer1_out[1394] | layer1_out[1395]);
     layer2_out[359] <= 1'b0;
     layer2_out[360] <= layer1_out[194] & ~layer1_out[195];
     layer2_out[361] <= ~(layer1_out[38] | layer1_out[39]);
     layer2_out[362] <= 1'b0;
     layer2_out[363] <= layer1_out[1451] & layer1_out[1452];
     layer2_out[364] <= 1'b1;
     layer2_out[365] <= 1'b0;
     layer2_out[366] <= ~layer1_out[1044] | layer1_out[1045];
     layer2_out[367] <= ~(layer1_out[474] & layer1_out[475]);
     layer2_out[368] <= layer1_out[40];
     layer2_out[369] <= layer1_out[1127] | layer1_out[1128];
     layer2_out[370] <= layer1_out[577];
     layer2_out[371] <= ~layer1_out[1053] | layer1_out[1052];
     layer2_out[372] <= ~layer1_out[1204] | layer1_out[1203];
     layer2_out[373] <= layer1_out[473];
     layer2_out[374] <= 1'b1;
     layer2_out[375] <= 1'b1;
     layer2_out[376] <= ~(layer1_out[1402] | layer1_out[1403]);
     layer2_out[377] <= layer1_out[989] | layer1_out[990];
     layer2_out[378] <= 1'b0;
     layer2_out[379] <= layer1_out[1014] | layer1_out[1015];
     layer2_out[380] <= ~layer1_out[614];
     layer2_out[381] <= ~layer1_out[1074];
     layer2_out[382] <= layer1_out[247] & layer1_out[248];
     layer2_out[383] <= 1'b1;
     layer2_out[384] <= 1'b0;
     layer2_out[385] <= 1'b0;
     layer2_out[386] <= ~(layer1_out[765] | layer1_out[766]);
     layer2_out[387] <= layer1_out[268] & layer1_out[269];
     layer2_out[388] <= layer1_out[1299] & ~layer1_out[1298];
     layer2_out[389] <= ~layer1_out[592] | layer1_out[591];
     layer2_out[390] <= ~layer1_out[536];
     layer2_out[391] <= layer1_out[702] | layer1_out[703];
     layer2_out[392] <= ~layer1_out[1462] | layer1_out[1461];
     layer2_out[393] <= 1'b1;
     layer2_out[394] <= ~layer1_out[854] | layer1_out[853];
     layer2_out[395] <= ~layer1_out[614];
     layer2_out[396] <= ~(layer1_out[985] & layer1_out[986]);
     layer2_out[397] <= layer1_out[214] & ~layer1_out[213];
     layer2_out[398] <= ~(layer1_out[279] ^ layer1_out[280]);
     layer2_out[399] <= layer1_out[1013] & ~layer1_out[1014];
     layer2_out[400] <= 1'b0;
     layer2_out[401] <= 1'b1;
     layer2_out[402] <= ~layer1_out[322];
     layer2_out[403] <= 1'b1;
     layer2_out[404] <= ~layer1_out[736] | layer1_out[735];
     layer2_out[405] <= layer1_out[743] & layer1_out[744];
     layer2_out[406] <= layer1_out[1157] ^ layer1_out[1158];
     layer2_out[407] <= layer1_out[423] | layer1_out[424];
     layer2_out[408] <= layer1_out[243] & layer1_out[244];
     layer2_out[409] <= ~(layer1_out[1427] | layer1_out[1428]);
     layer2_out[410] <= layer1_out[1243];
     layer2_out[411] <= ~layer1_out[721] | layer1_out[720];
     layer2_out[412] <= ~(layer1_out[970] & layer1_out[971]);
     layer2_out[413] <= 1'b1;
     layer2_out[414] <= ~layer1_out[72] | layer1_out[73];
     layer2_out[415] <= ~(layer1_out[307] & layer1_out[308]);
     layer2_out[416] <= 1'b0;
     layer2_out[417] <= ~layer1_out[804] | layer1_out[805];
     layer2_out[418] <= ~(layer1_out[583] | layer1_out[584]);
     layer2_out[419] <= 1'b1;
     layer2_out[420] <= ~layer1_out[387];
     layer2_out[421] <= ~layer1_out[632] | layer1_out[631];
     layer2_out[422] <= 1'b0;
     layer2_out[423] <= layer1_out[966];
     layer2_out[424] <= layer1_out[152];
     layer2_out[425] <= layer1_out[172];
     layer2_out[426] <= ~layer1_out[1491] | layer1_out[1490];
     layer2_out[427] <= ~layer1_out[306];
     layer2_out[428] <= layer1_out[888];
     layer2_out[429] <= 1'b1;
     layer2_out[430] <= 1'b0;
     layer2_out[431] <= layer1_out[1456] | layer1_out[1457];
     layer2_out[432] <= ~layer1_out[1277];
     layer2_out[433] <= layer1_out[297] & ~layer1_out[298];
     layer2_out[434] <= ~(layer1_out[549] & layer1_out[550]);
     layer2_out[435] <= layer1_out[783];
     layer2_out[436] <= 1'b1;
     layer2_out[437] <= layer1_out[413];
     layer2_out[438] <= 1'b1;
     layer2_out[439] <= ~(layer1_out[608] & layer1_out[609]);
     layer2_out[440] <= ~layer1_out[1405];
     layer2_out[441] <= layer1_out[413] & layer1_out[414];
     layer2_out[442] <= layer1_out[1122];
     layer2_out[443] <= layer1_out[464] & layer1_out[465];
     layer2_out[444] <= layer1_out[684] & layer1_out[685];
     layer2_out[445] <= ~(layer1_out[313] & layer1_out[314]);
     layer2_out[446] <= ~(layer1_out[35] | layer1_out[36]);
     layer2_out[447] <= ~(layer1_out[385] & layer1_out[386]);
     layer2_out[448] <= 1'b0;
     layer2_out[449] <= 1'b1;
     layer2_out[450] <= layer1_out[524] & ~layer1_out[523];
     layer2_out[451] <= ~(layer1_out[320] | layer1_out[321]);
     layer2_out[452] <= layer1_out[245] & ~layer1_out[246];
     layer2_out[453] <= ~(layer1_out[580] | layer1_out[581]);
     layer2_out[454] <= layer1_out[706] & ~layer1_out[707];
     layer2_out[455] <= layer1_out[817] & ~layer1_out[818];
     layer2_out[456] <= ~(layer1_out[58] & layer1_out[59]);
     layer2_out[457] <= ~(layer1_out[1114] | layer1_out[1115]);
     layer2_out[458] <= layer1_out[1086] | layer1_out[1087];
     layer2_out[459] <= layer1_out[545] & layer1_out[546];
     layer2_out[460] <= 1'b1;
     layer2_out[461] <= 1'b0;
     layer2_out[462] <= 1'b1;
     layer2_out[463] <= 1'b1;
     layer2_out[464] <= 1'b1;
     layer2_out[465] <= layer1_out[257] & layer1_out[258];
     layer2_out[466] <= ~layer1_out[1163];
     layer2_out[467] <= ~layer1_out[914] | layer1_out[913];
     layer2_out[468] <= ~layer1_out[1377];
     layer2_out[469] <= layer1_out[1226];
     layer2_out[470] <= layer1_out[896];
     layer2_out[471] <= ~(layer1_out[174] | layer1_out[175]);
     layer2_out[472] <= layer1_out[122] | layer1_out[123];
     layer2_out[473] <= ~(layer1_out[1182] & layer1_out[1183]);
     layer2_out[474] <= 1'b1;
     layer2_out[475] <= ~layer1_out[158] | layer1_out[159];
     layer2_out[476] <= layer1_out[141] & ~layer1_out[140];
     layer2_out[477] <= layer1_out[351] & ~layer1_out[350];
     layer2_out[478] <= layer1_out[1285] & ~layer1_out[1284];
     layer2_out[479] <= layer1_out[678] & ~layer1_out[677];
     layer2_out[480] <= ~layer1_out[852] | layer1_out[851];
     layer2_out[481] <= layer1_out[1450] ^ layer1_out[1451];
     layer2_out[482] <= ~layer1_out[661];
     layer2_out[483] <= 1'b0;
     layer2_out[484] <= ~(layer1_out[514] | layer1_out[515]);
     layer2_out[485] <= layer1_out[1139] & ~layer1_out[1140];
     layer2_out[486] <= ~(layer1_out[699] | layer1_out[700]);
     layer2_out[487] <= layer1_out[210] | layer1_out[211];
     layer2_out[488] <= ~layer1_out[1031] | layer1_out[1032];
     layer2_out[489] <= ~layer1_out[250];
     layer2_out[490] <= layer1_out[856] & layer1_out[857];
     layer2_out[491] <= ~(layer1_out[717] & layer1_out[718]);
     layer2_out[492] <= 1'b0;
     layer2_out[493] <= 1'b0;
     layer2_out[494] <= ~layer1_out[1002];
     layer2_out[495] <= 1'b0;
     layer2_out[496] <= layer1_out[145];
     layer2_out[497] <= 1'b1;
     layer2_out[498] <= layer1_out[1099];
     layer2_out[499] <= layer1_out[1278];
     layer2_out[500] <= layer1_out[551];
     layer2_out[501] <= ~layer1_out[1133];
     layer2_out[502] <= layer1_out[883];
     layer2_out[503] <= ~(layer1_out[1237] & layer1_out[1238]);
     layer2_out[504] <= layer1_out[143];
     layer2_out[505] <= layer1_out[824] & layer1_out[825];
     layer2_out[506] <= layer1_out[617] & ~layer1_out[616];
     layer2_out[507] <= layer1_out[34] | layer1_out[35];
     layer2_out[508] <= 1'b0;
     layer2_out[509] <= ~(layer1_out[603] | layer1_out[604]);
     layer2_out[510] <= 1'b1;
     layer2_out[511] <= 1'b0;
     layer2_out[512] <= 1'b1;
     layer2_out[513] <= ~layer1_out[112] | layer1_out[113];
     layer2_out[514] <= layer1_out[855] & ~layer1_out[856];
     layer2_out[515] <= layer1_out[1019];
     layer2_out[516] <= 1'b1;
     layer2_out[517] <= layer1_out[234];
     layer2_out[518] <= layer1_out[760] & ~layer1_out[761];
     layer2_out[519] <= layer1_out[365] & layer1_out[366];
     layer2_out[520] <= ~layer1_out[66] | layer1_out[67];
     layer2_out[521] <= layer1_out[816] & ~layer1_out[815];
     layer2_out[522] <= layer1_out[1301] & ~layer1_out[1302];
     layer2_out[523] <= layer1_out[1359] & ~layer1_out[1360];
     layer2_out[524] <= layer1_out[682] & ~layer1_out[683];
     layer2_out[525] <= ~layer1_out[338];
     layer2_out[526] <= layer1_out[187] & layer1_out[188];
     layer2_out[527] <= layer1_out[1138] & ~layer1_out[1137];
     layer2_out[528] <= 1'b1;
     layer2_out[529] <= layer1_out[495];
     layer2_out[530] <= ~layer1_out[28] | layer1_out[27];
     layer2_out[531] <= 1'b1;
     layer2_out[532] <= layer1_out[23];
     layer2_out[533] <= layer1_out[251] & layer1_out[252];
     layer2_out[534] <= ~layer1_out[1025];
     layer2_out[535] <= ~layer1_out[675];
     layer2_out[536] <= layer1_out[970] & ~layer1_out[969];
     layer2_out[537] <= ~(layer1_out[421] | layer1_out[422]);
     layer2_out[538] <= ~layer1_out[203];
     layer2_out[539] <= layer1_out[348] & ~layer1_out[349];
     layer2_out[540] <= ~(layer1_out[633] & layer1_out[634]);
     layer2_out[541] <= ~layer1_out[1339];
     layer2_out[542] <= ~layer1_out[419] | layer1_out[420];
     layer2_out[543] <= ~(layer1_out[414] & layer1_out[415]);
     layer2_out[544] <= ~layer1_out[829];
     layer2_out[545] <= layer1_out[1469] & ~layer1_out[1468];
     layer2_out[546] <= 1'b1;
     layer2_out[547] <= ~layer1_out[143] | layer1_out[142];
     layer2_out[548] <= layer1_out[791];
     layer2_out[549] <= layer1_out[149];
     layer2_out[550] <= layer1_out[280] & layer1_out[281];
     layer2_out[551] <= 1'b0;
     layer2_out[552] <= layer1_out[1042];
     layer2_out[553] <= layer1_out[1372] | layer1_out[1373];
     layer2_out[554] <= ~layer1_out[41] | layer1_out[42];
     layer2_out[555] <= layer1_out[915];
     layer2_out[556] <= layer1_out[955];
     layer2_out[557] <= layer1_out[298] | layer1_out[299];
     layer2_out[558] <= layer1_out[1022] & ~layer1_out[1021];
     layer2_out[559] <= ~layer1_out[65];
     layer2_out[560] <= layer1_out[141] & ~layer1_out[142];
     layer2_out[561] <= layer1_out[698] & ~layer1_out[699];
     layer2_out[562] <= layer1_out[98] | layer1_out[99];
     layer2_out[563] <= ~layer1_out[1104] | layer1_out[1103];
     layer2_out[564] <= ~layer1_out[1496] | layer1_out[1497];
     layer2_out[565] <= ~layer1_out[500] | layer1_out[501];
     layer2_out[566] <= layer1_out[1092] & ~layer1_out[1091];
     layer2_out[567] <= layer1_out[37] & ~layer1_out[38];
     layer2_out[568] <= layer1_out[734] & layer1_out[735];
     layer2_out[569] <= layer1_out[1089] & ~layer1_out[1090];
     layer2_out[570] <= ~layer1_out[668];
     layer2_out[571] <= ~(layer1_out[406] | layer1_out[407]);
     layer2_out[572] <= ~layer1_out[340] | layer1_out[341];
     layer2_out[573] <= ~layer1_out[488];
     layer2_out[574] <= layer1_out[927];
     layer2_out[575] <= layer1_out[1181] & layer1_out[1182];
     layer2_out[576] <= ~layer1_out[455] | layer1_out[454];
     layer2_out[577] <= layer1_out[866];
     layer2_out[578] <= layer1_out[723] & ~layer1_out[724];
     layer2_out[579] <= ~(layer1_out[1046] & layer1_out[1047]);
     layer2_out[580] <= layer1_out[1284];
     layer2_out[581] <= layer1_out[337] & ~layer1_out[336];
     layer2_out[582] <= layer1_out[1083];
     layer2_out[583] <= layer1_out[996] & ~layer1_out[995];
     layer2_out[584] <= 1'b0;
     layer2_out[585] <= layer1_out[1199] & layer1_out[1200];
     layer2_out[586] <= layer1_out[1369] & ~layer1_out[1368];
     layer2_out[587] <= ~(layer1_out[1485] | layer1_out[1486]);
     layer2_out[588] <= ~layer1_out[427];
     layer2_out[589] <= layer1_out[1084] & layer1_out[1085];
     layer2_out[590] <= layer1_out[1034] & ~layer1_out[1033];
     layer2_out[591] <= ~(layer1_out[1009] | layer1_out[1010]);
     layer2_out[592] <= ~layer1_out[1008] | layer1_out[1009];
     layer2_out[593] <= ~(layer1_out[46] & layer1_out[47]);
     layer2_out[594] <= ~layer1_out[528];
     layer2_out[595] <= layer1_out[947];
     layer2_out[596] <= layer1_out[839];
     layer2_out[597] <= 1'b0;
     layer2_out[598] <= ~layer1_out[1314] | layer1_out[1313];
     layer2_out[599] <= ~layer1_out[926];
     layer2_out[600] <= 1'b0;
     layer2_out[601] <= ~(layer1_out[1279] | layer1_out[1280]);
     layer2_out[602] <= ~layer1_out[903] | layer1_out[904];
     layer2_out[603] <= layer1_out[199];
     layer2_out[604] <= ~(layer1_out[89] | layer1_out[90]);
     layer2_out[605] <= ~(layer1_out[518] | layer1_out[519]);
     layer2_out[606] <= ~layer1_out[196] | layer1_out[197];
     layer2_out[607] <= ~(layer1_out[1253] | layer1_out[1254]);
     layer2_out[608] <= 1'b0;
     layer2_out[609] <= layer1_out[402] & layer1_out[403];
     layer2_out[610] <= 1'b1;
     layer2_out[611] <= ~layer1_out[903];
     layer2_out[612] <= ~layer1_out[540] | layer1_out[541];
     layer2_out[613] <= 1'b1;
     layer2_out[614] <= ~layer1_out[1208];
     layer2_out[615] <= 1'b1;
     layer2_out[616] <= layer1_out[1332] & layer1_out[1333];
     layer2_out[617] <= layer1_out[618] & ~layer1_out[617];
     layer2_out[618] <= 1'b0;
     layer2_out[619] <= 1'b1;
     layer2_out[620] <= layer1_out[1070] & ~layer1_out[1071];
     layer2_out[621] <= ~(layer1_out[1419] & layer1_out[1420]);
     layer2_out[622] <= layer1_out[770];
     layer2_out[623] <= ~layer1_out[1383];
     layer2_out[624] <= 1'b1;
     layer2_out[625] <= layer1_out[344];
     layer2_out[626] <= 1'b1;
     layer2_out[627] <= ~layer1_out[1056];
     layer2_out[628] <= ~layer1_out[62] | layer1_out[63];
     layer2_out[629] <= layer1_out[289] & ~layer1_out[290];
     layer2_out[630] <= layer1_out[1197] & layer1_out[1198];
     layer2_out[631] <= 1'b1;
     layer2_out[632] <= 1'b1;
     layer2_out[633] <= ~(layer1_out[75] | layer1_out[76]);
     layer2_out[634] <= ~layer1_out[1334] | layer1_out[1335];
     layer2_out[635] <= layer1_out[259];
     layer2_out[636] <= layer1_out[80] & ~layer1_out[79];
     layer2_out[637] <= ~layer1_out[14];
     layer2_out[638] <= layer1_out[31];
     layer2_out[639] <= layer1_out[560] ^ layer1_out[561];
     layer2_out[640] <= ~(layer1_out[1195] | layer1_out[1196]);
     layer2_out[641] <= ~(layer1_out[867] & layer1_out[868]);
     layer2_out[642] <= layer1_out[1439] | layer1_out[1440];
     layer2_out[643] <= 1'b0;
     layer2_out[644] <= 1'b1;
     layer2_out[645] <= 1'b1;
     layer2_out[646] <= layer1_out[789] | layer1_out[790];
     layer2_out[647] <= ~(layer1_out[1167] | layer1_out[1168]);
     layer2_out[648] <= layer1_out[576] & ~layer1_out[575];
     layer2_out[649] <= ~(layer1_out[949] & layer1_out[950]);
     layer2_out[650] <= ~(layer1_out[127] | layer1_out[128]);
     layer2_out[651] <= ~layer1_out[761];
     layer2_out[652] <= ~(layer1_out[1254] | layer1_out[1255]);
     layer2_out[653] <= ~(layer1_out[709] & layer1_out[710]);
     layer2_out[654] <= layer1_out[86] & ~layer1_out[85];
     layer2_out[655] <= 1'b1;
     layer2_out[656] <= layer1_out[1057] & ~layer1_out[1058];
     layer2_out[657] <= layer1_out[962] & layer1_out[963];
     layer2_out[658] <= ~(layer1_out[1169] & layer1_out[1170]);
     layer2_out[659] <= layer1_out[105] & layer1_out[106];
     layer2_out[660] <= ~layer1_out[449];
     layer2_out[661] <= ~(layer1_out[14] | layer1_out[15]);
     layer2_out[662] <= ~layer1_out[671];
     layer2_out[663] <= 1'b0;
     layer2_out[664] <= 1'b0;
     layer2_out[665] <= layer1_out[1387];
     layer2_out[666] <= ~(layer1_out[1492] | layer1_out[1493]);
     layer2_out[667] <= ~layer1_out[725] | layer1_out[724];
     layer2_out[668] <= ~layer1_out[1217];
     layer2_out[669] <= layer1_out[622] & layer1_out[623];
     layer2_out[670] <= 1'b0;
     layer2_out[671] <= ~layer1_out[278] | layer1_out[277];
     layer2_out[672] <= ~(layer1_out[1158] & layer1_out[1159]);
     layer2_out[673] <= 1'b0;
     layer2_out[674] <= layer1_out[1120] & ~layer1_out[1121];
     layer2_out[675] <= ~(layer1_out[912] & layer1_out[913]);
     layer2_out[676] <= ~layer1_out[1230] | layer1_out[1231];
     layer2_out[677] <= 1'b1;
     layer2_out[678] <= ~(layer1_out[1381] & layer1_out[1382]);
     layer2_out[679] <= ~layer1_out[1160] | layer1_out[1159];
     layer2_out[680] <= 1'b1;
     layer2_out[681] <= ~layer1_out[602];
     layer2_out[682] <= 1'b1;
     layer2_out[683] <= 1'b0;
     layer2_out[684] <= ~layer1_out[55] | layer1_out[54];
     layer2_out[685] <= layer1_out[958];
     layer2_out[686] <= layer1_out[836];
     layer2_out[687] <= 1'b0;
     layer2_out[688] <= ~(layer1_out[1333] & layer1_out[1334]);
     layer2_out[689] <= layer1_out[195] & layer1_out[196];
     layer2_out[690] <= ~layer1_out[716];
     layer2_out[691] <= ~(layer1_out[119] | layer1_out[120]);
     layer2_out[692] <= ~layer1_out[1263];
     layer2_out[693] <= ~layer1_out[539] | layer1_out[538];
     layer2_out[694] <= ~layer1_out[471];
     layer2_out[695] <= layer1_out[1041];
     layer2_out[696] <= 1'b0;
     layer2_out[697] <= layer1_out[706];
     layer2_out[698] <= layer1_out[929];
     layer2_out[699] <= layer1_out[645];
     layer2_out[700] <= ~layer1_out[667];
     layer2_out[701] <= ~layer1_out[905] | layer1_out[904];
     layer2_out[702] <= ~(layer1_out[349] | layer1_out[350]);
     layer2_out[703] <= 1'b0;
     layer2_out[704] <= ~layer1_out[1206];
     layer2_out[705] <= layer1_out[924];
     layer2_out[706] <= layer1_out[1233] & ~layer1_out[1232];
     layer2_out[707] <= 1'b1;
     layer2_out[708] <= layer1_out[843] & layer1_out[844];
     layer2_out[709] <= layer1_out[447];
     layer2_out[710] <= layer1_out[1116] & ~layer1_out[1117];
     layer2_out[711] <= ~layer1_out[893];
     layer2_out[712] <= layer1_out[1210] & ~layer1_out[1209];
     layer2_out[713] <= layer1_out[421] & ~layer1_out[420];
     layer2_out[714] <= layer1_out[1170];
     layer2_out[715] <= ~(layer1_out[814] & layer1_out[815]);
     layer2_out[716] <= 1'b1;
     layer2_out[717] <= layer1_out[1260] | layer1_out[1261];
     layer2_out[718] <= ~layer1_out[987];
     layer2_out[719] <= ~(layer1_out[778] | layer1_out[779]);
     layer2_out[720] <= layer1_out[1326];
     layer2_out[721] <= ~(layer1_out[861] & layer1_out[862]);
     layer2_out[722] <= ~layer1_out[1387];
     layer2_out[723] <= ~(layer1_out[672] & layer1_out[673]);
     layer2_out[724] <= ~layer1_out[1074];
     layer2_out[725] <= ~(layer1_out[811] ^ layer1_out[812]);
     layer2_out[726] <= layer1_out[1385] | layer1_out[1386];
     layer2_out[727] <= ~(layer1_out[791] & layer1_out[792]);
     layer2_out[728] <= ~(layer1_out[584] | layer1_out[585]);
     layer2_out[729] <= 1'b0;
     layer2_out[730] <= 1'b1;
     layer2_out[731] <= ~(layer1_out[462] & layer1_out[463]);
     layer2_out[732] <= ~layer1_out[1429] | layer1_out[1428];
     layer2_out[733] <= ~layer1_out[610] | layer1_out[611];
     layer2_out[734] <= layer1_out[1244] | layer1_out[1245];
     layer2_out[735] <= layer1_out[193] & ~layer1_out[192];
     layer2_out[736] <= layer1_out[19];
     layer2_out[737] <= ~(layer1_out[619] | layer1_out[620]);
     layer2_out[738] <= layer1_out[756];
     layer2_out[739] <= layer1_out[1210] | layer1_out[1211];
     layer2_out[740] <= 1'b0;
     layer2_out[741] <= ~layer1_out[531] | layer1_out[532];
     layer2_out[742] <= 1'b0;
     layer2_out[743] <= ~layer1_out[1141];
     layer2_out[744] <= 1'b0;
     layer2_out[745] <= 1'b1;
     layer2_out[746] <= layer1_out[373] & ~layer1_out[372];
     layer2_out[747] <= layer1_out[1154] & layer1_out[1155];
     layer2_out[748] <= ~layer1_out[87];
     layer2_out[749] <= layer1_out[1272] | layer1_out[1273];
     layer2_out[750] <= layer1_out[1132] & layer1_out[1133];
     layer2_out[751] <= layer1_out[319] & ~layer1_out[318];
     layer2_out[752] <= ~layer1_out[1081];
     layer2_out[753] <= layer1_out[1260] & ~layer1_out[1259];
     layer2_out[754] <= layer1_out[432] ^ layer1_out[433];
     layer2_out[755] <= layer1_out[444] & ~layer1_out[445];
     layer2_out[756] <= ~layer1_out[470];
     layer2_out[757] <= layer1_out[920] & ~layer1_out[921];
     layer2_out[758] <= layer1_out[751];
     layer2_out[759] <= layer1_out[433] | layer1_out[434];
     layer2_out[760] <= ~(layer1_out[1247] & layer1_out[1248]);
     layer2_out[761] <= ~layer1_out[752] | layer1_out[751];
     layer2_out[762] <= 1'b1;
     layer2_out[763] <= layer1_out[325] & ~layer1_out[324];
     layer2_out[764] <= ~(layer1_out[797] | layer1_out[798]);
     layer2_out[765] <= layer1_out[557] & ~layer1_out[558];
     layer2_out[766] <= ~layer1_out[991] | layer1_out[990];
     layer2_out[767] <= ~(layer1_out[343] | layer1_out[344]);
     layer2_out[768] <= layer1_out[457] | layer1_out[458];
     layer2_out[769] <= layer1_out[1328];
     layer2_out[770] <= layer1_out[303];
     layer2_out[771] <= 1'b1;
     layer2_out[772] <= 1'b0;
     layer2_out[773] <= 1'b1;
     layer2_out[774] <= layer1_out[435] & layer1_out[436];
     layer2_out[775] <= ~(layer1_out[301] | layer1_out[302]);
     layer2_out[776] <= ~layer1_out[19];
     layer2_out[777] <= layer1_out[1385];
     layer2_out[778] <= ~layer1_out[209] | layer1_out[208];
     layer2_out[779] <= ~(layer1_out[524] & layer1_out[525]);
     layer2_out[780] <= 1'b0;
     layer2_out[781] <= 1'b0;
     layer2_out[782] <= ~layer1_out[1013] | layer1_out[1012];
     layer2_out[783] <= ~(layer1_out[391] & layer1_out[392]);
     layer2_out[784] <= ~(layer1_out[1390] & layer1_out[1391]);
     layer2_out[785] <= layer1_out[857] & layer1_out[858];
     layer2_out[786] <= ~(layer1_out[377] ^ layer1_out[378]);
     layer2_out[787] <= 1'b0;
     layer2_out[788] <= layer1_out[1118];
     layer2_out[789] <= layer1_out[933] & ~layer1_out[932];
     layer2_out[790] <= layer1_out[1238] & ~layer1_out[1239];
     layer2_out[791] <= 1'b1;
     layer2_out[792] <= ~layer1_out[709] | layer1_out[708];
     layer2_out[793] <= ~layer1_out[330];
     layer2_out[794] <= ~(layer1_out[1340] | layer1_out[1341]);
     layer2_out[795] <= layer1_out[533] & ~layer1_out[534];
     layer2_out[796] <= ~(layer1_out[1039] | layer1_out[1040]);
     layer2_out[797] <= layer1_out[1319] & layer1_out[1320];
     layer2_out[798] <= layer1_out[1138];
     layer2_out[799] <= layer1_out[447] & ~layer1_out[448];
     layer2_out[800] <= layer1_out[230] | layer1_out[231];
     layer2_out[801] <= ~layer1_out[77] | layer1_out[76];
     layer2_out[802] <= ~layer1_out[441] | layer1_out[440];
     layer2_out[803] <= ~layer1_out[820];
     layer2_out[804] <= layer1_out[1166] & ~layer1_out[1165];
     layer2_out[805] <= layer1_out[1343] & layer1_out[1344];
     layer2_out[806] <= 1'b1;
     layer2_out[807] <= ~(layer1_out[805] | layer1_out[806]);
     layer2_out[808] <= ~(layer1_out[437] | layer1_out[438]);
     layer2_out[809] <= 1'b1;
     layer2_out[810] <= layer1_out[1106] | layer1_out[1107];
     layer2_out[811] <= layer1_out[927] & ~layer1_out[928];
     layer2_out[812] <= 1'b0;
     layer2_out[813] <= ~layer1_out[1028];
     layer2_out[814] <= layer1_out[1141] & layer1_out[1142];
     layer2_out[815] <= ~(layer1_out[1005] & layer1_out[1006]);
     layer2_out[816] <= layer1_out[1410];
     layer2_out[817] <= layer1_out[578] | layer1_out[579];
     layer2_out[818] <= layer1_out[274] & layer1_out[275];
     layer2_out[819] <= layer1_out[780] | layer1_out[781];
     layer2_out[820] <= layer1_out[921] & ~layer1_out[922];
     layer2_out[821] <= layer1_out[711] | layer1_out[712];
     layer2_out[822] <= ~layer1_out[1168];
     layer2_out[823] <= ~(layer1_out[944] | layer1_out[945]);
     layer2_out[824] <= layer1_out[1088];
     layer2_out[825] <= ~layer1_out[1290];
     layer2_out[826] <= layer1_out[964] | layer1_out[965];
     layer2_out[827] <= layer1_out[1415] & ~layer1_out[1414];
     layer2_out[828] <= layer1_out[317] & ~layer1_out[318];
     layer2_out[829] <= ~(layer1_out[907] & layer1_out[908]);
     layer2_out[830] <= layer1_out[137];
     layer2_out[831] <= layer1_out[222] & layer1_out[223];
     layer2_out[832] <= 1'b0;
     layer2_out[833] <= ~(layer1_out[968] & layer1_out[969]);
     layer2_out[834] <= layer1_out[275] | layer1_out[276];
     layer2_out[835] <= layer1_out[994];
     layer2_out[836] <= ~(layer1_out[637] | layer1_out[638]);
     layer2_out[837] <= ~(layer1_out[473] & layer1_out[474]);
     layer2_out[838] <= ~(layer1_out[785] & layer1_out[786]);
     layer2_out[839] <= layer1_out[1192];
     layer2_out[840] <= 1'b0;
     layer2_out[841] <= 1'b1;
     layer2_out[842] <= 1'b0;
     layer2_out[843] <= 1'b0;
     layer2_out[844] <= ~layer1_out[764];
     layer2_out[845] <= 1'b1;
     layer2_out[846] <= 1'b1;
     layer2_out[847] <= ~(layer1_out[266] & layer1_out[267]);
     layer2_out[848] <= 1'b0;
     layer2_out[849] <= ~layer1_out[1177];
     layer2_out[850] <= ~(layer1_out[770] & layer1_out[771]);
     layer2_out[851] <= 1'b0;
     layer2_out[852] <= 1'b1;
     layer2_out[853] <= layer1_out[950] & ~layer1_out[951];
     layer2_out[854] <= 1'b0;
     layer2_out[855] <= layer1_out[131] | layer1_out[132];
     layer2_out[856] <= 1'b1;
     layer2_out[857] <= layer1_out[772];
     layer2_out[858] <= 1'b1;
     layer2_out[859] <= layer1_out[1150];
     layer2_out[860] <= layer1_out[726];
     layer2_out[861] <= ~(layer1_out[910] ^ layer1_out[911]);
     layer2_out[862] <= layer1_out[1058] ^ layer1_out[1059];
     layer2_out[863] <= layer1_out[549] & ~layer1_out[548];
     layer2_out[864] <= ~(layer1_out[597] | layer1_out[598]);
     layer2_out[865] <= ~layer1_out[1095] | layer1_out[1094];
     layer2_out[866] <= ~layer1_out[436];
     layer2_out[867] <= ~layer1_out[207] | layer1_out[208];
     layer2_out[868] <= 1'b0;
     layer2_out[869] <= ~layer1_out[11] | layer1_out[10];
     layer2_out[870] <= 1'b0;
     layer2_out[871] <= layer1_out[398];
     layer2_out[872] <= layer1_out[315] & layer1_out[316];
     layer2_out[873] <= ~(layer1_out[1275] & layer1_out[1276]);
     layer2_out[874] <= layer1_out[638] | layer1_out[639];
     layer2_out[875] <= ~layer1_out[1411] | layer1_out[1410];
     layer2_out[876] <= ~layer1_out[1188] | layer1_out[1189];
     layer2_out[877] <= ~layer1_out[347] | layer1_out[346];
     layer2_out[878] <= ~layer1_out[1270];
     layer2_out[879] <= ~(layer1_out[306] ^ layer1_out[307]);
     layer2_out[880] <= ~layer1_out[287] | layer1_out[288];
     layer2_out[881] <= ~layer1_out[1236] | layer1_out[1235];
     layer2_out[882] <= ~layer1_out[975] | layer1_out[976];
     layer2_out[883] <= ~layer1_out[803];
     layer2_out[884] <= layer1_out[1208];
     layer2_out[885] <= layer1_out[942] & layer1_out[943];
     layer2_out[886] <= ~layer1_out[226] | layer1_out[225];
     layer2_out[887] <= layer1_out[381] & ~layer1_out[382];
     layer2_out[888] <= layer1_out[1224] & ~layer1_out[1225];
     layer2_out[889] <= layer1_out[849] & ~layer1_out[848];
     layer2_out[890] <= ~layer1_out[1371] | layer1_out[1372];
     layer2_out[891] <= layer1_out[897] | layer1_out[898];
     layer2_out[892] <= 1'b1;
     layer2_out[893] <= 1'b0;
     layer2_out[894] <= 1'b0;
     layer2_out[895] <= layer1_out[490] & ~layer1_out[489];
     layer2_out[896] <= ~layer1_out[73];
     layer2_out[897] <= 1'b0;
     layer2_out[898] <= layer1_out[826] & ~layer1_out[827];
     layer2_out[899] <= ~layer1_out[894];
     layer2_out[900] <= ~(layer1_out[1315] & layer1_out[1316]);
     layer2_out[901] <= layer1_out[9] & ~layer1_out[8];
     layer2_out[902] <= 1'b1;
     layer2_out[903] <= layer1_out[263] & ~layer1_out[262];
     layer2_out[904] <= layer1_out[1275] & ~layer1_out[1274];
     layer2_out[905] <= layer1_out[9] & ~layer1_out[10];
     layer2_out[906] <= ~layer1_out[408];
     layer2_out[907] <= ~(layer1_out[108] & layer1_out[109]);
     layer2_out[908] <= ~layer1_out[34];
     layer2_out[909] <= 1'b0;
     layer2_out[910] <= layer1_out[517] & layer1_out[518];
     layer2_out[911] <= layer1_out[451] & ~layer1_out[452];
     layer2_out[912] <= layer1_out[1035] & layer1_out[1036];
     layer2_out[913] <= layer1_out[81] & ~layer1_out[80];
     layer2_out[914] <= ~layer1_out[1283] | layer1_out[1282];
     layer2_out[915] <= layer1_out[267] & ~layer1_out[268];
     layer2_out[916] <= layer1_out[1203];
     layer2_out[917] <= layer1_out[650] | layer1_out[651];
     layer2_out[918] <= ~layer1_out[811] | layer1_out[810];
     layer2_out[919] <= layer1_out[981] & layer1_out[982];
     layer2_out[920] <= layer1_out[425] & layer1_out[426];
     layer2_out[921] <= layer1_out[1409] & ~layer1_out[1408];
     layer2_out[922] <= layer1_out[1302] & layer1_out[1303];
     layer2_out[923] <= ~(layer1_out[88] | layer1_out[89]);
     layer2_out[924] <= 1'b1;
     layer2_out[925] <= ~layer1_out[1240] | layer1_out[1241];
     layer2_out[926] <= ~(layer1_out[1454] | layer1_out[1455]);
     layer2_out[927] <= layer1_out[1290];
     layer2_out[928] <= 1'b1;
     layer2_out[929] <= 1'b0;
     layer2_out[930] <= ~layer1_out[872];
     layer2_out[931] <= 1'b0;
     layer2_out[932] <= ~layer1_out[87] | layer1_out[86];
     layer2_out[933] <= ~layer1_out[239];
     layer2_out[934] <= 1'b0;
     layer2_out[935] <= layer1_out[1051] & ~layer1_out[1050];
     layer2_out[936] <= layer1_out[996] & ~layer1_out[997];
     layer2_out[937] <= layer1_out[798] | layer1_out[799];
     layer2_out[938] <= ~layer1_out[1187];
     layer2_out[939] <= ~(layer1_out[1445] & layer1_out[1446]);
     layer2_out[940] <= ~(layer1_out[1025] & layer1_out[1026]);
     layer2_out[941] <= ~layer1_out[1328];
     layer2_out[942] <= layer1_out[862] | layer1_out[863];
     layer2_out[943] <= ~(layer1_out[209] | layer1_out[210]);
     layer2_out[944] <= layer1_out[389];
     layer2_out[945] <= ~(layer1_out[1077] & layer1_out[1078]);
     layer2_out[946] <= 1'b0;
     layer2_out[947] <= ~(layer1_out[155] ^ layer1_out[156]);
     layer2_out[948] <= 1'b0;
     layer2_out[949] <= ~layer1_out[505] | layer1_out[504];
     layer2_out[950] <= ~(layer1_out[829] | layer1_out[830]);
     layer2_out[951] <= layer1_out[443] ^ layer1_out[444];
     layer2_out[952] <= layer1_out[594] & layer1_out[595];
     layer2_out[953] <= layer1_out[760] & ~layer1_out[759];
     layer2_out[954] <= layer1_out[688] & layer1_out[689];
     layer2_out[955] <= layer1_out[775] | layer1_out[776];
     layer2_out[956] <= ~layer1_out[1234] | layer1_out[1233];
     layer2_out[957] <= ~layer1_out[509] | layer1_out[508];
     layer2_out[958] <= layer1_out[565] & layer1_out[566];
     layer2_out[959] <= layer1_out[467] & ~layer1_out[466];
     layer2_out[960] <= layer1_out[177] & ~layer1_out[176];
     layer2_out[961] <= layer1_out[1437];
     layer2_out[962] <= layer1_out[1071];
     layer2_out[963] <= ~layer1_out[882];
     layer2_out[964] <= layer1_out[285] & ~layer1_out[286];
     layer2_out[965] <= ~layer1_out[590] | layer1_out[589];
     layer2_out[966] <= 1'b1;
     layer2_out[967] <= ~layer1_out[789] | layer1_out[788];
     layer2_out[968] <= layer1_out[820] & ~layer1_out[819];
     layer2_out[969] <= ~(layer1_out[74] | layer1_out[75]);
     layer2_out[970] <= layer1_out[1011];
     layer2_out[971] <= layer1_out[395];
     layer2_out[972] <= ~(layer1_out[1226] | layer1_out[1227]);
     layer2_out[973] <= ~layer1_out[1127] | layer1_out[1126];
     layer2_out[974] <= 1'b1;
     layer2_out[975] <= layer1_out[503] & ~layer1_out[502];
     layer2_out[976] <= 1'b0;
     layer2_out[977] <= layer1_out[326];
     layer2_out[978] <= ~layer1_out[940];
     layer2_out[979] <= ~layer1_out[863] | layer1_out[864];
     layer2_out[980] <= ~(layer1_out[332] | layer1_out[333]);
     layer2_out[981] <= layer1_out[411] & ~layer1_out[412];
     layer2_out[982] <= layer1_out[291] | layer1_out[292];
     layer2_out[983] <= layer1_out[265] & layer1_out[266];
     layer2_out[984] <= 1'b1;
     layer2_out[985] <= layer1_out[1189] | layer1_out[1190];
     layer2_out[986] <= layer1_out[1442] & layer1_out[1443];
     layer2_out[987] <= ~layer1_out[710] | layer1_out[711];
     layer2_out[988] <= ~layer1_out[353] | layer1_out[354];
     layer2_out[989] <= layer1_out[782] & ~layer1_out[781];
     layer2_out[990] <= 1'b1;
     layer2_out[991] <= layer1_out[547] & layer1_out[548];
     layer2_out[992] <= ~layer1_out[640];
     layer2_out[993] <= layer1_out[264];
     layer2_out[994] <= ~layer1_out[1479] | layer1_out[1478];
     layer2_out[995] <= ~(layer1_out[1160] & layer1_out[1161]);
     layer2_out[996] <= ~(layer1_out[96] | layer1_out[97]);
     layer2_out[997] <= 1'b1;
     layer2_out[998] <= ~(layer1_out[1291] & layer1_out[1292]);
     layer2_out[999] <= layer1_out[730];
     layer2_out[1000] <= ~(layer1_out[1280] & layer1_out[1281]);
     layer2_out[1001] <= layer1_out[102];
     layer2_out[1002] <= layer1_out[588] & ~layer1_out[587];
     layer2_out[1003] <= ~(layer1_out[807] & layer1_out[808]);
     layer2_out[1004] <= 1'b1;
     layer2_out[1005] <= ~(layer1_out[539] | layer1_out[540]);
     layer2_out[1006] <= layer1_out[216] | layer1_out[217];
     layer2_out[1007] <= ~layer1_out[592];
     layer2_out[1008] <= layer1_out[57] | layer1_out[58];
     layer2_out[1009] <= ~layer1_out[432];
     layer2_out[1010] <= layer1_out[854];
     layer2_out[1011] <= 1'b0;
     layer2_out[1012] <= ~(layer1_out[1212] | layer1_out[1213]);
     layer2_out[1013] <= layer1_out[516];
     layer2_out[1014] <= ~(layer1_out[1349] & layer1_out[1350]);
     layer2_out[1015] <= 1'b1;
     layer2_out[1016] <= ~layer1_out[1172] | layer1_out[1171];
     layer2_out[1017] <= ~(layer1_out[685] & layer1_out[686]);
     layer2_out[1018] <= 1'b1;
     layer2_out[1019] <= layer1_out[335];
     layer2_out[1020] <= layer1_out[1305] & layer1_out[1306];
     layer2_out[1021] <= ~layer1_out[253] | layer1_out[254];
     layer2_out[1022] <= layer1_out[806] & layer1_out[807];
     layer2_out[1023] <= ~(layer1_out[546] | layer1_out[547]);
     layer2_out[1024] <= layer1_out[563] & ~layer1_out[564];
     layer2_out[1025] <= layer1_out[1483] & ~layer1_out[1482];
     layer2_out[1026] <= ~(layer1_out[675] & layer1_out[676]);
     layer2_out[1027] <= 1'b1;
     layer2_out[1028] <= layer1_out[373] & layer1_out[374];
     layer2_out[1029] <= ~layer1_out[1322];
     layer2_out[1030] <= 1'b0;
     layer2_out[1031] <= layer1_out[69] & layer1_out[70];
     layer2_out[1032] <= layer1_out[736] & layer1_out[737];
     layer2_out[1033] <= ~(layer1_out[417] | layer1_out[418]);
     layer2_out[1034] <= layer1_out[1433];
     layer2_out[1035] <= ~(layer1_out[859] | layer1_out[860]);
     layer2_out[1036] <= ~layer1_out[884];
     layer2_out[1037] <= 1'b0;
     layer2_out[1038] <= ~(layer1_out[1325] & layer1_out[1326]);
     layer2_out[1039] <= layer1_out[1366] & layer1_out[1367];
     layer2_out[1040] <= layer1_out[973] | layer1_out[974];
     layer2_out[1041] <= layer1_out[1061] & ~layer1_out[1060];
     layer2_out[1042] <= ~layer1_out[483] | layer1_out[484];
     layer2_out[1043] <= ~(layer1_out[776] | layer1_out[777]);
     layer2_out[1044] <= 1'b1;
     layer2_out[1045] <= layer1_out[1430];
     layer2_out[1046] <= 1'b1;
     layer2_out[1047] <= ~layer1_out[1476] | layer1_out[1477];
     layer2_out[1048] <= layer1_out[1053];
     layer2_out[1049] <= layer1_out[1360] | layer1_out[1361];
     layer2_out[1050] <= ~layer1_out[1097];
     layer2_out[1051] <= ~layer1_out[1113];
     layer2_out[1052] <= layer1_out[476] & layer1_out[477];
     layer2_out[1053] <= layer1_out[364];
     layer2_out[1054] <= ~layer1_out[353] | layer1_out[352];
     layer2_out[1055] <= layer1_out[647] & ~layer1_out[646];
     layer2_out[1056] <= layer1_out[733] & ~layer1_out[732];
     layer2_out[1057] <= ~layer1_out[1354];
     layer2_out[1058] <= ~layer1_out[133] | layer1_out[132];
     layer2_out[1059] <= layer1_out[1112];
     layer2_out[1060] <= ~(layer1_out[742] | layer1_out[743]);
     layer2_out[1061] <= ~(layer1_out[665] & layer1_out[666]);
     layer2_out[1062] <= layer1_out[300] | layer1_out[301];
     layer2_out[1063] <= ~(layer1_out[1216] | layer1_out[1217]);
     layer2_out[1064] <= ~layer1_out[190] | layer1_out[191];
     layer2_out[1065] <= layer1_out[1444] & layer1_out[1445];
     layer2_out[1066] <= layer1_out[1281] & layer1_out[1282];
     layer2_out[1067] <= layer1_out[422] | layer1_out[423];
     layer2_out[1068] <= ~(layer1_out[1047] & layer1_out[1048]);
     layer2_out[1069] <= layer1_out[93];
     layer2_out[1070] <= ~layer1_out[944];
     layer2_out[1071] <= 1'b1;
     layer2_out[1072] <= layer1_out[746] & ~layer1_out[745];
     layer2_out[1073] <= layer1_out[122] & ~layer1_out[121];
     layer2_out[1074] <= layer1_out[461] & layer1_out[462];
     layer2_out[1075] <= 1'b1;
     layer2_out[1076] <= ~(layer1_out[510] | layer1_out[511]);
     layer2_out[1077] <= layer1_out[607] & layer1_out[608];
     layer2_out[1078] <= ~layer1_out[27] | layer1_out[26];
     layer2_out[1079] <= 1'b1;
     layer2_out[1080] <= layer1_out[754] | layer1_out[755];
     layer2_out[1081] <= layer1_out[660];
     layer2_out[1082] <= 1'b1;
     layer2_out[1083] <= 1'b1;
     layer2_out[1084] <= layer1_out[295] & ~layer1_out[296];
     layer2_out[1085] <= ~(layer1_out[239] & layer1_out[240]);
     layer2_out[1086] <= layer1_out[485];
     layer2_out[1087] <= ~(layer1_out[1469] | layer1_out[1470]);
     layer2_out[1088] <= layer1_out[749] & ~layer1_out[750];
     layer2_out[1089] <= ~(layer1_out[477] | layer1_out[478]);
     layer2_out[1090] <= ~layer1_out[1297];
     layer2_out[1091] <= ~layer1_out[1162];
     layer2_out[1092] <= 1'b1;
     layer2_out[1093] <= ~layer1_out[91];
     layer2_out[1094] <= layer1_out[205] & layer1_out[206];
     layer2_out[1095] <= layer1_out[821] | layer1_out[822];
     layer2_out[1096] <= 1'b1;
     layer2_out[1097] <= ~layer1_out[1164] | layer1_out[1165];
     layer2_out[1098] <= 1'b0;
     layer2_out[1099] <= ~layer1_out[486];
     layer2_out[1100] <= 1'b0;
     layer2_out[1101] <= 1'b1;
     layer2_out[1102] <= layer1_out[842] & ~layer1_out[843];
     layer2_out[1103] <= ~(layer1_out[999] | layer1_out[1000]);
     layer2_out[1104] <= layer1_out[95] & ~layer1_out[94];
     layer2_out[1105] <= layer1_out[636] | layer1_out[637];
     layer2_out[1106] <= layer1_out[1488];
     layer2_out[1107] <= 1'b0;
     layer2_out[1108] <= ~(layer1_out[1404] & layer1_out[1405]);
     layer2_out[1109] <= 1'b0;
     layer2_out[1110] <= ~layer1_out[77];
     layer2_out[1111] <= 1'b0;
     layer2_out[1112] <= ~layer1_out[215];
     layer2_out[1113] <= layer1_out[479] & ~layer1_out[478];
     layer2_out[1114] <= layer1_out[1142] & ~layer1_out[1143];
     layer2_out[1115] <= layer1_out[499] | layer1_out[500];
     layer2_out[1116] <= ~layer1_out[224];
     layer2_out[1117] <= layer1_out[272] & layer1_out[273];
     layer2_out[1118] <= 1'b1;
     layer2_out[1119] <= layer1_out[70] & layer1_out[71];
     layer2_out[1120] <= ~layer1_out[45];
     layer2_out[1121] <= 1'b1;
     layer2_out[1122] <= layer1_out[15] & ~layer1_out[16];
     layer2_out[1123] <= 1'b0;
     layer2_out[1124] <= 1'b0;
     layer2_out[1125] <= layer1_out[290];
     layer2_out[1126] <= ~(layer1_out[931] | layer1_out[932]);
     layer2_out[1127] <= ~layer1_out[438];
     layer2_out[1128] <= ~(layer1_out[794] | layer1_out[795]);
     layer2_out[1129] <= ~layer1_out[1299];
     layer2_out[1130] <= ~(layer1_out[1110] | layer1_out[1111]);
     layer2_out[1131] <= layer1_out[405] & ~layer1_out[406];
     layer2_out[1132] <= layer1_out[630] & ~layer1_out[629];
     layer2_out[1133] <= 1'b1;
     layer2_out[1134] <= ~layer1_out[740] | layer1_out[739];
     layer2_out[1135] <= layer1_out[1128] & layer1_out[1129];
     layer2_out[1136] <= ~layer1_out[1195];
     layer2_out[1137] <= layer1_out[335] & ~layer1_out[334];
     layer2_out[1138] <= layer1_out[911] & layer1_out[912];
     layer2_out[1139] <= layer1_out[571];
     layer2_out[1140] <= layer1_out[1022];
     layer2_out[1141] <= layer1_out[941] & ~layer1_out[942];
     layer2_out[1142] <= layer1_out[920] & ~layer1_out[919];
     layer2_out[1143] <= layer1_out[533] & ~layer1_out[532];
     layer2_out[1144] <= layer1_out[270] | layer1_out[271];
     layer2_out[1145] <= 1'b1;
     layer2_out[1146] <= 1'b1;
     layer2_out[1147] <= ~layer1_out[980] | layer1_out[979];
     layer2_out[1148] <= 1'b1;
     layer2_out[1149] <= ~layer1_out[5];
     layer2_out[1150] <= 1'b0;
     layer2_out[1151] <= ~(layer1_out[201] & layer1_out[202]);
     layer2_out[1152] <= ~(layer1_out[1172] ^ layer1_out[1173]);
     layer2_out[1153] <= ~(layer1_out[526] & layer1_out[527]);
     layer2_out[1154] <= layer1_out[503];
     layer2_out[1155] <= layer1_out[1085];
     layer2_out[1156] <= ~(layer1_out[1082] | layer1_out[1083]);
     layer2_out[1157] <= 1'b1;
     layer2_out[1158] <= 1'b0;
     layer2_out[1159] <= ~layer1_out[404] | layer1_out[405];
     layer2_out[1160] <= layer1_out[493] & ~layer1_out[494];
     layer2_out[1161] <= ~layer1_out[1246] | layer1_out[1247];
     layer2_out[1162] <= 1'b1;
     layer2_out[1163] <= layer1_out[1042];
     layer2_out[1164] <= ~layer1_out[801];
     layer2_out[1165] <= 1'b1;
     layer2_out[1166] <= layer1_out[260] & ~layer1_out[261];
     layer2_out[1167] <= ~(layer1_out[718] | layer1_out[719]);
     layer2_out[1168] <= layer1_out[116] | layer1_out[117];
     layer2_out[1169] <= ~layer1_out[378];
     layer2_out[1170] <= ~(layer1_out[124] | layer1_out[125]);
     layer2_out[1171] <= layer1_out[1417] & ~layer1_out[1416];
     layer2_out[1172] <= ~(layer1_out[328] & layer1_out[329]);
     layer2_out[1173] <= layer1_out[345] & layer1_out[346];
     layer2_out[1174] <= ~layer1_out[364];
     layer2_out[1175] <= layer1_out[1144] & layer1_out[1145];
     layer2_out[1176] <= layer1_out[1037] & ~layer1_out[1036];
     layer2_out[1177] <= layer1_out[1198] & layer1_out[1199];
     layer2_out[1178] <= ~layer1_out[135] | layer1_out[136];
     layer2_out[1179] <= ~(layer1_out[316] & layer1_out[317]);
     layer2_out[1180] <= ~layer1_out[612] | layer1_out[613];
     layer2_out[1181] <= 1'b1;
     layer2_out[1182] <= ~(layer1_out[872] & layer1_out[873]);
     layer2_out[1183] <= 1'b0;
     layer2_out[1184] <= ~layer1_out[1049];
     layer2_out[1185] <= ~(layer1_out[1185] | layer1_out[1186]);
     layer2_out[1186] <= ~layer1_out[964] | layer1_out[963];
     layer2_out[1187] <= layer1_out[886];
     layer2_out[1188] <= 1'b1;
     layer2_out[1189] <= 1'b0;
     layer2_out[1190] <= layer1_out[740] & ~layer1_out[741];
     layer2_out[1191] <= layer1_out[1391] | layer1_out[1392];
     layer2_out[1192] <= 1'b1;
     layer2_out[1193] <= ~(layer1_out[530] & layer1_out[531]);
     layer2_out[1194] <= 1'b0;
     layer2_out[1195] <= 1'b0;
     layer2_out[1196] <= 1'b0;
     layer2_out[1197] <= ~(layer1_out[154] | layer1_out[155]);
     layer2_out[1198] <= layer1_out[712] | layer1_out[713];
     layer2_out[1199] <= 1'b0;
     layer2_out[1200] <= layer1_out[380] & ~layer1_out[379];
     layer2_out[1201] <= ~layer1_out[1393];
     layer2_out[1202] <= layer1_out[117] & ~layer1_out[118];
     layer2_out[1203] <= layer1_out[1249];
     layer2_out[1204] <= layer1_out[838];
     layer2_out[1205] <= layer1_out[1154] & ~layer1_out[1153];
     layer2_out[1206] <= layer1_out[355];
     layer2_out[1207] <= layer1_out[1034];
     layer2_out[1208] <= ~layer1_out[1426];
     layer2_out[1209] <= 1'b1;
     layer2_out[1210] <= 1'b0;
     layer2_out[1211] <= ~layer1_out[529] | layer1_out[528];
     layer2_out[1212] <= 1'b1;
     layer2_out[1213] <= layer1_out[1090] | layer1_out[1091];
     layer2_out[1214] <= layer1_out[279] & ~layer1_out[278];
     layer2_out[1215] <= ~(layer1_out[495] & layer1_out[496]);
     layer2_out[1216] <= ~layer1_out[1380] | layer1_out[1381];
     layer2_out[1217] <= layer1_out[1097] & ~layer1_out[1098];
     layer2_out[1218] <= 1'b1;
     layer2_out[1219] <= ~layer1_out[481];
     layer2_out[1220] <= layer1_out[1092] & ~layer1_out[1093];
     layer2_out[1221] <= ~layer1_out[831];
     layer2_out[1222] <= layer1_out[150] & ~layer1_out[151];
     layer2_out[1223] <= 1'b1;
     layer2_out[1224] <= 1'b0;
     layer2_out[1225] <= 1'b0;
     layer2_out[1226] <= 1'b0;
     layer2_out[1227] <= layer1_out[1403] & layer1_out[1404];
     layer2_out[1228] <= ~layer1_out[47] | layer1_out[48];
     layer2_out[1229] <= layer1_out[582] & ~layer1_out[581];
     layer2_out[1230] <= layer1_out[1471] & ~layer1_out[1472];
     layer2_out[1231] <= ~(layer1_out[82] | layer1_out[83]);
     layer2_out[1232] <= ~layer1_out[987] | layer1_out[988];
     layer2_out[1233] <= ~layer1_out[40] | layer1_out[39];
     layer2_out[1234] <= layer1_out[1078] | layer1_out[1079];
     layer2_out[1235] <= layer1_out[1466] & ~layer1_out[1467];
     layer2_out[1236] <= layer1_out[600] | layer1_out[601];
     layer2_out[1237] <= layer1_out[1109] | layer1_out[1110];
     layer2_out[1238] <= 1'b0;
     layer2_out[1239] <= 1'b0;
     layer2_out[1240] <= ~layer1_out[567] | layer1_out[566];
     layer2_out[1241] <= layer1_out[664] | layer1_out[665];
     layer2_out[1242] <= layer1_out[569] & ~layer1_out[568];
     layer2_out[1243] <= ~(layer1_out[416] | layer1_out[417]);
     layer2_out[1244] <= ~(layer1_out[390] & layer1_out[391]);
     layer2_out[1245] <= ~layer1_out[544];
     layer2_out[1246] <= 1'b0;
     layer2_out[1247] <= layer1_out[1101] & ~layer1_out[1102];
     layer2_out[1248] <= ~(layer1_out[1068] & layer1_out[1069]);
     layer2_out[1249] <= ~layer1_out[542] | layer1_out[541];
     layer2_out[1250] <= 1'b1;
     layer2_out[1251] <= 1'b0;
     layer2_out[1252] <= ~layer1_out[914] | layer1_out[915];
     layer2_out[1253] <= ~layer1_out[1346];
     layer2_out[1254] <= ~(layer1_out[1361] | layer1_out[1362]);
     layer2_out[1255] <= 1'b0;
     layer2_out[1256] <= 1'b0;
     layer2_out[1257] <= layer1_out[1354];
     layer2_out[1258] <= ~layer1_out[1249];
     layer2_out[1259] <= ~layer1_out[1298] | layer1_out[1297];
     layer2_out[1260] <= 1'b1;
     layer2_out[1261] <= layer1_out[204] & ~layer1_out[205];
     layer2_out[1262] <= layer1_out[1102] & layer1_out[1103];
     layer2_out[1263] <= layer1_out[355] ^ layer1_out[356];
     layer2_out[1264] <= layer1_out[983] & ~layer1_out[982];
     layer2_out[1265] <= 1'b0;
     layer2_out[1266] <= 1'b0;
     layer2_out[1267] <= layer1_out[878] & ~layer1_out[879];
     layer2_out[1268] <= layer1_out[1018] | layer1_out[1019];
     layer2_out[1269] <= ~(layer1_out[337] & layer1_out[338]);
     layer2_out[1270] <= ~layer1_out[1251] | layer1_out[1250];
     layer2_out[1271] <= layer1_out[905] & ~layer1_out[906];
     layer2_out[1272] <= ~layer1_out[1055];
     layer2_out[1273] <= layer1_out[1454] & ~layer1_out[1453];
     layer2_out[1274] <= layer1_out[1296] & ~layer1_out[1295];
     layer2_out[1275] <= ~layer1_out[1055];
     layer2_out[1276] <= layer1_out[84];
     layer2_out[1277] <= ~layer1_out[192] | layer1_out[191];
     layer2_out[1278] <= layer1_out[441] & layer1_out[442];
     layer2_out[1279] <= ~layer1_out[222] | layer1_out[221];
     layer2_out[1280] <= ~(layer1_out[1352] & layer1_out[1353]);
     layer2_out[1281] <= ~(layer1_out[123] | layer1_out[124]);
     layer2_out[1282] <= 1'b0;
     layer2_out[1283] <= ~layer1_out[110] | layer1_out[109];
     layer2_out[1284] <= ~(layer1_out[380] & layer1_out[381]);
     layer2_out[1285] <= ~layer1_out[1244];
     layer2_out[1286] <= ~layer1_out[1115];
     layer2_out[1287] <= ~layer1_out[612];
     layer2_out[1288] <= ~(layer1_out[21] | layer1_out[22]);
     layer2_out[1289] <= ~layer1_out[115] | layer1_out[116];
     layer2_out[1290] <= ~(layer1_out[1401] | layer1_out[1402]);
     layer2_out[1291] <= ~layer1_out[1076] | layer1_out[1075];
     layer2_out[1292] <= layer1_out[1462] & ~layer1_out[1463];
     layer2_out[1293] <= layer1_out[1432] ^ layer1_out[1433];
     layer2_out[1294] <= layer1_out[395] & ~layer1_out[394];
     layer2_out[1295] <= ~layer1_out[220] | layer1_out[221];
     layer2_out[1296] <= layer1_out[137];
     layer2_out[1297] <= ~layer1_out[1030] | layer1_out[1031];
     layer2_out[1298] <= ~(layer1_out[572] | layer1_out[573]);
     layer2_out[1299] <= ~layer1_out[1228] | layer1_out[1227];
     layer2_out[1300] <= layer1_out[1261] | layer1_out[1262];
     layer2_out[1301] <= layer1_out[874] & layer1_out[875];
     layer2_out[1302] <= layer1_out[662] & layer1_out[663];
     layer2_out[1303] <= layer1_out[1257];
     layer2_out[1304] <= 1'b1;
     layer2_out[1305] <= ~layer1_out[169];
     layer2_out[1306] <= ~layer1_out[197] | layer1_out[198];
     layer2_out[1307] <= 1'b0;
     layer2_out[1308] <= ~layer1_out[1] | layer1_out[0];
     layer2_out[1309] <= 1'b1;
     layer2_out[1310] <= layer1_out[1350] & ~layer1_out[1351];
     layer2_out[1311] <= ~layer1_out[899] | layer1_out[900];
     layer2_out[1312] <= 1'b0;
     layer2_out[1313] <= layer1_out[1363] | layer1_out[1364];
     layer2_out[1314] <= ~layer1_out[321];
     layer2_out[1315] <= 1'b1;
     layer2_out[1316] <= ~layer1_out[508];
     layer2_out[1317] <= layer1_out[360] & ~layer1_out[359];
     layer2_out[1318] <= ~layer1_out[325] | layer1_out[326];
     layer2_out[1319] <= layer1_out[43] & layer1_out[44];
     layer2_out[1320] <= ~layer1_out[1348];
     layer2_out[1321] <= layer1_out[3] & ~layer1_out[4];
     layer2_out[1322] <= ~layer1_out[1099];
     layer2_out[1323] <= 1'b0;
     layer2_out[1324] <= ~layer1_out[1436] | layer1_out[1435];
     layer2_out[1325] <= 1'b1;
     layer2_out[1326] <= layer1_out[703];
     layer2_out[1327] <= layer1_out[388] | layer1_out[389];
     layer2_out[1328] <= layer1_out[567] & ~layer1_out[568];
     layer2_out[1329] <= layer1_out[284] & ~layer1_out[283];
     layer2_out[1330] <= layer1_out[66] & ~layer1_out[65];
     layer2_out[1331] <= ~layer1_out[952] | layer1_out[951];
     layer2_out[1332] <= ~(layer1_out[1465] & layer1_out[1466]);
     layer2_out[1333] <= layer1_out[1043] & layer1_out[1044];
     layer2_out[1334] <= ~layer1_out[1240] | layer1_out[1239];
     layer2_out[1335] <= layer1_out[167];
     layer2_out[1336] <= ~(layer1_out[452] | layer1_out[453]);
     layer2_out[1337] <= ~layer1_out[193];
     layer2_out[1338] <= 1'b0;
     layer2_out[1339] <= ~layer1_out[369] | layer1_out[368];
     layer2_out[1340] <= ~layer1_out[834] | layer1_out[835];
     layer2_out[1341] <= ~layer1_out[721] | layer1_out[722];
     layer2_out[1342] <= 1'b1;
     layer2_out[1343] <= layer1_out[1065];
     layer2_out[1344] <= 1'b1;
     layer2_out[1345] <= 1'b1;
     layer2_out[1346] <= layer1_out[1342] & layer1_out[1343];
     layer2_out[1347] <= ~layer1_out[385] | layer1_out[384];
     layer2_out[1348] <= 1'b1;
     layer2_out[1349] <= ~(layer1_out[125] & layer1_out[126]);
     layer2_out[1350] <= ~layer1_out[884];
     layer2_out[1351] <= layer1_out[113] & layer1_out[114];
     layer2_out[1352] <= layer1_out[1320] & layer1_out[1321];
     layer2_out[1353] <= 1'b1;
     layer2_out[1354] <= layer1_out[1027] | layer1_out[1028];
     layer2_out[1355] <= 1'b0;
     layer2_out[1356] <= ~(layer1_out[1304] | layer1_out[1305]);
     layer2_out[1357] <= layer1_out[360] & ~layer1_out[361];
     layer2_out[1358] <= ~(layer1_out[160] | layer1_out[161]);
     layer2_out[1359] <= layer1_out[833];
     layer2_out[1360] <= 1'b0;
     layer2_out[1361] <= 1'b1;
     layer2_out[1362] <= ~layer1_out[1176] | layer1_out[1177];
     layer2_out[1363] <= ~layer1_out[826] | layer1_out[825];
     layer2_out[1364] <= ~(layer1_out[694] & layer1_out[695]);
     layer2_out[1365] <= layer1_out[808] & layer1_out[809];
     layer2_out[1366] <= ~(layer1_out[1341] ^ layer1_out[1342]);
     layer2_out[1367] <= layer1_out[1292];
     layer2_out[1368] <= ~(layer1_out[1001] & layer1_out[1002]);
     layer2_out[1369] <= layer1_out[615] | layer1_out[616];
     layer2_out[1370] <= ~layer1_out[1288] | layer1_out[1289];
     layer2_out[1371] <= ~layer1_out[1213] | layer1_out[1214];
     layer2_out[1372] <= ~layer1_out[476];
     layer2_out[1373] <= 1'b0;
     layer2_out[1374] <= 1'b1;
     layer2_out[1375] <= ~layer1_out[1176] | layer1_out[1175];
     layer2_out[1376] <= layer1_out[1264] & ~layer1_out[1265];
     layer2_out[1377] <= ~(layer1_out[410] & layer1_out[411]);
     layer2_out[1378] <= layer1_out[100];
     layer2_out[1379] <= layer1_out[876];
     layer2_out[1380] <= ~layer1_out[902];
     layer2_out[1381] <= 1'b0;
     layer2_out[1382] <= layer1_out[393] & ~layer1_out[394];
     layer2_out[1383] <= ~layer1_out[680] | layer1_out[681];
     layer2_out[1384] <= ~layer1_out[131];
     layer2_out[1385] <= 1'b1;
     layer2_out[1386] <= layer1_out[952] & ~layer1_out[953];
     layer2_out[1387] <= ~layer1_out[235] | layer1_out[236];
     layer2_out[1388] <= ~layer1_out[906] | layer1_out[907];
     layer2_out[1389] <= layer1_out[69] & ~layer1_out[68];
     layer2_out[1390] <= layer1_out[1374] | layer1_out[1375];
     layer2_out[1391] <= 1'b0;
     layer2_out[1392] <= 1'b0;
     layer2_out[1393] <= layer1_out[1345];
     layer2_out[1394] <= layer1_out[520] | layer1_out[521];
     layer2_out[1395] <= layer1_out[642];
     layer2_out[1396] <= layer1_out[687];
     layer2_out[1397] <= layer1_out[935];
     layer2_out[1398] <= ~layer1_out[1211] | layer1_out[1212];
     layer2_out[1399] <= ~(layer1_out[1263] | layer1_out[1264]);
     layer2_out[1400] <= ~(layer1_out[223] & layer1_out[224]);
     layer2_out[1401] <= ~layer1_out[657];
     layer2_out[1402] <= ~(layer1_out[731] & layer1_out[732]);
     layer2_out[1403] <= 1'b1;
     layer2_out[1404] <= ~(layer1_out[1048] & layer1_out[1049]);
     layer2_out[1405] <= ~layer1_out[233];
     layer2_out[1406] <= layer1_out[177];
     layer2_out[1407] <= layer1_out[606];
     layer2_out[1408] <= ~layer1_out[916] | layer1_out[917];
     layer2_out[1409] <= 1'b0;
     layer2_out[1410] <= layer1_out[619];
     layer2_out[1411] <= ~layer1_out[1441];
     layer2_out[1412] <= 1'b0;
     layer2_out[1413] <= 1'b0;
     layer2_out[1414] <= layer1_out[1294];
     layer2_out[1415] <= ~layer1_out[1352] | layer1_out[1351];
     layer2_out[1416] <= ~layer1_out[520];
     layer2_out[1417] <= ~layer1_out[1301] | layer1_out[1300];
     layer2_out[1418] <= ~layer1_out[589];
     layer2_out[1419] <= ~layer1_out[372];
     layer2_out[1420] <= ~layer1_out[254] | layer1_out[255];
     layer2_out[1421] <= ~(layer1_out[691] | layer1_out[692]);
     layer2_out[1422] <= layer1_out[654] | layer1_out[655];
     layer2_out[1423] <= ~(layer1_out[323] | layer1_out[324]);
     layer2_out[1424] <= ~layer1_out[1173] | layer1_out[1174];
     layer2_out[1425] <= 1'b0;
     layer2_out[1426] <= ~layer1_out[796];
     layer2_out[1427] <= ~(layer1_out[1397] | layer1_out[1398]);
     layer2_out[1428] <= ~(layer1_out[1411] & layer1_out[1412]);
     layer2_out[1429] <= 1'b0;
     layer2_out[1430] <= 1'b0;
     layer2_out[1431] <= layer1_out[510] & ~layer1_out[509];
     layer2_out[1432] <= layer1_out[1101] & ~layer1_out[1100];
     layer2_out[1433] <= layer1_out[553] & layer1_out[554];
     layer2_out[1434] <= ~layer1_out[282];
     layer2_out[1435] <= layer1_out[17] & ~layer1_out[18];
     layer2_out[1436] <= layer1_out[812];
     layer2_out[1437] <= layer1_out[1109];
     layer2_out[1438] <= layer1_out[1308] & ~layer1_out[1307];
     layer2_out[1439] <= 1'b0;
     layer2_out[1440] <= ~layer1_out[957];
     layer2_out[1441] <= ~layer1_out[1151] | layer1_out[1152];
     layer2_out[1442] <= layer1_out[182] & ~layer1_out[181];
     layer2_out[1443] <= layer1_out[845];
     layer2_out[1444] <= layer1_out[1396] | layer1_out[1397];
     layer2_out[1445] <= 1'b0;
     layer2_out[1446] <= layer1_out[642] & ~layer1_out[643];
     layer2_out[1447] <= ~layer1_out[649] | layer1_out[648];
     layer2_out[1448] <= ~layer1_out[659] | layer1_out[660];
     layer2_out[1449] <= 1'b0;
     layer2_out[1450] <= 1'b0;
     layer2_out[1451] <= 1'b1;
     layer2_out[1452] <= ~(layer1_out[1357] ^ layer1_out[1358]);
     layer2_out[1453] <= layer1_out[269] & ~layer1_out[270];
     layer2_out[1454] <= layer1_out[227];
     layer2_out[1455] <= ~layer1_out[794];
     layer2_out[1456] <= layer1_out[679] & ~layer1_out[678];
     layer2_out[1457] <= layer1_out[156];
     layer2_out[1458] <= layer1_out[1267] & ~layer1_out[1268];
     layer2_out[1459] <= layer1_out[1434] | layer1_out[1435];
     layer2_out[1460] <= 1'b1;
     layer2_out[1461] <= layer1_out[103] | layer1_out[104];
     layer2_out[1462] <= layer1_out[1464] & layer1_out[1465];
     layer2_out[1463] <= ~layer1_out[217];
     layer2_out[1464] <= ~layer1_out[865] | layer1_out[864];
     layer2_out[1465] <= ~layer1_out[256];
     layer2_out[1466] <= layer1_out[777] & ~layer1_out[778];
     layer2_out[1467] <= ~(layer1_out[100] | layer1_out[101]);
     layer2_out[1468] <= layer1_out[1309] | layer1_out[1310];
     layer2_out[1469] <= 1'b0;
     layer2_out[1470] <= 1'b1;
     layer2_out[1471] <= 1'b1;
     layer2_out[1472] <= ~layer1_out[1131] | layer1_out[1130];
     layer2_out[1473] <= 1'b0;
     layer2_out[1474] <= ~layer1_out[1388] | layer1_out[1389];
     layer2_out[1475] <= layer1_out[1193] & layer1_out[1194];
     layer2_out[1476] <= ~(layer1_out[673] & layer1_out[674]);
     layer2_out[1477] <= ~(layer1_out[852] & layer1_out[853]);
     layer2_out[1478] <= 1'b1;
     layer2_out[1479] <= layer1_out[460] & ~layer1_out[461];
     layer2_out[1480] <= ~layer1_out[909];
     layer2_out[1481] <= layer1_out[947] & ~layer1_out[948];
     layer2_out[1482] <= ~layer1_out[1191];
     layer2_out[1483] <= 1'b0;
     layer2_out[1484] <= layer1_out[594] & ~layer1_out[593];
     layer2_out[1485] <= 1'b0;
     layer2_out[1486] <= 1'b0;
     layer2_out[1487] <= ~layer1_out[20] | layer1_out[21];
     layer2_out[1488] <= layer1_out[327];
     layer2_out[1489] <= ~(layer1_out[97] | layer1_out[98]);
     layer2_out[1490] <= layer1_out[149] & ~layer1_out[148];
     layer2_out[1491] <= 1'b0;
     layer2_out[1492] <= ~layer1_out[628] | layer1_out[629];
     layer2_out[1493] <= ~layer1_out[1258];
     layer2_out[1494] <= layer1_out[1348];
     layer2_out[1495] <= layer1_out[924] | layer1_out[925];
     layer2_out[1496] <= 1'b1;
     layer2_out[1497] <= ~(layer1_out[1389] | layer1_out[1390]);
     layer2_out[1498] <= layer1_out[647] | layer1_out[648];
     layer2_out[1499] <= 1'b0;
     layer3_out[0] <= ~layer2_out[21] | layer2_out[20];
     layer3_out[1] <= layer2_out[1255] & layer2_out[1256];
     layer3_out[2] <= layer2_out[1311] & ~layer2_out[1312];
     layer3_out[3] <= layer2_out[1492] & layer2_out[1493];
     layer3_out[4] <= 1'b1;
     layer3_out[5] <= layer2_out[1426];
     layer3_out[6] <= ~layer2_out[762] | layer2_out[761];
     layer3_out[7] <= layer2_out[907];
     layer3_out[8] <= layer2_out[340] | layer2_out[341];
     layer3_out[9] <= ~layer2_out[452];
     layer3_out[10] <= 1'b0;
     layer3_out[11] <= ~(layer2_out[531] | layer2_out[532]);
     layer3_out[12] <= layer2_out[119];
     layer3_out[13] <= ~layer2_out[1213];
     layer3_out[14] <= ~layer2_out[1478];
     layer3_out[15] <= layer2_out[528] | layer2_out[529];
     layer3_out[16] <= layer2_out[683] | layer2_out[684];
     layer3_out[17] <= ~layer2_out[1081];
     layer3_out[18] <= layer2_out[675] & ~layer2_out[676];
     layer3_out[19] <= ~layer2_out[646] | layer2_out[645];
     layer3_out[20] <= ~layer2_out[137];
     layer3_out[21] <= layer2_out[1231];
     layer3_out[22] <= ~layer2_out[486] | layer2_out[487];
     layer3_out[23] <= ~(layer2_out[158] | layer2_out[159]);
     layer3_out[24] <= layer2_out[1254];
     layer3_out[25] <= ~(layer2_out[1383] & layer2_out[1384]);
     layer3_out[26] <= layer2_out[313];
     layer3_out[27] <= layer2_out[9] & ~layer2_out[8];
     layer3_out[28] <= ~(layer2_out[887] ^ layer2_out[888]);
     layer3_out[29] <= layer2_out[1107] & ~layer2_out[1108];
     layer3_out[30] <= layer2_out[470];
     layer3_out[31] <= layer2_out[830] & layer2_out[831];
     layer3_out[32] <= ~layer2_out[756];
     layer3_out[33] <= layer2_out[1106] & layer2_out[1107];
     layer3_out[34] <= ~layer2_out[1024] | layer2_out[1023];
     layer3_out[35] <= layer2_out[611];
     layer3_out[36] <= layer2_out[338] & layer2_out[339];
     layer3_out[37] <= layer2_out[1077] & ~layer2_out[1076];
     layer3_out[38] <= layer2_out[959];
     layer3_out[39] <= ~(layer2_out[939] | layer2_out[940]);
     layer3_out[40] <= 1'b1;
     layer3_out[41] <= layer2_out[13] | layer2_out[14];
     layer3_out[42] <= layer2_out[1176] & layer2_out[1177];
     layer3_out[43] <= ~(layer2_out[595] | layer2_out[596]);
     layer3_out[44] <= ~layer2_out[1047];
     layer3_out[45] <= ~layer2_out[1217] | layer2_out[1218];
     layer3_out[46] <= layer2_out[522] & layer2_out[523];
     layer3_out[47] <= layer2_out[250] & ~layer2_out[249];
     layer3_out[48] <= ~layer2_out[572] | layer2_out[571];
     layer3_out[49] <= ~(layer2_out[46] ^ layer2_out[47]);
     layer3_out[50] <= ~layer2_out[105] | layer2_out[106];
     layer3_out[51] <= layer2_out[108] & layer2_out[109];
     layer3_out[52] <= layer2_out[257];
     layer3_out[53] <= ~(layer2_out[59] & layer2_out[60]);
     layer3_out[54] <= 1'b0;
     layer3_out[55] <= layer2_out[314] & layer2_out[315];
     layer3_out[56] <= layer2_out[494];
     layer3_out[57] <= ~(layer2_out[913] | layer2_out[914]);
     layer3_out[58] <= ~layer2_out[1492] | layer2_out[1491];
     layer3_out[59] <= 1'b0;
     layer3_out[60] <= ~layer2_out[910];
     layer3_out[61] <= layer2_out[113] & layer2_out[114];
     layer3_out[62] <= layer2_out[832] & ~layer2_out[833];
     layer3_out[63] <= 1'b0;
     layer3_out[64] <= ~layer2_out[706] | layer2_out[705];
     layer3_out[65] <= ~layer2_out[590];
     layer3_out[66] <= layer2_out[576] & ~layer2_out[575];
     layer3_out[67] <= layer2_out[1384] & ~layer2_out[1385];
     layer3_out[68] <= layer2_out[851] & layer2_out[852];
     layer3_out[69] <= ~layer2_out[866];
     layer3_out[70] <= layer2_out[93] & ~layer2_out[92];
     layer3_out[71] <= ~layer2_out[261] | layer2_out[262];
     layer3_out[72] <= ~layer2_out[1283];
     layer3_out[73] <= ~(layer2_out[203] | layer2_out[204]);
     layer3_out[74] <= layer2_out[287] & layer2_out[288];
     layer3_out[75] <= layer2_out[1285];
     layer3_out[76] <= layer2_out[672];
     layer3_out[77] <= layer2_out[412];
     layer3_out[78] <= ~layer2_out[511] | layer2_out[512];
     layer3_out[79] <= ~layer2_out[369];
     layer3_out[80] <= 1'b1;
     layer3_out[81] <= layer2_out[172] & ~layer2_out[171];
     layer3_out[82] <= 1'b1;
     layer3_out[83] <= ~layer2_out[276] | layer2_out[277];
     layer3_out[84] <= ~layer2_out[1039];
     layer3_out[85] <= ~layer2_out[401];
     layer3_out[86] <= 1'b0;
     layer3_out[87] <= layer2_out[119] & ~layer2_out[118];
     layer3_out[88] <= layer2_out[209] & ~layer2_out[208];
     layer3_out[89] <= 1'b1;
     layer3_out[90] <= layer2_out[1431];
     layer3_out[91] <= layer2_out[879] | layer2_out[880];
     layer3_out[92] <= ~(layer2_out[1086] | layer2_out[1087]);
     layer3_out[93] <= ~layer2_out[1456];
     layer3_out[94] <= ~layer2_out[1429];
     layer3_out[95] <= layer2_out[533] & ~layer2_out[534];
     layer3_out[96] <= layer2_out[40];
     layer3_out[97] <= ~(layer2_out[335] | layer2_out[336]);
     layer3_out[98] <= layer2_out[534] & layer2_out[535];
     layer3_out[99] <= ~layer2_out[484];
     layer3_out[100] <= 1'b1;
     layer3_out[101] <= ~(layer2_out[1367] | layer2_out[1368]);
     layer3_out[102] <= layer2_out[78] & layer2_out[79];
     layer3_out[103] <= 1'b1;
     layer3_out[104] <= ~layer2_out[1077];
     layer3_out[105] <= layer2_out[717] & ~layer2_out[718];
     layer3_out[106] <= layer2_out[731];
     layer3_out[107] <= ~layer2_out[712];
     layer3_out[108] <= layer2_out[1377];
     layer3_out[109] <= ~layer2_out[0] | layer2_out[2];
     layer3_out[110] <= ~(layer2_out[91] & layer2_out[92]);
     layer3_out[111] <= ~layer2_out[539] | layer2_out[540];
     layer3_out[112] <= 1'b0;
     layer3_out[113] <= layer2_out[961] ^ layer2_out[962];
     layer3_out[114] <= layer2_out[1146];
     layer3_out[115] <= ~(layer2_out[845] | layer2_out[846]);
     layer3_out[116] <= layer2_out[278] & layer2_out[279];
     layer3_out[117] <= 1'b0;
     layer3_out[118] <= ~layer2_out[952] | layer2_out[951];
     layer3_out[119] <= ~layer2_out[1356];
     layer3_out[120] <= ~(layer2_out[501] & layer2_out[502]);
     layer3_out[121] <= 1'b1;
     layer3_out[122] <= ~layer2_out[1266];
     layer3_out[123] <= ~layer2_out[710] | layer2_out[709];
     layer3_out[124] <= 1'b0;
     layer3_out[125] <= layer2_out[475] & ~layer2_out[476];
     layer3_out[126] <= ~layer2_out[325];
     layer3_out[127] <= layer2_out[1421] & ~layer2_out[1420];
     layer3_out[128] <= ~layer2_out[1263];
     layer3_out[129] <= layer2_out[1063];
     layer3_out[130] <= ~layer2_out[896];
     layer3_out[131] <= layer2_out[978] | layer2_out[979];
     layer3_out[132] <= ~layer2_out[1129];
     layer3_out[133] <= ~(layer2_out[1480] | layer2_out[1481]);
     layer3_out[134] <= ~(layer2_out[1498] | layer2_out[1499]);
     layer3_out[135] <= 1'b1;
     layer3_out[136] <= 1'b0;
     layer3_out[137] <= layer2_out[1271] | layer2_out[1272];
     layer3_out[138] <= 1'b1;
     layer3_out[139] <= ~layer2_out[259];
     layer3_out[140] <= ~(layer2_out[711] & layer2_out[712]);
     layer3_out[141] <= layer2_out[935] & layer2_out[936];
     layer3_out[142] <= ~layer2_out[816] | layer2_out[817];
     layer3_out[143] <= 1'b0;
     layer3_out[144] <= layer2_out[236] & ~layer2_out[235];
     layer3_out[145] <= ~layer2_out[1291] | layer2_out[1290];
     layer3_out[146] <= ~layer2_out[885];
     layer3_out[147] <= layer2_out[689] & layer2_out[690];
     layer3_out[148] <= ~layer2_out[1372] | layer2_out[1373];
     layer3_out[149] <= layer2_out[844];
     layer3_out[150] <= ~(layer2_out[1211] | layer2_out[1212]);
     layer3_out[151] <= ~layer2_out[316] | layer2_out[315];
     layer3_out[152] <= layer2_out[1354];
     layer3_out[153] <= ~layer2_out[65] | layer2_out[66];
     layer3_out[154] <= layer2_out[808] & ~layer2_out[809];
     layer3_out[155] <= layer2_out[920];
     layer3_out[156] <= layer2_out[285] & ~layer2_out[286];
     layer3_out[157] <= ~(layer2_out[1308] | layer2_out[1309]);
     layer3_out[158] <= layer2_out[347];
     layer3_out[159] <= layer2_out[1399] & ~layer2_out[1398];
     layer3_out[160] <= 1'b1;
     layer3_out[161] <= ~layer2_out[140] | layer2_out[139];
     layer3_out[162] <= 1'b1;
     layer3_out[163] <= ~(layer2_out[716] | layer2_out[717]);
     layer3_out[164] <= layer2_out[251] & ~layer2_out[252];
     layer3_out[165] <= layer2_out[641] | layer2_out[642];
     layer3_out[166] <= layer2_out[279];
     layer3_out[167] <= layer2_out[1365] & layer2_out[1366];
     layer3_out[168] <= layer2_out[12] & ~layer2_out[11];
     layer3_out[169] <= ~layer2_out[196] | layer2_out[197];
     layer3_out[170] <= ~layer2_out[358] | layer2_out[357];
     layer3_out[171] <= ~layer2_out[300] | layer2_out[299];
     layer3_out[172] <= ~layer2_out[1104] | layer2_out[1105];
     layer3_out[173] <= 1'b1;
     layer3_out[174] <= 1'b0;
     layer3_out[175] <= 1'b1;
     layer3_out[176] <= layer2_out[549] & layer2_out[550];
     layer3_out[177] <= 1'b0;
     layer3_out[178] <= ~layer2_out[385] | layer2_out[386];
     layer3_out[179] <= 1'b1;
     layer3_out[180] <= layer2_out[1204] & ~layer2_out[1203];
     layer3_out[181] <= layer2_out[760];
     layer3_out[182] <= ~layer2_out[800] | layer2_out[799];
     layer3_out[183] <= layer2_out[420] & layer2_out[421];
     layer3_out[184] <= 1'b1;
     layer3_out[185] <= ~layer2_out[1354];
     layer3_out[186] <= 1'b1;
     layer3_out[187] <= layer2_out[838] & ~layer2_out[837];
     layer3_out[188] <= layer2_out[793] & layer2_out[794];
     layer3_out[189] <= layer2_out[28] & ~layer2_out[29];
     layer3_out[190] <= layer2_out[1090] | layer2_out[1091];
     layer3_out[191] <= ~(layer2_out[331] & layer2_out[332]);
     layer3_out[192] <= ~layer2_out[840] | layer2_out[841];
     layer3_out[193] <= ~layer2_out[212];
     layer3_out[194] <= layer2_out[881] | layer2_out[882];
     layer3_out[195] <= 1'b0;
     layer3_out[196] <= ~layer2_out[1380] | layer2_out[1379];
     layer3_out[197] <= layer2_out[726] | layer2_out[727];
     layer3_out[198] <= ~layer2_out[1136];
     layer3_out[199] <= ~layer2_out[1346] | layer2_out[1347];
     layer3_out[200] <= layer2_out[743] ^ layer2_out[744];
     layer3_out[201] <= layer2_out[423] | layer2_out[424];
     layer3_out[202] <= ~layer2_out[860] | layer2_out[861];
     layer3_out[203] <= ~layer2_out[152];
     layer3_out[204] <= layer2_out[999] | layer2_out[1000];
     layer3_out[205] <= layer2_out[1092] & ~layer2_out[1091];
     layer3_out[206] <= layer2_out[776];
     layer3_out[207] <= layer2_out[236];
     layer3_out[208] <= 1'b1;
     layer3_out[209] <= layer2_out[791] | layer2_out[792];
     layer3_out[210] <= layer2_out[1093] & layer2_out[1094];
     layer3_out[211] <= layer2_out[47];
     layer3_out[212] <= layer2_out[386] | layer2_out[387];
     layer3_out[213] <= ~layer2_out[628] | layer2_out[627];
     layer3_out[214] <= ~(layer2_out[1000] & layer2_out[1001]);
     layer3_out[215] <= ~layer2_out[139] | layer2_out[138];
     layer3_out[216] <= ~layer2_out[235] | layer2_out[234];
     layer3_out[217] <= 1'b0;
     layer3_out[218] <= ~layer2_out[593];
     layer3_out[219] <= layer2_out[244];
     layer3_out[220] <= 1'b1;
     layer3_out[221] <= layer2_out[27] | layer2_out[28];
     layer3_out[222] <= ~layer2_out[754];
     layer3_out[223] <= ~layer2_out[616];
     layer3_out[224] <= ~layer2_out[526] | layer2_out[527];
     layer3_out[225] <= layer2_out[1227] & ~layer2_out[1228];
     layer3_out[226] <= layer2_out[565];
     layer3_out[227] <= layer2_out[874] & ~layer2_out[873];
     layer3_out[228] <= layer2_out[1258] | layer2_out[1259];
     layer3_out[229] <= layer2_out[1101] | layer2_out[1102];
     layer3_out[230] <= layer2_out[899] ^ layer2_out[900];
     layer3_out[231] <= 1'b1;
     layer3_out[232] <= layer2_out[1200];
     layer3_out[233] <= layer2_out[1095] | layer2_out[1096];
     layer3_out[234] <= ~layer2_out[1009];
     layer3_out[235] <= ~layer2_out[174];
     layer3_out[236] <= ~layer2_out[986] | layer2_out[987];
     layer3_out[237] <= 1'b1;
     layer3_out[238] <= ~(layer2_out[1315] & layer2_out[1316]);
     layer3_out[239] <= ~layer2_out[1404];
     layer3_out[240] <= ~layer2_out[380];
     layer3_out[241] <= ~(layer2_out[871] & layer2_out[872]);
     layer3_out[242] <= 1'b0;
     layer3_out[243] <= ~layer2_out[1045] | layer2_out[1046];
     layer3_out[244] <= 1'b1;
     layer3_out[245] <= ~(layer2_out[1182] | layer2_out[1183]);
     layer3_out[246] <= layer2_out[1404];
     layer3_out[247] <= ~(layer2_out[545] & layer2_out[546]);
     layer3_out[248] <= ~(layer2_out[981] | layer2_out[982]);
     layer3_out[249] <= ~(layer2_out[770] | layer2_out[771]);
     layer3_out[250] <= 1'b1;
     layer3_out[251] <= layer2_out[1157];
     layer3_out[252] <= 1'b0;
     layer3_out[253] <= ~layer2_out[931] | layer2_out[930];
     layer3_out[254] <= ~(layer2_out[474] | layer2_out[475]);
     layer3_out[255] <= ~layer2_out[998] | layer2_out[999];
     layer3_out[256] <= layer2_out[499];
     layer3_out[257] <= ~layer2_out[1090];
     layer3_out[258] <= ~(layer2_out[572] & layer2_out[573]);
     layer3_out[259] <= 1'b1;
     layer3_out[260] <= ~layer2_out[954] | layer2_out[953];
     layer3_out[261] <= layer2_out[1166] & layer2_out[1167];
     layer3_out[262] <= layer2_out[1196] & ~layer2_out[1195];
     layer3_out[263] <= layer2_out[1280];
     layer3_out[264] <= layer2_out[214] & ~layer2_out[215];
     layer3_out[265] <= layer2_out[135];
     layer3_out[266] <= ~layer2_out[88];
     layer3_out[267] <= ~layer2_out[405] | layer2_out[404];
     layer3_out[268] <= ~(layer2_out[1154] & layer2_out[1155]);
     layer3_out[269] <= ~layer2_out[964] | layer2_out[965];
     layer3_out[270] <= 1'b1;
     layer3_out[271] <= ~layer2_out[1083];
     layer3_out[272] <= layer2_out[384] & ~layer2_out[383];
     layer3_out[273] <= layer2_out[1041] ^ layer2_out[1042];
     layer3_out[274] <= ~layer2_out[1261] | layer2_out[1260];
     layer3_out[275] <= ~layer2_out[430];
     layer3_out[276] <= ~layer2_out[1075];
     layer3_out[277] <= ~layer2_out[814];
     layer3_out[278] <= ~(layer2_out[566] | layer2_out[567]);
     layer3_out[279] <= layer2_out[148] & layer2_out[149];
     layer3_out[280] <= ~layer2_out[575] | layer2_out[574];
     layer3_out[281] <= ~(layer2_out[560] | layer2_out[561]);
     layer3_out[282] <= layer2_out[256] & ~layer2_out[255];
     layer3_out[283] <= layer2_out[94] & ~layer2_out[95];
     layer3_out[284] <= layer2_out[295] | layer2_out[296];
     layer3_out[285] <= 1'b0;
     layer3_out[286] <= ~layer2_out[359];
     layer3_out[287] <= layer2_out[1234];
     layer3_out[288] <= layer2_out[1419] & ~layer2_out[1418];
     layer3_out[289] <= ~(layer2_out[692] ^ layer2_out[693]);
     layer3_out[290] <= 1'b1;
     layer3_out[291] <= layer2_out[247] & ~layer2_out[248];
     layer3_out[292] <= 1'b0;
     layer3_out[293] <= layer2_out[1063] & ~layer2_out[1064];
     layer3_out[294] <= ~(layer2_out[954] | layer2_out[955]);
     layer3_out[295] <= layer2_out[111];
     layer3_out[296] <= 1'b0;
     layer3_out[297] <= ~(layer2_out[6] | layer2_out[7]);
     layer3_out[298] <= layer2_out[611];
     layer3_out[299] <= layer2_out[943] | layer2_out[944];
     layer3_out[300] <= ~layer2_out[245];
     layer3_out[301] <= 1'b1;
     layer3_out[302] <= 1'b0;
     layer3_out[303] <= ~layer2_out[1141];
     layer3_out[304] <= layer2_out[631];
     layer3_out[305] <= ~layer2_out[422];
     layer3_out[306] <= ~layer2_out[150];
     layer3_out[307] <= ~(layer2_out[1200] & layer2_out[1201]);
     layer3_out[308] <= layer2_out[687] & ~layer2_out[688];
     layer3_out[309] <= layer2_out[901] & ~layer2_out[900];
     layer3_out[310] <= ~layer2_out[672] | layer2_out[673];
     layer3_out[311] <= layer2_out[562];
     layer3_out[312] <= ~layer2_out[1037] | layer2_out[1038];
     layer3_out[313] <= layer2_out[169] & ~layer2_out[168];
     layer3_out[314] <= layer2_out[858] | layer2_out[859];
     layer3_out[315] <= ~(layer2_out[669] & layer2_out[670]);
     layer3_out[316] <= ~layer2_out[1108];
     layer3_out[317] <= ~(layer2_out[82] | layer2_out[83]);
     layer3_out[318] <= layer2_out[904] & layer2_out[905];
     layer3_out[319] <= 1'b1;
     layer3_out[320] <= layer2_out[765];
     layer3_out[321] <= layer2_out[1187];
     layer3_out[322] <= ~layer2_out[18] | layer2_out[17];
     layer3_out[323] <= 1'b0;
     layer3_out[324] <= ~layer2_out[568] | layer2_out[567];
     layer3_out[325] <= layer2_out[541] & layer2_out[542];
     layer3_out[326] <= layer2_out[1413] & layer2_out[1414];
     layer3_out[327] <= layer2_out[981] & ~layer2_out[980];
     layer3_out[328] <= ~layer2_out[737] | layer2_out[738];
     layer3_out[329] <= ~layer2_out[151];
     layer3_out[330] <= ~layer2_out[439];
     layer3_out[331] <= ~(layer2_out[416] | layer2_out[417]);
     layer3_out[332] <= ~(layer2_out[403] | layer2_out[404]);
     layer3_out[333] <= ~layer2_out[72] | layer2_out[73];
     layer3_out[334] <= 1'b0;
     layer3_out[335] <= layer2_out[1161] & layer2_out[1162];
     layer3_out[336] <= ~(layer2_out[306] & layer2_out[307]);
     layer3_out[337] <= ~layer2_out[844] | layer2_out[845];
     layer3_out[338] <= 1'b1;
     layer3_out[339] <= ~(layer2_out[1348] & layer2_out[1349]);
     layer3_out[340] <= ~layer2_out[585];
     layer3_out[341] <= ~layer2_out[656] | layer2_out[657];
     layer3_out[342] <= layer2_out[488] | layer2_out[489];
     layer3_out[343] <= layer2_out[399];
     layer3_out[344] <= ~layer2_out[1121] | layer2_out[1120];
     layer3_out[345] <= layer2_out[994];
     layer3_out[346] <= layer2_out[1333];
     layer3_out[347] <= layer2_out[1132];
     layer3_out[348] <= layer2_out[31];
     layer3_out[349] <= layer2_out[1380];
     layer3_out[350] <= layer2_out[746];
     layer3_out[351] <= ~layer2_out[1189] | layer2_out[1188];
     layer3_out[352] <= 1'b1;
     layer3_out[353] <= layer2_out[223] & ~layer2_out[222];
     layer3_out[354] <= layer2_out[418];
     layer3_out[355] <= layer2_out[874] & ~layer2_out[875];
     layer3_out[356] <= ~layer2_out[1136] | layer2_out[1137];
     layer3_out[357] <= ~layer2_out[1113];
     layer3_out[358] <= ~(layer2_out[352] | layer2_out[353]);
     layer3_out[359] <= ~layer2_out[509] | layer2_out[508];
     layer3_out[360] <= ~(layer2_out[43] & layer2_out[44]);
     layer3_out[361] <= layer2_out[700];
     layer3_out[362] <= ~layer2_out[216] | layer2_out[215];
     layer3_out[363] <= ~(layer2_out[1440] ^ layer2_out[1441]);
     layer3_out[364] <= layer2_out[53] | layer2_out[54];
     layer3_out[365] <= layer2_out[268] & ~layer2_out[269];
     layer3_out[366] <= ~(layer2_out[371] & layer2_out[372]);
     layer3_out[367] <= layer2_out[1439];
     layer3_out[368] <= layer2_out[790] & ~layer2_out[791];
     layer3_out[369] <= layer2_out[131] & layer2_out[132];
     layer3_out[370] <= layer2_out[260];
     layer3_out[371] <= layer2_out[523] & layer2_out[524];
     layer3_out[372] <= 1'b1;
     layer3_out[373] <= layer2_out[587] & ~layer2_out[586];
     layer3_out[374] <= layer2_out[923] | layer2_out[924];
     layer3_out[375] <= ~layer2_out[1254];
     layer3_out[376] <= layer2_out[1414] & ~layer2_out[1415];
     layer3_out[377] <= layer2_out[252];
     layer3_out[378] <= layer2_out[70] | layer2_out[71];
     layer3_out[379] <= ~layer2_out[137];
     layer3_out[380] <= 1'b0;
     layer3_out[381] <= ~(layer2_out[375] | layer2_out[376]);
     layer3_out[382] <= ~layer2_out[1043];
     layer3_out[383] <= layer2_out[661] & layer2_out[662];
     layer3_out[384] <= layer2_out[1028] & layer2_out[1029];
     layer3_out[385] <= layer2_out[821] | layer2_out[822];
     layer3_out[386] <= ~layer2_out[336];
     layer3_out[387] <= layer2_out[1134];
     layer3_out[388] <= ~(layer2_out[536] | layer2_out[537]);
     layer3_out[389] <= layer2_out[484] & ~layer2_out[485];
     layer3_out[390] <= 1'b0;
     layer3_out[391] <= layer2_out[238];
     layer3_out[392] <= layer2_out[1124];
     layer3_out[393] <= ~layer2_out[1031];
     layer3_out[394] <= ~layer2_out[477] | layer2_out[476];
     layer3_out[395] <= layer2_out[907] | layer2_out[908];
     layer3_out[396] <= layer2_out[937];
     layer3_out[397] <= layer2_out[1109] & ~layer2_out[1110];
     layer3_out[398] <= ~layer2_out[308];
     layer3_out[399] <= ~layer2_out[1358] | layer2_out[1359];
     layer3_out[400] <= ~layer2_out[461] | layer2_out[462];
     layer3_out[401] <= layer2_out[454];
     layer3_out[402] <= ~(layer2_out[1117] & layer2_out[1118]);
     layer3_out[403] <= ~layer2_out[1128] | layer2_out[1127];
     layer3_out[404] <= ~layer2_out[1378];
     layer3_out[405] <= ~layer2_out[88];
     layer3_out[406] <= layer2_out[736] & ~layer2_out[737];
     layer3_out[407] <= 1'b1;
     layer3_out[408] <= layer2_out[147];
     layer3_out[409] <= layer2_out[830];
     layer3_out[410] <= ~layer2_out[110];
     layer3_out[411] <= ~layer2_out[985];
     layer3_out[412] <= layer2_out[301] & ~layer2_out[302];
     layer3_out[413] <= layer2_out[1096] | layer2_out[1097];
     layer3_out[414] <= 1'b1;
     layer3_out[415] <= ~(layer2_out[1167] | layer2_out[1168]);
     layer3_out[416] <= ~layer2_out[629];
     layer3_out[417] <= ~layer2_out[186] | layer2_out[187];
     layer3_out[418] <= layer2_out[775];
     layer3_out[419] <= ~layer2_out[272];
     layer3_out[420] <= layer2_out[353] & ~layer2_out[354];
     layer3_out[421] <= ~layer2_out[648];
     layer3_out[422] <= layer2_out[1489] & ~layer2_out[1490];
     layer3_out[423] <= ~layer2_out[1366] | layer2_out[1367];
     layer3_out[424] <= ~layer2_out[414];
     layer3_out[425] <= ~layer2_out[714] | layer2_out[713];
     layer3_out[426] <= 1'b1;
     layer3_out[427] <= layer2_out[1305] | layer2_out[1306];
     layer3_out[428] <= ~layer2_out[552] | layer2_out[553];
     layer3_out[429] <= layer2_out[549] & ~layer2_out[548];
     layer3_out[430] <= layer2_out[1442] & ~layer2_out[1443];
     layer3_out[431] <= layer2_out[1036];
     layer3_out[432] <= 1'b0;
     layer3_out[433] <= ~layer2_out[1437] | layer2_out[1438];
     layer3_out[434] <= layer2_out[272] | layer2_out[273];
     layer3_out[435] <= ~layer2_out[1026];
     layer3_out[436] <= ~layer2_out[1335];
     layer3_out[437] <= layer2_out[71] & ~layer2_out[72];
     layer3_out[438] <= ~layer2_out[1013] | layer2_out[1014];
     layer3_out[439] <= ~(layer2_out[833] | layer2_out[834]);
     layer3_out[440] <= layer2_out[339] ^ layer2_out[340];
     layer3_out[441] <= layer2_out[159] & ~layer2_out[160];
     layer3_out[442] <= ~(layer2_out[973] | layer2_out[974]);
     layer3_out[443] <= 1'b0;
     layer3_out[444] <= layer2_out[910] & ~layer2_out[911];
     layer3_out[445] <= 1'b0;
     layer3_out[446] <= layer2_out[1349] & layer2_out[1350];
     layer3_out[447] <= ~layer2_out[32];
     layer3_out[448] <= layer2_out[1460] & ~layer2_out[1461];
     layer3_out[449] <= layer2_out[580];
     layer3_out[450] <= ~layer2_out[1171] | layer2_out[1170];
     layer3_out[451] <= layer2_out[1177] & layer2_out[1178];
     layer3_out[452] <= ~layer2_out[285];
     layer3_out[453] <= layer2_out[1444] | layer2_out[1445];
     layer3_out[454] <= layer2_out[932];
     layer3_out[455] <= ~layer2_out[603] | layer2_out[602];
     layer3_out[456] <= ~(layer2_out[1252] | layer2_out[1253]);
     layer3_out[457] <= 1'b0;
     layer3_out[458] <= 1'b1;
     layer3_out[459] <= ~(layer2_out[45] | layer2_out[46]);
     layer3_out[460] <= ~layer2_out[1475] | layer2_out[1474];
     layer3_out[461] <= layer2_out[1247] & ~layer2_out[1248];
     layer3_out[462] <= layer2_out[649];
     layer3_out[463] <= layer2_out[101] & layer2_out[102];
     layer3_out[464] <= 1'b1;
     layer3_out[465] <= layer2_out[287];
     layer3_out[466] <= ~(layer2_out[191] & layer2_out[192]);
     layer3_out[467] <= ~layer2_out[1276];
     layer3_out[468] <= layer2_out[1213] | layer2_out[1214];
     layer3_out[469] <= ~layer2_out[1099];
     layer3_out[470] <= ~layer2_out[606];
     layer3_out[471] <= layer2_out[1465] & layer2_out[1466];
     layer3_out[472] <= ~layer2_out[153];
     layer3_out[473] <= layer2_out[426];
     layer3_out[474] <= ~layer2_out[179] | layer2_out[180];
     layer3_out[475] <= layer2_out[15];
     layer3_out[476] <= layer2_out[1449];
     layer3_out[477] <= ~(layer2_out[1381] & layer2_out[1382]);
     layer3_out[478] <= layer2_out[428] & ~layer2_out[429];
     layer3_out[479] <= layer2_out[812];
     layer3_out[480] <= layer2_out[897] & layer2_out[898];
     layer3_out[481] <= layer2_out[938] & ~layer2_out[937];
     layer3_out[482] <= 1'b0;
     layer3_out[483] <= ~layer2_out[194];
     layer3_out[484] <= layer2_out[1181] | layer2_out[1182];
     layer3_out[485] <= layer2_out[1320];
     layer3_out[486] <= layer2_out[733];
     layer3_out[487] <= layer2_out[1406] & ~layer2_out[1407];
     layer3_out[488] <= ~(layer2_out[332] | layer2_out[333]);
     layer3_out[489] <= layer2_out[544];
     layer3_out[490] <= layer2_out[991] & ~layer2_out[992];
     layer3_out[491] <= ~(layer2_out[1229] & layer2_out[1230]);
     layer3_out[492] <= 1'b0;
     layer3_out[493] <= layer2_out[370];
     layer3_out[494] <= ~(layer2_out[399] & layer2_out[400]);
     layer3_out[495] <= 1'b0;
     layer3_out[496] <= layer2_out[1362] | layer2_out[1363];
     layer3_out[497] <= layer2_out[1125];
     layer3_out[498] <= ~layer2_out[826] | layer2_out[825];
     layer3_out[499] <= 1'b0;
     layer3_out[500] <= layer2_out[1030] & ~layer2_out[1029];
     layer3_out[501] <= ~(layer2_out[755] & layer2_out[756]);
     layer3_out[502] <= ~layer2_out[643];
     layer3_out[503] <= ~(layer2_out[1197] & layer2_out[1198]);
     layer3_out[504] <= ~layer2_out[389] | layer2_out[390];
     layer3_out[505] <= ~layer2_out[1457];
     layer3_out[506] <= layer2_out[792] | layer2_out[793];
     layer3_out[507] <= ~(layer2_out[1206] | layer2_out[1207]);
     layer3_out[508] <= layer2_out[1047];
     layer3_out[509] <= layer2_out[739] & layer2_out[740];
     layer3_out[510] <= ~(layer2_out[89] | layer2_out[90]);
     layer3_out[511] <= layer2_out[969];
     layer3_out[512] <= 1'b1;
     layer3_out[513] <= layer2_out[977] & layer2_out[978];
     layer3_out[514] <= layer2_out[688] | layer2_out[689];
     layer3_out[515] <= 1'b1;
     layer3_out[516] <= layer2_out[1242];
     layer3_out[517] <= layer2_out[1268] & layer2_out[1269];
     layer3_out[518] <= layer2_out[1453] & ~layer2_out[1452];
     layer3_out[519] <= layer2_out[316];
     layer3_out[520] <= layer2_out[887];
     layer3_out[521] <= ~(layer2_out[1232] | layer2_out[1233]);
     layer3_out[522] <= ~layer2_out[1056] | layer2_out[1055];
     layer3_out[523] <= ~(layer2_out[1292] & layer2_out[1293]);
     layer3_out[524] <= 1'b1;
     layer3_out[525] <= layer2_out[120] & ~layer2_out[121];
     layer3_out[526] <= layer2_out[184] & ~layer2_out[185];
     layer3_out[527] <= layer2_out[1332] & layer2_out[1333];
     layer3_out[528] <= layer2_out[823] & ~layer2_out[822];
     layer3_out[529] <= ~layer2_out[303];
     layer3_out[530] <= ~(layer2_out[1433] | layer2_out[1434]);
     layer3_out[531] <= ~(layer2_out[106] | layer2_out[107]);
     layer3_out[532] <= ~layer2_out[1265] | layer2_out[1264];
     layer3_out[533] <= 1'b0;
     layer3_out[534] <= ~layer2_out[896] | layer2_out[895];
     layer3_out[535] <= ~(layer2_out[621] | layer2_out[622]);
     layer3_out[536] <= layer2_out[1105] & layer2_out[1106];
     layer3_out[537] <= ~(layer2_out[750] & layer2_out[751]);
     layer3_out[538] <= ~layer2_out[1142] | layer2_out[1143];
     layer3_out[539] <= ~(layer2_out[392] & layer2_out[393]);
     layer3_out[540] <= ~layer2_out[1013] | layer2_out[1012];
     layer3_out[541] <= ~(layer2_out[1321] & layer2_out[1322]);
     layer3_out[542] <= 1'b1;
     layer3_out[543] <= ~(layer2_out[1375] | layer2_out[1376]);
     layer3_out[544] <= 1'b0;
     layer3_out[545] <= ~layer2_out[363] | layer2_out[364];
     layer3_out[546] <= layer2_out[623];
     layer3_out[547] <= 1'b0;
     layer3_out[548] <= ~layer2_out[662];
     layer3_out[549] <= layer2_out[665];
     layer3_out[550] <= ~layer2_out[620];
     layer3_out[551] <= ~(layer2_out[326] & layer2_out[327]);
     layer3_out[552] <= layer2_out[602] & ~layer2_out[601];
     layer3_out[553] <= 1'b1;
     layer3_out[554] <= ~layer2_out[248] | layer2_out[249];
     layer3_out[555] <= 1'b0;
     layer3_out[556] <= ~layer2_out[1370];
     layer3_out[557] <= ~(layer2_out[50] | layer2_out[51]);
     layer3_out[558] <= layer2_out[470] & ~layer2_out[471];
     layer3_out[559] <= ~layer2_out[1386] | layer2_out[1385];
     layer3_out[560] <= ~(layer2_out[551] & layer2_out[552]);
     layer3_out[561] <= ~layer2_out[698] | layer2_out[699];
     layer3_out[562] <= layer2_out[1296] & ~layer2_out[1295];
     layer3_out[563] <= 1'b0;
     layer3_out[564] <= ~layer2_out[441] | layer2_out[442];
     layer3_out[565] <= ~layer2_out[342];
     layer3_out[566] <= layer2_out[949];
     layer3_out[567] <= layer2_out[60] & layer2_out[61];
     layer3_out[568] <= layer2_out[100] & layer2_out[101];
     layer3_out[569] <= layer2_out[1276];
     layer3_out[570] <= 1'b1;
     layer3_out[571] <= ~layer2_out[1395] | layer2_out[1396];
     layer3_out[572] <= 1'b1;
     layer3_out[573] <= layer2_out[118];
     layer3_out[574] <= layer2_out[355] & layer2_out[356];
     layer3_out[575] <= layer2_out[146] & ~layer2_out[147];
     layer3_out[576] <= ~(layer2_out[524] & layer2_out[525]);
     layer3_out[577] <= layer2_out[376];
     layer3_out[578] <= layer2_out[1484];
     layer3_out[579] <= ~layer2_out[1158];
     layer3_out[580] <= layer2_out[632];
     layer3_out[581] <= layer2_out[1248] | layer2_out[1249];
     layer3_out[582] <= ~layer2_out[557];
     layer3_out[583] <= 1'b0;
     layer3_out[584] <= 1'b1;
     layer3_out[585] <= ~layer2_out[1307];
     layer3_out[586] <= layer2_out[97] & layer2_out[98];
     layer3_out[587] <= 1'b0;
     layer3_out[588] <= layer2_out[1402] & ~layer2_out[1401];
     layer3_out[589] <= 1'b0;
     layer3_out[590] <= 1'b0;
     layer3_out[591] <= ~layer2_out[656];
     layer3_out[592] <= 1'b0;
     layer3_out[593] <= layer2_out[1133] & ~layer2_out[1134];
     layer3_out[594] <= 1'b0;
     layer3_out[595] <= ~layer2_out[233] | layer2_out[232];
     layer3_out[596] <= layer2_out[503] & ~layer2_out[504];
     layer3_out[597] <= ~layer2_out[164] | layer2_out[165];
     layer3_out[598] <= layer2_out[32] | layer2_out[33];
     layer3_out[599] <= ~(layer2_out[988] | layer2_out[989]);
     layer3_out[600] <= 1'b1;
     layer3_out[601] <= ~layer2_out[371];
     layer3_out[602] <= ~(layer2_out[1419] | layer2_out[1420]);
     layer3_out[603] <= ~layer2_out[685];
     layer3_out[604] <= layer2_out[697] | layer2_out[698];
     layer3_out[605] <= ~layer2_out[377];
     layer3_out[606] <= 1'b1;
     layer3_out[607] <= ~layer2_out[2] | layer2_out[1];
     layer3_out[608] <= ~layer2_out[1174];
     layer3_out[609] <= ~(layer2_out[690] & layer2_out[691]);
     layer3_out[610] <= 1'b0;
     layer3_out[611] <= ~layer2_out[264];
     layer3_out[612] <= layer2_out[1119] | layer2_out[1120];
     layer3_out[613] <= ~(layer2_out[181] ^ layer2_out[182]);
     layer3_out[614] <= layer2_out[419] | layer2_out[420];
     layer3_out[615] <= ~layer2_out[891];
     layer3_out[616] <= layer2_out[98] ^ layer2_out[99];
     layer3_out[617] <= ~layer2_out[612];
     layer3_out[618] <= layer2_out[350] & ~layer2_out[349];
     layer3_out[619] <= 1'b1;
     layer3_out[620] <= ~(layer2_out[1482] & layer2_out[1483]);
     layer3_out[621] <= 1'b1;
     layer3_out[622] <= layer2_out[1389];
     layer3_out[623] <= layer2_out[903];
     layer3_out[624] <= 1'b0;
     layer3_out[625] <= ~layer2_out[1446];
     layer3_out[626] <= layer2_out[468] | layer2_out[469];
     layer3_out[627] <= layer2_out[1329] & ~layer2_out[1330];
     layer3_out[628] <= ~layer2_out[1169];
     layer3_out[629] <= layer2_out[457] | layer2_out[458];
     layer3_out[630] <= ~layer2_out[802];
     layer3_out[631] <= layer2_out[473] | layer2_out[474];
     layer3_out[632] <= ~layer2_out[1473] | layer2_out[1472];
     layer3_out[633] <= layer2_out[1351] & layer2_out[1352];
     layer3_out[634] <= ~layer2_out[1088] | layer2_out[1089];
     layer3_out[635] <= ~layer2_out[1401] | layer2_out[1400];
     layer3_out[636] <= 1'b0;
     layer3_out[637] <= ~layer2_out[207] | layer2_out[208];
     layer3_out[638] <= 1'b1;
     layer3_out[639] <= ~(layer2_out[608] & layer2_out[609]);
     layer3_out[640] <= ~layer2_out[254] | layer2_out[253];
     layer3_out[641] <= ~layer2_out[784];
     layer3_out[642] <= ~(layer2_out[933] | layer2_out[934]);
     layer3_out[643] <= layer2_out[1314];
     layer3_out[644] <= ~(layer2_out[1422] & layer2_out[1423]);
     layer3_out[645] <= 1'b0;
     layer3_out[646] <= layer2_out[1288] & ~layer2_out[1289];
     layer3_out[647] <= layer2_out[44] ^ layer2_out[45];
     layer3_out[648] <= ~layer2_out[408] | layer2_out[409];
     layer3_out[649] <= layer2_out[320] | layer2_out[321];
     layer3_out[650] <= layer2_out[223] | layer2_out[224];
     layer3_out[651] <= ~layer2_out[582];
     layer3_out[652] <= ~layer2_out[1428] | layer2_out[1427];
     layer3_out[653] <= ~layer2_out[1325];
     layer3_out[654] <= ~layer2_out[1070];
     layer3_out[655] <= 1'b0;
     layer3_out[656] <= layer2_out[259] & layer2_out[260];
     layer3_out[657] <= ~layer2_out[884];
     layer3_out[658] <= layer2_out[1157] & ~layer2_out[1156];
     layer3_out[659] <= ~layer2_out[1302];
     layer3_out[660] <= ~layer2_out[1197];
     layer3_out[661] <= ~layer2_out[774] | layer2_out[773];
     layer3_out[662] <= 1'b0;
     layer3_out[663] <= layer2_out[590] | layer2_out[591];
     layer3_out[664] <= layer2_out[1269] | layer2_out[1270];
     layer3_out[665] <= layer2_out[714] & layer2_out[715];
     layer3_out[666] <= layer2_out[233];
     layer3_out[667] <= layer2_out[351] | layer2_out[352];
     layer3_out[668] <= layer2_out[879] & ~layer2_out[878];
     layer3_out[669] <= 1'b0;
     layer3_out[670] <= ~(layer2_out[1165] | layer2_out[1166]);
     layer3_out[671] <= 1'b0;
     layer3_out[672] <= layer2_out[666] & ~layer2_out[665];
     layer3_out[673] <= ~layer2_out[709];
     layer3_out[674] <= 1'b1;
     layer3_out[675] <= layer2_out[938];
     layer3_out[676] <= ~layer2_out[1283];
     layer3_out[677] <= 1'b0;
     layer3_out[678] <= ~(layer2_out[216] & layer2_out[217]);
     layer3_out[679] <= 1'b1;
     layer3_out[680] <= 1'b0;
     layer3_out[681] <= layer2_out[1386] & layer2_out[1387];
     layer3_out[682] <= ~layer2_out[136] | layer2_out[135];
     layer3_out[683] <= ~(layer2_out[1466] & layer2_out[1467]);
     layer3_out[684] <= ~(layer2_out[1434] | layer2_out[1435]);
     layer3_out[685] <= ~layer2_out[427];
     layer3_out[686] <= layer2_out[361] & ~layer2_out[360];
     layer3_out[687] <= layer2_out[1163] & ~layer2_out[1162];
     layer3_out[688] <= ~(layer2_out[1493] & layer2_out[1494]);
     layer3_out[689] <= ~layer2_out[941];
     layer3_out[690] <= layer2_out[318] | layer2_out[319];
     layer3_out[691] <= ~(layer2_out[374] | layer2_out[375]);
     layer3_out[692] <= ~(layer2_out[1138] & layer2_out[1139]);
     layer3_out[693] <= ~layer2_out[1149] | layer2_out[1148];
     layer3_out[694] <= ~(layer2_out[921] & layer2_out[922]);
     layer3_out[695] <= 1'b1;
     layer3_out[696] <= layer2_out[414];
     layer3_out[697] <= 1'b1;
     layer3_out[698] <= 1'b0;
     layer3_out[699] <= ~layer2_out[839];
     layer3_out[700] <= 1'b1;
     layer3_out[701] <= layer2_out[405] & ~layer2_out[406];
     layer3_out[702] <= layer2_out[225] & ~layer2_out[224];
     layer3_out[703] <= ~(layer2_out[970] & layer2_out[971]);
     layer3_out[704] <= ~(layer2_out[785] & layer2_out[786]);
     layer3_out[705] <= ~layer2_out[1190] | layer2_out[1191];
     layer3_out[706] <= ~layer2_out[975];
     layer3_out[707] <= layer2_out[727] & ~layer2_out[728];
     layer3_out[708] <= layer2_out[242] & ~layer2_out[241];
     layer3_out[709] <= layer2_out[959];
     layer3_out[710] <= ~layer2_out[560];
     layer3_out[711] <= layer2_out[170] & ~layer2_out[171];
     layer3_out[712] <= ~layer2_out[1259];
     layer3_out[713] <= ~layer2_out[1084] | layer2_out[1083];
     layer3_out[714] <= ~(layer2_out[1320] | layer2_out[1321]);
     layer3_out[715] <= 1'b0;
     layer3_out[716] <= layer2_out[740] & ~layer2_out[741];
     layer3_out[717] <= ~layer2_out[1309];
     layer3_out[718] <= layer2_out[762] | layer2_out[763];
     layer3_out[719] <= ~(layer2_out[1032] & layer2_out[1033]);
     layer3_out[720] <= ~layer2_out[201];
     layer3_out[721] <= ~(layer2_out[52] | layer2_out[53]);
     layer3_out[722] <= layer2_out[221] & ~layer2_out[220];
     layer3_out[723] <= 1'b1;
     layer3_out[724] <= 1'b1;
     layer3_out[725] <= layer2_out[1084] & ~layer2_out[1085];
     layer3_out[726] <= layer2_out[205];
     layer3_out[727] <= layer2_out[983] | layer2_out[984];
     layer3_out[728] <= ~(layer2_out[348] & layer2_out[349]);
     layer3_out[729] <= ~layer2_out[290];
     layer3_out[730] <= ~layer2_out[707] | layer2_out[706];
     layer3_out[731] <= 1'b1;
     layer3_out[732] <= layer2_out[562] | layer2_out[563];
     layer3_out[733] <= ~(layer2_out[940] ^ layer2_out[941]);
     layer3_out[734] <= ~(layer2_out[1323] ^ layer2_out[1324]);
     layer3_out[735] <= ~(layer2_out[228] ^ layer2_out[229]);
     layer3_out[736] <= layer2_out[926] & ~layer2_out[925];
     layer3_out[737] <= ~layer2_out[472];
     layer3_out[738] <= ~(layer2_out[240] | layer2_out[241]);
     layer3_out[739] <= 1'b0;
     layer3_out[740] <= layer2_out[804];
     layer3_out[741] <= layer2_out[1019];
     layer3_out[742] <= ~(layer2_out[1017] ^ layer2_out[1018]);
     layer3_out[743] <= ~layer2_out[789];
     layer3_out[744] <= layer2_out[448] & ~layer2_out[449];
     layer3_out[745] <= ~(layer2_out[1397] | layer2_out[1398]);
     layer3_out[746] <= ~layer2_out[115] | layer2_out[116];
     layer3_out[747] <= layer2_out[903] & ~layer2_out[904];
     layer3_out[748] <= ~layer2_out[1003];
     layer3_out[749] <= ~(layer2_out[1285] | layer2_out[1286]);
     layer3_out[750] <= ~layer2_out[975];
     layer3_out[751] <= layer2_out[1336] & ~layer2_out[1337];
     layer3_out[752] <= layer2_out[1048] ^ layer2_out[1049];
     layer3_out[753] <= layer2_out[1393];
     layer3_out[754] <= 1'b0;
     layer3_out[755] <= ~layer2_out[1150] | layer2_out[1149];
     layer3_out[756] <= layer2_out[1355] & layer2_out[1356];
     layer3_out[757] <= layer2_out[592];
     layer3_out[758] <= layer2_out[1179];
     layer3_out[759] <= 1'b0;
     layer3_out[760] <= ~layer2_out[1040] | layer2_out[1039];
     layer3_out[761] <= 1'b1;
     layer3_out[762] <= ~(layer2_out[1244] & layer2_out[1245]);
     layer3_out[763] <= ~layer2_out[213] | layer2_out[214];
     layer3_out[764] <= ~layer2_out[1117];
     layer3_out[765] <= layer2_out[1327] | layer2_out[1328];
     layer3_out[766] <= ~(layer2_out[180] | layer2_out[181]);
     layer3_out[767] <= 1'b1;
     layer3_out[768] <= ~layer2_out[1497];
     layer3_out[769] <= layer2_out[41] & layer2_out[42];
     layer3_out[770] <= ~(layer2_out[588] | layer2_out[589]);
     layer3_out[771] <= layer2_out[8] & ~layer2_out[7];
     layer3_out[772] <= layer2_out[77] & ~layer2_out[78];
     layer3_out[773] <= ~(layer2_out[1131] & layer2_out[1132]);
     layer3_out[774] <= ~layer2_out[1017] | layer2_out[1016];
     layer3_out[775] <= 1'b0;
     layer3_out[776] <= layer2_out[182] & layer2_out[183];
     layer3_out[777] <= layer2_out[1069];
     layer3_out[778] <= layer2_out[516] ^ layer2_out[517];
     layer3_out[779] <= layer2_out[389] & ~layer2_out[388];
     layer3_out[780] <= layer2_out[299] & ~layer2_out[298];
     layer3_out[781] <= layer2_out[422] & layer2_out[423];
     layer3_out[782] <= ~(layer2_out[624] & layer2_out[625]);
     layer3_out[783] <= layer2_out[599] | layer2_out[600];
     layer3_out[784] <= layer2_out[1350];
     layer3_out[785] <= ~layer2_out[202];
     layer3_out[786] <= ~layer2_out[1325];
     layer3_out[787] <= ~(layer2_out[1238] & layer2_out[1239]);
     layer3_out[788] <= ~(layer2_out[280] | layer2_out[281]);
     layer3_out[789] <= ~layer2_out[749];
     layer3_out[790] <= 1'b0;
     layer3_out[791] <= layer2_out[1250];
     layer3_out[792] <= ~layer2_out[117] | layer2_out[116];
     layer3_out[793] <= layer2_out[934] | layer2_out[935];
     layer3_out[794] <= layer2_out[1065] & layer2_out[1066];
     layer3_out[795] <= ~layer2_out[1236];
     layer3_out[796] <= layer2_out[1394];
     layer3_out[797] <= layer2_out[1150] & ~layer2_out[1151];
     layer3_out[798] <= layer2_out[507];
     layer3_out[799] <= layer2_out[694];
     layer3_out[800] <= layer2_out[1216] & ~layer2_out[1217];
     layer3_out[801] <= layer2_out[200];
     layer3_out[802] <= ~layer2_out[390];
     layer3_out[803] <= 1'b1;
     layer3_out[804] <= ~layer2_out[373] | layer2_out[372];
     layer3_out[805] <= 1'b1;
     layer3_out[806] <= layer2_out[0];
     layer3_out[807] <= layer2_out[1364] | layer2_out[1365];
     layer3_out[808] <= ~layer2_out[564];
     layer3_out[809] <= ~(layer2_out[479] | layer2_out[480]);
     layer3_out[810] <= 1'b0;
     layer3_out[811] <= ~(layer2_out[485] & layer2_out[486]);
     layer3_out[812] <= layer2_out[128] & layer2_out[129];
     layer3_out[813] <= ~layer2_out[805];
     layer3_out[814] <= 1'b1;
     layer3_out[815] <= 1'b1;
     layer3_out[816] <= ~(layer2_out[1467] | layer2_out[1468]);
     layer3_out[817] <= layer2_out[190] & layer2_out[191];
     layer3_out[818] <= ~layer2_out[967];
     layer3_out[819] <= ~(layer2_out[492] & layer2_out[493]);
     layer3_out[820] <= ~layer2_out[1171] | layer2_out[1172];
     layer3_out[821] <= layer2_out[230];
     layer3_out[822] <= layer2_out[827] & ~layer2_out[826];
     layer3_out[823] <= ~layer2_out[18] | layer2_out[19];
     layer3_out[824] <= 1'b0;
     layer3_out[825] <= layer2_out[458];
     layer3_out[826] <= layer2_out[1152] & ~layer2_out[1153];
     layer3_out[827] <= 1'b0;
     layer3_out[828] <= ~(layer2_out[396] & layer2_out[397]);
     layer3_out[829] <= 1'b1;
     layer3_out[830] <= layer2_out[1179];
     layer3_out[831] <= layer2_out[104];
     layer3_out[832] <= 1'b1;
     layer3_out[833] <= ~layer2_out[723] | layer2_out[722];
     layer3_out[834] <= layer2_out[704];
     layer3_out[835] <= layer2_out[720] ^ layer2_out[721];
     layer3_out[836] <= ~layer2_out[1028] | layer2_out[1027];
     layer3_out[837] <= 1'b1;
     layer3_out[838] <= layer2_out[324] ^ layer2_out[325];
     layer3_out[839] <= ~(layer2_out[358] & layer2_out[359]);
     layer3_out[840] <= 1'b1;
     layer3_out[841] <= layer2_out[1472] & ~layer2_out[1471];
     layer3_out[842] <= 1'b1;
     layer3_out[843] <= 1'b0;
     layer3_out[844] <= ~(layer2_out[1470] | layer2_out[1471]);
     layer3_out[845] <= layer2_out[155] & ~layer2_out[156];
     layer3_out[846] <= layer2_out[547] | layer2_out[548];
     layer3_out[847] <= ~(layer2_out[304] | layer2_out[305]);
     layer3_out[848] <= ~layer2_out[765];
     layer3_out[849] <= layer2_out[270] & ~layer2_out[269];
     layer3_out[850] <= layer2_out[90] | layer2_out[91];
     layer3_out[851] <= ~(layer2_out[1335] | layer2_out[1336]);
     layer3_out[852] <= layer2_out[1139];
     layer3_out[853] <= ~layer2_out[438];
     layer3_out[854] <= layer2_out[891] | layer2_out[892];
     layer3_out[855] <= layer2_out[490] & ~layer2_out[491];
     layer3_out[856] <= layer2_out[860];
     layer3_out[857] <= ~(layer2_out[519] | layer2_out[520]);
     layer3_out[858] <= ~(layer2_out[412] | layer2_out[413]);
     layer3_out[859] <= ~layer2_out[79];
     layer3_out[860] <= layer2_out[1049];
     layer3_out[861] <= layer2_out[1204];
     layer3_out[862] <= ~layer2_out[228] | layer2_out[227];
     layer3_out[863] <= ~(layer2_out[1168] & layer2_out[1169]);
     layer3_out[864] <= ~(layer2_out[581] | layer2_out[582]);
     layer3_out[865] <= ~layer2_out[788];
     layer3_out[866] <= 1'b1;
     layer3_out[867] <= ~(layer2_out[1391] & layer2_out[1392]);
     layer3_out[868] <= layer2_out[556];
     layer3_out[869] <= 1'b0;
     layer3_out[870] <= ~layer2_out[1095] | layer2_out[1094];
     layer3_out[871] <= ~layer2_out[1271] | layer2_out[1270];
     layer3_out[872] <= ~(layer2_out[378] | layer2_out[379]);
     layer3_out[873] <= ~layer2_out[551] | layer2_out[550];
     layer3_out[874] <= ~layer2_out[759] | layer2_out[760];
     layer3_out[875] <= ~layer2_out[218];
     layer3_out[876] <= layer2_out[356] & ~layer2_out[357];
     layer3_out[877] <= 1'b1;
     layer3_out[878] <= 1'b1;
     layer3_out[879] <= ~layer2_out[554] | layer2_out[555];
     layer3_out[880] <= layer2_out[983] & ~layer2_out[982];
     layer3_out[881] <= layer2_out[1226] & ~layer2_out[1225];
     layer3_out[882] <= ~layer2_out[168];
     layer3_out[883] <= 1'b1;
     layer3_out[884] <= layer2_out[1314];
     layer3_out[885] <= layer2_out[188];
     layer3_out[886] <= ~layer2_out[1406] | layer2_out[1405];
     layer3_out[887] <= 1'b0;
     layer3_out[888] <= layer2_out[1001];
     layer3_out[889] <= ~(layer2_out[1185] & layer2_out[1186]);
     layer3_out[890] <= ~layer2_out[530] | layer2_out[529];
     layer3_out[891] <= ~(layer2_out[225] | layer2_out[226]);
     layer3_out[892] <= ~(layer2_out[204] | layer2_out[205]);
     layer3_out[893] <= layer2_out[211] & ~layer2_out[210];
     layer3_out[894] <= layer2_out[1208] & ~layer2_out[1209];
     layer3_out[895] <= layer2_out[963];
     layer3_out[896] <= 1'b0;
     layer3_out[897] <= ~(layer2_out[81] & layer2_out[82]);
     layer3_out[898] <= ~layer2_out[74];
     layer3_out[899] <= layer2_out[1374] | layer2_out[1375];
     layer3_out[900] <= ~layer2_out[1257];
     layer3_out[901] <= layer2_out[1052] & layer2_out[1053];
     layer3_out[902] <= ~(layer2_out[1299] | layer2_out[1300]);
     layer3_out[903] <= layer2_out[1458];
     layer3_out[904] <= layer2_out[1387] & layer2_out[1388];
     layer3_out[905] <= ~layer2_out[1210] | layer2_out[1211];
     layer3_out[906] <= ~layer2_out[124];
     layer3_out[907] <= layer2_out[908] ^ layer2_out[909];
     layer3_out[908] <= layer2_out[128] & ~layer2_out[127];
     layer3_out[909] <= ~(layer2_out[1257] & layer2_out[1258]);
     layer3_out[910] <= layer2_out[971];
     layer3_out[911] <= layer2_out[321] ^ layer2_out[322];
     layer3_out[912] <= ~(layer2_out[1236] & layer2_out[1237]);
     layer3_out[913] <= ~layer2_out[742] | layer2_out[741];
     layer3_out[914] <= ~layer2_out[343];
     layer3_out[915] <= layer2_out[1215];
     layer3_out[916] <= layer2_out[303];
     layer3_out[917] <= ~(layer2_out[802] ^ layer2_out[803]);
     layer3_out[918] <= layer2_out[681] & ~layer2_out[680];
     layer3_out[919] <= layer2_out[1229] & ~layer2_out[1228];
     layer3_out[920] <= layer2_out[1041];
     layer3_out[921] <= ~layer2_out[767];
     layer3_out[922] <= ~layer2_out[12] | layer2_out[13];
     layer3_out[923] <= layer2_out[380] & ~layer2_out[381];
     layer3_out[924] <= 1'b0;
     layer3_out[925] <= 1'b0;
     layer3_out[926] <= ~layer2_out[543] | layer2_out[544];
     layer3_out[927] <= layer2_out[218] | layer2_out[219];
     layer3_out[928] <= layer2_out[464] & ~layer2_out[465];
     layer3_out[929] <= 1'b1;
     layer3_out[930] <= layer2_out[758] & layer2_out[759];
     layer3_out[931] <= ~layer2_out[516] | layer2_out[515];
     layer3_out[932] <= ~layer2_out[1098] | layer2_out[1097];
     layer3_out[933] <= ~(layer2_out[1075] | layer2_out[1076]);
     layer3_out[934] <= layer2_out[1111] & ~layer2_out[1110];
     layer3_out[935] <= ~layer2_out[728];
     layer3_out[936] <= layer2_out[451];
     layer3_out[937] <= layer2_out[627];
     layer3_out[938] <= 1'b0;
     layer3_out[939] <= layer2_out[39];
     layer3_out[940] <= layer2_out[313] & ~layer2_out[314];
     layer3_out[941] <= layer2_out[724] & ~layer2_out[723];
     layer3_out[942] <= layer2_out[1436];
     layer3_out[943] <= ~(layer2_out[494] | layer2_out[495]);
     layer3_out[944] <= layer2_out[1044];
     layer3_out[945] <= ~(layer2_out[819] ^ layer2_out[820]);
     layer3_out[946] <= layer2_out[500];
     layer3_out[947] <= ~(layer2_out[409] & layer2_out[410]);
     layer3_out[948] <= layer2_out[1330];
     layer3_out[949] <= ~layer2_out[881] | layer2_out[880];
     layer3_out[950] <= layer2_out[659];
     layer3_out[951] <= layer2_out[197] | layer2_out[198];
     layer3_out[952] <= 1'b1;
     layer3_out[953] <= layer2_out[37];
     layer3_out[954] <= layer2_out[431];
     layer3_out[955] <= layer2_out[558] ^ layer2_out[559];
     layer3_out[956] <= 1'b0;
     layer3_out[957] <= ~layer2_out[772] | layer2_out[771];
     layer3_out[958] <= ~layer2_out[1346] | layer2_out[1345];
     layer3_out[959] <= layer2_out[735] & ~layer2_out[734];
     layer3_out[960] <= layer2_out[883] & ~layer2_out[882];
     layer3_out[961] <= ~layer2_out[1301] | layer2_out[1300];
     layer3_out[962] <= 1'b1;
     layer3_out[963] <= layer2_out[212];
     layer3_out[964] <= layer2_out[958] & ~layer2_out[957];
     layer3_out[965] <= ~(layer2_out[465] & layer2_out[466]);
     layer3_out[966] <= layer2_out[875] | layer2_out[876];
     layer3_out[967] <= layer2_out[221];
     layer3_out[968] <= layer2_out[957];
     layer3_out[969] <= ~(layer2_out[932] | layer2_out[933]);
     layer3_out[970] <= ~layer2_out[539] | layer2_out[538];
     layer3_out[971] <= ~layer2_out[1219];
     layer3_out[972] <= 1'b1;
     layer3_out[973] <= ~layer2_out[1007] | layer2_out[1008];
     layer3_out[974] <= ~layer2_out[1311];
     layer3_out[975] <= ~layer2_out[911];
     layer3_out[976] <= layer2_out[1261] & ~layer2_out[1262];
     layer3_out[977] <= ~(layer2_out[1289] & layer2_out[1290]);
     layer3_out[978] <= layer2_out[305] & ~layer2_out[306];
     layer3_out[979] <= ~layer2_out[668] | layer2_out[669];
     layer3_out[980] <= layer2_out[1115];
     layer3_out[981] <= ~layer2_out[74] | layer2_out[75];
     layer3_out[982] <= layer2_out[24] & ~layer2_out[23];
     layer3_out[983] <= ~(layer2_out[1274] ^ layer2_out[1275]);
     layer3_out[984] <= ~layer2_out[165];
     layer3_out[985] <= 1'b0;
     layer3_out[986] <= ~(layer2_out[989] & layer2_out[990]);
     layer3_out[987] <= ~(layer2_out[472] | layer2_out[473]);
     layer3_out[988] <= layer2_out[1059] | layer2_out[1060];
     layer3_out[989] <= layer2_out[140];
     layer3_out[990] <= ~layer2_out[668] | layer2_out[667];
     layer3_out[991] <= layer2_out[161] & ~layer2_out[160];
     layer3_out[992] <= layer2_out[1010];
     layer3_out[993] <= layer2_out[1235] & ~layer2_out[1234];
     layer3_out[994] <= layer2_out[1421] & layer2_out[1422];
     layer3_out[995] <= ~(layer2_out[1180] | layer2_out[1181]);
     layer3_out[996] <= layer2_out[1159] & ~layer2_out[1160];
     layer3_out[997] <= layer2_out[388];
     layer3_out[998] <= ~(layer2_out[1483] & layer2_out[1484]);
     layer3_out[999] <= layer2_out[506];
     layer3_out[1000] <= layer2_out[639];
     layer3_out[1001] <= layer2_out[443] & layer2_out[444];
     layer3_out[1002] <= layer2_out[55];
     layer3_out[1003] <= layer2_out[636] & ~layer2_out[635];
     layer3_out[1004] <= layer2_out[943];
     layer3_out[1005] <= 1'b0;
     layer3_out[1006] <= 1'b1;
     layer3_out[1007] <= ~layer2_out[1331];
     layer3_out[1008] <= layer2_out[194] & layer2_out[195];
     layer3_out[1009] <= ~(layer2_out[1224] & layer2_out[1225]);
     layer3_out[1010] <= layer2_out[25] & ~layer2_out[26];
     layer3_out[1011] <= ~(layer2_out[704] & layer2_out[705]);
     layer3_out[1012] <= ~layer2_out[1085];
     layer3_out[1013] <= layer2_out[767] & ~layer2_out[768];
     layer3_out[1014] <= ~layer2_out[961] | layer2_out[960];
     layer3_out[1015] <= layer2_out[1370];
     layer3_out[1016] <= ~layer2_out[1129];
     layer3_out[1017] <= ~(layer2_out[1410] | layer2_out[1411]);
     layer3_out[1018] <= ~layer2_out[1141] | layer2_out[1140];
     layer3_out[1019] <= layer2_out[1368] | layer2_out[1369];
     layer3_out[1020] <= 1'b0;
     layer3_out[1021] <= ~(layer2_out[1207] | layer2_out[1208]);
     layer3_out[1022] <= ~layer2_out[250];
     layer3_out[1023] <= ~(layer2_out[842] & layer2_out[843]);
     layer3_out[1024] <= ~layer2_out[142] | layer2_out[141];
     layer3_out[1025] <= ~layer2_out[1219];
     layer3_out[1026] <= layer2_out[748];
     layer3_out[1027] <= 1'b0;
     layer3_out[1028] <= layer2_out[782];
     layer3_out[1029] <= layer2_out[177] & layer2_out[178];
     layer3_out[1030] <= layer2_out[517] & ~layer2_out[518];
     layer3_out[1031] <= 1'b1;
     layer3_out[1032] <= layer2_out[1060] & ~layer2_out[1061];
     layer3_out[1033] <= ~layer2_out[1252];
     layer3_out[1034] <= layer2_out[804] & layer2_out[805];
     layer3_out[1035] <= ~layer2_out[1044] | layer2_out[1043];
     layer3_out[1036] <= ~layer2_out[594] | layer2_out[595];
     layer3_out[1037] <= layer2_out[866];
     layer3_out[1038] <= 1'b1;
     layer3_out[1039] <= layer2_out[1292] & ~layer2_out[1291];
     layer3_out[1040] <= ~layer2_out[607] | layer2_out[606];
     layer3_out[1041] <= layer2_out[175] & ~layer2_out[174];
     layer3_out[1042] <= layer2_out[454];
     layer3_out[1043] <= layer2_out[176];
     layer3_out[1044] <= layer2_out[748];
     layer3_out[1045] <= ~layer2_out[297];
     layer3_out[1046] <= layer2_out[823] | layer2_out[824];
     layer3_out[1047] <= ~(layer2_out[226] & layer2_out[227]);
     layer3_out[1048] <= layer2_out[699] & layer2_out[700];
     layer3_out[1049] <= 1'b0;
     layer3_out[1050] <= layer2_out[1125] & ~layer2_out[1126];
     layer3_out[1051] <= ~(layer2_out[1409] | layer2_out[1410]);
     layer3_out[1052] <= 1'b0;
     layer3_out[1053] <= layer2_out[726] & ~layer2_out[725];
     layer3_out[1054] <= layer2_out[818] & ~layer2_out[817];
     layer3_out[1055] <= layer2_out[1226] & ~layer2_out[1227];
     layer3_out[1056] <= layer2_out[820];
     layer3_out[1057] <= layer2_out[794] & layer2_out[795];
     layer3_out[1058] <= ~layer2_out[1215];
     layer3_out[1059] <= layer2_out[382] & ~layer2_out[381];
     layer3_out[1060] <= layer2_out[1067] | layer2_out[1068];
     layer3_out[1061] <= layer2_out[130] | layer2_out[131];
     layer3_out[1062] <= layer2_out[347];
     layer3_out[1063] <= layer2_out[825];
     layer3_out[1064] <= ~(layer2_out[603] & layer2_out[604]);
     layer3_out[1065] <= 1'b1;
     layer3_out[1066] <= layer2_out[239] & ~layer2_out[240];
     layer3_out[1067] <= layer2_out[1403];
     layer3_out[1068] <= ~layer2_out[828];
     layer3_out[1069] <= layer2_out[499];
     layer3_out[1070] <= layer2_out[107] & layer2_out[108];
     layer3_out[1071] <= layer2_out[555];
     layer3_out[1072] <= ~layer2_out[868] | layer2_out[867];
     layer3_out[1073] <= layer2_out[446];
     layer3_out[1074] <= ~(layer2_out[779] | layer2_out[780]);
     layer3_out[1075] <= layer2_out[1020] & layer2_out[1021];
     layer3_out[1076] <= ~layer2_out[468];
     layer3_out[1077] <= layer2_out[238] & ~layer2_out[239];
     layer3_out[1078] <= ~layer2_out[190] | layer2_out[189];
     layer3_out[1079] <= layer2_out[1357];
     layer3_out[1080] <= layer2_out[310] & ~layer2_out[311];
     layer3_out[1081] <= ~layer2_out[913] | layer2_out[912];
     layer3_out[1082] <= layer2_out[965] | layer2_out[966];
     layer3_out[1083] <= ~layer2_out[1099];
     layer3_out[1084] <= layer2_out[702] & layer2_out[703];
     layer3_out[1085] <= ~(layer2_out[1485] & layer2_out[1486]);
     layer3_out[1086] <= ~(layer2_out[1281] & layer2_out[1282]);
     layer3_out[1087] <= ~(layer2_out[778] | layer2_out[779]);
     layer3_out[1088] <= ~(layer2_out[658] & layer2_out[659]);
     layer3_out[1089] <= ~layer2_out[49];
     layer3_out[1090] <= ~(layer2_out[391] | layer2_out[392]);
     layer3_out[1091] <= 1'b1;
     layer3_out[1092] <= 1'b0;
     layer3_out[1093] <= 1'b0;
     layer3_out[1094] <= ~layer2_out[1488] | layer2_out[1487];
     layer3_out[1095] <= layer2_out[597] & ~layer2_out[596];
     layer3_out[1096] <= ~layer2_out[994];
     layer3_out[1097] <= ~layer2_out[633] | layer2_out[634];
     layer3_out[1098] <= ~(layer2_out[1294] | layer2_out[1295]);
     layer3_out[1099] <= layer2_out[63] & ~layer2_out[64];
     layer3_out[1100] <= layer2_out[1479] & ~layer2_out[1480];
     layer3_out[1101] <= layer2_out[478] & layer2_out[479];
     layer3_out[1102] <= layer2_out[553];
     layer3_out[1103] <= layer2_out[1249] | layer2_out[1250];
     layer3_out[1104] <= ~layer2_out[1416] | layer2_out[1417];
     layer3_out[1105] <= ~layer2_out[1007] | layer2_out[1006];
     layer3_out[1106] <= layer2_out[169];
     layer3_out[1107] <= ~(layer2_out[984] | layer2_out[985]);
     layer3_out[1108] <= ~layer2_out[588] | layer2_out[587];
     layer3_out[1109] <= layer2_out[926] & layer2_out[927];
     layer3_out[1110] <= layer2_out[1130] | layer2_out[1131];
     layer3_out[1111] <= layer2_out[1152] & ~layer2_out[1151];
     layer3_out[1112] <= ~layer2_out[569];
     layer3_out[1113] <= layer2_out[685];
     layer3_out[1114] <= ~(layer2_out[636] | layer2_out[637]);
     layer3_out[1115] <= ~layer2_out[1417] | layer2_out[1418];
     layer3_out[1116] <= 1'b0;
     layer3_out[1117] <= layer2_out[443] & ~layer2_out[442];
     layer3_out[1118] <= 1'b0;
     layer3_out[1119] <= ~layer2_out[1024];
     layer3_out[1120] <= ~layer2_out[195];
     layer3_out[1121] <= ~(layer2_out[1394] & layer2_out[1395]);
     layer3_out[1122] <= layer2_out[415];
     layer3_out[1123] <= layer2_out[674] & layer2_out[675];
     layer3_out[1124] <= layer2_out[451];
     layer3_out[1125] <= layer2_out[835];
     layer3_out[1126] <= layer2_out[916];
     layer3_out[1127] <= ~layer2_out[873];
     layer3_out[1128] <= layer2_out[1347] | layer2_out[1348];
     layer3_out[1129] <= ~layer2_out[184];
     layer3_out[1130] <= ~(layer2_out[254] & layer2_out[255]);
     layer3_out[1131] <= layer2_out[721] | layer2_out[722];
     layer3_out[1132] <= layer2_out[849] | layer2_out[850];
     layer3_out[1133] <= ~layer2_out[433];
     layer3_out[1134] <= ~layer2_out[490] | layer2_out[489];
     layer3_out[1135] <= layer2_out[435] & ~layer2_out[434];
     layer3_out[1136] <= ~(layer2_out[530] | layer2_out[531]);
     layer3_out[1137] <= ~layer2_out[123] | layer2_out[124];
     layer3_out[1138] <= layer2_out[541];
     layer3_out[1139] <= ~layer2_out[754];
     layer3_out[1140] <= layer2_out[1074] & ~layer2_out[1073];
     layer3_out[1141] <= layer2_out[1122] & layer2_out[1123];
     layer3_out[1142] <= layer2_out[1081];
     layer3_out[1143] <= layer2_out[1072];
     layer3_out[1144] <= ~layer2_out[1475] | layer2_out[1476];
     layer3_out[1145] <= ~layer2_out[338] | layer2_out[337];
     layer3_out[1146] <= layer2_out[1184] & ~layer2_out[1185];
     layer3_out[1147] <= 1'b0;
     layer3_out[1148] <= layer2_out[1273] & layer2_out[1274];
     layer3_out[1149] <= layer2_out[129] & ~layer2_out[130];
     layer3_out[1150] <= 1'b0;
     layer3_out[1151] <= layer2_out[846];
     layer3_out[1152] <= ~layer2_out[1222] | layer2_out[1221];
     layer3_out[1153] <= 1'b0;
     layer3_out[1154] <= layer2_out[67] & ~layer2_out[66];
     layer3_out[1155] <= layer2_out[37] & ~layer2_out[36];
     layer3_out[1156] <= layer2_out[81];
     layer3_out[1157] <= layer2_out[532] | layer2_out[533];
     layer3_out[1158] <= layer2_out[1030] & layer2_out[1031];
     layer3_out[1159] <= layer2_out[1022] & ~layer2_out[1023];
     layer3_out[1160] <= layer2_out[537] ^ layer2_out[538];
     layer3_out[1161] <= layer2_out[1066] | layer2_out[1067];
     layer3_out[1162] <= ~(layer2_out[1337] & layer2_out[1338]);
     layer3_out[1163] <= layer2_out[695] & layer2_out[696];
     layer3_out[1164] <= 1'b1;
     layer3_out[1165] <= 1'b0;
     layer3_out[1166] <= layer2_out[495] & ~layer2_out[496];
     layer3_out[1167] <= ~layer2_out[481] | layer2_out[480];
     layer3_out[1168] <= layer2_out[1494];
     layer3_out[1169] <= layer2_out[1281];
     layer3_out[1170] <= 1'b1;
     layer3_out[1171] <= layer2_out[920] | layer2_out[921];
     layer3_out[1172] <= layer2_out[1056] | layer2_out[1057];
     layer3_out[1173] <= layer2_out[809] | layer2_out[810];
     layer3_out[1174] <= ~layer2_out[1342] | layer2_out[1341];
     layer3_out[1175] <= 1'b1;
     layer3_out[1176] <= 1'b0;
     layer3_out[1177] <= layer2_out[408] & ~layer2_out[407];
     layer3_out[1178] <= ~layer2_out[1479];
     layer3_out[1179] <= ~layer2_out[1374];
     layer3_out[1180] <= ~(layer2_out[58] | layer2_out[59]);
     layer3_out[1181] <= layer2_out[282] & layer2_out[283];
     layer3_out[1182] <= 1'b1;
     layer3_out[1183] <= layer2_out[1036] & ~layer2_out[1035];
     layer3_out[1184] <= layer2_out[27] & ~layer2_out[26];
     layer3_out[1185] <= layer2_out[3];
     layer3_out[1186] <= ~(layer2_out[1342] | layer2_out[1343]);
     layer3_out[1187] <= layer2_out[153] & layer2_out[154];
     layer3_out[1188] <= 1'b1;
     layer3_out[1189] <= layer2_out[4];
     layer3_out[1190] <= ~(layer2_out[1053] & layer2_out[1054]);
     layer3_out[1191] <= ~layer2_out[426];
     layer3_out[1192] <= ~(layer2_out[143] & layer2_out[144]);
     layer3_out[1193] <= layer2_out[394] ^ layer2_out[395];
     layer3_out[1194] <= layer2_out[924] | layer2_out[925];
     layer3_out[1195] <= layer2_out[1008] & ~layer2_out[1009];
     layer3_out[1196] <= layer2_out[262];
     layer3_out[1197] <= layer2_out[432] | layer2_out[433];
     layer3_out[1198] <= ~layer2_out[96] | layer2_out[97];
     layer3_out[1199] <= ~(layer2_out[343] & layer2_out[344]);
     layer3_out[1200] <= layer2_out[1050] ^ layer2_out[1051];
     layer3_out[1201] <= layer2_out[1203];
     layer3_out[1202] <= 1'b1;
     layer3_out[1203] <= layer2_out[1449];
     layer3_out[1204] <= ~(layer2_out[22] ^ layer2_out[23]);
     layer3_out[1205] <= layer2_out[996];
     layer3_out[1206] <= 1'b1;
     layer3_out[1207] <= ~(layer2_out[637] & layer2_out[638]);
     layer3_out[1208] <= ~layer2_out[1172];
     layer3_out[1209] <= ~(layer2_out[1194] & layer2_out[1195]);
     layer3_out[1210] <= 1'b1;
     layer3_out[1211] <= ~layer2_out[1034] | layer2_out[1035];
     layer3_out[1212] <= layer2_out[946];
     layer3_out[1213] <= ~layer2_out[738] | layer2_out[739];
     layer3_out[1214] <= layer2_out[84] & ~layer2_out[83];
     layer3_out[1215] <= layer2_out[643];
     layer3_out[1216] <= ~layer2_out[836];
     layer3_out[1217] <= layer2_out[648] & layer2_out[649];
     layer3_out[1218] <= layer2_out[573] & layer2_out[574];
     layer3_out[1219] <= ~layer2_out[614];
     layer3_out[1220] <= 1'b1;
     layer3_out[1221] <= ~(layer2_out[1011] & layer2_out[1012]);
     layer3_out[1222] <= 1'b0;
     layer3_out[1223] <= ~layer2_out[431] | layer2_out[430];
     layer3_out[1224] <= ~layer2_out[839];
     layer3_out[1225] <= ~layer2_out[498];
     layer3_out[1226] <= layer2_out[1005] & layer2_out[1006];
     layer3_out[1227] <= ~(layer2_out[1443] & layer2_out[1444]);
     layer3_out[1228] <= ~layer2_out[143] | layer2_out[142];
     layer3_out[1229] <= layer2_out[294];
     layer3_out[1230] <= ~layer2_out[1278] | layer2_out[1279];
     layer3_out[1231] <= layer2_out[1473] & ~layer2_out[1474];
     layer3_out[1232] <= 1'b1;
     layer3_out[1233] <= layer2_out[103] & layer2_out[104];
     layer3_out[1234] <= layer2_out[789] & layer2_out[790];
     layer3_out[1235] <= ~(layer2_out[1051] & layer2_out[1052]);
     layer3_out[1236] <= layer2_out[456];
     layer3_out[1237] <= layer2_out[1240] & ~layer2_out[1241];
     layer3_out[1238] <= layer2_out[3] ^ layer2_out[4];
     layer3_out[1239] <= layer2_out[1423];
     layer3_out[1240] <= layer2_out[638] & layer2_out[639];
     layer3_out[1241] <= 1'b0;
     layer3_out[1242] <= layer2_out[172];
     layer3_out[1243] <= layer2_out[1459];
     layer3_out[1244] <= layer2_out[1457];
     layer3_out[1245] <= layer2_out[192] & layer2_out[193];
     layer3_out[1246] <= ~layer2_out[282] | layer2_out[281];
     layer3_out[1247] <= layer2_out[1014];
     layer3_out[1248] <= layer2_out[482];
     layer3_out[1249] <= layer2_out[477] & ~layer2_out[478];
     layer3_out[1250] <= ~layer2_out[17];
     layer3_out[1251] <= layer2_out[774] | layer2_out[775];
     layer3_out[1252] <= ~(layer2_out[604] | layer2_out[605]);
     layer3_out[1253] <= ~layer2_out[1065];
     layer3_out[1254] <= layer2_out[198] & ~layer2_out[199];
     layer3_out[1255] <= layer2_out[1372] & ~layer2_out[1371];
     layer3_out[1256] <= ~layer2_out[1464];
     layer3_out[1257] <= layer2_out[1453] | layer2_out[1454];
     layer3_out[1258] <= 1'b0;
     layer3_out[1259] <= ~(layer2_out[1415] & layer2_out[1416]);
     layer3_out[1260] <= layer2_out[888];
     layer3_out[1261] <= layer2_out[507] & ~layer2_out[506];
     layer3_out[1262] <= layer2_out[447];
     layer3_out[1263] <= layer2_out[617] ^ layer2_out[618];
     layer3_out[1264] <= 1'b0;
     layer3_out[1265] <= ~(layer2_out[283] & layer2_out[284]);
     layer3_out[1266] <= ~layer2_out[513];
     layer3_out[1267] <= ~layer2_out[157];
     layer3_out[1268] <= ~layer2_out[462];
     layer3_out[1269] <= ~layer2_out[1069] | layer2_out[1070];
     layer3_out[1270] <= ~(layer2_out[1488] & layer2_out[1489]);
     layer3_out[1271] <= ~layer2_out[801] | layer2_out[800];
     layer3_out[1272] <= layer2_out[1298];
     layer3_out[1273] <= ~layer2_out[652] | layer2_out[653];
     layer3_out[1274] <= ~(layer2_out[916] & layer2_out[917]);
     layer3_out[1275] <= layer2_out[1388] & layer2_out[1389];
     layer3_out[1276] <= 1'b1;
     layer3_out[1277] <= ~layer2_out[6] | layer2_out[5];
     layer3_out[1278] <= ~(layer2_out[35] & layer2_out[36]);
     layer3_out[1279] <= layer2_out[1087];
     layer3_out[1280] <= ~(layer2_out[1265] & layer2_out[1266]);
     layer3_out[1281] <= ~layer2_out[1413] | layer2_out[1412];
     layer3_out[1282] <= ~(layer2_out[769] | layer2_out[770]);
     layer3_out[1283] <= ~layer2_out[799];
     layer3_out[1284] <= ~layer2_out[57];
     layer3_out[1285] <= 1'b1;
     layer3_out[1286] <= layer2_out[889] & layer2_out[890];
     layer3_out[1287] <= 1'b0;
     layer3_out[1288] <= layer2_out[1361] & ~layer2_out[1362];
     layer3_out[1289] <= layer2_out[1360] & ~layer2_out[1361];
     layer3_out[1290] <= ~layer2_out[310];
     layer3_out[1291] <= 1'b0;
     layer3_out[1292] <= layer2_out[177] & ~layer2_out[176];
     layer3_out[1293] <= layer2_out[768] | layer2_out[769];
     layer3_out[1294] <= layer2_out[278];
     layer3_out[1295] <= layer2_out[265] & layer2_out[266];
     layer3_out[1296] <= layer2_out[670] & ~layer2_out[671];
     layer3_out[1297] <= 1'b0;
     layer3_out[1298] <= ~layer2_out[464] | layer2_out[463];
     layer3_out[1299] <= ~layer2_out[695];
     layer3_out[1300] <= layer2_out[50] & ~layer2_out[49];
     layer3_out[1301] <= ~layer2_out[585] | layer2_out[584];
     layer3_out[1302] <= ~(layer2_out[782] | layer2_out[783]);
     layer3_out[1303] <= layer2_out[993] & ~layer2_out[992];
     layer3_out[1304] <= 1'b0;
     layer3_out[1305] <= layer2_out[1222] & ~layer2_out[1223];
     layer3_out[1306] <= layer2_out[647] & ~layer2_out[646];
     layer3_out[1307] <= ~layer2_out[1312] | layer2_out[1313];
     layer3_out[1308] <= layer2_out[624] & ~layer2_out[623];
     layer3_out[1309] <= ~(layer2_out[513] | layer2_out[514]);
     layer3_out[1310] <= layer2_out[185];
     layer3_out[1311] <= ~(layer2_out[57] & layer2_out[58]);
     layer3_out[1312] <= layer2_out[857] & ~layer2_out[856];
     layer3_out[1313] <= layer2_out[497] & ~layer2_out[496];
     layer3_out[1314] <= ~(layer2_out[786] & layer2_out[787]);
     layer3_out[1315] <= 1'b0;
     layer3_out[1316] <= ~(layer2_out[361] & layer2_out[362]);
     layer3_out[1317] <= ~layer2_out[1302] | layer2_out[1301];
     layer3_out[1318] <= 1'b1;
     layer3_out[1319] <= layer2_out[1323] & ~layer2_out[1322];
     layer3_out[1320] <= ~layer2_out[65] | layer2_out[64];
     layer3_out[1321] <= layer2_out[742] & layer2_out[743];
     layer3_out[1322] <= layer2_out[1115];
     layer3_out[1323] <= ~(layer2_out[328] ^ layer2_out[329]);
     layer3_out[1324] <= layer2_out[459] & layer2_out[460];
     layer3_out[1325] <= 1'b0;
     layer3_out[1326] <= ~layer2_out[731];
     layer3_out[1327] <= layer2_out[440] & ~layer2_out[441];
     layer3_out[1328] <= ~layer2_out[868] | layer2_out[869];
     layer3_out[1329] <= ~layer2_out[635] | layer2_out[634];
     layer3_out[1330] <= 1'b1;
     layer3_out[1331] <= ~layer2_out[1426] | layer2_out[1427];
     layer3_out[1332] <= 1'b1;
     layer3_out[1333] <= layer2_out[263] & layer2_out[264];
     layer3_out[1334] <= layer2_out[1359] & layer2_out[1360];
     layer3_out[1335] <= ~(layer2_out[1277] | layer2_out[1278]);
     layer3_out[1336] <= layer2_out[641];
     layer3_out[1337] <= ~layer2_out[654] | layer2_out[655];
     layer3_out[1338] <= layer2_out[950] & ~layer2_out[951];
     layer3_out[1339] <= ~(layer2_out[1192] | layer2_out[1193]);
     layer3_out[1340] <= ~layer2_out[877];
     layer3_out[1341] <= ~layer2_out[1184];
     layer3_out[1342] <= 1'b0;
     layer3_out[1343] <= layer2_out[334] & ~layer2_out[335];
     layer3_out[1344] <= layer2_out[855] | layer2_out[856];
     layer3_out[1345] <= ~(layer2_out[987] & layer2_out[988]);
     layer3_out[1346] <= layer2_out[615] & ~layer2_out[614];
     layer3_out[1347] <= layer2_out[732] | layer2_out[733];
     layer3_out[1348] <= ~layer2_out[320];
     layer3_out[1349] <= layer2_out[1411] & ~layer2_out[1412];
     layer3_out[1350] <= layer2_out[1408] & layer2_out[1409];
     layer3_out[1351] <= 1'b1;
     layer3_out[1352] <= ~layer2_out[1145];
     layer3_out[1353] <= ~layer2_out[1469] | layer2_out[1470];
     layer3_out[1354] <= ~layer2_out[1018];
     layer3_out[1355] <= ~layer2_out[716];
     layer3_out[1356] <= layer2_out[397] & ~layer2_out[398];
     layer3_out[1357] <= ~layer2_out[1377];
     layer3_out[1358] <= ~layer2_out[1339] | layer2_out[1340];
     layer3_out[1359] <= ~layer2_out[446];
     layer3_out[1360] <= ~layer2_out[324];
     layer3_out[1361] <= 1'b1;
     layer3_out[1362] <= ~(layer2_out[362] & layer2_out[363]);
     layer3_out[1363] <= layer2_out[267] & ~layer2_out[268];
     layer3_out[1364] <= ~(layer2_out[1431] & layer2_out[1432]);
     layer3_out[1365] <= 1'b1;
     layer3_out[1366] <= layer2_out[1446] & layer2_out[1447];
     layer3_out[1367] <= ~layer2_out[1224];
     layer3_out[1368] <= layer2_out[710];
     layer3_out[1369] <= ~layer2_out[837];
     layer3_out[1370] <= 1'b0;
     layer3_out[1371] <= ~layer2_out[1119];
     layer3_out[1372] <= ~layer2_out[145];
     layer3_out[1373] <= layer2_out[719];
     layer3_out[1374] <= layer2_out[1399] & ~layer2_out[1400];
     layer3_out[1375] <= ~layer2_out[86];
     layer3_out[1376] <= layer2_out[1026] | layer2_out[1027];
     layer3_out[1377] <= layer2_out[679] & ~layer2_out[678];
     layer3_out[1378] <= ~layer2_out[863] | layer2_out[862];
     layer3_out[1379] <= ~layer2_out[9];
     layer3_out[1380] <= layer2_out[597] | layer2_out[598];
     layer3_out[1381] <= ~layer2_out[1352];
     layer3_out[1382] <= ~layer2_out[275] | layer2_out[274];
     layer3_out[1383] <= ~layer2_out[1477];
     layer3_out[1384] <= layer2_out[1055];
     layer3_out[1385] <= layer2_out[1194] & ~layer2_out[1193];
     layer3_out[1386] <= layer2_out[1238] & ~layer2_out[1237];
     layer3_out[1387] <= layer2_out[1112];
     layer3_out[1388] <= 1'b1;
     layer3_out[1389] <= 1'b1;
     layer3_out[1390] <= layer2_out[425] & ~layer2_out[424];
     layer3_out[1391] <= layer2_out[644] | layer2_out[645];
     layer3_out[1392] <= layer2_out[653];
     layer3_out[1393] <= ~layer2_out[780];
     layer3_out[1394] <= ~(layer2_out[1263] | layer2_out[1264]);
     layer3_out[1395] <= ~layer2_out[980] | layer2_out[979];
     layer3_out[1396] <= ~layer2_out[1433];
     layer3_out[1397] <= layer2_out[230];
     layer3_out[1398] <= layer2_out[997];
     layer3_out[1399] <= ~layer2_out[322];
     layer3_out[1400] <= ~(layer2_out[905] & layer2_out[906]);
     layer3_out[1401] <= ~layer2_out[696] | layer2_out[697];
     layer3_out[1402] <= layer2_out[1145] & ~layer2_out[1144];
     layer3_out[1403] <= layer2_out[827] & ~layer2_out[828];
     layer3_out[1404] <= layer2_out[29];
     layer3_out[1405] <= 1'b1;
     layer3_out[1406] <= layer2_out[1407] & ~layer2_out[1408];
     layer3_out[1407] <= ~(layer2_out[563] | layer2_out[564]);
     layer3_out[1408] <= ~layer2_out[729] | layer2_out[730];
     layer3_out[1409] <= ~layer2_out[854] | layer2_out[855];
     layer3_out[1410] <= 1'b0;
     layer3_out[1411] <= ~layer2_out[777];
     layer3_out[1412] <= ~layer2_out[1137];
     layer3_out[1413] <= 1'b1;
     layer3_out[1414] <= layer2_out[482];
     layer3_out[1415] <= layer2_out[577];
     layer3_out[1416] <= layer2_out[927] | layer2_out[928];
     layer3_out[1417] <= layer2_out[917] & ~layer2_out[918];
     layer3_out[1418] <= ~layer2_out[243] | layer2_out[242];
     layer3_out[1419] <= ~layer2_out[1317];
     layer3_out[1420] <= layer2_out[818];
     layer3_out[1421] <= ~layer2_out[1497] | layer2_out[1498];
     layer3_out[1422] <= layer2_out[763] & ~layer2_out[764];
     layer3_out[1423] <= ~layer2_out[189] | layer2_out[188];
     layer3_out[1424] <= ~(layer2_out[1003] | layer2_out[1004]);
     layer3_out[1425] <= ~layer2_out[1338];
     layer3_out[1426] <= layer2_out[848] & ~layer2_out[847];
     layer3_out[1427] <= layer2_out[1455];
     layer3_out[1428] <= ~(layer2_out[395] | layer2_out[396]);
     layer3_out[1429] <= ~layer2_out[111];
     layer3_out[1430] <= ~layer2_out[1316];
     layer3_out[1431] <= 1'b0;
     layer3_out[1432] <= ~layer2_out[1160];
     layer3_out[1433] <= ~(layer2_out[1267] | layer2_out[1268]);
     layer3_out[1434] <= ~layer2_out[417];
     layer3_out[1435] <= ~layer2_out[1298];
     layer3_out[1436] <= 1'b1;
     layer3_out[1437] <= ~(layer2_out[718] & layer2_out[719]);
     layer3_out[1438] <= layer2_out[199] & layer2_out[200];
     layer3_out[1439] <= 1'b1;
     layer3_out[1440] <= 1'b1;
     layer3_out[1441] <= ~(layer2_out[1071] & layer2_out[1072]);
     layer3_out[1442] <= ~(layer2_out[1173] | layer2_out[1174]);
     layer3_out[1443] <= ~(layer2_out[1111] ^ layer2_out[1112]);
     layer3_out[1444] <= 1'b1;
     layer3_out[1445] <= ~(layer2_out[144] | layer2_out[145]);
     layer3_out[1446] <= layer2_out[1061] & layer2_out[1062];
     layer3_out[1447] <= ~layer2_out[945] | layer2_out[944];
     layer3_out[1448] <= ~(layer2_out[615] & layer2_out[616]);
     layer3_out[1449] <= layer2_out[1486] | layer2_out[1487];
     layer3_out[1450] <= layer2_out[67] & ~layer2_out[68];
     layer3_out[1451] <= layer2_out[162] & ~layer2_out[161];
     layer3_out[1452] <= ~(layer2_out[745] | layer2_out[746]);
     layer3_out[1453] <= ~layer2_out[346] | layer2_out[345];
     layer3_out[1454] <= layer2_out[967];
     layer3_out[1455] <= ~layer2_out[520] | layer2_out[521];
     layer3_out[1456] <= ~(layer2_out[1451] & layer2_out[1452]);
     layer3_out[1457] <= ~(layer2_out[350] ^ layer2_out[351]);
     layer3_out[1458] <= ~layer2_out[1103] | layer2_out[1102];
     layer3_out[1459] <= layer2_out[521];
     layer3_out[1460] <= layer2_out[1191] & ~layer2_out[1192];
     layer3_out[1461] <= layer2_out[948] & ~layer2_out[947];
     layer3_out[1462] <= ~layer2_out[95];
     layer3_out[1463] <= ~(layer2_out[592] | layer2_out[593]);
     layer3_out[1464] <= layer2_out[751] & layer2_out[752];
     layer3_out[1465] <= layer2_out[1239] & ~layer2_out[1240];
     layer3_out[1466] <= 1'b1;
     layer3_out[1467] <= ~(layer2_out[33] | layer2_out[34]);
     layer3_out[1468] <= layer2_out[355];
     layer3_out[1469] <= ~layer2_out[209] | layer2_out[210];
     layer3_out[1470] <= 1'b1;
     layer3_out[1471] <= layer2_out[724];
     layer3_out[1472] <= ~(layer2_out[864] | layer2_out[865]);
     layer3_out[1473] <= layer2_out[811];
     layer3_out[1474] <= 1'b0;
     layer3_out[1475] <= layer2_out[666] & layer2_out[667];
     layer3_out[1476] <= ~layer2_out[1126] | layer2_out[1127];
     layer3_out[1477] <= layer2_out[1293];
     layer3_out[1478] <= ~layer2_out[995];
     layer3_out[1479] <= ~(layer2_out[61] & layer2_out[62]);
     layer3_out[1480] <= layer2_out[1318] | layer2_out[1319];
     layer3_out[1481] <= layer2_out[1155] | layer2_out[1156];
     layer3_out[1482] <= layer2_out[1220] & ~layer2_out[1221];
     layer3_out[1483] <= layer2_out[773];
     layer3_out[1484] <= layer2_out[811];
     layer3_out[1485] <= ~(layer2_out[1153] & layer2_out[1154]);
     layer3_out[1486] <= 1'b1;
     layer3_out[1487] <= ~layer2_out[365] | layer2_out[364];
     layer3_out[1488] <= 1'b0;
     layer3_out[1489] <= 1'b1;
     layer3_out[1490] <= layer2_out[366] & ~layer2_out[367];
     layer3_out[1491] <= ~layer2_out[1164] | layer2_out[1165];
     layer3_out[1492] <= layer2_out[157];
     layer3_out[1493] <= ~layer2_out[1205] | layer2_out[1206];
     layer3_out[1494] <= layer2_out[290] | layer2_out[291];
     layer3_out[1495] <= layer2_out[1464] & ~layer2_out[1463];
     layer3_out[1496] <= layer2_out[1343];
     layer3_out[1497] <= layer2_out[618];
     layer3_out[1498] <= ~layer2_out[373];
     layer3_out[1499] <= layer2_out[848] & layer2_out[849];
     layer4_out[0] <= ~layer3_out[34];
     layer4_out[1] <= layer3_out[643] & ~layer3_out[642];
     layer4_out[2] <= ~layer3_out[783] | layer3_out[784];
     layer4_out[3] <= ~(layer3_out[546] & layer3_out[547]);
     layer4_out[4] <= layer3_out[956] & ~layer3_out[955];
     layer4_out[5] <= layer3_out[931] | layer3_out[932];
     layer4_out[6] <= ~layer3_out[857];
     layer4_out[7] <= ~layer3_out[364];
     layer4_out[8] <= ~layer3_out[870] | layer3_out[869];
     layer4_out[9] <= 1'b0;
     layer4_out[10] <= layer3_out[1492];
     layer4_out[11] <= layer3_out[454] | layer3_out[455];
     layer4_out[12] <= ~(layer3_out[1161] & layer3_out[1162]);
     layer4_out[13] <= ~(layer3_out[1470] & layer3_out[1471]);
     layer4_out[14] <= layer3_out[3];
     layer4_out[15] <= layer3_out[518] & layer3_out[519];
     layer4_out[16] <= layer3_out[1238] | layer3_out[1239];
     layer4_out[17] <= layer3_out[11] & ~layer3_out[12];
     layer4_out[18] <= layer3_out[385];
     layer4_out[19] <= layer3_out[321] & ~layer3_out[322];
     layer4_out[20] <= ~(layer3_out[1295] ^ layer3_out[1296]);
     layer4_out[21] <= layer3_out[96] ^ layer3_out[97];
     layer4_out[22] <= layer3_out[1083];
     layer4_out[23] <= ~layer3_out[636] | layer3_out[635];
     layer4_out[24] <= layer3_out[1298] ^ layer3_out[1299];
     layer4_out[25] <= layer3_out[941] & ~layer3_out[940];
     layer4_out[26] <= layer3_out[899] & layer3_out[900];
     layer4_out[27] <= layer3_out[3];
     layer4_out[28] <= ~layer3_out[601] | layer3_out[600];
     layer4_out[29] <= ~(layer3_out[1290] | layer3_out[1291]);
     layer4_out[30] <= ~layer3_out[1490];
     layer4_out[31] <= ~layer3_out[1106];
     layer4_out[32] <= layer3_out[1286] & ~layer3_out[1285];
     layer4_out[33] <= layer3_out[117] & ~layer3_out[118];
     layer4_out[34] <= 1'b0;
     layer4_out[35] <= ~layer3_out[983];
     layer4_out[36] <= 1'b0;
     layer4_out[37] <= layer3_out[359] | layer3_out[360];
     layer4_out[38] <= layer3_out[868];
     layer4_out[39] <= layer3_out[1454];
     layer4_out[40] <= ~layer3_out[1074] | layer3_out[1075];
     layer4_out[41] <= layer3_out[588] & layer3_out[589];
     layer4_out[42] <= ~layer3_out[302] | layer3_out[301];
     layer4_out[43] <= layer3_out[818] & ~layer3_out[819];
     layer4_out[44] <= layer3_out[989] & layer3_out[990];
     layer4_out[45] <= layer3_out[519] & layer3_out[520];
     layer4_out[46] <= ~layer3_out[461] | layer3_out[460];
     layer4_out[47] <= ~layer3_out[1007] | layer3_out[1006];
     layer4_out[48] <= ~layer3_out[1462] | layer3_out[1463];
     layer4_out[49] <= ~layer3_out[792] | layer3_out[791];
     layer4_out[50] <= layer3_out[1257];
     layer4_out[51] <= layer3_out[628];
     layer4_out[52] <= layer3_out[1310] & ~layer3_out[1311];
     layer4_out[53] <= layer3_out[158] ^ layer3_out[159];
     layer4_out[54] <= ~layer3_out[822] | layer3_out[821];
     layer4_out[55] <= ~layer3_out[1077] | layer3_out[1076];
     layer4_out[56] <= ~(layer3_out[1174] | layer3_out[1175]);
     layer4_out[57] <= layer3_out[451];
     layer4_out[58] <= layer3_out[1085];
     layer4_out[59] <= ~(layer3_out[1013] | layer3_out[1014]);
     layer4_out[60] <= ~layer3_out[842];
     layer4_out[61] <= ~(layer3_out[999] & layer3_out[1000]);
     layer4_out[62] <= layer3_out[1175] & layer3_out[1176];
     layer4_out[63] <= ~layer3_out[1286];
     layer4_out[64] <= layer3_out[1437];
     layer4_out[65] <= ~layer3_out[1046];
     layer4_out[66] <= ~(layer3_out[967] | layer3_out[968]);
     layer4_out[67] <= layer3_out[1416];
     layer4_out[68] <= layer3_out[407] & ~layer3_out[408];
     layer4_out[69] <= ~(layer3_out[73] | layer3_out[74]);
     layer4_out[70] <= layer3_out[1180];
     layer4_out[71] <= ~(layer3_out[328] & layer3_out[329]);
     layer4_out[72] <= layer3_out[1197];
     layer4_out[73] <= layer3_out[110] ^ layer3_out[111];
     layer4_out[74] <= ~layer3_out[662];
     layer4_out[75] <= layer3_out[320] & layer3_out[321];
     layer4_out[76] <= layer3_out[535] & ~layer3_out[536];
     layer4_out[77] <= layer3_out[1269];
     layer4_out[78] <= layer3_out[732] & layer3_out[733];
     layer4_out[79] <= layer3_out[1307] & ~layer3_out[1308];
     layer4_out[80] <= ~layer3_out[1445] | layer3_out[1444];
     layer4_out[81] <= ~(layer3_out[1020] & layer3_out[1021]);
     layer4_out[82] <= 1'b0;
     layer4_out[83] <= 1'b0;
     layer4_out[84] <= ~(layer3_out[1357] ^ layer3_out[1358]);
     layer4_out[85] <= ~(layer3_out[1279] | layer3_out[1280]);
     layer4_out[86] <= layer3_out[276] & ~layer3_out[275];
     layer4_out[87] <= 1'b0;
     layer4_out[88] <= ~(layer3_out[424] & layer3_out[425]);
     layer4_out[89] <= 1'b0;
     layer4_out[90] <= ~layer3_out[1248];
     layer4_out[91] <= ~(layer3_out[651] | layer3_out[652]);
     layer4_out[92] <= layer3_out[918] & ~layer3_out[917];
     layer4_out[93] <= layer3_out[992];
     layer4_out[94] <= ~(layer3_out[665] | layer3_out[666]);
     layer4_out[95] <= layer3_out[198];
     layer4_out[96] <= ~layer3_out[733];
     layer4_out[97] <= layer3_out[1244] & layer3_out[1245];
     layer4_out[98] <= layer3_out[693] & ~layer3_out[692];
     layer4_out[99] <= ~(layer3_out[859] & layer3_out[860]);
     layer4_out[100] <= ~(layer3_out[28] ^ layer3_out[29]);
     layer4_out[101] <= layer3_out[774];
     layer4_out[102] <= layer3_out[1067];
     layer4_out[103] <= 1'b0;
     layer4_out[104] <= layer3_out[258] & ~layer3_out[259];
     layer4_out[105] <= ~(layer3_out[430] | layer3_out[431]);
     layer4_out[106] <= ~layer3_out[349];
     layer4_out[107] <= layer3_out[866] | layer3_out[867];
     layer4_out[108] <= ~layer3_out[1399];
     layer4_out[109] <= layer3_out[20];
     layer4_out[110] <= ~(layer3_out[927] & layer3_out[928]);
     layer4_out[111] <= ~(layer3_out[1246] | layer3_out[1247]);
     layer4_out[112] <= layer3_out[1419] ^ layer3_out[1420];
     layer4_out[113] <= ~(layer3_out[347] | layer3_out[348]);
     layer4_out[114] <= ~(layer3_out[1189] & layer3_out[1190]);
     layer4_out[115] <= layer3_out[304] & ~layer3_out[303];
     layer4_out[116] <= layer3_out[1465] & ~layer3_out[1466];
     layer4_out[117] <= layer3_out[909] & layer3_out[910];
     layer4_out[118] <= ~(layer3_out[91] | layer3_out[92]);
     layer4_out[119] <= layer3_out[36];
     layer4_out[120] <= layer3_out[450] & ~layer3_out[449];
     layer4_out[121] <= layer3_out[615] & layer3_out[616];
     layer4_out[122] <= 1'b0;
     layer4_out[123] <= 1'b1;
     layer4_out[124] <= ~layer3_out[1139];
     layer4_out[125] <= layer3_out[190] & layer3_out[191];
     layer4_out[126] <= ~layer3_out[162];
     layer4_out[127] <= layer3_out[354];
     layer4_out[128] <= ~(layer3_out[765] ^ layer3_out[766]);
     layer4_out[129] <= layer3_out[294] & layer3_out[295];
     layer4_out[130] <= ~layer3_out[1030];
     layer4_out[131] <= 1'b1;
     layer4_out[132] <= ~layer3_out[1005];
     layer4_out[133] <= layer3_out[710] & ~layer3_out[709];
     layer4_out[134] <= layer3_out[988] & ~layer3_out[989];
     layer4_out[135] <= ~(layer3_out[569] ^ layer3_out[570]);
     layer4_out[136] <= layer3_out[1079] & ~layer3_out[1078];
     layer4_out[137] <= layer3_out[1302] ^ layer3_out[1303];
     layer4_out[138] <= ~layer3_out[691];
     layer4_out[139] <= layer3_out[1056] & ~layer3_out[1055];
     layer4_out[140] <= ~layer3_out[1250];
     layer4_out[141] <= layer3_out[1058] & ~layer3_out[1057];
     layer4_out[142] <= layer3_out[1226] | layer3_out[1227];
     layer4_out[143] <= layer3_out[663];
     layer4_out[144] <= ~layer3_out[152];
     layer4_out[145] <= ~(layer3_out[1056] & layer3_out[1057]);
     layer4_out[146] <= layer3_out[1050] & ~layer3_out[1051];
     layer4_out[147] <= ~layer3_out[168];
     layer4_out[148] <= layer3_out[796] & ~layer3_out[795];
     layer4_out[149] <= ~(layer3_out[44] & layer3_out[45]);
     layer4_out[150] <= layer3_out[696] | layer3_out[697];
     layer4_out[151] <= layer3_out[1393] & ~layer3_out[1394];
     layer4_out[152] <= ~layer3_out[1193] | layer3_out[1194];
     layer4_out[153] <= 1'b0;
     layer4_out[154] <= ~layer3_out[849];
     layer4_out[155] <= ~(layer3_out[695] ^ layer3_out[696]);
     layer4_out[156] <= layer3_out[247] & layer3_out[248];
     layer4_out[157] <= layer3_out[1009];
     layer4_out[158] <= 1'b1;
     layer4_out[159] <= layer3_out[1123] ^ layer3_out[1124];
     layer4_out[160] <= layer3_out[1186] & layer3_out[1187];
     layer4_out[161] <= layer3_out[69] & ~layer3_out[70];
     layer4_out[162] <= layer3_out[1461] & ~layer3_out[1460];
     layer4_out[163] <= ~(layer3_out[653] ^ layer3_out[654]);
     layer4_out[164] <= ~layer3_out[285] | layer3_out[286];
     layer4_out[165] <= layer3_out[830];
     layer4_out[166] <= ~layer3_out[604];
     layer4_out[167] <= layer3_out[750];
     layer4_out[168] <= layer3_out[893] & layer3_out[894];
     layer4_out[169] <= layer3_out[322];
     layer4_out[170] <= ~(layer3_out[704] | layer3_out[705]);
     layer4_out[171] <= layer3_out[1456] | layer3_out[1457];
     layer4_out[172] <= ~layer3_out[1271] | layer3_out[1272];
     layer4_out[173] <= ~(layer3_out[1039] | layer3_out[1040]);
     layer4_out[174] <= ~layer3_out[522];
     layer4_out[175] <= ~layer3_out[13] | layer3_out[14];
     layer4_out[176] <= ~layer3_out[960];
     layer4_out[177] <= layer3_out[1344] | layer3_out[1345];
     layer4_out[178] <= layer3_out[554] & ~layer3_out[555];
     layer4_out[179] <= ~layer3_out[1356];
     layer4_out[180] <= ~(layer3_out[926] ^ layer3_out[927]);
     layer4_out[181] <= ~(layer3_out[1180] & layer3_out[1181]);
     layer4_out[182] <= ~layer3_out[560];
     layer4_out[183] <= layer3_out[671];
     layer4_out[184] <= ~(layer3_out[1483] & layer3_out[1484]);
     layer4_out[185] <= layer3_out[500] & ~layer3_out[501];
     layer4_out[186] <= ~(layer3_out[1404] & layer3_out[1405]);
     layer4_out[187] <= layer3_out[1252] & ~layer3_out[1253];
     layer4_out[188] <= ~layer3_out[333];
     layer4_out[189] <= layer3_out[469];
     layer4_out[190] <= layer3_out[711];
     layer4_out[191] <= ~(layer3_out[340] & layer3_out[341]);
     layer4_out[192] <= ~layer3_out[1014];
     layer4_out[193] <= layer3_out[1118] | layer3_out[1119];
     layer4_out[194] <= ~(layer3_out[529] ^ layer3_out[530]);
     layer4_out[195] <= layer3_out[416];
     layer4_out[196] <= ~(layer3_out[339] | layer3_out[340]);
     layer4_out[197] <= layer3_out[1032];
     layer4_out[198] <= layer3_out[299] | layer3_out[300];
     layer4_out[199] <= layer3_out[1450];
     layer4_out[200] <= layer3_out[1316] ^ layer3_out[1317];
     layer4_out[201] <= ~layer3_out[42] | layer3_out[41];
     layer4_out[202] <= layer3_out[1017] | layer3_out[1018];
     layer4_out[203] <= ~(layer3_out[155] & layer3_out[156]);
     layer4_out[204] <= 1'b0;
     layer4_out[205] <= ~layer3_out[1382];
     layer4_out[206] <= ~layer3_out[464] | layer3_out[463];
     layer4_out[207] <= layer3_out[472] & ~layer3_out[473];
     layer4_out[208] <= ~layer3_out[396];
     layer4_out[209] <= layer3_out[144] & layer3_out[145];
     layer4_out[210] <= layer3_out[1431] & ~layer3_out[1430];
     layer4_out[211] <= ~layer3_out[1135] | layer3_out[1134];
     layer4_out[212] <= ~layer3_out[190] | layer3_out[189];
     layer4_out[213] <= layer3_out[136];
     layer4_out[214] <= ~layer3_out[1080] | layer3_out[1081];
     layer4_out[215] <= ~layer3_out[691];
     layer4_out[216] <= ~(layer3_out[1378] | layer3_out[1379]);
     layer4_out[217] <= ~layer3_out[806];
     layer4_out[218] <= ~layer3_out[526] | layer3_out[527];
     layer4_out[219] <= layer3_out[1222] & ~layer3_out[1221];
     layer4_out[220] <= layer3_out[1154];
     layer4_out[221] <= 1'b1;
     layer4_out[222] <= 1'b1;
     layer4_out[223] <= 1'b0;
     layer4_out[224] <= layer3_out[942] ^ layer3_out[943];
     layer4_out[225] <= layer3_out[1480] ^ layer3_out[1481];
     layer4_out[226] <= ~layer3_out[196];
     layer4_out[227] <= ~(layer3_out[465] ^ layer3_out[466]);
     layer4_out[228] <= 1'b1;
     layer4_out[229] <= layer3_out[1122] & ~layer3_out[1121];
     layer4_out[230] <= ~layer3_out[1417];
     layer4_out[231] <= ~layer3_out[76] | layer3_out[77];
     layer4_out[232] <= layer3_out[825];
     layer4_out[233] <= layer3_out[862];
     layer4_out[234] <= ~layer3_out[436];
     layer4_out[235] <= layer3_out[853] & ~layer3_out[854];
     layer4_out[236] <= ~layer3_out[827];
     layer4_out[237] <= ~layer3_out[540];
     layer4_out[238] <= 1'b1;
     layer4_out[239] <= ~layer3_out[543];
     layer4_out[240] <= layer3_out[1016] | layer3_out[1017];
     layer4_out[241] <= ~(layer3_out[478] & layer3_out[479]);
     layer4_out[242] <= layer3_out[667] & ~layer3_out[666];
     layer4_out[243] <= ~layer3_out[934];
     layer4_out[244] <= ~layer3_out[49] | layer3_out[50];
     layer4_out[245] <= ~(layer3_out[194] | layer3_out[195]);
     layer4_out[246] <= ~layer3_out[352];
     layer4_out[247] <= ~layer3_out[1402];
     layer4_out[248] <= layer3_out[421];
     layer4_out[249] <= layer3_out[426] & ~layer3_out[425];
     layer4_out[250] <= layer3_out[24] | layer3_out[25];
     layer4_out[251] <= ~layer3_out[830];
     layer4_out[252] <= ~layer3_out[264];
     layer4_out[253] <= 1'b1;
     layer4_out[254] <= ~layer3_out[912];
     layer4_out[255] <= layer3_out[994];
     layer4_out[256] <= ~layer3_out[1498];
     layer4_out[257] <= layer3_out[12] | layer3_out[13];
     layer4_out[258] <= ~layer3_out[416];
     layer4_out[259] <= ~(layer3_out[317] & layer3_out[318]);
     layer4_out[260] <= ~layer3_out[1223];
     layer4_out[261] <= layer3_out[1424] & ~layer3_out[1423];
     layer4_out[262] <= ~layer3_out[1427] | layer3_out[1426];
     layer4_out[263] <= ~(layer3_out[5] ^ layer3_out[6]);
     layer4_out[264] <= layer3_out[1209];
     layer4_out[265] <= layer3_out[987] & ~layer3_out[986];
     layer4_out[266] <= layer3_out[498];
     layer4_out[267] <= layer3_out[1371];
     layer4_out[268] <= layer3_out[770];
     layer4_out[269] <= 1'b0;
     layer4_out[270] <= ~(layer3_out[934] ^ layer3_out[935]);
     layer4_out[271] <= ~(layer3_out[1276] | layer3_out[1277]);
     layer4_out[272] <= layer3_out[227];
     layer4_out[273] <= layer3_out[239] | layer3_out[240];
     layer4_out[274] <= layer3_out[990] & layer3_out[991];
     layer4_out[275] <= ~(layer3_out[823] ^ layer3_out[824]);
     layer4_out[276] <= layer3_out[1382];
     layer4_out[277] <= ~layer3_out[278];
     layer4_out[278] <= layer3_out[530] & ~layer3_out[531];
     layer4_out[279] <= ~layer3_out[627] | layer3_out[626];
     layer4_out[280] <= layer3_out[246];
     layer4_out[281] <= ~(layer3_out[295] & layer3_out[296]);
     layer4_out[282] <= layer3_out[1297] & ~layer3_out[1298];
     layer4_out[283] <= ~(layer3_out[1100] & layer3_out[1101]);
     layer4_out[284] <= layer3_out[1397];
     layer4_out[285] <= ~(layer3_out[367] & layer3_out[368]);
     layer4_out[286] <= ~layer3_out[508];
     layer4_out[287] <= layer3_out[1434] & ~layer3_out[1435];
     layer4_out[288] <= layer3_out[1115] | layer3_out[1116];
     layer4_out[289] <= layer3_out[816];
     layer4_out[290] <= layer3_out[748] & ~layer3_out[749];
     layer4_out[291] <= layer3_out[946] & ~layer3_out[947];
     layer4_out[292] <= layer3_out[810] | layer3_out[811];
     layer4_out[293] <= layer3_out[1040];
     layer4_out[294] <= ~(layer3_out[718] | layer3_out[719]);
     layer4_out[295] <= layer3_out[1206] | layer3_out[1207];
     layer4_out[296] <= ~layer3_out[169] | layer3_out[170];
     layer4_out[297] <= ~layer3_out[1007];
     layer4_out[298] <= ~layer3_out[146];
     layer4_out[299] <= ~(layer3_out[657] & layer3_out[658]);
     layer4_out[300] <= ~layer3_out[837] | layer3_out[836];
     layer4_out[301] <= layer3_out[497] & ~layer3_out[496];
     layer4_out[302] <= layer3_out[349] | layer3_out[350];
     layer4_out[303] <= layer3_out[767];
     layer4_out[304] <= layer3_out[23] | layer3_out[24];
     layer4_out[305] <= ~layer3_out[354] | layer3_out[353];
     layer4_out[306] <= ~layer3_out[1266] | layer3_out[1265];
     layer4_out[307] <= layer3_out[707] & ~layer3_out[708];
     layer4_out[308] <= ~layer3_out[507];
     layer4_out[309] <= 1'b1;
     layer4_out[310] <= ~(layer3_out[170] ^ layer3_out[171]);
     layer4_out[311] <= ~layer3_out[1233] | layer3_out[1234];
     layer4_out[312] <= layer3_out[1425] & layer3_out[1426];
     layer4_out[313] <= ~(layer3_out[1379] | layer3_out[1380]);
     layer4_out[314] <= layer3_out[619] | layer3_out[620];
     layer4_out[315] <= layer3_out[1365];
     layer4_out[316] <= layer3_out[508] & ~layer3_out[507];
     layer4_out[317] <= layer3_out[648];
     layer4_out[318] <= ~layer3_out[489];
     layer4_out[319] <= layer3_out[1166] & ~layer3_out[1167];
     layer4_out[320] <= ~layer3_out[344];
     layer4_out[321] <= 1'b0;
     layer4_out[322] <= 1'b1;
     layer4_out[323] <= layer3_out[1331];
     layer4_out[324] <= layer3_out[181] ^ layer3_out[182];
     layer4_out[325] <= layer3_out[475] & ~layer3_out[474];
     layer4_out[326] <= ~layer3_out[62];
     layer4_out[327] <= ~layer3_out[1394];
     layer4_out[328] <= layer3_out[504] & ~layer3_out[505];
     layer4_out[329] <= layer3_out[550];
     layer4_out[330] <= ~(layer3_out[186] & layer3_out[187]);
     layer4_out[331] <= ~layer3_out[1413] | layer3_out[1412];
     layer4_out[332] <= layer3_out[879];
     layer4_out[333] <= ~layer3_out[561] | layer3_out[562];
     layer4_out[334] <= layer3_out[1132] & ~layer3_out[1131];
     layer4_out[335] <= layer3_out[668];
     layer4_out[336] <= layer3_out[252] & ~layer3_out[253];
     layer4_out[337] <= layer3_out[1112];
     layer4_out[338] <= ~(layer3_out[520] & layer3_out[521]);
     layer4_out[339] <= ~layer3_out[1476];
     layer4_out[340] <= layer3_out[487] & layer3_out[488];
     layer4_out[341] <= ~(layer3_out[499] & layer3_out[500]);
     layer4_out[342] <= ~layer3_out[478] | layer3_out[477];
     layer4_out[343] <= layer3_out[429];
     layer4_out[344] <= ~layer3_out[777];
     layer4_out[345] <= ~layer3_out[1352] | layer3_out[1353];
     layer4_out[346] <= ~layer3_out[937] | layer3_out[938];
     layer4_out[347] <= ~(layer3_out[1242] & layer3_out[1243]);
     layer4_out[348] <= ~layer3_out[746];
     layer4_out[349] <= ~layer3_out[639] | layer3_out[640];
     layer4_out[350] <= ~layer3_out[441] | layer3_out[440];
     layer4_out[351] <= layer3_out[580] | layer3_out[581];
     layer4_out[352] <= layer3_out[613] & ~layer3_out[614];
     layer4_out[353] <= layer3_out[415] & ~layer3_out[414];
     layer4_out[354] <= layer3_out[945];
     layer4_out[355] <= layer3_out[267] & layer3_out[268];
     layer4_out[356] <= ~(layer3_out[1002] ^ layer3_out[1003]);
     layer4_out[357] <= layer3_out[719];
     layer4_out[358] <= ~(layer3_out[121] | layer3_out[122]);
     layer4_out[359] <= ~layer3_out[187] | layer3_out[188];
     layer4_out[360] <= layer3_out[721] | layer3_out[722];
     layer4_out[361] <= ~layer3_out[1455] | layer3_out[1456];
     layer4_out[362] <= layer3_out[99] ^ layer3_out[100];
     layer4_out[363] <= ~layer3_out[1408];
     layer4_out[364] <= ~layer3_out[642] | layer3_out[641];
     layer4_out[365] <= ~layer3_out[898] | layer3_out[897];
     layer4_out[366] <= layer3_out[1277] & ~layer3_out[1278];
     layer4_out[367] <= layer3_out[1095] & layer3_out[1096];
     layer4_out[368] <= layer3_out[90] & ~layer3_out[89];
     layer4_out[369] <= layer3_out[1058] | layer3_out[1059];
     layer4_out[370] <= ~layer3_out[680];
     layer4_out[371] <= ~layer3_out[902];
     layer4_out[372] <= ~layer3_out[335];
     layer4_out[373] <= 1'b1;
     layer4_out[374] <= layer3_out[60] | layer3_out[61];
     layer4_out[375] <= layer3_out[289];
     layer4_out[376] <= ~(layer3_out[1140] & layer3_out[1141]);
     layer4_out[377] <= layer3_out[1235];
     layer4_out[378] <= ~layer3_out[602] | layer3_out[603];
     layer4_out[379] <= layer3_out[32];
     layer4_out[380] <= layer3_out[1494] & layer3_out[1495];
     layer4_out[381] <= ~layer3_out[261] | layer3_out[260];
     layer4_out[382] <= ~layer3_out[1390] | layer3_out[1391];
     layer4_out[383] <= layer3_out[865] & ~layer3_out[866];
     layer4_out[384] <= layer3_out[933] & ~layer3_out[932];
     layer4_out[385] <= layer3_out[361];
     layer4_out[386] <= 1'b0;
     layer4_out[387] <= ~layer3_out[265];
     layer4_out[388] <= ~(layer3_out[62] & layer3_out[63]);
     layer4_out[389] <= ~layer3_out[456];
     layer4_out[390] <= ~(layer3_out[634] | layer3_out[635]);
     layer4_out[391] <= layer3_out[279] & layer3_out[280];
     layer4_out[392] <= ~layer3_out[481] | layer3_out[480];
     layer4_out[393] <= ~(layer3_out[0] & layer3_out[2]);
     layer4_out[394] <= layer3_out[161];
     layer4_out[395] <= ~layer3_out[521] | layer3_out[522];
     layer4_out[396] <= ~layer3_out[1038];
     layer4_out[397] <= ~(layer3_out[1171] | layer3_out[1172]);
     layer4_out[398] <= ~(layer3_out[1420] | layer3_out[1421]);
     layer4_out[399] <= ~(layer3_out[1051] & layer3_out[1052]);
     layer4_out[400] <= layer3_out[831];
     layer4_out[401] <= layer3_out[404];
     layer4_out[402] <= ~layer3_out[812] | layer3_out[813];
     layer4_out[403] <= layer3_out[1264] & ~layer3_out[1265];
     layer4_out[404] <= layer3_out[1437];
     layer4_out[405] <= layer3_out[485];
     layer4_out[406] <= layer3_out[281];
     layer4_out[407] <= ~layer3_out[660];
     layer4_out[408] <= layer3_out[1003] | layer3_out[1004];
     layer4_out[409] <= layer3_out[84];
     layer4_out[410] <= layer3_out[880];
     layer4_out[411] <= layer3_out[1114] & ~layer3_out[1113];
     layer4_out[412] <= layer3_out[323] & layer3_out[324];
     layer4_out[413] <= 1'b0;
     layer4_out[414] <= ~(layer3_out[584] | layer3_out[585]);
     layer4_out[415] <= layer3_out[104] & layer3_out[105];
     layer4_out[416] <= layer3_out[1209];
     layer4_out[417] <= ~layer3_out[177] | layer3_out[178];
     layer4_out[418] <= ~(layer3_out[107] & layer3_out[108]);
     layer4_out[419] <= layer3_out[365] & ~layer3_out[364];
     layer4_out[420] <= layer3_out[660] | layer3_out[661];
     layer4_out[421] <= ~layer3_out[971];
     layer4_out[422] <= ~layer3_out[1148];
     layer4_out[423] <= ~(layer3_out[380] & layer3_out[381]);
     layer4_out[424] <= layer3_out[1110];
     layer4_out[425] <= ~(layer3_out[1054] & layer3_out[1055]);
     layer4_out[426] <= ~layer3_out[734];
     layer4_out[427] <= layer3_out[112] & ~layer3_out[111];
     layer4_out[428] <= layer3_out[92];
     layer4_out[429] <= ~layer3_out[292];
     layer4_out[430] <= ~layer3_out[231];
     layer4_out[431] <= ~(layer3_out[687] | layer3_out[688]);
     layer4_out[432] <= layer3_out[325] | layer3_out[326];
     layer4_out[433] <= layer3_out[369] | layer3_out[370];
     layer4_out[434] <= layer3_out[610] & layer3_out[611];
     layer4_out[435] <= layer3_out[1374] & ~layer3_out[1375];
     layer4_out[436] <= ~layer3_out[1128] | layer3_out[1129];
     layer4_out[437] <= 1'b1;
     layer4_out[438] <= layer3_out[1424] ^ layer3_out[1425];
     layer4_out[439] <= 1'b1;
     layer4_out[440] <= layer3_out[1153] & ~layer3_out[1152];
     layer4_out[441] <= ~layer3_out[446];
     layer4_out[442] <= layer3_out[762] & layer3_out[763];
     layer4_out[443] <= layer3_out[395] & ~layer3_out[394];
     layer4_out[444] <= ~layer3_out[282] | layer3_out[283];
     layer4_out[445] <= ~layer3_out[787];
     layer4_out[446] <= layer3_out[1192];
     layer4_out[447] <= layer3_out[1350] | layer3_out[1351];
     layer4_out[448] <= layer3_out[10] & layer3_out[11];
     layer4_out[449] <= ~layer3_out[722] | layer3_out[723];
     layer4_out[450] <= layer3_out[1173];
     layer4_out[451] <= ~layer3_out[694];
     layer4_out[452] <= ~layer3_out[973] | layer3_out[972];
     layer4_out[453] <= ~layer3_out[21];
     layer4_out[454] <= layer3_out[317] & ~layer3_out[316];
     layer4_out[455] <= layer3_out[701];
     layer4_out[456] <= ~(layer3_out[913] | layer3_out[914]);
     layer4_out[457] <= ~layer3_out[1139] | layer3_out[1140];
     layer4_out[458] <= ~layer3_out[238];
     layer4_out[459] <= ~(layer3_out[148] & layer3_out[149]);
     layer4_out[460] <= ~(layer3_out[670] & layer3_out[671]);
     layer4_out[461] <= ~(layer3_out[139] | layer3_out[140]);
     layer4_out[462] <= ~(layer3_out[1144] | layer3_out[1145]);
     layer4_out[463] <= ~layer3_out[1368] | layer3_out[1367];
     layer4_out[464] <= layer3_out[751];
     layer4_out[465] <= layer3_out[138] | layer3_out[139];
     layer4_out[466] <= 1'b1;
     layer4_out[467] <= ~layer3_out[741] | layer3_out[742];
     layer4_out[468] <= ~(layer3_out[393] | layer3_out[394]);
     layer4_out[469] <= layer3_out[954];
     layer4_out[470] <= layer3_out[882];
     layer4_out[471] <= layer3_out[164];
     layer4_out[472] <= ~(layer3_out[1348] & layer3_out[1349]);
     layer4_out[473] <= ~layer3_out[626] | layer3_out[625];
     layer4_out[474] <= ~(layer3_out[156] & layer3_out[157]);
     layer4_out[475] <= ~(layer3_out[1428] | layer3_out[1429]);
     layer4_out[476] <= layer3_out[94];
     layer4_out[477] <= ~(layer3_out[564] | layer3_out[565]);
     layer4_out[478] <= layer3_out[614] & ~layer3_out[615];
     layer4_out[479] <= ~layer3_out[176] | layer3_out[177];
     layer4_out[480] <= layer3_out[299];
     layer4_out[481] <= 1'b0;
     layer4_out[482] <= layer3_out[593] ^ layer3_out[594];
     layer4_out[483] <= 1'b0;
     layer4_out[484] <= layer3_out[1044];
     layer4_out[485] <= layer3_out[1301] | layer3_out[1302];
     layer4_out[486] <= layer3_out[504] & ~layer3_out[503];
     layer4_out[487] <= layer3_out[213] & ~layer3_out[214];
     layer4_out[488] <= layer3_out[1340] | layer3_out[1341];
     layer4_out[489] <= ~layer3_out[1411];
     layer4_out[490] <= ~layer3_out[1253] | layer3_out[1254];
     layer4_out[491] <= 1'b1;
     layer4_out[492] <= layer3_out[254] & ~layer3_out[253];
     layer4_out[493] <= ~layer3_out[390] | layer3_out[389];
     layer4_out[494] <= layer3_out[1377] | layer3_out[1378];
     layer4_out[495] <= layer3_out[1027] & ~layer3_out[1028];
     layer4_out[496] <= layer3_out[578] & ~layer3_out[577];
     layer4_out[497] <= 1'b1;
     layer4_out[498] <= ~layer3_out[1346] | layer3_out[1345];
     layer4_out[499] <= layer3_out[330];
     layer4_out[500] <= ~layer3_out[754];
     layer4_out[501] <= layer3_out[153] & ~layer3_out[152];
     layer4_out[502] <= layer3_out[1268] & ~layer3_out[1267];
     layer4_out[503] <= ~layer3_out[985] | layer3_out[984];
     layer4_out[504] <= ~(layer3_out[490] | layer3_out[491]);
     layer4_out[505] <= layer3_out[115] | layer3_out[116];
     layer4_out[506] <= ~(layer3_out[1104] & layer3_out[1105]);
     layer4_out[507] <= ~layer3_out[398];
     layer4_out[508] <= layer3_out[1171] & ~layer3_out[1170];
     layer4_out[509] <= layer3_out[401];
     layer4_out[510] <= layer3_out[1359] & layer3_out[1360];
     layer4_out[511] <= ~layer3_out[344] | layer3_out[345];
     layer4_out[512] <= ~layer3_out[30];
     layer4_out[513] <= layer3_out[1230];
     layer4_out[514] <= ~layer3_out[1236];
     layer4_out[515] <= ~layer3_out[379] | layer3_out[380];
     layer4_out[516] <= ~layer3_out[725] | layer3_out[726];
     layer4_out[517] <= ~layer3_out[841] | layer3_out[840];
     layer4_out[518] <= ~layer3_out[884];
     layer4_out[519] <= ~layer3_out[438];
     layer4_out[520] <= layer3_out[1284] ^ layer3_out[1285];
     layer4_out[521] <= ~(layer3_out[858] & layer3_out[859]);
     layer4_out[522] <= ~(layer3_out[327] | layer3_out[328]);
     layer4_out[523] <= ~layer3_out[1238] | layer3_out[1237];
     layer4_out[524] <= layer3_out[1085];
     layer4_out[525] <= ~layer3_out[1354];
     layer4_out[526] <= ~layer3_out[1244];
     layer4_out[527] <= layer3_out[716] & layer3_out[717];
     layer4_out[528] <= layer3_out[307];
     layer4_out[529] <= layer3_out[228];
     layer4_out[530] <= layer3_out[208] | layer3_out[209];
     layer4_out[531] <= ~layer3_out[131] | layer3_out[132];
     layer4_out[532] <= ~(layer3_out[452] | layer3_out[453]);
     layer4_out[533] <= ~layer3_out[1250];
     layer4_out[534] <= ~(layer3_out[596] & layer3_out[597]);
     layer4_out[535] <= layer3_out[78];
     layer4_out[536] <= layer3_out[305];
     layer4_out[537] <= ~(layer3_out[204] | layer3_out[205]);
     layer4_out[538] <= ~layer3_out[572] | layer3_out[573];
     layer4_out[539] <= ~layer3_out[214];
     layer4_out[540] <= layer3_out[809] & ~layer3_out[810];
     layer4_out[541] <= ~layer3_out[358];
     layer4_out[542] <= 1'b0;
     layer4_out[543] <= layer3_out[785];
     layer4_out[544] <= ~layer3_out[428];
     layer4_out[545] <= layer3_out[976] | layer3_out[977];
     layer4_out[546] <= ~layer3_out[361];
     layer4_out[547] <= layer3_out[1033] | layer3_out[1034];
     layer4_out[548] <= ~(layer3_out[180] & layer3_out[181]);
     layer4_out[549] <= ~layer3_out[1313] | layer3_out[1312];
     layer4_out[550] <= layer3_out[336] | layer3_out[337];
     layer4_out[551] <= layer3_out[581];
     layer4_out[552] <= 1'b1;
     layer4_out[553] <= ~(layer3_out[541] ^ layer3_out[542]);
     layer4_out[554] <= layer3_out[1478];
     layer4_out[555] <= ~(layer3_out[742] & layer3_out[743]);
     layer4_out[556] <= ~(layer3_out[549] & layer3_out[550]);
     layer4_out[557] <= ~(layer3_out[220] & layer3_out[221]);
     layer4_out[558] <= ~layer3_out[1399];
     layer4_out[559] <= ~(layer3_out[775] & layer3_out[776]);
     layer4_out[560] <= layer3_out[1192] & layer3_out[1193];
     layer4_out[561] <= ~(layer3_out[895] | layer3_out[896]);
     layer4_out[562] <= layer3_out[623] & ~layer3_out[622];
     layer4_out[563] <= layer3_out[1386] & layer3_out[1387];
     layer4_out[564] <= ~(layer3_out[806] & layer3_out[807]);
     layer4_out[565] <= layer3_out[1471] & ~layer3_out[1472];
     layer4_out[566] <= ~(layer3_out[514] | layer3_out[515]);
     layer4_out[567] <= layer3_out[496] & ~layer3_out[495];
     layer4_out[568] <= 1'b1;
     layer4_out[569] <= layer3_out[173];
     layer4_out[570] <= ~(layer3_out[1473] | layer3_out[1474]);
     layer4_out[571] <= layer3_out[1155] | layer3_out[1156];
     layer4_out[572] <= ~layer3_out[982] | layer3_out[981];
     layer4_out[573] <= layer3_out[72] | layer3_out[73];
     layer4_out[574] <= 1'b1;
     layer4_out[575] <= layer3_out[650];
     layer4_out[576] <= layer3_out[376] ^ layer3_out[377];
     layer4_out[577] <= ~(layer3_out[974] & layer3_out[975]);
     layer4_out[578] <= layer3_out[410];
     layer4_out[579] <= ~(layer3_out[646] & layer3_out[647]);
     layer4_out[580] <= layer3_out[1261] & ~layer3_out[1262];
     layer4_out[581] <= layer3_out[1317] & layer3_out[1318];
     layer4_out[582] <= ~layer3_out[1242];
     layer4_out[583] <= layer3_out[74];
     layer4_out[584] <= layer3_out[1073] & layer3_out[1074];
     layer4_out[585] <= layer3_out[1495];
     layer4_out[586] <= ~(layer3_out[669] & layer3_out[670]);
     layer4_out[587] <= layer3_out[826] & ~layer3_out[827];
     layer4_out[588] <= ~layer3_out[1103] | layer3_out[1104];
     layer4_out[589] <= ~layer3_out[1216];
     layer4_out[590] <= layer3_out[1341];
     layer4_out[591] <= layer3_out[417] & layer3_out[418];
     layer4_out[592] <= layer3_out[492] ^ layer3_out[493];
     layer4_out[593] <= ~layer3_out[96];
     layer4_out[594] <= ~layer3_out[618] | layer3_out[619];
     layer4_out[595] <= ~layer3_out[235] | layer3_out[236];
     layer4_out[596] <= ~layer3_out[128] | layer3_out[129];
     layer4_out[597] <= layer3_out[137];
     layer4_out[598] <= layer3_out[81] & ~layer3_out[82];
     layer4_out[599] <= layer3_out[652] & layer3_out[653];
     layer4_out[600] <= ~layer3_out[375] | layer3_out[376];
     layer4_out[601] <= layer3_out[312] & layer3_out[313];
     layer4_out[602] <= ~layer3_out[1373];
     layer4_out[603] <= 1'b1;
     layer4_out[604] <= layer3_out[552];
     layer4_out[605] <= ~layer3_out[729] | layer3_out[730];
     layer4_out[606] <= ~layer3_out[433];
     layer4_out[607] <= layer3_out[26] & ~layer3_out[27];
     layer4_out[608] <= ~layer3_out[790] | layer3_out[791];
     layer4_out[609] <= ~layer3_out[786] | layer3_out[787];
     layer4_out[610] <= 1'b1;
     layer4_out[611] <= layer3_out[538];
     layer4_out[612] <= ~(layer3_out[819] | layer3_out[820]);
     layer4_out[613] <= layer3_out[1019];
     layer4_out[614] <= layer3_out[744];
     layer4_out[615] <= layer3_out[1343] & ~layer3_out[1344];
     layer4_out[616] <= layer3_out[405] | layer3_out[406];
     layer4_out[617] <= layer3_out[747];
     layer4_out[618] <= ~layer3_out[59] | layer3_out[58];
     layer4_out[619] <= layer3_out[1381];
     layer4_out[620] <= ~layer3_out[964];
     layer4_out[621] <= ~layer3_out[281] | layer3_out[280];
     layer4_out[622] <= 1'b0;
     layer4_out[623] <= layer3_out[345] | layer3_out[346];
     layer4_out[624] <= ~layer3_out[1099];
     layer4_out[625] <= layer3_out[1127];
     layer4_out[626] <= layer3_out[285] & ~layer3_out[284];
     layer4_out[627] <= ~layer3_out[937] | layer3_out[936];
     layer4_out[628] <= ~layer3_out[711];
     layer4_out[629] <= ~layer3_out[1177] | layer3_out[1178];
     layer4_out[630] <= layer3_out[1459] & layer3_out[1460];
     layer4_out[631] <= ~layer3_out[1475] | layer3_out[1476];
     layer4_out[632] <= ~layer3_out[807] | layer3_out[808];
     layer4_out[633] <= layer3_out[911] | layer3_out[912];
     layer4_out[634] <= ~layer3_out[1063];
     layer4_out[635] <= layer3_out[1090] & ~layer3_out[1091];
     layer4_out[636] <= layer3_out[288] & ~layer3_out[287];
     layer4_out[637] <= ~layer3_out[358] | layer3_out[359];
     layer4_out[638] <= layer3_out[777] | layer3_out[778];
     layer4_out[639] <= 1'b1;
     layer4_out[640] <= ~layer3_out[1462];
     layer4_out[641] <= layer3_out[890];
     layer4_out[642] <= ~layer3_out[1087];
     layer4_out[643] <= ~(layer3_out[1450] | layer3_out[1451]);
     layer4_out[644] <= layer3_out[103];
     layer4_out[645] <= layer3_out[1408] | layer3_out[1409];
     layer4_out[646] <= layer3_out[15] | layer3_out[16];
     layer4_out[647] <= layer3_out[792] & layer3_out[793];
     layer4_out[648] <= ~layer3_out[409] | layer3_out[408];
     layer4_out[649] <= 1'b0;
     layer4_out[650] <= ~layer3_out[1212] | layer3_out[1213];
     layer4_out[651] <= 1'b1;
     layer4_out[652] <= layer3_out[541];
     layer4_out[653] <= layer3_out[1290];
     layer4_out[654] <= ~layer3_out[707];
     layer4_out[655] <= ~layer3_out[622] | layer3_out[621];
     layer4_out[656] <= 1'b0;
     layer4_out[657] <= layer3_out[314] | layer3_out[315];
     layer4_out[658] <= layer3_out[712];
     layer4_out[659] <= ~layer3_out[953];
     layer4_out[660] <= ~layer3_out[1053];
     layer4_out[661] <= ~(layer3_out[534] & layer3_out[535]);
     layer4_out[662] <= layer3_out[223] & ~layer3_out[224];
     layer4_out[663] <= layer3_out[55];
     layer4_out[664] <= ~layer3_out[71] | layer3_out[72];
     layer4_out[665] <= layer3_out[1275] & layer3_out[1276];
     layer4_out[666] <= ~(layer3_out[770] & layer3_out[771]);
     layer4_out[667] <= ~(layer3_out[1278] | layer3_out[1279]);
     layer4_out[668] <= ~layer3_out[144];
     layer4_out[669] <= ~(layer3_out[701] | layer3_out[702]);
     layer4_out[670] <= ~layer3_out[1217];
     layer4_out[671] <= layer3_out[241];
     layer4_out[672] <= ~layer3_out[714];
     layer4_out[673] <= layer3_out[1485] & layer3_out[1486];
     layer4_out[674] <= ~layer3_out[1410];
     layer4_out[675] <= layer3_out[462] ^ layer3_out[463];
     layer4_out[676] <= ~layer3_out[1466];
     layer4_out[677] <= layer3_out[703] & ~layer3_out[704];
     layer4_out[678] <= ~layer3_out[679];
     layer4_out[679] <= layer3_out[637] | layer3_out[638];
     layer4_out[680] <= layer3_out[876];
     layer4_out[681] <= ~layer3_out[9];
     layer4_out[682] <= ~(layer3_out[185] & layer3_out[186]);
     layer4_out[683] <= layer3_out[812] & ~layer3_out[811];
     layer4_out[684] <= ~layer3_out[115] | layer3_out[114];
     layer4_out[685] <= ~layer3_out[183];
     layer4_out[686] <= layer3_out[1105] ^ layer3_out[1106];
     layer4_out[687] <= ~layer3_out[503];
     layer4_out[688] <= layer3_out[166] & layer3_out[167];
     layer4_out[689] <= layer3_out[1004] ^ layer3_out[1005];
     layer4_out[690] <= ~layer3_out[727] | layer3_out[728];
     layer4_out[691] <= layer3_out[316] & ~layer3_out[315];
     layer4_out[692] <= 1'b1;
     layer4_out[693] <= 1'b1;
     layer4_out[694] <= ~layer3_out[401];
     layer4_out[695] <= layer3_out[684] & layer3_out[685];
     layer4_out[696] <= ~layer3_out[1414];
     layer4_out[697] <= ~layer3_out[531];
     layer4_out[698] <= layer3_out[857] & layer3_out[858];
     layer4_out[699] <= ~layer3_out[1343];
     layer4_out[700] <= ~(layer3_out[929] | layer3_out[930]);
     layer4_out[701] <= ~layer3_out[291];
     layer4_out[702] <= ~(layer3_out[1070] | layer3_out[1071]);
     layer4_out[703] <= ~layer3_out[680] | layer3_out[681];
     layer4_out[704] <= ~layer3_out[1433];
     layer4_out[705] <= layer3_out[1468] | layer3_out[1469];
     layer4_out[706] <= layer3_out[682] | layer3_out[683];
     layer4_out[707] <= layer3_out[760];
     layer4_out[708] <= layer3_out[393];
     layer4_out[709] <= layer3_out[421] & layer3_out[422];
     layer4_out[710] <= layer3_out[864] & ~layer3_out[865];
     layer4_out[711] <= ~layer3_out[621];
     layer4_out[712] <= ~(layer3_out[1092] & layer3_out[1093]);
     layer4_out[713] <= layer3_out[210] & ~layer3_out[209];
     layer4_out[714] <= layer3_out[80];
     layer4_out[715] <= ~layer3_out[412] | layer3_out[411];
     layer4_out[716] <= ~(layer3_out[1035] & layer3_out[1036]);
     layer4_out[717] <= ~layer3_out[893];
     layer4_out[718] <= ~layer3_out[41];
     layer4_out[719] <= layer3_out[479] & layer3_out[480];
     layer4_out[720] <= ~layer3_out[1142];
     layer4_out[721] <= ~(layer3_out[98] | layer3_out[99]);
     layer4_out[722] <= layer3_out[391] & ~layer3_out[392];
     layer4_out[723] <= layer3_out[148];
     layer4_out[724] <= ~(layer3_out[1474] & layer3_out[1475]);
     layer4_out[725] <= ~layer3_out[835] | layer3_out[834];
     layer4_out[726] <= layer3_out[605];
     layer4_out[727] <= layer3_out[273];
     layer4_out[728] <= 1'b1;
     layer4_out[729] <= ~layer3_out[406];
     layer4_out[730] <= ~layer3_out[779];
     layer4_out[731] <= ~layer3_out[752] | layer3_out[751];
     layer4_out[732] <= layer3_out[1047];
     layer4_out[733] <= layer3_out[788];
     layer4_out[734] <= ~layer3_out[818] | layer3_out[817];
     layer4_out[735] <= ~layer3_out[1030] | layer3_out[1029];
     layer4_out[736] <= layer3_out[1348] & ~layer3_out[1347];
     layer4_out[737] <= layer3_out[828];
     layer4_out[738] <= layer3_out[1165] & layer3_out[1166];
     layer4_out[739] <= 1'b1;
     layer4_out[740] <= layer3_out[1002];
     layer4_out[741] <= layer3_out[165];
     layer4_out[742] <= ~(layer3_out[266] ^ layer3_out[267]);
     layer4_out[743] <= layer3_out[1155] & ~layer3_out[1154];
     layer4_out[744] <= layer3_out[1203] & ~layer3_out[1204];
     layer4_out[745] <= layer3_out[1107] & layer3_out[1108];
     layer4_out[746] <= ~layer3_out[962];
     layer4_out[747] <= ~layer3_out[457];
     layer4_out[748] <= layer3_out[212];
     layer4_out[749] <= ~layer3_out[678];
     layer4_out[750] <= layer3_out[1366];
     layer4_out[751] <= ~layer3_out[249] | layer3_out[250];
     layer4_out[752] <= 1'b0;
     layer4_out[753] <= ~layer3_out[481];
     layer4_out[754] <= ~layer3_out[242];
     layer4_out[755] <= ~layer3_out[1309];
     layer4_out[756] <= ~layer3_out[268];
     layer4_out[757] <= layer3_out[22] & layer3_out[23];
     layer4_out[758] <= ~layer3_out[1097];
     layer4_out[759] <= ~(layer3_out[616] & layer3_out[617]);
     layer4_out[760] <= ~layer3_out[1142];
     layer4_out[761] <= 1'b0;
     layer4_out[762] <= 1'b1;
     layer4_out[763] <= ~layer3_out[747];
     layer4_out[764] <= ~(layer3_out[1291] & layer3_out[1292]);
     layer4_out[765] <= ~layer3_out[956] | layer3_out[957];
     layer4_out[766] <= layer3_out[1446] | layer3_out[1447];
     layer4_out[767] <= ~(layer3_out[1172] & layer3_out[1173]);
     layer4_out[768] <= ~layer3_out[87];
     layer4_out[769] <= layer3_out[1103];
     layer4_out[770] <= ~layer3_out[1320];
     layer4_out[771] <= ~layer3_out[1264];
     layer4_out[772] <= ~layer3_out[185] | layer3_out[184];
     layer4_out[773] <= ~layer3_out[215] | layer3_out[216];
     layer4_out[774] <= layer3_out[275];
     layer4_out[775] <= layer3_out[887];
     layer4_out[776] <= ~layer3_out[577] | layer3_out[576];
     layer4_out[777] <= layer3_out[224];
     layer4_out[778] <= ~layer3_out[65];
     layer4_out[779] <= ~(layer3_out[154] | layer3_out[155]);
     layer4_out[780] <= layer3_out[1334] & layer3_out[1335];
     layer4_out[781] <= layer3_out[1484] & ~layer3_out[1485];
     layer4_out[782] <= ~(layer3_out[935] & layer3_out[936]);
     layer4_out[783] <= layer3_out[543] & ~layer3_out[542];
     layer4_out[784] <= layer3_out[1093] & ~layer3_out[1094];
     layer4_out[785] <= layer3_out[1369];
     layer4_out[786] <= 1'b1;
     layer4_out[787] <= ~(layer3_out[164] & layer3_out[165]);
     layer4_out[788] <= layer3_out[497] & layer3_out[498];
     layer4_out[789] <= ~layer3_out[402] | layer3_out[403];
     layer4_out[790] <= layer3_out[241];
     layer4_out[791] <= ~layer3_out[534];
     layer4_out[792] <= ~layer3_out[1066];
     layer4_out[793] <= ~layer3_out[251];
     layer4_out[794] <= layer3_out[1331] ^ layer3_out[1332];
     layer4_out[795] <= layer3_out[1066] & ~layer3_out[1065];
     layer4_out[796] <= layer3_out[82] & layer3_out[83];
     layer4_out[797] <= layer3_out[101] & layer3_out[102];
     layer4_out[798] <= layer3_out[1288] ^ layer3_out[1289];
     layer4_out[799] <= ~(layer3_out[1024] & layer3_out[1025]);
     layer4_out[800] <= layer3_out[557];
     layer4_out[801] <= layer3_out[1263];
     layer4_out[802] <= layer3_out[1211] & ~layer3_out[1210];
     layer4_out[803] <= layer3_out[48] & ~layer3_out[47];
     layer4_out[804] <= ~layer3_out[234];
     layer4_out[805] <= layer3_out[591];
     layer4_out[806] <= layer3_out[198];
     layer4_out[807] <= layer3_out[663];
     layer4_out[808] <= ~(layer3_out[1062] & layer3_out[1063]);
     layer4_out[809] <= layer3_out[687];
     layer4_out[810] <= ~layer3_out[804];
     layer4_out[811] <= layer3_out[1026];
     layer4_out[812] <= layer3_out[1383] | layer3_out[1384];
     layer4_out[813] <= layer3_out[880] & layer3_out[881];
     layer4_out[814] <= layer3_out[451] & ~layer3_out[452];
     layer4_out[815] <= ~(layer3_out[802] & layer3_out[803]);
     layer4_out[816] <= ~layer3_out[765];
     layer4_out[817] <= 1'b0;
     layer4_out[818] <= layer3_out[1001];
     layer4_out[819] <= layer3_out[485];
     layer4_out[820] <= layer3_out[1122] & layer3_out[1123];
     layer4_out[821] <= ~layer3_out[1384];
     layer4_out[822] <= ~layer3_out[919] | layer3_out[920];
     layer4_out[823] <= layer3_out[578];
     layer4_out[824] <= ~layer3_out[125] | layer3_out[126];
     layer4_out[825] <= ~(layer3_out[27] | layer3_out[28]);
     layer4_out[826] <= ~layer3_out[35];
     layer4_out[827] <= ~(layer3_out[199] | layer3_out[200]);
     layer4_out[828] <= layer3_out[1112];
     layer4_out[829] <= ~layer3_out[781] | layer3_out[782];
     layer4_out[830] <= layer3_out[795];
     layer4_out[831] <= layer3_out[178] | layer3_out[179];
     layer4_out[832] <= ~layer3_out[1323];
     layer4_out[833] <= 1'b1;
     layer4_out[834] <= ~layer3_out[175] | layer3_out[174];
     layer4_out[835] <= ~layer3_out[676];
     layer4_out[836] <= layer3_out[1167] | layer3_out[1168];
     layer4_out[837] <= layer3_out[685];
     layer4_out[838] <= layer3_out[758];
     layer4_out[839] <= layer3_out[950] & ~layer3_out[949];
     layer4_out[840] <= layer3_out[1087];
     layer4_out[841] <= ~layer3_out[1488] | layer3_out[1487];
     layer4_out[842] <= ~(layer3_out[1431] | layer3_out[1432]);
     layer4_out[843] <= layer3_out[623];
     layer4_out[844] <= ~(layer3_out[1088] | layer3_out[1089]);
     layer4_out[845] <= ~layer3_out[1185] | layer3_out[1184];
     layer4_out[846] <= layer3_out[900];
     layer4_out[847] <= ~layer3_out[42];
     layer4_out[848] <= ~(layer3_out[977] | layer3_out[978]);
     layer4_out[849] <= layer3_out[1333];
     layer4_out[850] <= ~(layer3_out[1355] & layer3_out[1356]);
     layer4_out[851] <= ~layer3_out[1151];
     layer4_out[852] <= 1'b0;
     layer4_out[853] <= ~layer3_out[1114];
     layer4_out[854] <= layer3_out[996];
     layer4_out[855] <= ~(layer3_out[1126] | layer3_out[1127]);
     layer4_out[856] <= layer3_out[906] & layer3_out[907];
     layer4_out[857] <= 1'b0;
     layer4_out[858] <= layer3_out[985] ^ layer3_out[986];
     layer4_out[859] <= ~layer3_out[1470] | layer3_out[1469];
     layer4_out[860] <= ~layer3_out[396];
     layer4_out[861] <= layer3_out[633] | layer3_out[634];
     layer4_out[862] <= layer3_out[603] & layer3_out[604];
     layer4_out[863] <= ~(layer3_out[873] | layer3_out[874]);
     layer4_out[864] <= layer3_out[1008];
     layer4_out[865] <= layer3_out[730] | layer3_out[731];
     layer4_out[866] <= ~(layer3_out[1403] & layer3_out[1404]);
     layer4_out[867] <= ~layer3_out[228];
     layer4_out[868] <= layer3_out[910];
     layer4_out[869] <= ~layer3_out[856] | layer3_out[855];
     layer4_out[870] <= layer3_out[471];
     layer4_out[871] <= 1'b0;
     layer4_out[872] <= ~layer3_out[675];
     layer4_out[873] <= layer3_out[1467];
     layer4_out[874] <= ~layer3_out[217];
     layer4_out[875] <= layer3_out[419] & ~layer3_out[418];
     layer4_out[876] <= ~layer3_out[1069] | layer3_out[1068];
     layer4_out[877] <= ~layer3_out[703] | layer3_out[702];
     layer4_out[878] <= 1'b0;
     layer4_out[879] <= layer3_out[17];
     layer4_out[880] <= ~layer3_out[904];
     layer4_out[881] <= ~(layer3_out[365] & layer3_out[366]);
     layer4_out[882] <= layer3_out[1272];
     layer4_out[883] <= layer3_out[426] | layer3_out[427];
     layer4_out[884] <= layer3_out[630];
     layer4_out[885] <= ~(layer3_out[793] & layer3_out[794]);
     layer4_out[886] <= layer3_out[206];
     layer4_out[887] <= layer3_out[465] & ~layer3_out[464];
     layer4_out[888] <= layer3_out[1200];
     layer4_out[889] <= ~(layer3_out[839] | layer3_out[840]);
     layer4_out[890] <= layer3_out[1293] ^ layer3_out[1294];
     layer4_out[891] <= ~layer3_out[1363];
     layer4_out[892] <= layer3_out[1158] & layer3_out[1159];
     layer4_out[893] <= 1'b1;
     layer4_out[894] <= ~layer3_out[1212] | layer3_out[1211];
     layer4_out[895] <= ~(layer3_out[1417] & layer3_out[1418]);
     layer4_out[896] <= layer3_out[905] ^ layer3_out[906];
     layer4_out[897] <= ~(layer3_out[739] & layer3_out[740]);
     layer4_out[898] <= layer3_out[970] & ~layer3_out[969];
     layer4_out[899] <= layer3_out[951];
     layer4_out[900] <= ~layer3_out[561];
     layer4_out[901] <= layer3_out[1022];
     layer4_out[902] <= ~layer3_out[127] | layer3_out[126];
     layer4_out[903] <= layer3_out[1050];
     layer4_out[904] <= layer3_out[725] & ~layer3_out[724];
     layer4_out[905] <= ~(layer3_out[297] & layer3_out[298]);
     layer4_out[906] <= layer3_out[456] & ~layer3_out[457];
     layer4_out[907] <= ~layer3_out[648];
     layer4_out[908] <= layer3_out[1133] & ~layer3_out[1134];
     layer4_out[909] <= ~(layer3_out[924] & layer3_out[925]);
     layer4_out[910] <= ~layer3_out[1143];
     layer4_out[911] <= layer3_out[355] | layer3_out[356];
     layer4_out[912] <= ~(layer3_out[106] | layer3_out[107]);
     layer4_out[913] <= ~layer3_out[644] | layer3_out[643];
     layer4_out[914] <= ~layer3_out[124];
     layer4_out[915] <= layer3_out[196];
     layer4_out[916] <= 1'b1;
     layer4_out[917] <= layer3_out[436] & ~layer3_out[435];
     layer4_out[918] <= ~layer3_out[1195] | layer3_out[1194];
     layer4_out[919] <= ~layer3_out[1071];
     layer4_out[920] <= ~layer3_out[1214] | layer3_out[1215];
     layer4_out[921] <= ~(layer3_out[305] | layer3_out[306]);
     layer4_out[922] <= ~layer3_out[803] | layer3_out[804];
     layer4_out[923] <= 1'b0;
     layer4_out[924] <= 1'b0;
     layer4_out[925] <= ~layer3_out[193];
     layer4_out[926] <= ~layer3_out[245];
     layer4_out[927] <= layer3_out[681] | layer3_out[682];
     layer4_out[928] <= layer3_out[66] & ~layer3_out[65];
     layer4_out[929] <= 1'b1;
     layer4_out[930] <= ~layer3_out[721];
     layer4_out[931] <= ~(layer3_out[938] ^ layer3_out[939]);
     layer4_out[932] <= ~layer3_out[174];
     layer4_out[933] <= layer3_out[252] & ~layer3_out[251];
     layer4_out[934] <= layer3_out[264] & ~layer3_out[263];
     layer4_out[935] <= layer3_out[1392] ^ layer3_out[1393];
     layer4_out[936] <= ~layer3_out[1390];
     layer4_out[937] <= ~(layer3_out[510] & layer3_out[511]);
     layer4_out[938] <= ~(layer3_out[715] & layer3_out[716]);
     layer4_out[939] <= ~layer3_out[219] | layer3_out[218];
     layer4_out[940] <= ~layer3_out[1387];
     layer4_out[941] <= 1'b1;
     layer4_out[942] <= ~(layer3_out[921] | layer3_out[922]);
     layer4_out[943] <= ~(layer3_out[1413] | layer3_out[1414]);
     layer4_out[944] <= layer3_out[200] & ~layer3_out[201];
     layer4_out[945] <= layer3_out[1223] & ~layer3_out[1222];
     layer4_out[946] <= layer3_out[113];
     layer4_out[947] <= ~layer3_out[1373];
     layer4_out[948] <= layer3_out[1096];
     layer4_out[949] <= layer3_out[310] | layer3_out[311];
     layer4_out[950] <= ~layer3_out[639];
     layer4_out[951] <= layer3_out[551] | layer3_out[552];
     layer4_out[952] <= layer3_out[1190] & layer3_out[1191];
     layer4_out[953] <= layer3_out[86];
     layer4_out[954] <= layer3_out[518] & ~layer3_out[517];
     layer4_out[955] <= ~layer3_out[785] | layer3_out[784];
     layer4_out[956] <= layer3_out[1035];
     layer4_out[957] <= ~layer3_out[494] | layer3_out[493];
     layer4_out[958] <= ~(layer3_out[851] | layer3_out[852]);
     layer4_out[959] <= layer3_out[592] & ~layer3_out[591];
     layer4_out[960] <= ~(layer3_out[419] | layer3_out[420]);
     layer4_out[961] <= ~layer3_out[636] | layer3_out[637];
     layer4_out[962] <= ~layer3_out[189];
     layer4_out[963] <= ~layer3_out[1016];
     layer4_out[964] <= layer3_out[1170] & ~layer3_out[1169];
     layer4_out[965] <= 1'b0;
     layer4_out[966] <= ~layer3_out[547];
     layer4_out[967] <= layer3_out[257] | layer3_out[258];
     layer4_out[968] <= layer3_out[1270];
     layer4_out[969] <= ~layer3_out[1183];
     layer4_out[970] <= layer3_out[772] & ~layer3_out[771];
     layer4_out[971] <= layer3_out[423] & ~layer3_out[422];
     layer4_out[972] <= ~layer3_out[30];
     layer4_out[973] <= ~layer3_out[1303];
     layer4_out[974] <= ~layer3_out[1070];
     layer4_out[975] <= ~layer3_out[176];
     layer4_out[976] <= ~layer3_out[1133] | layer3_out[1132];
     layer4_out[977] <= layer3_out[855];
     layer4_out[978] <= ~layer3_out[586];
     layer4_out[979] <= ~layer3_out[573] | layer3_out[574];
     layer4_out[980] <= ~layer3_out[987] | layer3_out[988];
     layer4_out[981] <= ~layer3_out[255] | layer3_out[256];
     layer4_out[982] <= layer3_out[846];
     layer4_out[983] <= ~layer3_out[945];
     layer4_out[984] <= ~(layer3_out[799] & layer3_out[800]);
     layer4_out[985] <= layer3_out[592] & layer3_out[593];
     layer4_out[986] <= layer3_out[439] & ~layer3_out[440];
     layer4_out[987] <= layer3_out[1195] & layer3_out[1196];
     layer4_out[988] <= layer3_out[566] & ~layer3_out[567];
     layer4_out[989] <= layer3_out[1449];
     layer4_out[990] <= layer3_out[236] | layer3_out[237];
     layer4_out[991] <= 1'b0;
     layer4_out[992] <= ~layer3_out[1231] | layer3_out[1230];
     layer4_out[993] <= ~layer3_out[832] | layer3_out[833];
     layer4_out[994] <= 1'b1;
     layer4_out[995] <= ~layer3_out[895];
     layer4_out[996] <= layer3_out[1218] | layer3_out[1219];
     layer4_out[997] <= layer3_out[796] | layer3_out[797];
     layer4_out[998] <= layer3_out[553] & layer3_out[554];
     layer4_out[999] <= layer3_out[350] & ~layer3_out[351];
     layer4_out[1000] <= 1'b0;
     layer4_out[1001] <= layer3_out[1422] | layer3_out[1423];
     layer4_out[1002] <= layer3_out[958];
     layer4_out[1003] <= ~layer3_out[971];
     layer4_out[1004] <= layer3_out[1309] & layer3_out[1310];
     layer4_out[1005] <= ~(layer3_out[608] & layer3_out[609]);
     layer4_out[1006] <= layer3_out[1151] ^ layer3_out[1152];
     layer4_out[1007] <= layer3_out[1292];
     layer4_out[1008] <= layer3_out[332] & ~layer3_out[333];
     layer4_out[1009] <= ~(layer3_out[736] | layer3_out[737]);
     layer4_out[1010] <= layer3_out[410] ^ layer3_out[411];
     layer4_out[1011] <= layer3_out[1080];
     layer4_out[1012] <= ~(layer3_out[763] & layer3_out[764]);
     layer4_out[1013] <= ~layer3_out[150];
     layer4_out[1014] <= 1'b0;
     layer4_out[1015] <= layer3_out[249];
     layer4_out[1016] <= layer3_out[869] & ~layer3_out[868];
     layer4_out[1017] <= ~(layer3_out[567] & layer3_out[568]);
     layer4_out[1018] <= ~layer3_out[1145] | layer3_out[1146];
     layer4_out[1019] <= layer3_out[238] | layer3_out[239];
     layer4_out[1020] <= ~layer3_out[536];
     layer4_out[1021] <= 1'b0;
     layer4_out[1022] <= ~layer3_out[150];
     layer4_out[1023] <= ~layer3_out[1202];
     layer4_out[1024] <= ~(layer3_out[269] | layer3_out[270]);
     layer4_out[1025] <= layer3_out[1216] | layer3_out[1217];
     layer4_out[1026] <= ~layer3_out[1121];
     layer4_out[1027] <= layer3_out[461] & ~layer3_out[462];
     layer4_out[1028] <= layer3_out[991] & ~layer3_out[992];
     layer4_out[1029] <= ~(layer3_out[1245] & layer3_out[1246]);
     layer4_out[1030] <= layer3_out[576];
     layer4_out[1031] <= ~layer3_out[1327];
     layer4_out[1032] <= layer3_out[838] & ~layer3_out[839];
     layer4_out[1033] <= ~layer3_out[816] | layer3_out[815];
     layer4_out[1034] <= layer3_out[272];
     layer4_out[1035] <= layer3_out[923];
     layer4_out[1036] <= ~layer3_out[50];
     layer4_out[1037] <= layer3_out[207] & ~layer3_out[206];
     layer4_out[1038] <= ~layer3_out[39] | layer3_out[40];
     layer4_out[1039] <= layer3_out[1119] & layer3_out[1120];
     layer4_out[1040] <= ~layer3_out[210];
     layer4_out[1041] <= ~(layer3_out[1294] | layer3_out[1295]);
     layer4_out[1042] <= layer3_out[1280] | layer3_out[1281];
     layer4_out[1043] <= ~layer3_out[35];
     layer4_out[1044] <= 1'b1;
     layer4_out[1045] <= ~layer3_out[140];
     layer4_out[1046] <= ~(layer3_out[1328] | layer3_out[1329]);
     layer4_out[1047] <= ~(layer3_out[862] & layer3_out[863]);
     layer4_out[1048] <= ~layer3_out[194] | layer3_out[193];
     layer4_out[1049] <= ~layer3_out[1241];
     layer4_out[1050] <= ~layer3_out[1229];
     layer4_out[1051] <= ~(layer3_out[963] & layer3_out[964]);
     layer4_out[1052] <= layer3_out[1032] | layer3_out[1033];
     layer4_out[1053] <= layer3_out[1282];
     layer4_out[1054] <= layer3_out[1095];
     layer4_out[1055] <= ~layer3_out[1463];
     layer4_out[1056] <= ~layer3_out[1367];
     layer4_out[1057] <= ~layer3_out[18];
     layer4_out[1058] <= layer3_out[1108];
     layer4_out[1059] <= 1'b1;
     layer4_out[1060] <= layer3_out[326] & ~layer3_out[327];
     layer4_out[1061] <= layer3_out[1100];
     layer4_out[1062] <= 1'b0;
     layer4_out[1063] <= layer3_out[337];
     layer4_out[1064] <= layer3_out[1083] | layer3_out[1084];
     layer4_out[1065] <= layer3_out[979];
     layer4_out[1066] <= 1'b1;
     layer4_out[1067] <= layer3_out[217] & ~layer3_out[216];
     layer4_out[1068] <= ~(layer3_out[1457] ^ layer3_out[1458]);
     layer4_out[1069] <= layer3_out[1200] & layer3_out[1201];
     layer4_out[1070] <= layer3_out[386] & layer3_out[387];
     layer4_out[1071] <= layer3_out[761] | layer3_out[762];
     layer4_out[1072] <= layer3_out[201] & ~layer3_out[202];
     layer4_out[1073] <= ~layer3_out[124] | layer3_out[123];
     layer4_out[1074] <= layer3_out[797] & ~layer3_out[798];
     layer4_out[1075] <= ~layer3_out[1161];
     layer4_out[1076] <= layer3_out[545] ^ layer3_out[546];
     layer4_out[1077] <= layer3_out[1256];
     layer4_out[1078] <= layer3_out[234] | layer3_out[235];
     layer4_out[1079] <= layer3_out[32];
     layer4_out[1080] <= layer3_out[448] | layer3_out[449];
     layer4_out[1081] <= layer3_out[468] & ~layer3_out[469];
     layer4_out[1082] <= layer3_out[1028];
     layer4_out[1083] <= ~layer3_out[886];
     layer4_out[1084] <= ~layer3_out[325] | layer3_out[324];
     layer4_out[1085] <= ~(layer3_out[1375] | layer3_out[1376]);
     layer4_out[1086] <= layer3_out[302] | layer3_out[303];
     layer4_out[1087] <= ~layer3_out[143] | layer3_out[142];
     layer4_out[1088] <= layer3_out[825] | layer3_out[826];
     layer4_out[1089] <= layer3_out[1260] & ~layer3_out[1261];
     layer4_out[1090] <= ~layer3_out[586] | layer3_out[587];
     layer4_out[1091] <= ~layer3_out[511] | layer3_out[512];
     layer4_out[1092] <= ~layer3_out[1473] | layer3_out[1472];
     layer4_out[1093] <= layer3_out[47];
     layer4_out[1094] <= layer3_out[232] & ~layer3_out[233];
     layer4_out[1095] <= ~layer3_out[467];
     layer4_out[1096] <= layer3_out[382] | layer3_out[383];
     layer4_out[1097] <= layer3_out[1477] & layer3_out[1478];
     layer4_out[1098] <= ~layer3_out[1441];
     layer4_out[1099] <= layer3_out[54] & ~layer3_out[53];
     layer4_out[1100] <= ~(layer3_out[630] & layer3_out[631]);
     layer4_out[1101] <= ~layer3_out[447];
     layer4_out[1102] <= layer3_out[625];
     layer4_out[1103] <= layer3_out[1407];
     layer4_out[1104] <= layer3_out[568] | layer3_out[569];
     layer4_out[1105] <= ~layer3_out[45] | layer3_out[46];
     layer4_out[1106] <= ~(layer3_out[1447] | layer3_out[1448]);
     layer4_out[1107] <= ~layer3_out[798];
     layer4_out[1108] <= ~layer3_out[596] | layer3_out[595];
     layer4_out[1109] <= ~layer3_out[1232] | layer3_out[1233];
     layer4_out[1110] <= ~(layer3_out[1391] | layer3_out[1392]);
     layer4_out[1111] <= ~layer3_out[1220];
     layer4_out[1112] <= layer3_out[724];
     layer4_out[1113] <= layer3_out[1397];
     layer4_out[1114] <= ~layer3_out[1494];
     layer4_out[1115] <= ~(layer3_out[1213] ^ layer3_out[1214]);
     layer4_out[1116] <= layer3_out[529];
     layer4_out[1117] <= layer3_out[726] & layer3_out[727];
     layer4_out[1118] <= ~layer3_out[808];
     layer4_out[1119] <= ~layer3_out[371];
     layer4_out[1120] <= layer3_out[848];
     layer4_out[1121] <= layer3_out[1442];
     layer4_out[1122] <= ~layer3_out[1136] | layer3_out[1137];
     layer4_out[1123] <= ~layer3_out[975];
     layer4_out[1124] <= ~(layer3_out[1] | layer3_out[2]);
     layer4_out[1125] <= ~layer3_out[246];
     layer4_out[1126] <= ~layer3_out[852];
     layer4_out[1127] <= layer3_out[532];
     layer4_out[1128] <= layer3_out[231];
     layer4_out[1129] <= layer3_out[470] & layer3_out[471];
     layer4_out[1130] <= ~layer3_out[278];
     layer4_out[1131] <= layer3_out[203] & ~layer3_out[204];
     layer4_out[1132] <= ~layer3_out[1301] | layer3_out[1300];
     layer4_out[1133] <= layer3_out[948] & layer3_out[949];
     layer4_out[1134] <= ~layer3_out[159] | layer3_out[160];
     layer4_out[1135] <= 1'b1;
     layer4_out[1136] <= ~(layer3_out[597] | layer3_out[598]);
     layer4_out[1137] <= ~layer3_out[1319] | layer3_out[1318];
     layer4_out[1138] <= layer3_out[713] ^ layer3_out[714];
     layer4_out[1139] <= ~layer3_out[684] | layer3_out[683];
     layer4_out[1140] <= ~layer3_out[525] | layer3_out[524];
     layer4_out[1141] <= ~(layer3_out[1385] & layer3_out[1386]);
     layer4_out[1142] <= layer3_out[161];
     layer4_out[1143] <= layer3_out[1137] & layer3_out[1138];
     layer4_out[1144] <= layer3_out[844];
     layer4_out[1145] <= ~layer3_out[916];
     layer4_out[1146] <= layer3_out[287];
     layer4_out[1147] <= ~layer3_out[137];
     layer4_out[1148] <= ~(layer3_out[501] | layer3_out[502]);
     layer4_out[1149] <= layer3_out[1239] | layer3_out[1240];
     layer4_out[1150] <= layer3_out[672];
     layer4_out[1151] <= layer3_out[775];
     layer4_out[1152] <= layer3_out[388];
     layer4_out[1153] <= layer3_out[1482] & ~layer3_out[1483];
     layer4_out[1154] <= layer3_out[475] & layer3_out[476];
     layer4_out[1155] <= layer3_out[778] & layer3_out[779];
     layer4_out[1156] <= ~layer3_out[342];
     layer4_out[1157] <= layer3_out[658] & ~layer3_out[659];
     layer4_out[1158] <= layer3_out[837] & layer3_out[838];
     layer4_out[1159] <= ~(layer3_out[1418] & layer3_out[1419]);
     layer4_out[1160] <= layer3_out[1019] | layer3_out[1020];
     layer4_out[1161] <= layer3_out[1149] & layer3_out[1150];
     layer4_out[1162] <= ~(layer3_out[1299] | layer3_out[1300]);
     layer4_out[1163] <= layer3_out[1042] ^ layer3_out[1043];
     layer4_out[1164] <= layer3_out[119] & ~layer3_out[120];
     layer4_out[1165] <= layer3_out[847] & ~layer3_out[848];
     layer4_out[1166] <= 1'b1;
     layer4_out[1167] <= layer3_out[1311] & ~layer3_out[1312];
     layer4_out[1168] <= layer3_out[861];
     layer4_out[1169] <= layer3_out[1042];
     layer4_out[1170] <= layer3_out[939] & ~layer3_out[940];
     layer4_out[1171] <= ~(layer3_out[14] | layer3_out[15]);
     layer4_out[1172] <= ~layer3_out[1164];
     layer4_out[1173] <= layer3_out[1231] & layer3_out[1232];
     layer4_out[1174] <= ~layer3_out[311];
     layer4_out[1175] <= ~layer3_out[371] | layer3_out[372];
     layer4_out[1176] <= ~(layer3_out[55] & layer3_out[56]);
     layer4_out[1177] <= layer3_out[644];
     layer4_out[1178] <= ~layer3_out[823];
     layer4_out[1179] <= layer3_out[356];
     layer4_out[1180] <= layer3_out[1315] & ~layer3_out[1316];
     layer4_out[1181] <= ~layer3_out[454] | layer3_out[453];
     layer4_out[1182] <= ~(layer3_out[134] & layer3_out[135]);
     layer4_out[1183] <= layer3_out[974];
     layer4_out[1184] <= 1'b1;
     layer4_out[1185] <= ~layer3_out[631];
     layer4_out[1186] <= ~layer3_out[9];
     layer4_out[1187] <= layer3_out[67] & ~layer3_out[68];
     layer4_out[1188] <= ~layer3_out[583] | layer3_out[584];
     layer4_out[1189] <= ~(layer3_out[146] & layer3_out[147]);
     layer4_out[1190] <= layer3_out[813];
     layer4_out[1191] <= ~layer3_out[951];
     layer4_out[1192] <= ~(layer3_out[261] ^ layer3_out[262]);
     layer4_out[1193] <= ~layer3_out[442] | layer3_out[443];
     layer4_out[1194] <= ~layer3_out[1073];
     layer4_out[1195] <= 1'b1;
     layer4_out[1196] <= layer3_out[1236] & ~layer3_out[1235];
     layer4_out[1197] <= layer3_out[960] & layer3_out[961];
     layer4_out[1198] <= 1'b0;
     layer4_out[1199] <= layer3_out[372] & ~layer3_out[373];
     layer4_out[1200] <= layer3_out[588];
     layer4_out[1201] <= ~layer3_out[1324];
     layer4_out[1202] <= layer3_out[347] & ~layer3_out[346];
     layer4_out[1203] <= layer3_out[76] & ~layer3_out[75];
     layer4_out[1204] <= ~(layer3_out[38] | layer3_out[39]);
     layer4_out[1205] <= layer3_out[1060] | layer3_out[1061];
     layer4_out[1206] <= ~layer3_out[87];
     layer4_out[1207] <= layer3_out[699];
     layer4_out[1208] <= layer3_out[226];
     layer4_out[1209] <= layer3_out[431];
     layer4_out[1210] <= layer3_out[695] & ~layer3_out[694];
     layer4_out[1211] <= ~layer3_out[90] | layer3_out[91];
     layer4_out[1212] <= layer3_out[1335];
     layer4_out[1213] <= ~layer3_out[1208] | layer3_out[1207];
     layer4_out[1214] <= layer3_out[1037];
     layer4_out[1215] <= layer3_out[1296] & layer3_out[1297];
     layer4_out[1216] <= layer3_out[294];
     layer4_out[1217] <= ~layer3_out[958];
     layer4_out[1218] <= layer3_out[1059] & layer3_out[1060];
     layer4_out[1219] <= layer3_out[289];
     layer4_out[1220] <= layer3_out[891] | layer3_out[892];
     layer4_out[1221] <= layer3_out[1026] & ~layer3_out[1027];
     layer4_out[1222] <= layer3_out[513] & ~layer3_out[514];
     layer4_out[1223] <= layer3_out[690];
     layer4_out[1224] <= ~layer3_out[1062];
     layer4_out[1225] <= ~(layer3_out[645] & layer3_out[646]);
     layer4_out[1226] <= ~layer3_out[1388];
     layer4_out[1227] <= ~layer3_out[773];
     layer4_out[1228] <= layer3_out[1227] & ~layer3_out[1228];
     layer4_out[1229] <= ~layer3_out[1497] | layer3_out[1496];
     layer4_out[1230] <= ~layer3_out[270];
     layer4_out[1231] <= layer3_out[931];
     layer4_out[1232] <= layer3_out[571] ^ layer3_out[572];
     layer4_out[1233] <= 1'b1;
     layer4_out[1234] <= ~layer3_out[769] | layer3_out[768];
     layer4_out[1235] <= ~layer3_out[728] | layer3_out[729];
     layer4_out[1236] <= layer3_out[1224] & layer3_out[1225];
     layer4_out[1237] <= layer3_out[699];
     layer4_out[1238] <= ~(layer3_out[1064] | layer3_out[1065]);
     layer4_out[1239] <= layer3_out[759] | layer3_out[760];
     layer4_out[1240] <= layer3_out[1492];
     layer4_out[1241] <= layer3_out[1410] & ~layer3_out[1411];
     layer4_out[1242] <= layer3_out[994] | layer3_out[995];
     layer4_out[1243] <= ~(layer3_out[109] & layer3_out[110]);
     layer4_out[1244] <= ~(layer3_out[1346] ^ layer3_out[1347]);
     layer4_out[1245] <= ~(layer3_out[1101] & layer3_out[1102]);
     layer4_out[1246] <= 1'b0;
     layer4_out[1247] <= ~(layer3_out[262] & layer3_out[263]);
     layer4_out[1248] <= layer3_out[1187];
     layer4_out[1249] <= layer3_out[1183] | layer3_out[1184];
     layer4_out[1250] <= 1'b1;
     layer4_out[1251] <= layer3_out[0] ^ layer3_out[1];
     layer4_out[1252] <= layer3_out[628] | layer3_out[629];
     layer4_out[1253] <= 1'b0;
     layer4_out[1254] <= ~layer3_out[908];
     layer4_out[1255] <= ~(layer3_out[916] | layer3_out[917]);
     layer4_out[1256] <= layer3_out[7];
     layer4_out[1257] <= 1'b1;
     layer4_out[1258] <= layer3_out[929];
     layer4_out[1259] <= layer3_out[25];
     layer4_out[1260] <= layer3_out[202] & layer3_out[203];
     layer4_out[1261] <= layer3_out[901];
     layer4_out[1262] <= ~layer3_out[601];
     layer4_out[1263] <= layer3_out[171];
     layer4_out[1264] <= layer3_out[606] | layer3_out[607];
     layer4_out[1265] <= ~layer3_out[1435];
     layer4_out[1266] <= layer3_out[997];
     layer4_out[1267] <= ~(layer3_out[833] | layer3_out[834]);
     layer4_out[1268] <= ~layer3_out[872] | layer3_out[871];
     layer4_out[1269] <= layer3_out[429] | layer3_out[430];
     layer4_out[1270] <= ~(layer3_out[1427] | layer3_out[1428]);
     layer4_out[1271] <= ~layer3_out[382];
     layer4_out[1272] <= layer3_out[1090];
     layer4_out[1273] <= layer3_out[1188];
     layer4_out[1274] <= layer3_out[562] & ~layer3_out[563];
     layer4_out[1275] <= layer3_out[444];
     layer4_out[1276] <= ~layer3_out[1053] | layer3_out[1054];
     layer4_out[1277] <= ~layer3_out[610] | layer3_out[609];
     layer4_out[1278] <= layer3_out[914] & layer3_out[915];
     layer4_out[1279] <= layer3_out[736] & ~layer3_out[735];
     layer4_out[1280] <= layer3_out[1159] ^ layer3_out[1160];
     layer4_out[1281] <= layer3_out[516] & layer3_out[517];
     layer4_out[1282] <= layer3_out[1147] & layer3_out[1148];
     layer4_out[1283] <= ~layer3_out[459];
     layer4_out[1284] <= ~(layer3_out[874] ^ layer3_out[875]);
     layer4_out[1285] <= layer3_out[1130] & ~layer3_out[1129];
     layer4_out[1286] <= ~(layer3_out[904] | layer3_out[905]);
     layer4_out[1287] <= ~layer3_out[1125] | layer3_out[1124];
     layer4_out[1288] <= ~layer3_out[1441] | layer3_out[1442];
     layer4_out[1289] <= layer3_out[132] & layer3_out[133];
     layer4_out[1290] <= layer3_out[77];
     layer4_out[1291] <= ~layer3_out[717] | layer3_out[718];
     layer4_out[1292] <= ~layer3_out[756] | layer3_out[755];
     layer4_out[1293] <= ~layer3_out[998];
     layer4_out[1294] <= layer3_out[1023] ^ layer3_out[1024];
     layer4_out[1295] <= layer3_out[657];
     layer4_out[1296] <= layer3_out[594] & ~layer3_out[595];
     layer4_out[1297] <= ~layer3_out[1048];
     layer4_out[1298] <= layer3_out[1157];
     layer4_out[1299] <= ~layer3_out[222];
     layer4_out[1300] <= layer3_out[1304] & layer3_out[1305];
     layer4_out[1301] <= ~(layer3_out[920] | layer3_out[921]);
     layer4_out[1302] <= ~(layer3_out[390] & layer3_out[391]);
     layer4_out[1303] <= ~layer3_out[548];
     layer4_out[1304] <= layer3_out[907] & ~layer3_out[908];
     layer4_out[1305] <= layer3_out[708] | layer3_out[709];
     layer4_out[1306] <= 1'b1;
     layer4_out[1307] <= ~layer3_out[93];
     layer4_out[1308] <= layer3_out[8] & ~layer3_out[7];
     layer4_out[1309] <= ~layer3_out[439] | layer3_out[438];
     layer4_out[1310] <= layer3_out[1091];
     layer4_out[1311] <= ~layer3_out[510];
     layer4_out[1312] <= ~layer3_out[60] | layer3_out[59];
     layer4_out[1313] <= ~(layer3_out[1022] ^ layer3_out[1023]);
     layer4_out[1314] <= ~(layer3_out[863] | layer3_out[864]);
     layer4_out[1315] <= layer3_out[982] & ~layer3_out[983];
     layer4_out[1316] <= layer3_out[996] & ~layer3_out[997];
     layer4_out[1317] <= layer3_out[884];
     layer4_out[1318] <= layer3_out[154] & ~layer3_out[153];
     layer4_out[1319] <= layer3_out[53] & ~layer3_out[52];
     layer4_out[1320] <= layer3_out[1438];
     layer4_out[1321] <= layer3_out[133] & layer3_out[134];
     layer4_out[1322] <= layer3_out[308] & layer3_out[309];
     layer4_out[1323] <= layer3_out[21] & ~layer3_out[20];
     layer4_out[1324] <= layer3_out[898] | layer3_out[899];
     layer4_out[1325] <= ~layer3_out[1337] | layer3_out[1336];
     layer4_out[1326] <= layer3_out[375];
     layer4_out[1327] <= ~(layer3_out[640] | layer3_out[641]);
     layer4_out[1328] <= ~layer3_out[388];
     layer4_out[1329] <= ~layer3_out[618];
     layer4_out[1330] <= ~layer3_out[1352] | layer3_out[1351];
     layer4_out[1331] <= 1'b1;
     layer4_out[1332] <= layer3_out[1012] | layer3_out[1013];
     layer4_out[1333] <= ~(layer3_out[743] ^ layer3_out[744]);
     layer4_out[1334] <= 1'b1;
     layer4_out[1335] <= layer3_out[38] & ~layer3_out[37];
     layer4_out[1336] <= layer3_out[1339] | layer3_out[1340];
     layer4_out[1337] <= ~(layer3_out[120] | layer3_out[121]);
     layer4_out[1338] <= layer3_out[487];
     layer4_out[1339] <= layer3_out[1443];
     layer4_out[1340] <= layer3_out[1077] | layer3_out[1078];
     layer4_out[1341] <= layer3_out[70];
     layer4_out[1342] <= 1'b0;
     layer4_out[1343] <= ~layer3_out[923];
     layer4_out[1344] <= ~layer3_out[119] | layer3_out[118];
     layer4_out[1345] <= layer3_out[435] & ~layer3_out[434];
     layer4_out[1346] <= layer3_out[1371] | layer3_out[1372];
     layer4_out[1347] <= 1'b0;
     layer4_out[1348] <= layer3_out[192];
     layer4_out[1349] <= layer3_out[67];
     layer4_out[1350] <= ~layer3_out[753];
     layer4_out[1351] <= layer3_out[590];
     layer4_out[1352] <= ~(layer3_out[1011] | layer3_out[1012]);
     layer4_out[1353] <= ~(layer3_out[844] | layer3_out[845]);
     layer4_out[1354] <= ~(layer3_out[157] | layer3_out[158]);
     layer4_out[1355] <= ~layer3_out[870] | layer3_out[871];
     layer4_out[1356] <= ~layer3_out[1196];
     layer4_out[1357] <= layer3_out[1395] & layer3_out[1396];
     layer4_out[1358] <= ~layer3_out[1117] | layer3_out[1116];
     layer4_out[1359] <= layer3_out[309] & ~layer3_out[310];
     layer4_out[1360] <= layer3_out[1339];
     layer4_out[1361] <= ~layer3_out[1185];
     layer4_out[1362] <= layer3_out[180];
     layer4_out[1363] <= layer3_out[1359];
     layer4_out[1364] <= ~(layer3_out[1268] | layer3_out[1269]);
     layer4_out[1365] <= layer3_out[141];
     layer4_out[1366] <= layer3_out[308];
     layer4_out[1367] <= 1'b0;
     layer4_out[1368] <= layer3_out[574] & ~layer3_out[575];
     layer4_out[1369] <= layer3_out[888] & ~layer3_out[889];
     layer4_out[1370] <= layer3_out[342] | layer3_out[343];
     layer4_out[1371] <= ~(layer3_out[1329] | layer3_out[1330]);
     layer4_out[1372] <= ~layer3_out[1458] | layer3_out[1459];
     layer4_out[1373] <= ~layer3_out[319];
     layer4_out[1374] <= ~layer3_out[1147];
     layer4_out[1375] <= ~layer3_out[1165] | layer3_out[1164];
     layer4_out[1376] <= ~(layer3_out[398] & layer3_out[399]);
     layer4_out[1377] <= layer3_out[1333];
     layer4_out[1378] <= 1'b1;
     layer4_out[1379] <= ~layer3_out[1323];
     layer4_out[1380] <= ~layer3_out[331];
     layer4_out[1381] <= ~layer3_out[841] | layer3_out[842];
     layer4_out[1382] <= layer3_out[665] & ~layer3_out[664];
     layer4_out[1383] <= layer3_out[1081];
     layer4_out[1384] <= ~(layer3_out[300] | layer3_out[301]);
     layer4_out[1385] <= layer3_out[489] | layer3_out[490];
     layer4_out[1386] <= layer3_out[1405];
     layer4_out[1387] <= layer3_out[168] & ~layer3_out[169];
     layer4_out[1388] <= 1'b0;
     layer4_out[1389] <= layer3_out[128];
     layer4_out[1390] <= ~layer3_out[1338] | layer3_out[1337];
     layer4_out[1391] <= layer3_out[948] & ~layer3_out[947];
     layer4_out[1392] <= 1'b0;
     layer4_out[1393] <= layer3_out[51] | layer3_out[52];
     layer4_out[1394] <= layer3_out[1275] & ~layer3_out[1274];
     layer4_out[1395] <= layer3_out[373] & ~layer3_out[374];
     layer4_out[1396] <= 1'b1;
     layer4_out[1397] <= layer3_out[403] & layer3_out[404];
     layer4_out[1398] <= layer3_out[476] & ~layer3_out[477];
     layer4_out[1399] <= ~layer3_out[926] | layer3_out[925];
     layer4_out[1400] <= ~layer3_out[256] | layer3_out[257];
     layer4_out[1401] <= ~(layer3_out[1305] & layer3_out[1306]);
     layer4_out[1402] <= ~layer3_out[836];
     layer4_out[1403] <= ~layer3_out[1313];
     layer4_out[1404] <= ~layer3_out[1204] | layer3_out[1205];
     layer4_out[1405] <= ~layer3_out[942];
     layer4_out[1406] <= ~(layer3_out[738] & layer3_out[739]);
     layer4_out[1407] <= ~(layer3_out[1168] | layer3_out[1169]);
     layer4_out[1408] <= layer3_out[688] & layer3_out[689];
     layer4_out[1409] <= ~(layer3_out[1109] | layer3_out[1110]);
     layer4_out[1410] <= 1'b0;
     layer4_out[1411] <= ~layer3_out[446] | layer3_out[445];
     layer4_out[1412] <= layer3_out[130];
     layer4_out[1413] <= ~layer3_out[423];
     layer4_out[1414] <= layer3_out[1125];
     layer4_out[1415] <= ~(layer3_out[259] | layer3_out[260]);
     layer4_out[1416] <= ~layer3_out[1490] | layer3_out[1489];
     layer4_out[1417] <= layer3_out[1258] | layer3_out[1259];
     layer4_out[1418] <= layer3_out[1117] & layer3_out[1118];
     layer4_out[1419] <= ~layer3_out[213] | layer3_out[212];
     layer4_out[1420] <= ~(layer3_out[1043] & layer3_out[1044]);
     layer4_out[1421] <= layer3_out[1451] & ~layer3_out[1452];
     layer4_out[1422] <= layer3_out[1283];
     layer4_out[1423] <= ~(layer3_out[57] & layer3_out[58]);
     layer4_out[1424] <= ~layer3_out[103];
     layer4_out[1425] <= layer3_out[740] & layer3_out[741];
     layer4_out[1426] <= ~layer3_out[1445] | layer3_out[1446];
     layer4_out[1427] <= layer3_out[754] | layer3_out[755];
     layer4_out[1428] <= layer3_out[1287] & layer3_out[1288];
     layer4_out[1429] <= ~(layer3_out[1010] | layer3_out[1011]);
     layer4_out[1430] <= layer3_out[1361] | layer3_out[1362];
     layer4_out[1431] <= ~layer3_out[106] | layer3_out[105];
     layer4_out[1432] <= layer3_out[1259];
     layer4_out[1433] <= layer3_out[1283];
     layer4_out[1434] <= layer3_out[801] & layer3_out[802];
     layer4_out[1435] <= layer3_out[1455];
     layer4_out[1436] <= layer3_out[674] & ~layer3_out[673];
     layer4_out[1437] <= ~(layer3_out[1429] & layer3_out[1430]);
     layer4_out[1438] <= ~layer3_out[81];
     layer4_out[1439] <= ~layer3_out[1047];
     layer4_out[1440] <= layer3_out[383];
     layer4_out[1441] <= layer3_out[254] & ~layer3_out[255];
     layer4_out[1442] <= ~layer3_out[555];
     layer4_out[1443] <= ~layer3_out[738];
     layer4_out[1444] <= layer3_out[1464] & layer3_out[1465];
     layer4_out[1445] <= layer3_out[820] & layer3_out[821];
     layer4_out[1446] <= layer3_out[654] & layer3_out[655];
     layer4_out[1447] <= layer3_out[545];
     layer4_out[1448] <= layer3_out[782];
     layer4_out[1449] <= layer3_out[1307];
     layer4_out[1450] <= layer3_out[1486] | layer3_out[1487];
     layer4_out[1451] <= ~layer3_out[63] | layer3_out[64];
     layer4_out[1452] <= layer3_out[571] & ~layer3_out[570];
     layer4_out[1453] <= layer3_out[183];
     layer4_out[1454] <= ~layer3_out[505];
     layer4_out[1455] <= layer3_out[116] & ~layer3_out[117];
     layer4_out[1456] <= ~layer3_out[56] | layer3_out[57];
     layer4_out[1457] <= ~layer3_out[109];
     layer4_out[1458] <= ~(layer3_out[579] | layer3_out[580]);
     layer4_out[1459] <= layer3_out[633];
     layer4_out[1460] <= 1'b1;
     layer4_out[1461] <= ~(layer3_out[766] & layer3_out[767]);
     layer4_out[1462] <= ~(layer3_out[962] ^ layer3_out[963]);
     layer4_out[1463] <= layer3_out[352];
     layer4_out[1464] <= layer3_out[980] | layer3_out[981];
     layer4_out[1465] <= ~layer3_out[1376];
     layer4_out[1466] <= ~(layer3_out[1225] & layer3_out[1226]);
     layer4_out[1467] <= ~layer3_out[412] | layer3_out[413];
     layer4_out[1468] <= layer3_out[483] & ~layer3_out[484];
     layer4_out[1469] <= layer3_out[1479] & ~layer3_out[1480];
     layer4_out[1470] <= ~layer3_out[846];
     layer4_out[1471] <= ~(layer3_out[1251] | layer3_out[1252]);
     layer4_out[1472] <= ~layer3_out[757] | layer3_out[758];
     layer4_out[1473] <= ~layer3_out[1481];
     layer4_out[1474] <= layer3_out[467] & layer3_out[468];
     layer4_out[1475] <= layer3_out[44] & ~layer3_out[43];
     layer4_out[1476] <= layer3_out[1258];
     layer4_out[1477] <= layer3_out[1182];
     layer4_out[1478] <= layer3_out[877] | layer3_out[878];
     layer4_out[1479] <= layer3_out[608] & ~layer3_out[607];
     layer4_out[1480] <= layer3_out[697] ^ layer3_out[698];
     layer4_out[1481] <= layer3_out[801] & ~layer3_out[800];
     layer4_out[1482] <= ~(layer3_out[978] ^ layer3_out[979]);
     layer4_out[1483] <= layer3_out[319] & layer3_out[320];
     layer4_out[1484] <= ~layer3_out[1354] | layer3_out[1353];
     layer4_out[1485] <= ~(layer3_out[4] | layer3_out[5]);
     layer4_out[1486] <= layer3_out[1163] & ~layer3_out[1162];
     layer4_out[1487] <= ~layer3_out[385];
     layer4_out[1488] <= ~layer3_out[897];
     layer4_out[1489] <= ~layer3_out[131] | layer3_out[130];
     layer4_out[1490] <= layer3_out[525] ^ layer3_out[526];
     layer4_out[1491] <= layer3_out[1266];
     layer4_out[1492] <= layer3_out[68] | layer3_out[69];
     layer4_out[1493] <= ~layer3_out[851];
     layer4_out[1494] <= layer3_out[97];
     layer4_out[1495] <= 1'b1;
     layer4_out[1496] <= layer3_out[706] & ~layer3_out[705];
     layer4_out[1497] <= ~(layer3_out[378] & layer3_out[379]);
     layer4_out[1498] <= layer3_out[1037];
     layer4_out[1499] <= ~layer3_out[613] | layer3_out[612];
     layer5_out[0] <= layer4_out[411];
     layer5_out[1] <= ~(layer4_out[980] | layer4_out[981]);
     layer5_out[2] <= layer4_out[1098];
     layer5_out[3] <= ~layer4_out[354] | layer4_out[353];
     layer5_out[4] <= layer4_out[428];
     layer5_out[5] <= ~layer4_out[280];
     layer5_out[6] <= layer4_out[305];
     layer5_out[7] <= ~(layer4_out[427] ^ layer4_out[428]);
     layer5_out[8] <= layer4_out[25];
     layer5_out[9] <= ~(layer4_out[1435] | layer4_out[1436]);
     layer5_out[10] <= ~layer4_out[504] | layer4_out[503];
     layer5_out[11] <= layer4_out[100] & ~layer4_out[101];
     layer5_out[12] <= layer4_out[1161];
     layer5_out[13] <= ~(layer4_out[1120] ^ layer4_out[1121]);
     layer5_out[14] <= ~(layer4_out[1083] | layer4_out[1084]);
     layer5_out[15] <= ~layer4_out[1076] | layer4_out[1077];
     layer5_out[16] <= ~(layer4_out[552] ^ layer4_out[553]);
     layer5_out[17] <= layer4_out[1129];
     layer5_out[18] <= layer4_out[892];
     layer5_out[19] <= ~layer4_out[1385];
     layer5_out[20] <= layer4_out[205] & ~layer4_out[206];
     layer5_out[21] <= ~(layer4_out[1293] ^ layer4_out[1294]);
     layer5_out[22] <= ~(layer4_out[247] & layer4_out[248]);
     layer5_out[23] <= ~(layer4_out[701] ^ layer4_out[702]);
     layer5_out[24] <= layer4_out[1290];
     layer5_out[25] <= layer4_out[1472] & ~layer4_out[1473];
     layer5_out[26] <= ~(layer4_out[243] | layer4_out[244]);
     layer5_out[27] <= layer4_out[137];
     layer5_out[28] <= ~layer4_out[789];
     layer5_out[29] <= ~layer4_out[552];
     layer5_out[30] <= ~layer4_out[201] | layer4_out[200];
     layer5_out[31] <= layer4_out[95] ^ layer4_out[96];
     layer5_out[32] <= ~layer4_out[151];
     layer5_out[33] <= layer4_out[210] & ~layer4_out[211];
     layer5_out[34] <= ~layer4_out[645];
     layer5_out[35] <= layer4_out[482] & ~layer4_out[483];
     layer5_out[36] <= ~layer4_out[816];
     layer5_out[37] <= layer4_out[964];
     layer5_out[38] <= layer4_out[1051];
     layer5_out[39] <= layer4_out[1143];
     layer5_out[40] <= layer4_out[354] & layer4_out[355];
     layer5_out[41] <= ~layer4_out[1416];
     layer5_out[42] <= layer4_out[1279] ^ layer4_out[1280];
     layer5_out[43] <= ~layer4_out[835];
     layer5_out[44] <= ~layer4_out[793];
     layer5_out[45] <= layer4_out[734] & ~layer4_out[735];
     layer5_out[46] <= 1'b0;
     layer5_out[47] <= layer4_out[697] & ~layer4_out[698];
     layer5_out[48] <= layer4_out[631];
     layer5_out[49] <= ~layer4_out[1267] | layer4_out[1266];
     layer5_out[50] <= layer4_out[905] & ~layer4_out[904];
     layer5_out[51] <= layer4_out[299] & layer4_out[300];
     layer5_out[52] <= layer4_out[1390];
     layer5_out[53] <= ~(layer4_out[1282] ^ layer4_out[1283]);
     layer5_out[54] <= layer4_out[969] & ~layer4_out[970];
     layer5_out[55] <= ~layer4_out[273];
     layer5_out[56] <= layer4_out[331] | layer4_out[332];
     layer5_out[57] <= ~layer4_out[866] | layer4_out[867];
     layer5_out[58] <= ~layer4_out[494];
     layer5_out[59] <= layer4_out[442] & layer4_out[443];
     layer5_out[60] <= layer4_out[900];
     layer5_out[61] <= ~layer4_out[326] | layer4_out[327];
     layer5_out[62] <= ~layer4_out[45];
     layer5_out[63] <= layer4_out[121] & ~layer4_out[120];
     layer5_out[64] <= layer4_out[1430];
     layer5_out[65] <= ~layer4_out[1463];
     layer5_out[66] <= layer4_out[739] & layer4_out[740];
     layer5_out[67] <= ~layer4_out[493] | layer4_out[492];
     layer5_out[68] <= layer4_out[1088];
     layer5_out[69] <= layer4_out[524] | layer4_out[525];
     layer5_out[70] <= layer4_out[1332] & ~layer4_out[1333];
     layer5_out[71] <= layer4_out[1187] & ~layer4_out[1188];
     layer5_out[72] <= layer4_out[1483];
     layer5_out[73] <= ~(layer4_out[239] & layer4_out[240]);
     layer5_out[74] <= layer4_out[1350];
     layer5_out[75] <= layer4_out[653];
     layer5_out[76] <= layer4_out[521];
     layer5_out[77] <= ~(layer4_out[659] ^ layer4_out[660]);
     layer5_out[78] <= layer4_out[963];
     layer5_out[79] <= layer4_out[1086] | layer4_out[1087];
     layer5_out[80] <= layer4_out[528];
     layer5_out[81] <= ~layer4_out[433];
     layer5_out[82] <= ~layer4_out[351];
     layer5_out[83] <= layer4_out[578];
     layer5_out[84] <= ~layer4_out[712];
     layer5_out[85] <= ~layer4_out[161];
     layer5_out[86] <= ~(layer4_out[1283] & layer4_out[1284]);
     layer5_out[87] <= ~layer4_out[1204] | layer4_out[1203];
     layer5_out[88] <= ~layer4_out[1036] | layer4_out[1037];
     layer5_out[89] <= layer4_out[1117] & ~layer4_out[1118];
     layer5_out[90] <= ~layer4_out[518];
     layer5_out[91] <= 1'b1;
     layer5_out[92] <= layer4_out[543] ^ layer4_out[544];
     layer5_out[93] <= ~layer4_out[925];
     layer5_out[94] <= layer4_out[1372];
     layer5_out[95] <= layer4_out[1389];
     layer5_out[96] <= ~(layer4_out[1483] & layer4_out[1484]);
     layer5_out[97] <= ~layer4_out[918] | layer4_out[917];
     layer5_out[98] <= ~layer4_out[773];
     layer5_out[99] <= ~layer4_out[623];
     layer5_out[100] <= layer4_out[246] & ~layer4_out[245];
     layer5_out[101] <= ~layer4_out[59];
     layer5_out[102] <= ~layer4_out[886];
     layer5_out[103] <= layer4_out[494];
     layer5_out[104] <= layer4_out[212];
     layer5_out[105] <= ~(layer4_out[860] & layer4_out[861]);
     layer5_out[106] <= ~layer4_out[1165] | layer4_out[1166];
     layer5_out[107] <= ~(layer4_out[374] ^ layer4_out[375]);
     layer5_out[108] <= layer4_out[1420];
     layer5_out[109] <= layer4_out[1172] | layer4_out[1173];
     layer5_out[110] <= layer4_out[1303] ^ layer4_out[1304];
     layer5_out[111] <= ~layer4_out[1424];
     layer5_out[112] <= layer4_out[214];
     layer5_out[113] <= layer4_out[173];
     layer5_out[114] <= layer4_out[892] & ~layer4_out[893];
     layer5_out[115] <= layer4_out[803] & layer4_out[804];
     layer5_out[116] <= ~layer4_out[175];
     layer5_out[117] <= ~layer4_out[801] | layer4_out[802];
     layer5_out[118] <= layer4_out[495] & layer4_out[496];
     layer5_out[119] <= layer4_out[283] & ~layer4_out[284];
     layer5_out[120] <= ~layer4_out[1197] | layer4_out[1196];
     layer5_out[121] <= ~(layer4_out[1134] ^ layer4_out[1135]);
     layer5_out[122] <= ~(layer4_out[857] ^ layer4_out[858]);
     layer5_out[123] <= layer4_out[1007];
     layer5_out[124] <= layer4_out[1454];
     layer5_out[125] <= layer4_out[1075];
     layer5_out[126] <= ~(layer4_out[670] & layer4_out[671]);
     layer5_out[127] <= layer4_out[918] ^ layer4_out[919];
     layer5_out[128] <= ~layer4_out[1024] | layer4_out[1023];
     layer5_out[129] <= layer4_out[1034] & ~layer4_out[1033];
     layer5_out[130] <= ~(layer4_out[1287] & layer4_out[1288]);
     layer5_out[131] <= ~layer4_out[80] | layer4_out[79];
     layer5_out[132] <= ~layer4_out[521];
     layer5_out[133] <= ~layer4_out[90] | layer4_out[89];
     layer5_out[134] <= layer4_out[298];
     layer5_out[135] <= ~(layer4_out[1255] & layer4_out[1256]);
     layer5_out[136] <= ~layer4_out[779] | layer4_out[778];
     layer5_out[137] <= ~layer4_out[1020];
     layer5_out[138] <= layer4_out[225] & ~layer4_out[224];
     layer5_out[139] <= layer4_out[430] & ~layer4_out[429];
     layer5_out[140] <= layer4_out[1068] | layer4_out[1069];
     layer5_out[141] <= layer4_out[397] ^ layer4_out[398];
     layer5_out[142] <= layer4_out[421] ^ layer4_out[422];
     layer5_out[143] <= layer4_out[220] & layer4_out[221];
     layer5_out[144] <= layer4_out[683];
     layer5_out[145] <= ~layer4_out[714] | layer4_out[715];
     layer5_out[146] <= ~layer4_out[215] | layer4_out[214];
     layer5_out[147] <= layer4_out[218] & ~layer4_out[219];
     layer5_out[148] <= ~layer4_out[1023] | layer4_out[1022];
     layer5_out[149] <= ~layer4_out[1024];
     layer5_out[150] <= layer4_out[262];
     layer5_out[151] <= layer4_out[438] | layer4_out[439];
     layer5_out[152] <= ~(layer4_out[458] ^ layer4_out[459]);
     layer5_out[153] <= layer4_out[464];
     layer5_out[154] <= ~layer4_out[600] | layer4_out[599];
     layer5_out[155] <= layer4_out[423];
     layer5_out[156] <= layer4_out[743];
     layer5_out[157] <= ~layer4_out[1133];
     layer5_out[158] <= ~layer4_out[903];
     layer5_out[159] <= layer4_out[1064] & layer4_out[1065];
     layer5_out[160] <= ~layer4_out[235] | layer4_out[236];
     layer5_out[161] <= ~layer4_out[437];
     layer5_out[162] <= layer4_out[854] & ~layer4_out[855];
     layer5_out[163] <= layer4_out[744] & layer4_out[745];
     layer5_out[164] <= layer4_out[623] & ~layer4_out[622];
     layer5_out[165] <= ~layer4_out[431];
     layer5_out[166] <= ~layer4_out[546];
     layer5_out[167] <= layer4_out[166];
     layer5_out[168] <= ~layer4_out[737];
     layer5_out[169] <= layer4_out[370];
     layer5_out[170] <= ~layer4_out[1104] | layer4_out[1103];
     layer5_out[171] <= ~(layer4_out[837] & layer4_out[838]);
     layer5_out[172] <= layer4_out[1149];
     layer5_out[173] <= ~layer4_out[822];
     layer5_out[174] <= ~layer4_out[629] | layer4_out[628];
     layer5_out[175] <= layer4_out[1082] & ~layer4_out[1083];
     layer5_out[176] <= layer4_out[1031];
     layer5_out[177] <= layer4_out[567];
     layer5_out[178] <= ~layer4_out[1398];
     layer5_out[179] <= ~(layer4_out[179] & layer4_out[180]);
     layer5_out[180] <= ~layer4_out[1056] | layer4_out[1055];
     layer5_out[181] <= ~(layer4_out[359] & layer4_out[360]);
     layer5_out[182] <= layer4_out[516];
     layer5_out[183] <= layer4_out[408];
     layer5_out[184] <= layer4_out[713] & ~layer4_out[714];
     layer5_out[185] <= layer4_out[824] & layer4_out[825];
     layer5_out[186] <= layer4_out[1361];
     layer5_out[187] <= layer4_out[523];
     layer5_out[188] <= ~layer4_out[1054] | layer4_out[1055];
     layer5_out[189] <= layer4_out[346];
     layer5_out[190] <= ~(layer4_out[488] & layer4_out[489]);
     layer5_out[191] <= layer4_out[1142];
     layer5_out[192] <= ~layer4_out[770] | layer4_out[771];
     layer5_out[193] <= layer4_out[781] | layer4_out[782];
     layer5_out[194] <= layer4_out[1107];
     layer5_out[195] <= ~layer4_out[1064];
     layer5_out[196] <= ~layer4_out[591];
     layer5_out[197] <= layer4_out[153];
     layer5_out[198] <= ~(layer4_out[1154] ^ layer4_out[1155]);
     layer5_out[199] <= layer4_out[1412] & layer4_out[1413];
     layer5_out[200] <= layer4_out[531];
     layer5_out[201] <= ~(layer4_out[1485] & layer4_out[1486]);
     layer5_out[202] <= ~(layer4_out[229] & layer4_out[230]);
     layer5_out[203] <= layer4_out[250];
     layer5_out[204] <= layer4_out[346];
     layer5_out[205] <= layer4_out[1043];
     layer5_out[206] <= layer4_out[652];
     layer5_out[207] <= ~layer4_out[1494];
     layer5_out[208] <= 1'b1;
     layer5_out[209] <= layer4_out[304];
     layer5_out[210] <= 1'b0;
     layer5_out[211] <= ~layer4_out[389];
     layer5_out[212] <= ~(layer4_out[240] ^ layer4_out[241]);
     layer5_out[213] <= ~(layer4_out[414] ^ layer4_out[415]);
     layer5_out[214] <= layer4_out[944];
     layer5_out[215] <= layer4_out[615] ^ layer4_out[616];
     layer5_out[216] <= ~(layer4_out[87] | layer4_out[88]);
     layer5_out[217] <= layer4_out[823] & layer4_out[824];
     layer5_out[218] <= ~layer4_out[790] | layer4_out[791];
     layer5_out[219] <= ~(layer4_out[664] | layer4_out[665]);
     layer5_out[220] <= layer4_out[364] & ~layer4_out[365];
     layer5_out[221] <= layer4_out[942];
     layer5_out[222] <= ~layer4_out[1240] | layer4_out[1241];
     layer5_out[223] <= layer4_out[526];
     layer5_out[224] <= layer4_out[1381];
     layer5_out[225] <= layer4_out[934];
     layer5_out[226] <= ~layer4_out[827] | layer4_out[828];
     layer5_out[227] <= layer4_out[876] & ~layer4_out[875];
     layer5_out[228] <= ~layer4_out[256];
     layer5_out[229] <= layer4_out[1014] & ~layer4_out[1013];
     layer5_out[230] <= layer4_out[120];
     layer5_out[231] <= layer4_out[1052] ^ layer4_out[1053];
     layer5_out[232] <= layer4_out[681] ^ layer4_out[682];
     layer5_out[233] <= ~layer4_out[1140];
     layer5_out[234] <= ~(layer4_out[413] & layer4_out[414]);
     layer5_out[235] <= layer4_out[457];
     layer5_out[236] <= layer4_out[187] & layer4_out[188];
     layer5_out[237] <= ~layer4_out[1231];
     layer5_out[238] <= ~layer4_out[1006];
     layer5_out[239] <= ~layer4_out[441] | layer4_out[442];
     layer5_out[240] <= layer4_out[877];
     layer5_out[241] <= ~layer4_out[512];
     layer5_out[242] <= ~layer4_out[1199] | layer4_out[1200];
     layer5_out[243] <= ~layer4_out[1060];
     layer5_out[244] <= ~(layer4_out[953] & layer4_out[954]);
     layer5_out[245] <= layer4_out[1375];
     layer5_out[246] <= ~layer4_out[1434];
     layer5_out[247] <= layer4_out[636];
     layer5_out[248] <= ~layer4_out[1012];
     layer5_out[249] <= ~(layer4_out[985] & layer4_out[986]);
     layer5_out[250] <= layer4_out[1453];
     layer5_out[251] <= layer4_out[931] & ~layer4_out[932];
     layer5_out[252] <= ~layer4_out[1125];
     layer5_out[253] <= layer4_out[1428] | layer4_out[1429];
     layer5_out[254] <= ~layer4_out[1057];
     layer5_out[255] <= layer4_out[1237] & layer4_out[1238];
     layer5_out[256] <= layer4_out[627] & ~layer4_out[628];
     layer5_out[257] <= ~layer4_out[57];
     layer5_out[258] <= ~(layer4_out[27] ^ layer4_out[28]);
     layer5_out[259] <= ~layer4_out[407] | layer4_out[406];
     layer5_out[260] <= ~layer4_out[1087] | layer4_out[1088];
     layer5_out[261] <= layer4_out[803];
     layer5_out[262] <= ~(layer4_out[535] | layer4_out[536]);
     layer5_out[263] <= layer4_out[1133] & ~layer4_out[1134];
     layer5_out[264] <= ~layer4_out[529];
     layer5_out[265] <= ~(layer4_out[499] & layer4_out[500]);
     layer5_out[266] <= layer4_out[342];
     layer5_out[267] <= layer4_out[1048] & ~layer4_out[1047];
     layer5_out[268] <= layer4_out[1188] ^ layer4_out[1189];
     layer5_out[269] <= layer4_out[1311];
     layer5_out[270] <= layer4_out[951];
     layer5_out[271] <= layer4_out[971];
     layer5_out[272] <= layer4_out[1163] | layer4_out[1164];
     layer5_out[273] <= layer4_out[1169] & ~layer4_out[1168];
     layer5_out[274] <= layer4_out[172] & layer4_out[173];
     layer5_out[275] <= ~(layer4_out[592] & layer4_out[593]);
     layer5_out[276] <= 1'b1;
     layer5_out[277] <= layer4_out[1040];
     layer5_out[278] <= layer4_out[1193] & ~layer4_out[1194];
     layer5_out[279] <= ~(layer4_out[322] ^ layer4_out[323]);
     layer5_out[280] <= layer4_out[555] ^ layer4_out[556];
     layer5_out[281] <= 1'b0;
     layer5_out[282] <= ~layer4_out[640];
     layer5_out[283] <= ~layer4_out[369];
     layer5_out[284] <= ~layer4_out[265] | layer4_out[266];
     layer5_out[285] <= ~layer4_out[1170] | layer4_out[1169];
     layer5_out[286] <= ~layer4_out[180];
     layer5_out[287] <= layer4_out[246] ^ layer4_out[247];
     layer5_out[288] <= ~(layer4_out[1269] & layer4_out[1270]);
     layer5_out[289] <= ~(layer4_out[381] ^ layer4_out[382]);
     layer5_out[290] <= ~layer4_out[427];
     layer5_out[291] <= ~(layer4_out[608] | layer4_out[609]);
     layer5_out[292] <= layer4_out[1150] & layer4_out[1151];
     layer5_out[293] <= ~layer4_out[1356];
     layer5_out[294] <= layer4_out[1387];
     layer5_out[295] <= ~(layer4_out[1179] ^ layer4_out[1180]);
     layer5_out[296] <= 1'b0;
     layer5_out[297] <= layer4_out[1383];
     layer5_out[298] <= layer4_out[545];
     layer5_out[299] <= 1'b0;
     layer5_out[300] <= ~layer4_out[588] | layer4_out[589];
     layer5_out[301] <= ~layer4_out[1371] | layer4_out[1370];
     layer5_out[302] <= layer4_out[1493] | layer4_out[1494];
     layer5_out[303] <= ~layer4_out[46];
     layer5_out[304] <= layer4_out[1030] & ~layer4_out[1029];
     layer5_out[305] <= ~layer4_out[1295];
     layer5_out[306] <= layer4_out[914] ^ layer4_out[915];
     layer5_out[307] <= ~layer4_out[655];
     layer5_out[308] <= layer4_out[1356] & layer4_out[1357];
     layer5_out[309] <= layer4_out[1205] & ~layer4_out[1206];
     layer5_out[310] <= layer4_out[41] & ~layer4_out[42];
     layer5_out[311] <= ~(layer4_out[107] ^ layer4_out[108]);
     layer5_out[312] <= ~layer4_out[1277] | layer4_out[1276];
     layer5_out[313] <= ~layer4_out[777];
     layer5_out[314] <= ~(layer4_out[151] ^ layer4_out[152]);
     layer5_out[315] <= ~layer4_out[1286];
     layer5_out[316] <= layer4_out[1003] | layer4_out[1004];
     layer5_out[317] <= layer4_out[436] & layer4_out[437];
     layer5_out[318] <= layer4_out[3];
     layer5_out[319] <= ~layer4_out[746] | layer4_out[747];
     layer5_out[320] <= ~layer4_out[348] | layer4_out[349];
     layer5_out[321] <= ~(layer4_out[417] ^ layer4_out[418]);
     layer5_out[322] <= ~layer4_out[686];
     layer5_out[323] <= layer4_out[732] & ~layer4_out[731];
     layer5_out[324] <= layer4_out[888];
     layer5_out[325] <= 1'b1;
     layer5_out[326] <= layer4_out[1365];
     layer5_out[327] <= layer4_out[291] & ~layer4_out[290];
     layer5_out[328] <= layer4_out[1058] ^ layer4_out[1059];
     layer5_out[329] <= layer4_out[82];
     layer5_out[330] <= ~(layer4_out[570] & layer4_out[571]);
     layer5_out[331] <= ~(layer4_out[1444] ^ layer4_out[1445]);
     layer5_out[332] <= layer4_out[112];
     layer5_out[333] <= ~layer4_out[1050] | layer4_out[1051];
     layer5_out[334] <= layer4_out[359];
     layer5_out[335] <= ~layer4_out[764];
     layer5_out[336] <= layer4_out[618];
     layer5_out[337] <= layer4_out[78] | layer4_out[79];
     layer5_out[338] <= ~layer4_out[1015];
     layer5_out[339] <= layer4_out[696] | layer4_out[697];
     layer5_out[340] <= layer4_out[1346];
     layer5_out[341] <= ~layer4_out[448];
     layer5_out[342] <= ~layer4_out[864];
     layer5_out[343] <= ~(layer4_out[1398] | layer4_out[1399]);
     layer5_out[344] <= layer4_out[434] & layer4_out[435];
     layer5_out[345] <= ~layer4_out[1148];
     layer5_out[346] <= ~layer4_out[314];
     layer5_out[347] <= ~layer4_out[890];
     layer5_out[348] <= ~(layer4_out[500] & layer4_out[501]);
     layer5_out[349] <= ~(layer4_out[129] & layer4_out[130]);
     layer5_out[350] <= ~layer4_out[70];
     layer5_out[351] <= layer4_out[543];
     layer5_out[352] <= ~layer4_out[1228] | layer4_out[1229];
     layer5_out[353] <= layer4_out[949] & ~layer4_out[948];
     layer5_out[354] <= 1'b0;
     layer5_out[355] <= layer4_out[771] | layer4_out[772];
     layer5_out[356] <= ~layer4_out[1247];
     layer5_out[357] <= ~layer4_out[604];
     layer5_out[358] <= ~layer4_out[1452];
     layer5_out[359] <= layer4_out[748];
     layer5_out[360] <= layer4_out[1226] & ~layer4_out[1225];
     layer5_out[361] <= ~layer4_out[1126];
     layer5_out[362] <= layer4_out[1164] & layer4_out[1165];
     layer5_out[363] <= ~layer4_out[1158] | layer4_out[1159];
     layer5_out[364] <= layer4_out[378] & ~layer4_out[377];
     layer5_out[365] <= ~(layer4_out[404] & layer4_out[405]);
     layer5_out[366] <= ~layer4_out[357] | layer4_out[356];
     layer5_out[367] <= layer4_out[1216];
     layer5_out[368] <= ~layer4_out[1161] | layer4_out[1160];
     layer5_out[369] <= layer4_out[692];
     layer5_out[370] <= ~layer4_out[745];
     layer5_out[371] <= ~(layer4_out[420] ^ layer4_out[421]);
     layer5_out[372] <= ~(layer4_out[91] & layer4_out[92]);
     layer5_out[373] <= ~layer4_out[978] | layer4_out[977];
     layer5_out[374] <= ~(layer4_out[858] | layer4_out[859]);
     layer5_out[375] <= ~layer4_out[975];
     layer5_out[376] <= layer4_out[1370];
     layer5_out[377] <= layer4_out[1456] | layer4_out[1457];
     layer5_out[378] <= ~layer4_out[343];
     layer5_out[379] <= ~(layer4_out[516] | layer4_out[517]);
     layer5_out[380] <= ~layer4_out[1457];
     layer5_out[381] <= layer4_out[105];
     layer5_out[382] <= ~layer4_out[227];
     layer5_out[383] <= layer4_out[801];
     layer5_out[384] <= ~layer4_out[748];
     layer5_out[385] <= ~(layer4_out[1462] ^ layer4_out[1463]);
     layer5_out[386] <= ~layer4_out[35];
     layer5_out[387] <= ~layer4_out[921];
     layer5_out[388] <= ~layer4_out[580] | layer4_out[579];
     layer5_out[389] <= ~layer4_out[1043];
     layer5_out[390] <= 1'b0;
     layer5_out[391] <= layer4_out[767] & ~layer4_out[768];
     layer5_out[392] <= layer4_out[189] & ~layer4_out[188];
     layer5_out[393] <= layer4_out[1346];
     layer5_out[394] <= ~(layer4_out[533] & layer4_out[534]);
     layer5_out[395] <= ~layer4_out[274] | layer4_out[275];
     layer5_out[396] <= ~(layer4_out[258] & layer4_out[259]);
     layer5_out[397] <= layer4_out[103] & layer4_out[104];
     layer5_out[398] <= ~layer4_out[369];
     layer5_out[399] <= ~(layer4_out[1001] ^ layer4_out[1002]);
     layer5_out[400] <= ~(layer4_out[1159] & layer4_out[1160]);
     layer5_out[401] <= ~layer4_out[675];
     layer5_out[402] <= ~(layer4_out[1004] ^ layer4_out[1005]);
     layer5_out[403] <= layer4_out[1096] & ~layer4_out[1097];
     layer5_out[404] <= ~layer4_out[74];
     layer5_out[405] <= layer4_out[1309];
     layer5_out[406] <= 1'b1;
     layer5_out[407] <= layer4_out[39] & ~layer4_out[38];
     layer5_out[408] <= layer4_out[947];
     layer5_out[409] <= ~layer4_out[1414];
     layer5_out[410] <= layer4_out[387] ^ layer4_out[388];
     layer5_out[411] <= ~(layer4_out[909] & layer4_out[910]);
     layer5_out[412] <= ~layer4_out[467];
     layer5_out[413] <= layer4_out[601];
     layer5_out[414] <= layer4_out[1082] & ~layer4_out[1081];
     layer5_out[415] <= ~(layer4_out[1184] & layer4_out[1185]);
     layer5_out[416] <= ~layer4_out[538];
     layer5_out[417] <= layer4_out[738];
     layer5_out[418] <= layer4_out[1236] | layer4_out[1237];
     layer5_out[419] <= ~(layer4_out[636] & layer4_out[637]);
     layer5_out[420] <= ~layer4_out[967];
     layer5_out[421] <= layer4_out[1316] & layer4_out[1317];
     layer5_out[422] <= layer4_out[508] & layer4_out[509];
     layer5_out[423] <= layer4_out[137];
     layer5_out[424] <= layer4_out[594] & ~layer4_out[593];
     layer5_out[425] <= layer4_out[37] ^ layer4_out[38];
     layer5_out[426] <= ~layer4_out[1336] | layer4_out[1335];
     layer5_out[427] <= ~(layer4_out[658] & layer4_out[659]);
     layer5_out[428] <= ~layer4_out[1280];
     layer5_out[429] <= ~layer4_out[264] | layer4_out[263];
     layer5_out[430] <= layer4_out[641] & ~layer4_out[640];
     layer5_out[431] <= layer4_out[273] & ~layer4_out[274];
     layer5_out[432] <= layer4_out[550] | layer4_out[551];
     layer5_out[433] <= layer4_out[709] | layer4_out[710];
     layer5_out[434] <= layer4_out[71] & layer4_out[72];
     layer5_out[435] <= ~layer4_out[478] | layer4_out[479];
     layer5_out[436] <= 1'b1;
     layer5_out[437] <= ~layer4_out[1084];
     layer5_out[438] <= layer4_out[1335] & ~layer4_out[1334];
     layer5_out[439] <= layer4_out[1489] & ~layer4_out[1488];
     layer5_out[440] <= layer4_out[1208] & layer4_out[1209];
     layer5_out[441] <= layer4_out[266] & layer4_out[267];
     layer5_out[442] <= layer4_out[1034] | layer4_out[1035];
     layer5_out[443] <= ~layer4_out[1009];
     layer5_out[444] <= ~layer4_out[145];
     layer5_out[445] <= layer4_out[257] & ~layer4_out[258];
     layer5_out[446] <= ~layer4_out[424];
     layer5_out[447] <= ~(layer4_out[926] | layer4_out[927]);
     layer5_out[448] <= ~(layer4_out[1265] | layer4_out[1266]);
     layer5_out[449] <= ~(layer4_out[1497] | layer4_out[1498]);
     layer5_out[450] <= layer4_out[984];
     layer5_out[451] <= ~layer4_out[508];
     layer5_out[452] <= layer4_out[1433] | layer4_out[1434];
     layer5_out[453] <= layer4_out[1492];
     layer5_out[454] <= ~layer4_out[1305];
     layer5_out[455] <= layer4_out[448] & ~layer4_out[449];
     layer5_out[456] <= layer4_out[63];
     layer5_out[457] <= ~layer4_out[398] | layer4_out[399];
     layer5_out[458] <= layer4_out[1260];
     layer5_out[459] <= layer4_out[879] & layer4_out[880];
     layer5_out[460] <= layer4_out[12] & layer4_out[13];
     layer5_out[461] <= layer4_out[1476];
     layer5_out[462] <= layer4_out[1143];
     layer5_out[463] <= ~layer4_out[686] | layer4_out[687];
     layer5_out[464] <= ~layer4_out[952];
     layer5_out[465] <= layer4_out[836] & layer4_out[837];
     layer5_out[466] <= layer4_out[1182];
     layer5_out[467] <= ~(layer4_out[446] ^ layer4_out[447]);
     layer5_out[468] <= ~layer4_out[1315];
     layer5_out[469] <= layer4_out[1328];
     layer5_out[470] <= layer4_out[1110];
     layer5_out[471] <= ~(layer4_out[719] ^ layer4_out[720]);
     layer5_out[472] <= ~layer4_out[1219] | layer4_out[1218];
     layer5_out[473] <= layer4_out[238] & ~layer4_out[239];
     layer5_out[474] <= layer4_out[567];
     layer5_out[475] <= ~(layer4_out[317] & layer4_out[318]);
     layer5_out[476] <= ~(layer4_out[992] ^ layer4_out[993]);
     layer5_out[477] <= ~layer4_out[762];
     layer5_out[478] <= ~layer4_out[1254] | layer4_out[1255];
     layer5_out[479] <= layer4_out[484] & layer4_out[485];
     layer5_out[480] <= layer4_out[1230] & ~layer4_out[1229];
     layer5_out[481] <= ~(layer4_out[1201] ^ layer4_out[1202]);
     layer5_out[482] <= layer4_out[487];
     layer5_out[483] <= layer4_out[583] ^ layer4_out[584];
     layer5_out[484] <= layer4_out[186] ^ layer4_out[187];
     layer5_out[485] <= layer4_out[1074];
     layer5_out[486] <= ~layer4_out[218];
     layer5_out[487] <= ~layer4_out[363] | layer4_out[364];
     layer5_out[488] <= ~layer4_out[1186];
     layer5_out[489] <= layer4_out[755];
     layer5_out[490] <= ~layer4_out[97];
     layer5_out[491] <= layer4_out[937] | layer4_out[938];
     layer5_out[492] <= layer4_out[158] ^ layer4_out[159];
     layer5_out[493] <= layer4_out[256] & layer4_out[257];
     layer5_out[494] <= layer4_out[1186];
     layer5_out[495] <= ~layer4_out[1392] | layer4_out[1393];
     layer5_out[496] <= layer4_out[1471];
     layer5_out[497] <= layer4_out[960];
     layer5_out[498] <= ~(layer4_out[564] | layer4_out[565]);
     layer5_out[499] <= layer4_out[270] & ~layer4_out[269];
     layer5_out[500] <= ~(layer4_out[455] ^ layer4_out[456]);
     layer5_out[501] <= layer4_out[1461];
     layer5_out[502] <= ~layer4_out[308];
     layer5_out[503] <= ~layer4_out[632] | layer4_out[631];
     layer5_out[504] <= ~layer4_out[139] | layer4_out[138];
     layer5_out[505] <= ~layer4_out[1354];
     layer5_out[506] <= layer4_out[1144] | layer4_out[1145];
     layer5_out[507] <= layer4_out[114] & layer4_out[115];
     layer5_out[508] <= layer4_out[142];
     layer5_out[509] <= ~(layer4_out[961] & layer4_out[962]);
     layer5_out[510] <= layer4_out[455];
     layer5_out[511] <= layer4_out[1312] & ~layer4_out[1311];
     layer5_out[512] <= ~layer4_out[1419] | layer4_out[1420];
     layer5_out[513] <= layer4_out[1440];
     layer5_out[514] <= ~(layer4_out[9] ^ layer4_out[10]);
     layer5_out[515] <= layer4_out[470] & ~layer4_out[471];
     layer5_out[516] <= layer4_out[813] & layer4_out[814];
     layer5_out[517] <= ~(layer4_out[444] ^ layer4_out[445]);
     layer5_out[518] <= ~layer4_out[705];
     layer5_out[519] <= layer4_out[16];
     layer5_out[520] <= ~layer4_out[440];
     layer5_out[521] <= ~layer4_out[177];
     layer5_out[522] <= layer4_out[1181];
     layer5_out[523] <= ~layer4_out[167];
     layer5_out[524] <= ~layer4_out[1017];
     layer5_out[525] <= ~layer4_out[1090] | layer4_out[1089];
     layer5_out[526] <= layer4_out[505];
     layer5_out[527] <= layer4_out[971] & ~layer4_out[972];
     layer5_out[528] <= ~layer4_out[1325];
     layer5_out[529] <= ~(layer4_out[469] | layer4_out[470]);
     layer5_out[530] <= ~layer4_out[734];
     layer5_out[531] <= layer4_out[881];
     layer5_out[532] <= ~(layer4_out[171] | layer4_out[172]);
     layer5_out[533] <= ~layer4_out[1232];
     layer5_out[534] <= layer4_out[722] & layer4_out[723];
     layer5_out[535] <= layer4_out[598] & layer4_out[599];
     layer5_out[536] <= layer4_out[996] ^ layer4_out[997];
     layer5_out[537] <= ~layer4_out[1047];
     layer5_out[538] <= ~layer4_out[838];
     layer5_out[539] <= ~layer4_out[1278];
     layer5_out[540] <= ~layer4_out[1383] | layer4_out[1382];
     layer5_out[541] <= ~layer4_out[620];
     layer5_out[542] <= ~layer4_out[694];
     layer5_out[543] <= ~(layer4_out[942] & layer4_out[943]);
     layer5_out[544] <= layer4_out[386];
     layer5_out[545] <= ~layer4_out[1321];
     layer5_out[546] <= ~layer4_out[1382];
     layer5_out[547] <= ~(layer4_out[1425] & layer4_out[1426]);
     layer5_out[548] <= layer4_out[69] & ~layer4_out[68];
     layer5_out[549] <= layer4_out[724] & ~layer4_out[723];
     layer5_out[550] <= ~layer4_out[583];
     layer5_out[551] <= ~(layer4_out[1093] ^ layer4_out[1094]);
     layer5_out[552] <= layer4_out[702] | layer4_out[703];
     layer5_out[553] <= ~layer4_out[492];
     layer5_out[554] <= ~(layer4_out[935] | layer4_out[936]);
     layer5_out[555] <= layer4_out[1117] & ~layer4_out[1116];
     layer5_out[556] <= ~(layer4_out[910] | layer4_out[911]);
     layer5_out[557] <= layer4_out[609];
     layer5_out[558] <= layer4_out[282] & ~layer4_out[281];
     layer5_out[559] <= layer4_out[401] & ~layer4_out[402];
     layer5_out[560] <= ~(layer4_out[453] | layer4_out[454]);
     layer5_out[561] <= ~(layer4_out[1239] & layer4_out[1240]);
     layer5_out[562] <= layer4_out[1308] ^ layer4_out[1309];
     layer5_out[563] <= layer4_out[1329];
     layer5_out[564] <= layer4_out[768];
     layer5_out[565] <= layer4_out[1062] | layer4_out[1063];
     layer5_out[566] <= ~(layer4_out[840] ^ layer4_out[841]);
     layer5_out[567] <= ~(layer4_out[479] ^ layer4_out[480]);
     layer5_out[568] <= ~layer4_out[540] | layer4_out[541];
     layer5_out[569] <= ~(layer4_out[204] & layer4_out[205]);
     layer5_out[570] <= layer4_out[1408] | layer4_out[1409];
     layer5_out[571] <= layer4_out[1014] & layer4_out[1015];
     layer5_out[572] <= ~layer4_out[487] | layer4_out[486];
     layer5_out[573] <= layer4_out[716] & layer4_out[717];
     layer5_out[574] <= ~(layer4_out[999] ^ layer4_out[1000]);
     layer5_out[575] <= layer4_out[350];
     layer5_out[576] <= ~(layer4_out[1407] & layer4_out[1408]);
     layer5_out[577] <= ~(layer4_out[452] | layer4_out[453]);
     layer5_out[578] <= ~layer4_out[955] | layer4_out[956];
     layer5_out[579] <= ~layer4_out[277] | layer4_out[276];
     layer5_out[580] <= ~layer4_out[1411];
     layer5_out[581] <= layer4_out[1177] & layer4_out[1178];
     layer5_out[582] <= ~layer4_out[1323];
     layer5_out[583] <= ~layer4_out[784] | layer4_out[783];
     layer5_out[584] <= ~layer4_out[718];
     layer5_out[585] <= layer4_out[3] | layer4_out[4];
     layer5_out[586] <= ~(layer4_out[451] ^ layer4_out[452]);
     layer5_out[587] <= layer4_out[48];
     layer5_out[588] <= layer4_out[877];
     layer5_out[589] <= layer4_out[1158];
     layer5_out[590] <= ~layer4_out[375];
     layer5_out[591] <= ~(layer4_out[1118] & layer4_out[1119]);
     layer5_out[592] <= layer4_out[742] ^ layer4_out[743];
     layer5_out[593] <= ~layer4_out[700];
     layer5_out[594] <= ~layer4_out[895] | layer4_out[896];
     layer5_out[595] <= layer4_out[826];
     layer5_out[596] <= ~(layer4_out[1424] ^ layer4_out[1425]);
     layer5_out[597] <= layer4_out[22];
     layer5_out[598] <= layer4_out[949];
     layer5_out[599] <= ~layer4_out[475];
     layer5_out[600] <= ~(layer4_out[1216] ^ layer4_out[1217]);
     layer5_out[601] <= ~(layer4_out[357] ^ layer4_out[358]);
     layer5_out[602] <= ~(layer4_out[908] | layer4_out[909]);
     layer5_out[603] <= ~layer4_out[844];
     layer5_out[604] <= layer4_out[547];
     layer5_out[605] <= ~layer4_out[413] | layer4_out[412];
     layer5_out[606] <= ~(layer4_out[275] | layer4_out[276]);
     layer5_out[607] <= ~layer4_out[51];
     layer5_out[608] <= layer4_out[505];
     layer5_out[609] <= ~layer4_out[1005];
     layer5_out[610] <= ~layer4_out[267] | layer4_out[268];
     layer5_out[611] <= ~layer4_out[1247];
     layer5_out[612] <= layer4_out[766] & layer4_out[767];
     layer5_out[613] <= ~layer4_out[787] | layer4_out[788];
     layer5_out[614] <= ~layer4_out[850];
     layer5_out[615] <= layer4_out[537];
     layer5_out[616] <= ~(layer4_out[897] | layer4_out[898]);
     layer5_out[617] <= ~layer4_out[797];
     layer5_out[618] <= ~(layer4_out[254] | layer4_out[255]);
     layer5_out[619] <= layer4_out[849];
     layer5_out[620] <= layer4_out[531] & ~layer4_out[532];
     layer5_out[621] <= ~layer4_out[794];
     layer5_out[622] <= ~(layer4_out[1409] & layer4_out[1410]);
     layer5_out[623] <= layer4_out[664];
     layer5_out[624] <= ~(layer4_out[154] & layer4_out[155]);
     layer5_out[625] <= layer4_out[339];
     layer5_out[626] <= ~layer4_out[1067];
     layer5_out[627] <= layer4_out[896] ^ layer4_out[897];
     layer5_out[628] <= layer4_out[929] & ~layer4_out[930];
     layer5_out[629] <= ~layer4_out[846] | layer4_out[847];
     layer5_out[630] <= layer4_out[1100] & ~layer4_out[1101];
     layer5_out[631] <= layer4_out[700] & ~layer4_out[701];
     layer5_out[632] <= ~layer4_out[471];
     layer5_out[633] <= ~(layer4_out[692] | layer4_out[693]);
     layer5_out[634] <= ~layer4_out[394] | layer4_out[393];
     layer5_out[635] <= ~layer4_out[1331];
     layer5_out[636] <= layer4_out[1085] | layer4_out[1086];
     layer5_out[637] <= ~layer4_out[648];
     layer5_out[638] <= ~layer4_out[55];
     layer5_out[639] <= ~(layer4_out[987] | layer4_out[988]);
     layer5_out[640] <= ~(layer4_out[869] ^ layer4_out[870]);
     layer5_out[641] <= layer4_out[480];
     layer5_out[642] <= ~layer4_out[644] | layer4_out[643];
     layer5_out[643] <= layer4_out[54] & layer4_out[55];
     layer5_out[644] <= layer4_out[18];
     layer5_out[645] <= layer4_out[555] & ~layer4_out[554];
     layer5_out[646] <= layer4_out[391];
     layer5_out[647] <= ~layer4_out[403];
     layer5_out[648] <= 1'b0;
     layer5_out[649] <= ~layer4_out[232];
     layer5_out[650] <= ~layer4_out[40];
     layer5_out[651] <= ~(layer4_out[720] | layer4_out[721]);
     layer5_out[652] <= layer4_out[1477] & ~layer4_out[1478];
     layer5_out[653] <= layer4_out[681] & ~layer4_out[680];
     layer5_out[654] <= layer4_out[709];
     layer5_out[655] <= ~layer4_out[163];
     layer5_out[656] <= ~layer4_out[989];
     layer5_out[657] <= layer4_out[586];
     layer5_out[658] <= layer4_out[1458] & layer4_out[1459];
     layer5_out[659] <= ~layer4_out[1256];
     layer5_out[660] <= layer4_out[185] | layer4_out[186];
     layer5_out[661] <= layer4_out[871] & layer4_out[872];
     layer5_out[662] <= layer4_out[133];
     layer5_out[663] <= layer4_out[1372];
     layer5_out[664] <= layer4_out[367] & layer4_out[368];
     layer5_out[665] <= layer4_out[740];
     layer5_out[666] <= ~layer4_out[1397];
     layer5_out[667] <= ~layer4_out[1190] | layer4_out[1189];
     layer5_out[668] <= layer4_out[1422] & ~layer4_out[1423];
     layer5_out[669] <= layer4_out[182] & layer4_out[183];
     layer5_out[670] <= layer4_out[549];
     layer5_out[671] <= ~layer4_out[815];
     layer5_out[672] <= layer4_out[1027] | layer4_out[1028];
     layer5_out[673] <= layer4_out[582];
     layer5_out[674] <= ~layer4_out[109];
     layer5_out[675] <= layer4_out[689];
     layer5_out[676] <= ~(layer4_out[572] ^ layer4_out[573]);
     layer5_out[677] <= ~layer4_out[629];
     layer5_out[678] <= ~layer4_out[1414];
     layer5_out[679] <= ~layer4_out[1124] | layer4_out[1123];
     layer5_out[680] <= ~(layer4_out[795] ^ layer4_out[796]);
     layer5_out[681] <= ~(layer4_out[118] & layer4_out[119]);
     layer5_out[682] <= layer4_out[1222];
     layer5_out[683] <= layer4_out[753];
     layer5_out[684] <= ~layer4_out[401];
     layer5_out[685] <= ~layer4_out[341];
     layer5_out[686] <= layer4_out[148];
     layer5_out[687] <= layer4_out[1009] & ~layer4_out[1010];
     layer5_out[688] <= ~layer4_out[434];
     layer5_out[689] <= layer4_out[565] ^ layer4_out[566];
     layer5_out[690] <= ~layer4_out[855];
     layer5_out[691] <= ~(layer4_out[76] | layer4_out[77]);
     layer5_out[692] <= layer4_out[915];
     layer5_out[693] <= layer4_out[672] & ~layer4_out[673];
     layer5_out[694] <= ~layer4_out[294] | layer4_out[295];
     layer5_out[695] <= layer4_out[875];
     layer5_out[696] <= ~layer4_out[348];
     layer5_out[697] <= layer4_out[326] & ~layer4_out[325];
     layer5_out[698] <= 1'b0;
     layer5_out[699] <= ~layer4_out[1113] | layer4_out[1114];
     layer5_out[700] <= ~layer4_out[1045];
     layer5_out[701] <= ~layer4_out[1340];
     layer5_out[702] <= layer4_out[821];
     layer5_out[703] <= ~layer4_out[340];
     layer5_out[704] <= layer4_out[1281] ^ layer4_out[1282];
     layer5_out[705] <= ~layer4_out[1019];
     layer5_out[706] <= ~layer4_out[1029] | layer4_out[1028];
     layer5_out[707] <= 1'b1;
     layer5_out[708] <= ~layer4_out[1238] | layer4_out[1239];
     layer5_out[709] <= layer4_out[1011];
     layer5_out[710] <= ~(layer4_out[1432] & layer4_out[1433]);
     layer5_out[711] <= ~layer4_out[614];
     layer5_out[712] <= layer4_out[1081];
     layer5_out[713] <= layer4_out[724] ^ layer4_out[725];
     layer5_out[714] <= ~layer4_out[12];
     layer5_out[715] <= layer4_out[1395];
     layer5_out[716] <= ~layer4_out[1478];
     layer5_out[717] <= ~(layer4_out[973] ^ layer4_out[974]);
     layer5_out[718] <= ~layer4_out[538] | layer4_out[539];
     layer5_out[719] <= layer4_out[867] | layer4_out[868];
     layer5_out[720] <= ~layer4_out[1123] | layer4_out[1122];
     layer5_out[721] <= ~layer4_out[1466];
     layer5_out[722] <= layer4_out[1212];
     layer5_out[723] <= layer4_out[373];
     layer5_out[724] <= ~(layer4_out[919] | layer4_out[920]);
     layer5_out[725] <= 1'b0;
     layer5_out[726] <= ~layer4_out[1148];
     layer5_out[727] <= layer4_out[798] | layer4_out[799];
     layer5_out[728] <= ~layer4_out[353];
     layer5_out[729] <= ~layer4_out[197];
     layer5_out[730] <= ~layer4_out[1337];
     layer5_out[731] <= ~(layer4_out[1220] & layer4_out[1221]);
     layer5_out[732] <= 1'b1;
     layer5_out[733] <= ~layer4_out[143] | layer4_out[142];
     layer5_out[734] <= ~(layer4_out[386] & layer4_out[387]);
     layer5_out[735] <= layer4_out[146];
     layer5_out[736] <= layer4_out[660] & layer4_out[661];
     layer5_out[737] <= 1'b1;
     layer5_out[738] <= ~layer4_out[1139];
     layer5_out[739] <= ~(layer4_out[1366] & layer4_out[1367]);
     layer5_out[740] <= layer4_out[1175] | layer4_out[1176];
     layer5_out[741] <= layer4_out[1207];
     layer5_out[742] <= layer4_out[415];
     layer5_out[743] <= ~layer4_out[529];
     layer5_out[744] <= layer4_out[431] | layer4_out[432];
     layer5_out[745] <= layer4_out[1202] | layer4_out[1203];
     layer5_out[746] <= ~(layer4_out[48] | layer4_out[49]);
     layer5_out[747] <= ~(layer4_out[882] ^ layer4_out[883]);
     layer5_out[748] <= ~(layer4_out[514] & layer4_out[515]);
     layer5_out[749] <= layer4_out[853];
     layer5_out[750] <= ~layer4_out[921] | layer4_out[922];
     layer5_out[751] <= ~layer4_out[496];
     layer5_out[752] <= layer4_out[775];
     layer5_out[753] <= layer4_out[761] & ~layer4_out[760];
     layer5_out[754] <= ~layer4_out[1479] | layer4_out[1480];
     layer5_out[755] <= ~layer4_out[1305];
     layer5_out[756] <= ~layer4_out[787];
     layer5_out[757] <= ~layer4_out[1354] | layer4_out[1353];
     layer5_out[758] <= 1'b0;
     layer5_out[759] <= ~layer4_out[832];
     layer5_out[760] <= layer4_out[196] & layer4_out[197];
     layer5_out[761] <= ~(layer4_out[819] | layer4_out[820]);
     layer5_out[762] <= ~layer4_out[1116];
     layer5_out[763] <= layer4_out[1049] & ~layer4_out[1048];
     layer5_out[764] <= layer4_out[153];
     layer5_out[765] <= ~layer4_out[984];
     layer5_out[766] <= ~(layer4_out[1399] | layer4_out[1400]);
     layer5_out[767] <= ~layer4_out[192];
     layer5_out[768] <= ~layer4_out[591];
     layer5_out[769] <= layer4_out[924];
     layer5_out[770] <= ~(layer4_out[1437] & layer4_out[1438]);
     layer5_out[771] <= layer4_out[886];
     layer5_out[772] <= ~layer4_out[991];
     layer5_out[773] <= layer4_out[558] ^ layer4_out[559];
     layer5_out[774] <= layer4_out[1447];
     layer5_out[775] <= layer4_out[426] & ~layer4_out[425];
     layer5_out[776] <= 1'b0;
     layer5_out[777] <= ~layer4_out[322];
     layer5_out[778] <= ~layer4_out[655] | layer4_out[654];
     layer5_out[779] <= layer4_out[64] & layer4_out[65];
     layer5_out[780] <= layer4_out[127];
     layer5_out[781] <= layer4_out[826] & layer4_out[827];
     layer5_out[782] <= ~layer4_out[82] | layer4_out[81];
     layer5_out[783] <= layer4_out[1323] & ~layer4_out[1324];
     layer5_out[784] <= ~layer4_out[464] | layer4_out[463];
     layer5_out[785] <= layer4_out[633] & ~layer4_out[634];
     layer5_out[786] <= ~layer4_out[1107];
     layer5_out[787] <= layer4_out[589] & ~layer4_out[590];
     layer5_out[788] <= ~(layer4_out[391] | layer4_out[392]);
     layer5_out[789] <= layer4_out[840];
     layer5_out[790] <= ~layer4_out[1220] | layer4_out[1219];
     layer5_out[791] <= ~layer4_out[316];
     layer5_out[792] <= ~layer4_out[366];
     layer5_out[793] <= layer4_out[934];
     layer5_out[794] <= layer4_out[1347] & ~layer4_out[1348];
     layer5_out[795] <= layer4_out[1377] ^ layer4_out[1378];
     layer5_out[796] <= layer4_out[585];
     layer5_out[797] <= ~layer4_out[789] | layer4_out[788];
     layer5_out[798] <= layer4_out[641];
     layer5_out[799] <= layer4_out[1242] & layer4_out[1243];
     layer5_out[800] <= layer4_out[937] & ~layer4_out[936];
     layer5_out[801] <= ~(layer4_out[26] | layer4_out[27]);
     layer5_out[802] <= ~(layer4_out[83] ^ layer4_out[84]);
     layer5_out[803] <= 1'b0;
     layer5_out[804] <= ~layer4_out[381] | layer4_out[380];
     layer5_out[805] <= ~layer4_out[1249];
     layer5_out[806] <= layer4_out[815];
     layer5_out[807] <= ~(layer4_out[203] | layer4_out[204]);
     layer5_out[808] <= layer4_out[1438] & ~layer4_out[1439];
     layer5_out[809] <= ~layer4_out[106] | layer4_out[105];
     layer5_out[810] <= ~(layer4_out[862] & layer4_out[863]);
     layer5_out[811] <= ~layer4_out[1407];
     layer5_out[812] <= ~layer4_out[1441] | layer4_out[1442];
     layer5_out[813] <= layer4_out[234];
     layer5_out[814] <= layer4_out[272] & ~layer4_out[271];
     layer5_out[815] <= ~layer4_out[1058] | layer4_out[1057];
     layer5_out[816] <= layer4_out[6];
     layer5_out[817] <= layer4_out[594] & ~layer4_out[595];
     layer5_out[818] <= layer4_out[930] & layer4_out[931];
     layer5_out[819] <= ~(layer4_out[199] | layer4_out[200]);
     layer5_out[820] <= ~layer4_out[1295];
     layer5_out[821] <= layer4_out[1145] & layer4_out[1146];
     layer5_out[822] <= layer4_out[687];
     layer5_out[823] <= layer4_out[1411] & layer4_out[1412];
     layer5_out[824] <= ~(layer4_out[568] | layer4_out[569]);
     layer5_out[825] <= layer4_out[518];
     layer5_out[826] <= ~layer4_out[907];
     layer5_out[827] <= ~(layer4_out[1333] ^ layer4_out[1334]);
     layer5_out[828] <= ~layer4_out[663];
     layer5_out[829] <= ~(layer4_out[306] ^ layer4_out[307]);
     layer5_out[830] <= layer4_out[845] & ~layer4_out[844];
     layer5_out[831] <= ~(layer4_out[1261] | layer4_out[1262]);
     layer5_out[832] <= layer4_out[403] ^ layer4_out[404];
     layer5_out[833] <= ~layer4_out[1138];
     layer5_out[834] <= layer4_out[1498];
     layer5_out[835] <= ~layer4_out[1461];
     layer5_out[836] <= ~layer4_out[1298] | layer4_out[1299];
     layer5_out[837] <= ~layer4_out[374];
     layer5_out[838] <= layer4_out[1453] & ~layer4_out[1452];
     layer5_out[839] <= layer4_out[1387] & layer4_out[1388];
     layer5_out[840] <= ~(layer4_out[893] | layer4_out[894]);
     layer5_out[841] <= layer4_out[603] & ~layer4_out[602];
     layer5_out[842] <= layer4_out[117];
     layer5_out[843] <= layer4_out[14] & layer4_out[15];
     layer5_out[844] <= ~(layer4_out[1487] | layer4_out[1488]);
     layer5_out[845] <= layer4_out[1011];
     layer5_out[846] <= ~(layer4_out[1320] | layer4_out[1321]);
     layer5_out[847] <= layer4_out[1061] & ~layer4_out[1062];
     layer5_out[848] <= layer4_out[1459];
     layer5_out[849] <= ~layer4_out[1069];
     layer5_out[850] <= layer4_out[420];
     layer5_out[851] <= ~layer4_out[327];
     layer5_out[852] <= ~layer4_out[84] | layer4_out[85];
     layer5_out[853] <= ~layer4_out[195];
     layer5_out[854] <= ~layer4_out[80];
     layer5_out[855] <= layer4_out[1301];
     layer5_out[856] <= layer4_out[607];
     layer5_out[857] <= ~layer4_out[1095];
     layer5_out[858] <= ~layer4_out[1183];
     layer5_out[859] <= layer4_out[287];
     layer5_out[860] <= layer4_out[1495];
     layer5_out[861] <= layer4_out[457];
     layer5_out[862] <= ~(layer4_out[809] ^ layer4_out[810]);
     layer5_out[863] <= layer4_out[314] ^ layer4_out[315];
     layer5_out[864] <= ~layer4_out[99] | layer4_out[100];
     layer5_out[865] <= layer4_out[1442] ^ layer4_out[1443];
     layer5_out[866] <= layer4_out[14];
     layer5_out[867] <= layer4_out[122] | layer4_out[123];
     layer5_out[868] <= ~layer4_out[510] | layer4_out[509];
     layer5_out[869] <= ~(layer4_out[1352] | layer4_out[1353]);
     layer5_out[870] <= layer4_out[335] & ~layer4_out[334];
     layer5_out[871] <= layer4_out[140] & layer4_out[141];
     layer5_out[872] <= ~(layer4_out[7] ^ layer4_out[8]);
     layer5_out[873] <= layer4_out[328] & layer4_out[329];
     layer5_out[874] <= layer4_out[298];
     layer5_out[875] <= layer4_out[950] & ~layer4_out[951];
     layer5_out[876] <= ~layer4_out[905] | layer4_out[906];
     layer5_out[877] <= layer4_out[756] & ~layer4_out[757];
     layer5_out[878] <= ~layer4_out[1303] | layer4_out[1302];
     layer5_out[879] <= ~layer4_out[766];
     layer5_out[880] <= layer4_out[8];
     layer5_out[881] <= layer4_out[210];
     layer5_out[882] <= layer4_out[979];
     layer5_out[883] <= ~layer4_out[674];
     layer5_out[884] <= layer4_out[668];
     layer5_out[885] <= layer4_out[1253] ^ layer4_out[1254];
     layer5_out[886] <= ~(layer4_out[1190] | layer4_out[1191]);
     layer5_out[887] <= 1'b1;
     layer5_out[888] <= ~layer4_out[960];
     layer5_out[889] <= ~(layer4_out[730] | layer4_out[731]);
     layer5_out[890] <= ~(layer4_out[133] & layer4_out[134]);
     layer5_out[891] <= ~layer4_out[585];
     layer5_out[892] <= layer4_out[1343];
     layer5_out[893] <= ~(layer4_out[383] & layer4_out[384]);
     layer5_out[894] <= ~(layer4_out[1417] | layer4_out[1418]);
     layer5_out[895] <= layer4_out[928];
     layer5_out[896] <= ~(layer4_out[139] & layer4_out[140]);
     layer5_out[897] <= layer4_out[1405];
     layer5_out[898] <= ~layer4_out[1224] | layer4_out[1225];
     layer5_out[899] <= ~layer4_out[65];
     layer5_out[900] <= layer4_out[75];
     layer5_out[901] <= layer4_out[418];
     layer5_out[902] <= layer4_out[443];
     layer5_out[903] <= layer4_out[223];
     layer5_out[904] <= ~(layer4_out[307] & layer4_out[308]);
     layer5_out[905] <= ~layer4_out[396] | layer4_out[397];
     layer5_out[906] <= layer4_out[376];
     layer5_out[907] <= ~(layer4_out[1078] & layer4_out[1079]);
     layer5_out[908] <= layer4_out[1194];
     layer5_out[909] <= layer4_out[1357] ^ layer4_out[1358];
     layer5_out[910] <= ~layer4_out[939];
     layer5_out[911] <= layer4_out[1318] & layer4_out[1319];
     layer5_out[912] <= ~(layer4_out[333] | layer4_out[334]);
     layer5_out[913] <= layer4_out[498];
     layer5_out[914] <= ~layer4_out[792];
     layer5_out[915] <= ~(layer4_out[912] | layer4_out[913]);
     layer5_out[916] <= ~layer4_out[411];
     layer5_out[917] <= ~layer4_out[1363] | layer4_out[1364];
     layer5_out[918] <= layer4_out[436];
     layer5_out[919] <= ~layer4_out[725];
     layer5_out[920] <= layer4_out[30];
     layer5_out[921] <= layer4_out[221] ^ layer4_out[222];
     layer5_out[922] <= ~layer4_out[1167];
     layer5_out[923] <= ~layer4_out[639];
     layer5_out[924] <= layer4_out[103] & ~layer4_out[102];
     layer5_out[925] <= ~layer4_out[1192];
     layer5_out[926] <= ~layer4_out[1390];
     layer5_out[927] <= ~layer4_out[280];
     layer5_out[928] <= ~layer4_out[829];
     layer5_out[929] <= ~(layer4_out[1473] & layer4_out[1474]);
     layer5_out[930] <= layer4_out[1373];
     layer5_out[931] <= layer4_out[212];
     layer5_out[932] <= layer4_out[1001];
     layer5_out[933] <= ~layer4_out[812];
     layer5_out[934] <= layer4_out[773];
     layer5_out[935] <= layer4_out[1270] | layer4_out[1271];
     layer5_out[936] <= layer4_out[1293];
     layer5_out[937] <= ~layer4_out[1467];
     layer5_out[938] <= ~layer4_out[1470];
     layer5_out[939] <= ~(layer4_out[559] ^ layer4_out[560]);
     layer5_out[940] <= ~layer4_out[248] | layer4_out[249];
     layer5_out[941] <= ~layer4_out[611];
     layer5_out[942] <= ~(layer4_out[1097] | layer4_out[1098]);
     layer5_out[943] <= ~layer4_out[388] | layer4_out[389];
     layer5_out[944] <= ~layer4_out[1455];
     layer5_out[945] <= layer4_out[384] & layer4_out[385];
     layer5_out[946] <= ~layer4_out[982];
     layer5_out[947] <= ~layer4_out[1261] | layer4_out[1260];
     layer5_out[948] <= ~layer4_out[808];
     layer5_out[949] <= ~layer4_out[711] | layer4_out[712];
     layer5_out[950] <= ~layer4_out[832];
     layer5_out[951] <= layer4_out[940];
     layer5_out[952] <= layer4_out[669] | layer4_out[670];
     layer5_out[953] <= layer4_out[1244] & layer4_out[1245];
     layer5_out[954] <= ~layer4_out[562];
     layer5_out[955] <= ~layer4_out[922];
     layer5_out[956] <= layer4_out[1003];
     layer5_out[957] <= ~(layer4_out[160] | layer4_out[161]);
     layer5_out[958] <= layer4_out[1496] & ~layer4_out[1497];
     layer5_out[959] <= ~(layer4_out[43] ^ layer4_out[44]);
     layer5_out[960] <= layer4_out[318];
     layer5_out[961] <= layer4_out[1349] & ~layer4_out[1348];
     layer5_out[962] <= ~(layer4_out[1198] | layer4_out[1199]);
     layer5_out[963] <= layer4_out[124] | layer4_out[125];
     layer5_out[964] <= layer4_out[1060];
     layer5_out[965] <= ~layer4_out[1122];
     layer5_out[966] <= ~layer4_out[722] | layer4_out[721];
     layer5_out[967] <= layer4_out[534];
     layer5_out[968] <= layer4_out[1287];
     layer5_out[969] <= layer4_out[1224];
     layer5_out[970] <= ~layer4_out[843];
     layer5_out[971] <= ~layer4_out[683] | layer4_out[684];
     layer5_out[972] <= ~layer4_out[1271];
     layer5_out[973] <= layer4_out[351];
     layer5_out[974] <= ~(layer4_out[362] & layer4_out[363]);
     layer5_out[975] <= ~layer4_out[633] | layer4_out[632];
     layer5_out[976] <= layer4_out[136];
     layer5_out[977] <= layer4_out[968] & ~layer4_out[969];
     layer5_out[978] <= layer4_out[532];
     layer5_out[979] <= ~(layer4_out[44] | layer4_out[45]);
     layer5_out[980] <= ~layer4_out[291];
     layer5_out[981] <= layer4_out[845] ^ layer4_out[846];
     layer5_out[982] <= 1'b1;
     layer5_out[983] <= ~layer4_out[806];
     layer5_out[984] <= ~layer4_out[88] | layer4_out[89];
     layer5_out[985] <= layer4_out[680];
     layer5_out[986] <= layer4_out[847] & layer4_out[848];
     layer5_out[987] <= layer4_out[501];
     layer5_out[988] <= layer4_out[780] | layer4_out[781];
     layer5_out[989] <= ~layer4_out[237];
     layer5_out[990] <= layer4_out[1313] & ~layer4_out[1312];
     layer5_out[991] <= layer4_out[1402] & ~layer4_out[1401];
     layer5_out[992] <= ~layer4_out[514];
     layer5_out[993] <= layer4_out[1218];
     layer5_out[994] <= layer4_out[337];
     layer5_out[995] <= layer4_out[903];
     layer5_out[996] <= layer4_out[763];
     layer5_out[997] <= ~layer4_out[321];
     layer5_out[998] <= ~layer4_out[1264] | layer4_out[1263];
     layer5_out[999] <= layer4_out[819] & ~layer4_out[818];
     layer5_out[1000] <= layer4_out[287] ^ layer4_out[288];
     layer5_out[1001] <= ~(layer4_out[626] ^ layer4_out[627]);
     layer5_out[1002] <= layer4_out[763] ^ layer4_out[764];
     layer5_out[1003] <= ~layer4_out[657] | layer4_out[658];
     layer5_out[1004] <= ~layer4_out[1091] | layer4_out[1090];
     layer5_out[1005] <= layer4_out[1179] & ~layer4_out[1178];
     layer5_out[1006] <= layer4_out[110];
     layer5_out[1007] <= ~layer4_out[301];
     layer5_out[1008] <= ~layer4_out[1026];
     layer5_out[1009] <= ~layer4_out[1352] | layer4_out[1351];
     layer5_out[1010] <= ~(layer4_out[66] & layer4_out[67]);
     layer5_out[1011] <= ~(layer4_out[1153] & layer4_out[1154]);
     layer5_out[1012] <= ~(layer4_out[1376] & layer4_out[1377]);
     layer5_out[1013] <= layer4_out[1359] & ~layer4_out[1358];
     layer5_out[1014] <= ~layer4_out[653];
     layer5_out[1015] <= ~layer4_out[1428];
     layer5_out[1016] <= layer4_out[184] & ~layer4_out[183];
     layer5_out[1017] <= layer4_out[946] & ~layer4_out[945];
     layer5_out[1018] <= layer4_out[226];
     layer5_out[1019] <= ~(layer4_out[34] ^ layer4_out[35]);
     layer5_out[1020] <= layer4_out[736] & ~layer4_out[735];
     layer5_out[1021] <= ~layer4_out[296];
     layer5_out[1022] <= layer4_out[1152];
     layer5_out[1023] <= ~layer4_out[198];
     layer5_out[1024] <= layer4_out[979];
     layer5_out[1025] <= ~layer4_out[1041];
     layer5_out[1026] <= ~layer4_out[292];
     layer5_out[1027] <= layer4_out[1300] | layer4_out[1301];
     layer5_out[1028] <= layer4_out[916] ^ layer4_out[917];
     layer5_out[1029] <= ~layer4_out[93];
     layer5_out[1030] <= layer4_out[95] & ~layer4_out[94];
     layer5_out[1031] <= layer4_out[605] & ~layer4_out[606];
     layer5_out[1032] <= ~layer4_out[576];
     layer5_out[1033] <= layer4_out[611];
     layer5_out[1034] <= ~(layer4_out[1340] | layer4_out[1341]);
     layer5_out[1035] <= layer4_out[755] & layer4_out[756];
     layer5_out[1036] <= ~layer4_out[278];
     layer5_out[1037] <= layer4_out[704] ^ layer4_out[705];
     layer5_out[1038] <= ~(layer4_out[732] | layer4_out[733]);
     layer5_out[1039] <= ~layer4_out[190] | layer4_out[191];
     layer5_out[1040] <= ~layer4_out[782];
     layer5_out[1041] <= layer4_out[865] | layer4_out[866];
     layer5_out[1042] <= ~(layer4_out[1439] | layer4_out[1440]);
     layer5_out[1043] <= layer4_out[842];
     layer5_out[1044] <= ~layer4_out[1297];
     layer5_out[1045] <= ~layer4_out[1132];
     layer5_out[1046] <= layer4_out[1138];
     layer5_out[1047] <= layer4_out[679];
     layer5_out[1048] <= layer4_out[332] | layer4_out[333];
     layer5_out[1049] <= ~layer4_out[1276];
     layer5_out[1050] <= layer4_out[365];
     layer5_out[1051] <= ~layer4_out[1376] | layer4_out[1375];
     layer5_out[1052] <= ~layer4_out[806] | layer4_out[807];
     layer5_out[1053] <= ~(layer4_out[898] | layer4_out[899]);
     layer5_out[1054] <= ~layer4_out[1265];
     layer5_out[1055] <= layer4_out[1045];
     layer5_out[1056] <= ~(layer4_out[90] | layer4_out[91]);
     layer5_out[1057] <= ~layer4_out[1269];
     layer5_out[1058] <= layer4_out[1072] ^ layer4_out[1073];
     layer5_out[1059] <= layer4_out[168];
     layer5_out[1060] <= layer4_out[129];
     layer5_out[1061] <= ~layer4_out[736] | layer4_out[737];
     layer5_out[1062] <= layer4_out[868] & ~layer4_out[869];
     layer5_out[1063] <= ~layer4_out[1018];
     layer5_out[1064] <= layer4_out[1246];
     layer5_out[1065] <= layer4_out[1128];
     layer5_out[1066] <= ~layer4_out[263];
     layer5_out[1067] <= ~(layer4_out[1039] & layer4_out[1040]);
     layer5_out[1068] <= ~layer4_out[578];
     layer5_out[1069] <= layer4_out[1474] | layer4_out[1475];
     layer5_out[1070] <= ~(layer4_out[625] & layer4_out[626]);
     layer5_out[1071] <= ~layer4_out[617];
     layer5_out[1072] <= layer4_out[1234] & ~layer4_out[1233];
     layer5_out[1073] <= layer4_out[302];
     layer5_out[1074] <= ~(layer4_out[1136] | layer4_out[1137]);
     layer5_out[1075] <= layer4_out[243];
     layer5_out[1076] <= ~layer4_out[58] | layer4_out[57];
     layer5_out[1077] <= layer4_out[1101] & ~layer4_out[1102];
     layer5_out[1078] <= layer4_out[548] & layer4_out[549];
     layer5_out[1079] <= layer4_out[604];
     layer5_out[1080] <= ~(layer4_out[1443] ^ layer4_out[1444]);
     layer5_out[1081] <= ~(layer4_out[490] & layer4_out[491]);
     layer5_out[1082] <= layer4_out[625];
     layer5_out[1083] <= layer4_out[650];
     layer5_out[1084] <= layer4_out[108] | layer4_out[109];
     layer5_out[1085] <= 1'b1;
     layer5_out[1086] <= ~layer4_out[1108] | layer4_out[1109];
     layer5_out[1087] <= ~(layer4_out[440] ^ layer4_out[441]);
     layer5_out[1088] <= ~(layer4_out[157] | layer4_out[158]);
     layer5_out[1089] <= layer4_out[1299] & ~layer4_out[1300];
     layer5_out[1090] <= layer4_out[715] & ~layer4_out[716];
     layer5_out[1091] <= layer4_out[581];
     layer5_out[1092] <= ~layer4_out[489];
     layer5_out[1093] <= layer4_out[1486] & layer4_out[1487];
     layer5_out[1094] <= ~layer4_out[59];
     layer5_out[1095] <= layer4_out[92] & layer4_out[93];
     layer5_out[1096] <= ~(layer4_out[244] | layer4_out[245]);
     layer5_out[1097] <= layer4_out[1445];
     layer5_out[1098] <= layer4_out[1016] & ~layer4_out[1017];
     layer5_out[1099] <= layer4_out[1242];
     layer5_out[1100] <= layer4_out[1021] & ~layer4_out[1022];
     layer5_out[1101] <= ~(layer4_out[394] ^ layer4_out[395]);
     layer5_out[1102] <= layer4_out[203];
     layer5_out[1103] <= layer4_out[717];
     layer5_out[1104] <= layer4_out[997] & layer4_out[998];
     layer5_out[1105] <= layer4_out[1437] & ~layer4_out[1436];
     layer5_out[1106] <= ~(layer4_out[449] | layer4_out[450]);
     layer5_out[1107] <= ~layer4_out[1448];
     layer5_out[1108] <= layer4_out[546] & ~layer4_out[547];
     layer5_out[1109] <= ~layer4_out[684] | layer4_out[685];
     layer5_out[1110] <= layer4_out[2] & ~layer4_out[0];
     layer5_out[1111] <= layer4_out[1080];
     layer5_out[1112] <= ~(layer4_out[553] ^ layer4_out[554]);
     layer5_out[1113] <= layer4_out[975];
     layer5_out[1114] <= ~layer4_out[16];
     layer5_out[1115] <= layer4_out[1342] ^ layer4_out[1343];
     layer5_out[1116] <= layer4_out[101] | layer4_out[102];
     layer5_out[1117] <= layer4_out[779] | layer4_out[780];
     layer5_out[1118] <= layer4_out[1078] & ~layer4_out[1077];
     layer5_out[1119] <= ~(layer4_out[848] | layer4_out[849]);
     layer5_out[1120] <= layer4_out[270] | layer4_out[271];
     layer5_out[1121] <= layer4_out[268];
     layer5_out[1122] <= layer4_out[695] | layer4_out[696];
     layer5_out[1123] <= ~layer4_out[215];
     layer5_out[1124] <= ~layer4_out[149] | layer4_out[150];
     layer5_out[1125] <= layer4_out[1147];
     layer5_out[1126] <= layer4_out[1213];
     layer5_out[1127] <= ~layer4_out[690];
     layer5_out[1128] <= layer4_out[560] & layer4_out[561];
     layer5_out[1129] <= layer4_out[957];
     layer5_out[1130] <= layer4_out[176] | layer4_out[177];
     layer5_out[1131] <= ~(layer4_out[1243] ^ layer4_out[1244]);
     layer5_out[1132] <= layer4_out[1209];
     layer5_out[1133] <= ~layer4_out[220] | layer4_out[219];
     layer5_out[1134] <= ~layer4_out[53] | layer4_out[52];
     layer5_out[1135] <= ~layer4_out[477];
     layer5_out[1136] <= layer4_out[343] & layer4_out[344];
     layer5_out[1137] <= ~layer4_out[1228];
     layer5_out[1138] <= layer4_out[260] & ~layer4_out[259];
     layer5_out[1139] <= layer4_out[1450];
     layer5_out[1140] <= ~(layer4_out[665] ^ layer4_out[666]);
     layer5_out[1141] <= layer4_out[726] | layer4_out[727];
     layer5_out[1142] <= layer4_out[1249];
     layer5_out[1143] <= layer4_out[1201] & ~layer4_out[1200];
     layer5_out[1144] <= ~layer4_out[958];
     layer5_out[1145] <= ~(layer4_out[690] | layer4_out[691]);
     layer5_out[1146] <= layer4_out[596] & ~layer4_out[595];
     layer5_out[1147] <= ~layer4_out[1035] | layer4_out[1036];
     layer5_out[1148] <= ~(layer4_out[106] ^ layer4_out[107]);
     layer5_out[1149] <= ~layer4_out[1039];
     layer5_out[1150] <= ~(layer4_out[1257] | layer4_out[1258]);
     layer5_out[1151] <= layer4_out[965] & ~layer4_out[966];
     layer5_out[1152] <= ~(layer4_out[1070] ^ layer4_out[1071]);
     layer5_out[1153] <= ~layer4_out[622];
     layer5_out[1154] <= ~layer4_out[170];
     layer5_out[1155] <= layer4_out[355];
     layer5_out[1156] <= ~layer4_out[944];
     layer5_out[1157] <= ~layer4_out[223];
     layer5_out[1158] <= ~layer4_out[1394];
     layer5_out[1159] <= ~layer4_out[10];
     layer5_out[1160] <= layer4_out[574] ^ layer4_out[575];
     layer5_out[1161] <= layer4_out[541] | layer4_out[542];
     layer5_out[1162] <= layer4_out[1172];
     layer5_out[1163] <= ~(layer4_out[646] ^ layer4_out[647]);
     layer5_out[1164] <= ~(layer4_out[1466] ^ layer4_out[1467]);
     layer5_out[1165] <= ~(layer4_out[1341] & layer4_out[1342]);
     layer5_out[1166] <= ~(layer4_out[671] & layer4_out[672]);
     layer5_out[1167] <= 1'b1;
     layer5_out[1168] <= ~layer4_out[1175] | layer4_out[1174];
     layer5_out[1169] <= ~layer4_out[1091];
     layer5_out[1170] <= ~layer4_out[856];
     layer5_out[1171] <= layer4_out[901] & layer4_out[902];
     layer5_out[1172] <= ~layer4_out[1156];
     layer5_out[1173] <= ~layer4_out[1093];
     layer5_out[1174] <= layer4_out[752] ^ layer4_out[753];
     layer5_out[1175] <= layer4_out[1105] & layer4_out[1106];
     layer5_out[1176] <= ~layer4_out[1361] | layer4_out[1362];
     layer5_out[1177] <= layer4_out[98];
     layer5_out[1178] <= ~(layer4_out[116] ^ layer4_out[117]);
     layer5_out[1179] <= ~layer4_out[207] | layer4_out[206];
     layer5_out[1180] <= ~layer4_out[873];
     layer5_out[1181] <= ~layer4_out[498];
     layer5_out[1182] <= layer4_out[1365] | layer4_out[1366];
     layer5_out[1183] <= ~layer4_out[40];
     layer5_out[1184] <= layer4_out[360] & ~layer4_out[361];
     layer5_out[1185] <= layer4_out[468] | layer4_out[469];
     layer5_out[1186] <= layer4_out[1096];
     layer5_out[1187] <= ~layer4_out[208] | layer4_out[207];
     layer5_out[1188] <= ~(layer4_out[260] & layer4_out[261]);
     layer5_out[1189] <= ~layer4_out[115];
     layer5_out[1190] <= ~layer4_out[1211];
     layer5_out[1191] <= ~(layer4_out[1221] | layer4_out[1222]);
     layer5_out[1192] <= layer4_out[938];
     layer5_out[1193] <= layer4_out[805] & ~layer4_out[804];
     layer5_out[1194] <= ~layer4_out[955];
     layer5_out[1195] <= layer4_out[707];
     layer5_out[1196] <= layer4_out[1368] & layer4_out[1369];
     layer5_out[1197] <= layer4_out[462] & ~layer4_out[463];
     layer5_out[1198] <= layer4_out[22];
     layer5_out[1199] <= ~(layer4_out[963] | layer4_out[964]);
     layer5_out[1200] <= layer4_out[399] & ~layer4_out[400];
     layer5_out[1201] <= ~layer4_out[201];
     layer5_out[1202] <= 1'b0;
     layer5_out[1203] <= ~(layer4_out[694] | layer4_out[695]);
     layer5_out[1204] <= ~(layer4_out[1492] & layer4_out[1493]);
     layer5_out[1205] <= layer4_out[730];
     layer5_out[1206] <= ~layer4_out[283];
     layer5_out[1207] <= layer4_out[895] & ~layer4_out[894];
     layer5_out[1208] <= layer4_out[309] ^ layer4_out[310];
     layer5_out[1209] <= ~(layer4_out[1421] | layer4_out[1422]);
     layer5_out[1210] <= layer4_out[799];
     layer5_out[1211] <= layer4_out[933] & ~layer4_out[932];
     layer5_out[1212] <= layer4_out[124];
     layer5_out[1213] <= layer4_out[676] & ~layer4_out[677];
     layer5_out[1214] <= layer4_out[777] | layer4_out[778];
     layer5_out[1215] <= ~layer4_out[643];
     layer5_out[1216] <= layer4_out[285] & layer4_out[286];
     layer5_out[1217] <= layer4_out[143] | layer4_out[144];
     layer5_out[1218] <= ~layer4_out[121];
     layer5_out[1219] <= layer4_out[812];
     layer5_out[1220] <= ~layer4_out[409];
     layer5_out[1221] <= ~(layer4_out[637] & layer4_out[638]);
     layer5_out[1222] <= ~(layer4_out[241] ^ layer4_out[242]);
     layer5_out[1223] <= layer4_out[1065];
     layer5_out[1224] <= layer4_out[710] ^ layer4_out[711];
     layer5_out[1225] <= ~(layer4_out[1074] ^ layer4_out[1075]);
     layer5_out[1226] <= layer4_out[1485];
     layer5_out[1227] <= layer4_out[1328];
     layer5_out[1228] <= ~layer4_out[362] | layer4_out[361];
     layer5_out[1229] <= ~layer4_out[1111] | layer4_out[1112];
     layer5_out[1230] <= ~layer4_out[699];
     layer5_out[1231] <= layer4_out[1100];
     layer5_out[1232] <= ~(layer4_out[1181] & layer4_out[1182]);
     layer5_out[1233] <= layer4_out[20] & ~layer4_out[19];
     layer5_out[1234] <= ~layer4_out[249] | layer4_out[250];
     layer5_out[1235] <= layer4_out[1251] & ~layer4_out[1252];
     layer5_out[1236] <= layer4_out[994];
     layer5_out[1237] <= layer4_out[99];
     layer5_out[1238] <= ~(layer4_out[1480] & layer4_out[1481]);
     layer5_out[1239] <= layer4_out[228];
     layer5_out[1240] <= ~layer4_out[24];
     layer5_out[1241] <= layer4_out[294];
     layer5_out[1242] <= ~layer4_out[395];
     layer5_out[1243] <= ~layer4_out[1170];
     layer5_out[1244] <= ~(layer4_out[1325] & layer4_out[1326]);
     layer5_out[1245] <= ~layer4_out[526];
     layer5_out[1246] <= ~layer4_out[912];
     layer5_out[1247] <= layer4_out[884];
     layer5_out[1248] <= layer4_out[1468];
     layer5_out[1249] <= ~layer4_out[159] | layer4_out[160];
     layer5_out[1250] <= ~layer4_out[776];
     layer5_out[1251] <= layer4_out[1232];
     layer5_out[1252] <= layer4_out[729];
     layer5_out[1253] <= ~layer4_out[182] | layer4_out[181];
     layer5_out[1254] <= layer4_out[475];
     layer5_out[1255] <= 1'b0;
     layer5_out[1256] <= layer4_out[992];
     layer5_out[1257] <= ~(layer4_out[1104] & layer4_out[1105]);
     layer5_out[1258] <= layer4_out[1174];
     layer5_out[1259] <= layer4_out[30] & ~layer4_out[29];
     layer5_out[1260] <= layer4_out[229];
     layer5_out[1261] <= layer4_out[1214];
     layer5_out[1262] <= layer4_out[1379];
     layer5_out[1263] <= ~layer4_out[1128];
     layer5_out[1264] <= ~(layer4_out[33] & layer4_out[34]);
     layer5_out[1265] <= ~(layer4_out[833] & layer4_out[834]);
     layer5_out[1266] <= layer4_out[674] ^ layer4_out[675];
     layer5_out[1267] <= ~layer4_out[1395] | layer4_out[1396];
     layer5_out[1268] <= ~layer4_out[382];
     layer5_out[1269] <= ~layer4_out[539] | layer4_out[540];
     layer5_out[1270] <= ~layer4_out[1368];
     layer5_out[1271] <= ~layer4_out[1235] | layer4_out[1236];
     layer5_out[1272] <= ~layer4_out[372];
     layer5_out[1273] <= layer4_out[678];
     layer5_out[1274] <= ~layer4_out[859] | layer4_out[860];
     layer5_out[1275] <= layer4_out[1391] & layer4_out[1392];
     layer5_out[1276] <= ~layer4_out[597];
     layer5_out[1277] <= ~layer4_out[927];
     layer5_out[1278] <= ~(layer4_out[1226] ^ layer4_out[1227]);
     layer5_out[1279] <= ~layer4_out[166];
     layer5_out[1280] <= ~layer4_out[1290];
     layer5_out[1281] <= ~layer4_out[750];
     layer5_out[1282] <= ~layer4_out[1447];
     layer5_out[1283] <= layer4_out[617];
     layer5_out[1284] <= ~(layer4_out[556] | layer4_out[557]);
     layer5_out[1285] <= layer4_out[1278] | layer4_out[1279];
     layer5_out[1286] <= ~layer4_out[1470];
     layer5_out[1287] <= ~layer4_out[335];
     layer5_out[1288] <= layer4_out[1112] & layer4_out[1113];
     layer5_out[1289] <= layer4_out[461];
     layer5_out[1290] <= layer4_out[208] & ~layer4_out[209];
     layer5_out[1291] <= layer4_out[165];
     layer5_out[1292] <= ~layer4_out[1157] | layer4_out[1156];
     layer5_out[1293] <= layer4_out[656];
     layer5_out[1294] <= ~layer4_out[252] | layer4_out[251];
     layer5_out[1295] <= layer4_out[1267] ^ layer4_out[1268];
     layer5_out[1296] <= layer4_out[156] | layer4_out[157];
     layer5_out[1297] <= ~layer4_out[316];
     layer5_out[1298] <= ~layer4_out[862];
     layer5_out[1299] <= ~layer4_out[149] | layer4_out[148];
     layer5_out[1300] <= layer4_out[1272] & ~layer4_out[1273];
     layer5_out[1301] <= ~(layer4_out[563] | layer4_out[564]);
     layer5_out[1302] <= ~(layer4_out[1338] | layer4_out[1339]);
     layer5_out[1303] <= ~layer4_out[43];
     layer5_out[1304] <= ~(layer4_out[319] ^ layer4_out[320]);
     layer5_out[1305] <= ~layer4_out[1320];
     layer5_out[1306] <= ~layer4_out[76] | layer4_out[75];
     layer5_out[1307] <= layer4_out[337] | layer4_out[338];
     layer5_out[1308] <= layer4_out[1313] | layer4_out[1314];
     layer5_out[1309] <= ~layer4_out[667] | layer4_out[666];
     layer5_out[1310] <= ~layer4_out[29];
     layer5_out[1311] <= layer4_out[1481] | layer4_out[1482];
     layer5_out[1312] <= layer4_out[1115];
     layer5_out[1313] <= ~layer4_out[50];
     layer5_out[1314] <= layer4_out[1326];
     layer5_out[1315] <= layer4_out[612];
     layer5_out[1316] <= layer4_out[606] | layer4_out[607];
     layer5_out[1317] <= layer4_out[1037] ^ layer4_out[1038];
     layer5_out[1318] <= layer4_out[830];
     layer5_out[1319] <= layer4_out[820];
     layer5_out[1320] <= layer4_out[323] | layer4_out[324];
     layer5_out[1321] <= ~layer4_out[1362];
     layer5_out[1322] <= ~layer4_out[1259];
     layer5_out[1323] <= ~layer4_out[1360];
     layer5_out[1324] <= ~(layer4_out[86] & layer4_out[87]);
     layer5_out[1325] <= layer4_out[155] | layer4_out[156];
     layer5_out[1326] <= layer4_out[176] & ~layer4_out[175];
     layer5_out[1327] <= layer4_out[769];
     layer5_out[1328] <= ~(layer4_out[727] & layer4_out[728]);
     layer5_out[1329] <= ~layer4_out[1206];
     layer5_out[1330] <= layer4_out[63] & ~layer4_out[64];
     layer5_out[1331] <= layer4_out[645];
     layer5_out[1332] <= layer4_out[571] ^ layer4_out[572];
     layer5_out[1333] <= layer4_out[1168] & ~layer4_out[1167];
     layer5_out[1334] <= ~layer4_out[232];
     layer5_out[1335] <= layer4_out[19] & ~layer4_out[18];
     layer5_out[1336] <= layer4_out[946];
     layer5_out[1337] <= ~layer4_out[61];
     layer5_out[1338] <= ~layer4_out[1330];
     layer5_out[1339] <= ~layer4_out[61];
     layer5_out[1340] <= ~layer4_out[620];
     layer5_out[1341] <= 1'b0;
     layer5_out[1342] <= layer4_out[1297] & layer4_out[1298];
     layer5_out[1343] <= layer4_out[131] & ~layer4_out[130];
     layer5_out[1344] <= ~(layer4_out[1464] ^ layer4_out[1465]);
     layer5_out[1345] <= ~(layer4_out[195] | layer4_out[196]);
     layer5_out[1346] <= layer4_out[1262];
     layer5_out[1347] <= ~layer4_out[472] | layer4_out[473];
     layer5_out[1348] <= ~layer4_out[68];
     layer5_out[1349] <= layer4_out[345];
     layer5_out[1350] <= ~layer4_out[265];
     layer5_out[1351] <= ~(layer4_out[1] & layer4_out[2]);
     layer5_out[1352] <= layer4_out[1102] ^ layer4_out[1103];
     layer5_out[1353] <= ~layer4_out[445] | layer4_out[446];
     layer5_out[1354] <= layer4_out[993] ^ layer4_out[994];
     layer5_out[1355] <= layer4_out[668];
     layer5_out[1356] <= ~(layer4_out[127] | layer4_out[128]);
     layer5_out[1357] <= layer4_out[295] | layer4_out[296];
     layer5_out[1358] <= ~layer4_out[520];
     layer5_out[1359] <= ~layer4_out[1337];
     layer5_out[1360] <= ~layer4_out[577];
     layer5_out[1361] <= ~layer4_out[184] | layer4_out[185];
     layer5_out[1362] <= layer4_out[5];
     layer5_out[1363] <= ~layer4_out[750];
     layer5_out[1364] <= layer4_out[797] & ~layer4_out[798];
     layer5_out[1365] <= ~layer4_out[925];
     layer5_out[1366] <= ~layer4_out[828];
     layer5_out[1367] <= layer4_out[1308];
     layer5_out[1368] <= ~layer4_out[879];
     layer5_out[1369] <= ~layer4_out[378];
     layer5_out[1370] <= ~layer4_out[741] | layer4_out[742];
     layer5_out[1371] <= layer4_out[1418] | layer4_out[1419];
     layer5_out[1372] <= ~(layer4_out[1274] ^ layer4_out[1275]);
     layer5_out[1373] <= ~(layer4_out[1431] & layer4_out[1432]);
     layer5_out[1374] <= ~(layer4_out[465] | layer4_out[466]);
     layer5_out[1375] <= ~(layer4_out[1291] | layer4_out[1292]);
     layer5_out[1376] <= ~layer4_out[234];
     layer5_out[1377] <= ~(layer4_out[1197] & layer4_out[1198]);
     layer5_out[1378] <= layer4_out[1033];
     layer5_out[1379] <= ~(layer4_out[906] | layer4_out[907]);
     layer5_out[1380] <= ~layer4_out[811] | layer4_out[810];
     layer5_out[1381] <= ~(layer4_out[817] ^ layer4_out[818]);
     layer5_out[1382] <= ~layer4_out[1404] | layer4_out[1405];
     layer5_out[1383] <= layer4_out[1288] | layer4_out[1289];
     layer5_out[1384] <= ~(layer4_out[1252] ^ layer4_out[1253]);
     layer5_out[1385] <= ~layer4_out[111] | layer4_out[112];
     layer5_out[1386] <= ~(layer4_out[329] & layer4_out[330]);
     layer5_out[1387] <= layer4_out[379] & ~layer4_out[380];
     layer5_out[1388] <= ~(layer4_out[31] | layer4_out[32]);
     layer5_out[1389] <= layer4_out[587];
     layer5_out[1390] <= ~layer4_out[998];
     layer5_out[1391] <= ~layer4_out[888];
     layer5_out[1392] <= ~layer4_out[1402];
     layer5_out[1393] <= ~(layer4_out[884] & layer4_out[885]);
     layer5_out[1394] <= ~layer4_out[313];
     layer5_out[1395] <= layer4_out[189] & layer4_out[190];
     layer5_out[1396] <= layer4_out[557];
     layer5_out[1397] <= layer4_out[1450];
     layer5_out[1398] <= layer4_out[284] & layer4_out[285];
     layer5_out[1399] <= ~(layer4_out[981] & layer4_out[982]);
     layer5_out[1400] <= layer4_out[1316];
     layer5_out[1401] <= ~layer4_out[634];
     layer5_out[1402] <= layer4_out[1489] & layer4_out[1490];
     layer5_out[1403] <= ~layer4_out[192] | layer4_out[193];
     layer5_out[1404] <= layer4_out[613];
     layer5_out[1405] <= ~(layer4_out[311] ^ layer4_out[312]);
     layer5_out[1406] <= ~(layer4_out[506] | layer4_out[507]);
     layer5_out[1407] <= layer4_out[253];
     layer5_out[1408] <= ~layer4_out[649];
     layer5_out[1409] <= ~(layer4_out[1124] & layer4_out[1125]);
     layer5_out[1410] <= layer4_out[466] & ~layer4_out[467];
     layer5_out[1411] <= layer4_out[193];
     layer5_out[1412] <= layer4_out[988] & ~layer4_out[989];
     layer5_out[1413] <= layer4_out[408] & layer4_out[409];
     layer5_out[1414] <= ~layer4_out[392];
     layer5_out[1415] <= ~layer4_out[1];
     layer5_out[1416] <= layer4_out[1031];
     layer5_out[1417] <= layer4_out[278] & ~layer4_out[279];
     layer5_out[1418] <= ~(layer4_out[483] ^ layer4_out[484]);
     layer5_out[1419] <= layer4_out[424];
     layer5_out[1420] <= ~layer4_out[405];
     layer5_out[1421] <= layer4_out[913];
     layer5_out[1422] <= layer4_out[134] | layer4_out[135];
     layer5_out[1423] <= ~layer4_out[1285] | layer4_out[1284];
     layer5_out[1424] <= layer4_out[459];
     layer5_out[1425] <= layer4_out[52];
     layer5_out[1426] <= ~layer4_out[972];
     layer5_out[1427] <= ~layer4_out[474];
     layer5_out[1428] <= layer4_out[880] & layer4_out[881];
     layer5_out[1429] <= ~layer4_out[236];
     layer5_out[1430] <= layer4_out[324];
     layer5_out[1431] <= layer4_out[1317];
     layer5_out[1432] <= ~layer4_out[707];
     layer5_out[1433] <= layer4_out[113];
     layer5_out[1434] <= ~layer4_out[1196];
     layer5_out[1435] <= layer4_out[78];
     layer5_out[1436] <= layer4_out[976];
     layer5_out[1437] <= ~layer4_out[1109] | layer4_out[1110];
     layer5_out[1438] <= layer4_out[785] & ~layer4_out[784];
     layer5_out[1439] <= layer4_out[289] & ~layer4_out[288];
     layer5_out[1440] <= layer4_out[1213];
     layer5_out[1441] <= layer4_out[889] ^ layer4_out[890];
     layer5_out[1442] <= layer4_out[301] ^ layer4_out[302];
     layer5_out[1443] <= layer4_out[760];
     layer5_out[1444] <= layer4_out[1307];
     layer5_out[1445] <= ~layer4_out[481] | layer4_out[482];
     layer5_out[1446] <= ~layer4_out[1192] | layer4_out[1193];
     layer5_out[1447] <= layer4_out[870];
     layer5_out[1448] <= layer4_out[986];
     layer5_out[1449] <= layer4_out[254];
     layer5_out[1450] <= ~layer4_out[37];
     layer5_out[1451] <= ~layer4_out[1475];
     layer5_out[1452] <= ~layer4_out[1072];
     layer5_out[1453] <= ~layer4_out[704];
     layer5_out[1454] <= ~(layer4_out[1025] & layer4_out[1026]);
     layer5_out[1455] <= ~layer4_out[1274];
     layer5_out[1456] <= ~(layer4_out[573] ^ layer4_out[574]);
     layer5_out[1457] <= ~layer4_out[1177];
     layer5_out[1458] <= layer4_out[807] | layer4_out[808];
     layer5_out[1459] <= layer4_out[649] & ~layer4_out[650];
     layer5_out[1460] <= ~layer4_out[597];
     layer5_out[1461] <= layer4_out[874];
     layer5_out[1462] <= ~(layer4_out[1234] | layer4_out[1235]);
     layer5_out[1463] <= ~(layer4_out[835] | layer4_out[836]);
     layer5_out[1464] <= layer4_out[416];
     layer5_out[1465] <= ~(layer4_out[600] | layer4_out[601]);
     layer5_out[1466] <= layer4_out[785];
     layer5_out[1467] <= layer4_out[1251];
     layer5_out[1468] <= ~layer4_out[1135];
     layer5_out[1469] <= layer4_out[901];
     layer5_out[1470] <= ~layer4_out[1350];
     layer5_out[1471] <= layer4_out[20] & ~layer4_out[21];
     layer5_out[1472] <= ~layer4_out[522];
     layer5_out[1473] <= layer4_out[216] ^ layer4_out[217];
     layer5_out[1474] <= ~(layer4_out[131] | layer4_out[132]);
     layer5_out[1475] <= ~layer4_out[968] | layer4_out[967];
     layer5_out[1476] <= ~layer4_out[32];
     layer5_out[1477] <= ~layer4_out[1379];
     layer5_out[1478] <= layer4_out[25] & layer4_out[26];
     layer5_out[1479] <= ~(layer4_out[995] & layer4_out[996]);
     layer5_out[1480] <= ~layer4_out[1417];
     layer5_out[1481] <= ~(layer4_out[289] | layer4_out[290]);
     layer5_out[1482] <= ~layer4_out[486];
     layer5_out[1483] <= ~layer4_out[1204];
     layer5_out[1484] <= 1'b1;
     layer5_out[1485] <= ~layer4_out[231];
     layer5_out[1486] <= layer4_out[311] & ~layer4_out[310];
     layer5_out[1487] <= ~(layer4_out[1162] | layer4_out[1163]);
     layer5_out[1488] <= ~layer4_out[511];
     layer5_out[1489] <= ~layer4_out[561] | layer4_out[562];
     layer5_out[1490] <= layer4_out[1053];
     layer5_out[1491] <= layer4_out[71];
     layer5_out[1492] <= ~layer4_out[502];
     layer5_out[1493] <= layer4_out[1119] & ~layer4_out[1120];
     layer5_out[1494] <= layer4_out[661] & ~layer4_out[662];
     layer5_out[1495] <= ~layer4_out[1386] | layer4_out[1385];
     layer5_out[1496] <= ~(layer4_out[304] | layer4_out[305]);
     layer5_out[1497] <= layer4_out[1490];
     layer5_out[1498] <= layer4_out[85] & layer4_out[86];
     layer5_out[1499] <= ~(layer4_out[1403] & layer4_out[1404]);
     layer6_out[0] <= layer5_out[460];
     layer6_out[1] <= ~(layer5_out[1413] | layer5_out[1414]);
     layer6_out[2] <= 1'b0;
     layer6_out[3] <= ~(layer5_out[32] ^ layer5_out[33]);
     layer6_out[4] <= ~(layer5_out[1460] ^ layer5_out[1461]);
     layer6_out[5] <= ~layer5_out[104];
     layer6_out[6] <= layer5_out[236] ^ layer5_out[237];
     layer6_out[7] <= layer5_out[1067];
     layer6_out[8] <= layer5_out[789] | layer5_out[790];
     layer6_out[9] <= ~layer5_out[914] | layer5_out[915];
     layer6_out[10] <= ~layer5_out[942];
     layer6_out[11] <= ~layer5_out[43];
     layer6_out[12] <= layer5_out[429];
     layer6_out[13] <= ~layer5_out[506] | layer5_out[507];
     layer6_out[14] <= layer5_out[1092];
     layer6_out[15] <= ~layer5_out[492];
     layer6_out[16] <= layer5_out[720] & ~layer5_out[719];
     layer6_out[17] <= ~(layer5_out[463] | layer5_out[464]);
     layer6_out[18] <= ~layer5_out[736];
     layer6_out[19] <= layer5_out[1029];
     layer6_out[20] <= ~layer5_out[148];
     layer6_out[21] <= layer5_out[1112];
     layer6_out[22] <= ~layer5_out[802];
     layer6_out[23] <= layer5_out[910];
     layer6_out[24] <= layer5_out[114] ^ layer5_out[115];
     layer6_out[25] <= ~layer5_out[627] | layer5_out[626];
     layer6_out[26] <= layer5_out[196] & ~layer5_out[195];
     layer6_out[27] <= layer5_out[647] & layer5_out[648];
     layer6_out[28] <= layer5_out[466] & layer5_out[467];
     layer6_out[29] <= ~(layer5_out[1189] | layer5_out[1190]);
     layer6_out[30] <= ~layer5_out[347];
     layer6_out[31] <= ~layer5_out[1202];
     layer6_out[32] <= layer5_out[1419] ^ layer5_out[1420];
     layer6_out[33] <= ~layer5_out[1309] | layer5_out[1308];
     layer6_out[34] <= ~layer5_out[508];
     layer6_out[35] <= layer5_out[1406];
     layer6_out[36] <= ~layer5_out[385];
     layer6_out[37] <= layer5_out[462] | layer5_out[463];
     layer6_out[38] <= layer5_out[583];
     layer6_out[39] <= layer5_out[645];
     layer6_out[40] <= ~layer5_out[378] | layer5_out[379];
     layer6_out[41] <= 1'b0;
     layer6_out[42] <= ~layer5_out[1411] | layer5_out[1412];
     layer6_out[43] <= ~layer5_out[750];
     layer6_out[44] <= ~layer5_out[632];
     layer6_out[45] <= ~layer5_out[841] | layer5_out[842];
     layer6_out[46] <= ~(layer5_out[285] | layer5_out[286]);
     layer6_out[47] <= ~layer5_out[1413];
     layer6_out[48] <= ~layer5_out[47];
     layer6_out[49] <= ~(layer5_out[96] | layer5_out[97]);
     layer6_out[50] <= layer5_out[27];
     layer6_out[51] <= layer5_out[411];
     layer6_out[52] <= ~(layer5_out[517] ^ layer5_out[518]);
     layer6_out[53] <= layer5_out[945] & layer5_out[946];
     layer6_out[54] <= layer5_out[1084] ^ layer5_out[1085];
     layer6_out[55] <= layer5_out[739] ^ layer5_out[740];
     layer6_out[56] <= ~layer5_out[1318];
     layer6_out[57] <= layer5_out[322];
     layer6_out[58] <= ~(layer5_out[1011] ^ layer5_out[1012]);
     layer6_out[59] <= layer5_out[667] & ~layer5_out[666];
     layer6_out[60] <= layer5_out[526];
     layer6_out[61] <= ~layer5_out[249] | layer5_out[250];
     layer6_out[62] <= ~layer5_out[1164];
     layer6_out[63] <= ~layer5_out[71];
     layer6_out[64] <= layer5_out[785];
     layer6_out[65] <= ~layer5_out[698];
     layer6_out[66] <= layer5_out[582] ^ layer5_out[583];
     layer6_out[67] <= layer5_out[491] & ~layer5_out[490];
     layer6_out[68] <= layer5_out[330] & ~layer5_out[331];
     layer6_out[69] <= 1'b1;
     layer6_out[70] <= layer5_out[468] & ~layer5_out[467];
     layer6_out[71] <= ~(layer5_out[324] & layer5_out[325]);
     layer6_out[72] <= ~layer5_out[70];
     layer6_out[73] <= ~(layer5_out[777] ^ layer5_out[778]);
     layer6_out[74] <= layer5_out[1122] & ~layer5_out[1123];
     layer6_out[75] <= layer5_out[1176] & ~layer5_out[1177];
     layer6_out[76] <= ~layer5_out[979];
     layer6_out[77] <= layer5_out[1488] & ~layer5_out[1487];
     layer6_out[78] <= layer5_out[362] & layer5_out[363];
     layer6_out[79] <= layer5_out[221] ^ layer5_out[222];
     layer6_out[80] <= layer5_out[311] | layer5_out[312];
     layer6_out[81] <= ~layer5_out[966] | layer5_out[967];
     layer6_out[82] <= ~layer5_out[117] | layer5_out[116];
     layer6_out[83] <= ~layer5_out[784];
     layer6_out[84] <= layer5_out[612] ^ layer5_out[613];
     layer6_out[85] <= ~layer5_out[813];
     layer6_out[86] <= ~layer5_out[1024] | layer5_out[1023];
     layer6_out[87] <= ~layer5_out[47];
     layer6_out[88] <= layer5_out[1278];
     layer6_out[89] <= layer5_out[321];
     layer6_out[90] <= layer5_out[1365];
     layer6_out[91] <= ~layer5_out[1231] | layer5_out[1232];
     layer6_out[92] <= ~(layer5_out[575] ^ layer5_out[576]);
     layer6_out[93] <= layer5_out[89] | layer5_out[90];
     layer6_out[94] <= layer5_out[140];
     layer6_out[95] <= layer5_out[1166] ^ layer5_out[1167];
     layer6_out[96] <= layer5_out[187] | layer5_out[188];
     layer6_out[97] <= layer5_out[416];
     layer6_out[98] <= layer5_out[1182];
     layer6_out[99] <= ~layer5_out[427] | layer5_out[428];
     layer6_out[100] <= ~layer5_out[1008];
     layer6_out[101] <= ~layer5_out[1062] | layer5_out[1063];
     layer6_out[102] <= ~layer5_out[1022] | layer5_out[1023];
     layer6_out[103] <= layer5_out[1238];
     layer6_out[104] <= layer5_out[1330] ^ layer5_out[1331];
     layer6_out[105] <= layer5_out[1438];
     layer6_out[106] <= layer5_out[1454] & layer5_out[1455];
     layer6_out[107] <= layer5_out[646];
     layer6_out[108] <= layer5_out[1493];
     layer6_out[109] <= layer5_out[383];
     layer6_out[110] <= layer5_out[1151];
     layer6_out[111] <= ~layer5_out[456];
     layer6_out[112] <= ~layer5_out[1073];
     layer6_out[113] <= ~layer5_out[683];
     layer6_out[114] <= layer5_out[759] ^ layer5_out[760];
     layer6_out[115] <= layer5_out[1430];
     layer6_out[116] <= layer5_out[553] & ~layer5_out[554];
     layer6_out[117] <= layer5_out[724];
     layer6_out[118] <= ~(layer5_out[97] | layer5_out[98]);
     layer6_out[119] <= layer5_out[1016] & ~layer5_out[1017];
     layer6_out[120] <= ~layer5_out[972];
     layer6_out[121] <= layer5_out[0] & ~layer5_out[2];
     layer6_out[122] <= layer5_out[758] | layer5_out[759];
     layer6_out[123] <= layer5_out[623];
     layer6_out[124] <= ~layer5_out[782];
     layer6_out[125] <= layer5_out[1246] & layer5_out[1247];
     layer6_out[126] <= layer5_out[602];
     layer6_out[127] <= layer5_out[931];
     layer6_out[128] <= layer5_out[239] | layer5_out[240];
     layer6_out[129] <= 1'b0;
     layer6_out[130] <= layer5_out[955] | layer5_out[956];
     layer6_out[131] <= ~(layer5_out[1496] | layer5_out[1497]);
     layer6_out[132] <= layer5_out[419];
     layer6_out[133] <= layer5_out[613];
     layer6_out[134] <= layer5_out[379] & layer5_out[380];
     layer6_out[135] <= ~layer5_out[838];
     layer6_out[136] <= ~layer5_out[972];
     layer6_out[137] <= ~layer5_out[1251] | layer5_out[1250];
     layer6_out[138] <= layer5_out[660] & ~layer5_out[659];
     layer6_out[139] <= ~(layer5_out[1270] ^ layer5_out[1271]);
     layer6_out[140] <= ~layer5_out[792] | layer5_out[791];
     layer6_out[141] <= layer5_out[1379];
     layer6_out[142] <= layer5_out[180] & ~layer5_out[179];
     layer6_out[143] <= ~layer5_out[1212];
     layer6_out[144] <= layer5_out[929];
     layer6_out[145] <= layer5_out[425] | layer5_out[426];
     layer6_out[146] <= 1'b1;
     layer6_out[147] <= layer5_out[711] ^ layer5_out[712];
     layer6_out[148] <= ~layer5_out[306];
     layer6_out[149] <= layer5_out[1276];
     layer6_out[150] <= layer5_out[1382] ^ layer5_out[1383];
     layer6_out[151] <= ~layer5_out[1280] | layer5_out[1281];
     layer6_out[152] <= layer5_out[712];
     layer6_out[153] <= ~layer5_out[804] | layer5_out[805];
     layer6_out[154] <= ~layer5_out[1237] | layer5_out[1236];
     layer6_out[155] <= ~layer5_out[1030] | layer5_out[1031];
     layer6_out[156] <= layer5_out[1351];
     layer6_out[157] <= layer5_out[1003] & ~layer5_out[1002];
     layer6_out[158] <= ~layer5_out[1064] | layer5_out[1065];
     layer6_out[159] <= ~layer5_out[1060];
     layer6_out[160] <= ~(layer5_out[1381] ^ layer5_out[1382]);
     layer6_out[161] <= ~layer5_out[535];
     layer6_out[162] <= layer5_out[234] ^ layer5_out[235];
     layer6_out[163] <= ~(layer5_out[1129] & layer5_out[1130]);
     layer6_out[164] <= layer5_out[686];
     layer6_out[165] <= ~layer5_out[207];
     layer6_out[166] <= layer5_out[554] | layer5_out[555];
     layer6_out[167] <= layer5_out[1297];
     layer6_out[168] <= ~layer5_out[464] | layer5_out[465];
     layer6_out[169] <= layer5_out[952];
     layer6_out[170] <= layer5_out[1025];
     layer6_out[171] <= ~layer5_out[258] | layer5_out[259];
     layer6_out[172] <= ~(layer5_out[198] | layer5_out[199]);
     layer6_out[173] <= ~(layer5_out[890] | layer5_out[891]);
     layer6_out[174] <= ~layer5_out[1314] | layer5_out[1313];
     layer6_out[175] <= layer5_out[1489] & ~layer5_out[1488];
     layer6_out[176] <= ~layer5_out[494];
     layer6_out[177] <= ~layer5_out[1341];
     layer6_out[178] <= layer5_out[257] & ~layer5_out[256];
     layer6_out[179] <= ~layer5_out[1241];
     layer6_out[180] <= layer5_out[826] & ~layer5_out[825];
     layer6_out[181] <= ~layer5_out[1168];
     layer6_out[182] <= ~layer5_out[1294];
     layer6_out[183] <= ~(layer5_out[1086] | layer5_out[1087]);
     layer6_out[184] <= layer5_out[1384];
     layer6_out[185] <= layer5_out[62];
     layer6_out[186] <= ~layer5_out[418];
     layer6_out[187] <= ~layer5_out[963];
     layer6_out[188] <= layer5_out[611] ^ layer5_out[612];
     layer6_out[189] <= layer5_out[794];
     layer6_out[190] <= ~layer5_out[437];
     layer6_out[191] <= ~(layer5_out[713] | layer5_out[714]);
     layer6_out[192] <= layer5_out[805] & layer5_out[806];
     layer6_out[193] <= ~layer5_out[984] | layer5_out[983];
     layer6_out[194] <= ~layer5_out[526];
     layer6_out[195] <= layer5_out[710];
     layer6_out[196] <= ~layer5_out[907];
     layer6_out[197] <= ~(layer5_out[894] | layer5_out[895]);
     layer6_out[198] <= ~layer5_out[684];
     layer6_out[199] <= ~(layer5_out[247] ^ layer5_out[248]);
     layer6_out[200] <= layer5_out[1298] & layer5_out[1299];
     layer6_out[201] <= layer5_out[300] ^ layer5_out[301];
     layer6_out[202] <= ~layer5_out[552];
     layer6_out[203] <= ~layer5_out[1426];
     layer6_out[204] <= layer5_out[1125];
     layer6_out[205] <= 1'b1;
     layer6_out[206] <= ~layer5_out[218];
     layer6_out[207] <= layer5_out[843] & ~layer5_out[842];
     layer6_out[208] <= layer5_out[1400] | layer5_out[1401];
     layer6_out[209] <= ~layer5_out[1079];
     layer6_out[210] <= ~layer5_out[359];
     layer6_out[211] <= ~layer5_out[798] | layer5_out[799];
     layer6_out[212] <= ~layer5_out[859] | layer5_out[860];
     layer6_out[213] <= ~layer5_out[761] | layer5_out[762];
     layer6_out[214] <= layer5_out[690];
     layer6_out[215] <= layer5_out[989];
     layer6_out[216] <= layer5_out[777];
     layer6_out[217] <= ~(layer5_out[555] | layer5_out[556]);
     layer6_out[218] <= ~(layer5_out[87] & layer5_out[88]);
     layer6_out[219] <= layer5_out[1165] ^ layer5_out[1166];
     layer6_out[220] <= layer5_out[1155];
     layer6_out[221] <= layer5_out[780];
     layer6_out[222] <= layer5_out[731] & layer5_out[732];
     layer6_out[223] <= layer5_out[75] ^ layer5_out[76];
     layer6_out[224] <= ~layer5_out[73];
     layer6_out[225] <= ~layer5_out[429] | layer5_out[430];
     layer6_out[226] <= ~layer5_out[519];
     layer6_out[227] <= layer5_out[402] & ~layer5_out[401];
     layer6_out[228] <= layer5_out[836];
     layer6_out[229] <= layer5_out[908];
     layer6_out[230] <= ~(layer5_out[590] | layer5_out[591]);
     layer6_out[231] <= layer5_out[1314];
     layer6_out[232] <= layer5_out[244];
     layer6_out[233] <= layer5_out[749] ^ layer5_out[750];
     layer6_out[234] <= layer5_out[643];
     layer6_out[235] <= layer5_out[93];
     layer6_out[236] <= ~layer5_out[160];
     layer6_out[237] <= layer5_out[367];
     layer6_out[238] <= layer5_out[1233] & layer5_out[1234];
     layer6_out[239] <= layer5_out[1303] ^ layer5_out[1304];
     layer6_out[240] <= layer5_out[1200] & ~layer5_out[1199];
     layer6_out[241] <= layer5_out[741];
     layer6_out[242] <= layer5_out[1179];
     layer6_out[243] <= layer5_out[136] & ~layer5_out[135];
     layer6_out[244] <= layer5_out[803] | layer5_out[804];
     layer6_out[245] <= layer5_out[431] & ~layer5_out[432];
     layer6_out[246] <= ~layer5_out[531];
     layer6_out[247] <= layer5_out[1329] & ~layer5_out[1328];
     layer6_out[248] <= layer5_out[640];
     layer6_out[249] <= layer5_out[150];
     layer6_out[250] <= layer5_out[967] | layer5_out[968];
     layer6_out[251] <= layer5_out[744];
     layer6_out[252] <= layer5_out[1464];
     layer6_out[253] <= ~(layer5_out[940] | layer5_out[941]);
     layer6_out[254] <= layer5_out[262] ^ layer5_out[263];
     layer6_out[255] <= ~layer5_out[1086];
     layer6_out[256] <= ~(layer5_out[86] & layer5_out[87]);
     layer6_out[257] <= ~(layer5_out[1269] | layer5_out[1270]);
     layer6_out[258] <= ~layer5_out[1063];
     layer6_out[259] <= ~layer5_out[572];
     layer6_out[260] <= layer5_out[439] & ~layer5_out[440];
     layer6_out[261] <= 1'b0;
     layer6_out[262] <= ~layer5_out[808];
     layer6_out[263] <= layer5_out[1225];
     layer6_out[264] <= ~(layer5_out[856] | layer5_out[857]);
     layer6_out[265] <= layer5_out[12];
     layer6_out[266] <= ~layer5_out[1428];
     layer6_out[267] <= ~layer5_out[532];
     layer6_out[268] <= ~(layer5_out[716] ^ layer5_out[717]);
     layer6_out[269] <= ~layer5_out[110];
     layer6_out[270] <= ~(layer5_out[1200] ^ layer5_out[1201]);
     layer6_out[271] <= ~layer5_out[131];
     layer6_out[272] <= layer5_out[919] & ~layer5_out[918];
     layer6_out[273] <= layer5_out[974] & ~layer5_out[975];
     layer6_out[274] <= ~layer5_out[277] | layer5_out[278];
     layer6_out[275] <= layer5_out[1261];
     layer6_out[276] <= ~(layer5_out[950] & layer5_out[951]);
     layer6_out[277] <= ~(layer5_out[465] | layer5_out[466]);
     layer6_out[278] <= ~(layer5_out[237] ^ layer5_out[238]);
     layer6_out[279] <= ~layer5_out[1456] | layer5_out[1457];
     layer6_out[280] <= ~layer5_out[371];
     layer6_out[281] <= ~layer5_out[948];
     layer6_out[282] <= layer5_out[670] ^ layer5_out[671];
     layer6_out[283] <= layer5_out[1388];
     layer6_out[284] <= layer5_out[1008] ^ layer5_out[1009];
     layer6_out[285] <= 1'b1;
     layer6_out[286] <= layer5_out[408] & ~layer5_out[407];
     layer6_out[287] <= ~layer5_out[901] | layer5_out[900];
     layer6_out[288] <= ~layer5_out[1479];
     layer6_out[289] <= ~(layer5_out[899] | layer5_out[900]);
     layer6_out[290] <= layer5_out[728] | layer5_out[729];
     layer6_out[291] <= layer5_out[1360];
     layer6_out[292] <= ~layer5_out[970];
     layer6_out[293] <= ~layer5_out[174];
     layer6_out[294] <= layer5_out[994] & ~layer5_out[993];
     layer6_out[295] <= ~(layer5_out[399] & layer5_out[400]);
     layer6_out[296] <= ~(layer5_out[1478] & layer5_out[1479]);
     layer6_out[297] <= layer5_out[304];
     layer6_out[298] <= ~layer5_out[917] | layer5_out[918];
     layer6_out[299] <= layer5_out[1184] | layer5_out[1185];
     layer6_out[300] <= layer5_out[844];
     layer6_out[301] <= ~layer5_out[1227];
     layer6_out[302] <= layer5_out[904];
     layer6_out[303] <= layer5_out[1409] & ~layer5_out[1410];
     layer6_out[304] <= layer5_out[204] | layer5_out[205];
     layer6_out[305] <= ~(layer5_out[298] ^ layer5_out[299]);
     layer6_out[306] <= ~(layer5_out[1160] & layer5_out[1161]);
     layer6_out[307] <= layer5_out[603] & layer5_out[604];
     layer6_out[308] <= layer5_out[291] & ~layer5_out[290];
     layer6_out[309] <= layer5_out[1489] & ~layer5_out[1490];
     layer6_out[310] <= 1'b1;
     layer6_out[311] <= ~layer5_out[1485];
     layer6_out[312] <= ~layer5_out[365];
     layer6_out[313] <= layer5_out[325];
     layer6_out[314] <= layer5_out[1052];
     layer6_out[315] <= layer5_out[1465] | layer5_out[1466];
     layer6_out[316] <= ~(layer5_out[305] & layer5_out[306]);
     layer6_out[317] <= ~(layer5_out[1010] ^ layer5_out[1011]);
     layer6_out[318] <= ~layer5_out[1305];
     layer6_out[319] <= layer5_out[461] & layer5_out[462];
     layer6_out[320] <= ~layer5_out[135] | layer5_out[134];
     layer6_out[321] <= layer5_out[558] & layer5_out[559];
     layer6_out[322] <= layer5_out[317] ^ layer5_out[318];
     layer6_out[323] <= ~layer5_out[299];
     layer6_out[324] <= layer5_out[232];
     layer6_out[325] <= layer5_out[1094];
     layer6_out[326] <= layer5_out[231] & ~layer5_out[230];
     layer6_out[327] <= ~layer5_out[954];
     layer6_out[328] <= layer5_out[1260] & ~layer5_out[1259];
     layer6_out[329] <= layer5_out[342];
     layer6_out[330] <= layer5_out[137];
     layer6_out[331] <= layer5_out[1335] ^ layer5_out[1336];
     layer6_out[332] <= layer5_out[394];
     layer6_out[333] <= ~layer5_out[851];
     layer6_out[334] <= ~layer5_out[231];
     layer6_out[335] <= 1'b0;
     layer6_out[336] <= layer5_out[548] | layer5_out[549];
     layer6_out[337] <= layer5_out[1060];
     layer6_out[338] <= ~layer5_out[1242];
     layer6_out[339] <= layer5_out[407];
     layer6_out[340] <= layer5_out[690] & ~layer5_out[691];
     layer6_out[341] <= layer5_out[1193] & ~layer5_out[1192];
     layer6_out[342] <= ~layer5_out[108];
     layer6_out[343] <= layer5_out[523];
     layer6_out[344] <= layer5_out[16];
     layer6_out[345] <= layer5_out[197];
     layer6_out[346] <= ~(layer5_out[951] & layer5_out[952]);
     layer6_out[347] <= ~(layer5_out[591] | layer5_out[592]);
     layer6_out[348] <= layer5_out[692];
     layer6_out[349] <= ~layer5_out[354];
     layer6_out[350] <= layer5_out[505];
     layer6_out[351] <= 1'b0;
     layer6_out[352] <= layer5_out[431] & ~layer5_out[430];
     layer6_out[353] <= ~layer5_out[269];
     layer6_out[354] <= layer5_out[1393] & layer5_out[1394];
     layer6_out[355] <= ~layer5_out[142] | layer5_out[143];
     layer6_out[356] <= layer5_out[353];
     layer6_out[357] <= layer5_out[610];
     layer6_out[358] <= ~layer5_out[332];
     layer6_out[359] <= layer5_out[1336];
     layer6_out[360] <= ~(layer5_out[809] & layer5_out[810]);
     layer6_out[361] <= ~layer5_out[183];
     layer6_out[362] <= ~(layer5_out[589] ^ layer5_out[590]);
     layer6_out[363] <= 1'b1;
     layer6_out[364] <= ~layer5_out[765];
     layer6_out[365] <= layer5_out[1353];
     layer6_out[366] <= layer5_out[314];
     layer6_out[367] <= layer5_out[5];
     layer6_out[368] <= ~layer5_out[211] | layer5_out[212];
     layer6_out[369] <= layer5_out[1475];
     layer6_out[370] <= ~layer5_out[403];
     layer6_out[371] <= ~layer5_out[1268];
     layer6_out[372] <= layer5_out[227];
     layer6_out[373] <= layer5_out[268];
     layer6_out[374] <= layer5_out[819] & ~layer5_out[818];
     layer6_out[375] <= ~(layer5_out[113] | layer5_out[114]);
     layer6_out[376] <= layer5_out[770];
     layer6_out[377] <= layer5_out[1250] & ~layer5_out[1249];
     layer6_out[378] <= ~layer5_out[892];
     layer6_out[379] <= ~layer5_out[1073];
     layer6_out[380] <= ~layer5_out[1271];
     layer6_out[381] <= ~layer5_out[1317];
     layer6_out[382] <= ~layer5_out[472] | layer5_out[473];
     layer6_out[383] <= layer5_out[1070] & ~layer5_out[1071];
     layer6_out[384] <= layer5_out[1343];
     layer6_out[385] <= layer5_out[1155];
     layer6_out[386] <= layer5_out[240] | layer5_out[241];
     layer6_out[387] <= layer5_out[1295];
     layer6_out[388] <= ~layer5_out[435] | layer5_out[434];
     layer6_out[389] <= layer5_out[228] ^ layer5_out[229];
     layer6_out[390] <= layer5_out[593];
     layer6_out[391] <= ~layer5_out[1149];
     layer6_out[392] <= layer5_out[877];
     layer6_out[393] <= layer5_out[1175] ^ layer5_out[1176];
     layer6_out[394] <= ~(layer5_out[1347] & layer5_out[1348]);
     layer6_out[395] <= layer5_out[168] ^ layer5_out[169];
     layer6_out[396] <= layer5_out[1121] | layer5_out[1122];
     layer6_out[397] <= layer5_out[1120] & ~layer5_out[1121];
     layer6_out[398] <= layer5_out[58] & layer5_out[59];
     layer6_out[399] <= ~(layer5_out[1253] ^ layer5_out[1254]);
     layer6_out[400] <= layer5_out[319];
     layer6_out[401] <= layer5_out[279];
     layer6_out[402] <= layer5_out[1481] & ~layer5_out[1480];
     layer6_out[403] <= layer5_out[199] | layer5_out[200];
     layer6_out[404] <= ~layer5_out[996];
     layer6_out[405] <= ~layer5_out[1075];
     layer6_out[406] <= ~layer5_out[1195] | layer5_out[1196];
     layer6_out[407] <= ~layer5_out[992];
     layer6_out[408] <= layer5_out[193] ^ layer5_out[194];
     layer6_out[409] <= layer5_out[1077] ^ layer5_out[1078];
     layer6_out[410] <= layer5_out[1483] & ~layer5_out[1484];
     layer6_out[411] <= layer5_out[415] & ~layer5_out[416];
     layer6_out[412] <= layer5_out[214] ^ layer5_out[215];
     layer6_out[413] <= ~layer5_out[987];
     layer6_out[414] <= ~layer5_out[819];
     layer6_out[415] <= ~(layer5_out[1416] ^ layer5_out[1417]);
     layer6_out[416] <= ~layer5_out[157];
     layer6_out[417] <= layer5_out[1349] & ~layer5_out[1348];
     layer6_out[418] <= ~layer5_out[999] | layer5_out[998];
     layer6_out[419] <= ~layer5_out[825];
     layer6_out[420] <= layer5_out[671] | layer5_out[672];
     layer6_out[421] <= ~(layer5_out[81] ^ layer5_out[82]);
     layer6_out[422] <= ~layer5_out[630];
     layer6_out[423] <= layer5_out[1376] & layer5_out[1377];
     layer6_out[424] <= 1'b0;
     layer6_out[425] <= ~(layer5_out[834] | layer5_out[835]);
     layer6_out[426] <= layer5_out[1300] | layer5_out[1301];
     layer6_out[427] <= layer5_out[68];
     layer6_out[428] <= layer5_out[1163];
     layer6_out[429] <= layer5_out[239];
     layer6_out[430] <= ~layer5_out[83];
     layer6_out[431] <= layer5_out[1031];
     layer6_out[432] <= ~layer5_out[985];
     layer6_out[433] <= ~(layer5_out[1096] | layer5_out[1097]);
     layer6_out[434] <= ~(layer5_out[1194] | layer5_out[1195]);
     layer6_out[435] <= layer5_out[316] & ~layer5_out[315];
     layer6_out[436] <= layer5_out[499];
     layer6_out[437] <= layer5_out[45];
     layer6_out[438] <= ~(layer5_out[395] & layer5_out[396]);
     layer6_out[439] <= ~layer5_out[1226];
     layer6_out[440] <= layer5_out[1324] ^ layer5_out[1325];
     layer6_out[441] <= ~layer5_out[1152];
     layer6_out[442] <= layer5_out[550] & layer5_out[551];
     layer6_out[443] <= layer5_out[23] & ~layer5_out[22];
     layer6_out[444] <= layer5_out[18];
     layer6_out[445] <= layer5_out[56] & ~layer5_out[57];
     layer6_out[446] <= ~layer5_out[830];
     layer6_out[447] <= layer5_out[986] ^ layer5_out[987];
     layer6_out[448] <= layer5_out[420];
     layer6_out[449] <= layer5_out[252];
     layer6_out[450] <= layer5_out[375] & ~layer5_out[374];
     layer6_out[451] <= ~layer5_out[969];
     layer6_out[452] <= layer5_out[1286] & layer5_out[1287];
     layer6_out[453] <= ~layer5_out[178];
     layer6_out[454] <= layer5_out[1451] & layer5_out[1452];
     layer6_out[455] <= layer5_out[265] | layer5_out[266];
     layer6_out[456] <= layer5_out[1055];
     layer6_out[457] <= layer5_out[30];
     layer6_out[458] <= ~layer5_out[1262] | layer5_out[1261];
     layer6_out[459] <= ~(layer5_out[527] ^ layer5_out[528]);
     layer6_out[460] <= layer5_out[1133] & ~layer5_out[1134];
     layer6_out[461] <= ~layer5_out[377] | layer5_out[378];
     layer6_out[462] <= ~layer5_out[476];
     layer6_out[463] <= layer5_out[828] ^ layer5_out[829];
     layer6_out[464] <= layer5_out[599];
     layer6_out[465] <= ~layer5_out[272];
     layer6_out[466] <= layer5_out[639];
     layer6_out[467] <= ~layer5_out[655] | layer5_out[656];
     layer6_out[468] <= layer5_out[1256] | layer5_out[1257];
     layer6_out[469] <= layer5_out[699] & layer5_out[700];
     layer6_out[470] <= layer5_out[129];
     layer6_out[471] <= ~layer5_out[108] | layer5_out[107];
     layer6_out[472] <= ~layer5_out[1168];
     layer6_out[473] <= layer5_out[488];
     layer6_out[474] <= ~(layer5_out[1349] & layer5_out[1350]);
     layer6_out[475] <= ~layer5_out[165];
     layer6_out[476] <= ~layer5_out[1459];
     layer6_out[477] <= layer5_out[864] | layer5_out[865];
     layer6_out[478] <= ~(layer5_out[1427] | layer5_out[1428]);
     layer6_out[479] <= layer5_out[944] & ~layer5_out[945];
     layer6_out[480] <= layer5_out[145];
     layer6_out[481] <= layer5_out[328];
     layer6_out[482] <= ~layer5_out[1065];
     layer6_out[483] <= ~layer5_out[1140];
     layer6_out[484] <= ~layer5_out[1403] | layer5_out[1402];
     layer6_out[485] <= ~(layer5_out[166] ^ layer5_out[167]);
     layer6_out[486] <= ~layer5_out[9];
     layer6_out[487] <= ~layer5_out[653] | layer5_out[654];
     layer6_out[488] <= layer5_out[487] & ~layer5_out[486];
     layer6_out[489] <= layer5_out[565];
     layer6_out[490] <= layer5_out[882];
     layer6_out[491] <= layer5_out[162];
     layer6_out[492] <= ~(layer5_out[1375] | layer5_out[1376]);
     layer6_out[493] <= layer5_out[1441] & ~layer5_out[1442];
     layer6_out[494] <= layer5_out[632];
     layer6_out[495] <= ~(layer5_out[847] & layer5_out[848]);
     layer6_out[496] <= layer5_out[96] & ~layer5_out[95];
     layer6_out[497] <= ~layer5_out[1231] | layer5_out[1230];
     layer6_out[498] <= layer5_out[133] ^ layer5_out[134];
     layer6_out[499] <= ~layer5_out[1374];
     layer6_out[500] <= ~layer5_out[187] | layer5_out[186];
     layer6_out[501] <= layer5_out[186];
     layer6_out[502] <= ~(layer5_out[994] | layer5_out[995]);
     layer6_out[503] <= ~layer5_out[1391] | layer5_out[1390];
     layer6_out[504] <= ~layer5_out[766];
     layer6_out[505] <= ~(layer5_out[1049] | layer5_out[1050]);
     layer6_out[506] <= ~layer5_out[1183];
     layer6_out[507] <= layer5_out[522];
     layer6_out[508] <= layer5_out[1225] & ~layer5_out[1224];
     layer6_out[509] <= ~layer5_out[706];
     layer6_out[510] <= ~(layer5_out[1493] | layer5_out[1494]);
     layer6_out[511] <= ~layer5_out[521] | layer5_out[520];
     layer6_out[512] <= ~layer5_out[620] | layer5_out[621];
     layer6_out[513] <= ~layer5_out[77];
     layer6_out[514] <= ~layer5_out[1084] | layer5_out[1083];
     layer6_out[515] <= ~(layer5_out[1274] ^ layer5_out[1275]);
     layer6_out[516] <= layer5_out[722];
     layer6_out[517] <= layer5_out[424] & ~layer5_out[425];
     layer6_out[518] <= layer5_out[1342] & ~layer5_out[1341];
     layer6_out[519] <= ~layer5_out[664];
     layer6_out[520] <= ~layer5_out[1129];
     layer6_out[521] <= layer5_out[1306] & ~layer5_out[1305];
     layer6_out[522] <= ~layer5_out[1036] | layer5_out[1035];
     layer6_out[523] <= layer5_out[31] & ~layer5_out[32];
     layer6_out[524] <= layer5_out[709] | layer5_out[710];
     layer6_out[525] <= layer5_out[235];
     layer6_out[526] <= ~layer5_out[211];
     layer6_out[527] <= layer5_out[1358];
     layer6_out[528] <= ~layer5_out[531];
     layer6_out[529] <= layer5_out[1418];
     layer6_out[530] <= layer5_out[1198] & ~layer5_out[1199];
     layer6_out[531] <= layer5_out[369] | layer5_out[370];
     layer6_out[532] <= ~(layer5_out[946] & layer5_out[947]);
     layer6_out[533] <= layer5_out[499];
     layer6_out[534] <= ~(layer5_out[1440] & layer5_out[1441]);
     layer6_out[535] <= ~layer5_out[782];
     layer6_out[536] <= ~layer5_out[120] | layer5_out[119];
     layer6_out[537] <= layer5_out[530];
     layer6_out[538] <= ~layer5_out[154];
     layer6_out[539] <= layer5_out[508];
     layer6_out[540] <= ~layer5_out[478];
     layer6_out[541] <= ~layer5_out[287] | layer5_out[286];
     layer6_out[542] <= layer5_out[171] & ~layer5_out[170];
     layer6_out[543] <= ~layer5_out[53];
     layer6_out[544] <= layer5_out[1138];
     layer6_out[545] <= layer5_out[382] & ~layer5_out[381];
     layer6_out[546] <= layer5_out[743] & ~layer5_out[742];
     layer6_out[547] <= layer5_out[1323] | layer5_out[1324];
     layer6_out[548] <= layer5_out[450];
     layer6_out[549] <= layer5_out[1387] | layer5_out[1388];
     layer6_out[550] <= ~layer5_out[35] | layer5_out[36];
     layer6_out[551] <= ~layer5_out[1136];
     layer6_out[552] <= ~layer5_out[719];
     layer6_out[553] <= layer5_out[422] ^ layer5_out[423];
     layer6_out[554] <= layer5_out[984] ^ layer5_out[985];
     layer6_out[555] <= layer5_out[1450] & ~layer5_out[1451];
     layer6_out[556] <= ~layer5_out[920];
     layer6_out[557] <= layer5_out[293] & layer5_out[294];
     layer6_out[558] <= ~layer5_out[837];
     layer6_out[559] <= layer5_out[699];
     layer6_out[560] <= ~layer5_out[1283];
     layer6_out[561] <= layer5_out[752];
     layer6_out[562] <= layer5_out[1346];
     layer6_out[563] <= ~(layer5_out[976] | layer5_out[977]);
     layer6_out[564] <= layer5_out[45] & ~layer5_out[46];
     layer6_out[565] <= ~layer5_out[419] | layer5_out[420];
     layer6_out[566] <= layer5_out[868];
     layer6_out[567] <= ~(layer5_out[512] | layer5_out[513]);
     layer6_out[568] <= layer5_out[1043];
     layer6_out[569] <= ~(layer5_out[259] & layer5_out[260]);
     layer6_out[570] <= layer5_out[1137] ^ layer5_out[1138];
     layer6_out[571] <= ~(layer5_out[1332] | layer5_out[1333]);
     layer6_out[572] <= layer5_out[91] | layer5_out[92];
     layer6_out[573] <= layer5_out[846] ^ layer5_out[847];
     layer6_out[574] <= ~layer5_out[679];
     layer6_out[575] <= layer5_out[393];
     layer6_out[576] <= ~(layer5_out[1089] | layer5_out[1090]);
     layer6_out[577] <= layer5_out[880];
     layer6_out[578] <= ~(layer5_out[714] ^ layer5_out[715]);
     layer6_out[579] <= ~(layer5_out[1202] | layer5_out[1203]);
     layer6_out[580] <= ~layer5_out[722];
     layer6_out[581] <= ~(layer5_out[939] | layer5_out[940]);
     layer6_out[582] <= ~layer5_out[659] | layer5_out[658];
     layer6_out[583] <= ~(layer5_out[1119] ^ layer5_out[1120]);
     layer6_out[584] <= ~layer5_out[734];
     layer6_out[585] <= layer5_out[1147];
     layer6_out[586] <= ~(layer5_out[801] ^ layer5_out[802]);
     layer6_out[587] <= layer5_out[695] & layer5_out[696];
     layer6_out[588] <= ~(layer5_out[1445] | layer5_out[1446]);
     layer6_out[589] <= layer5_out[410];
     layer6_out[590] <= ~(layer5_out[849] ^ layer5_out[850]);
     layer6_out[591] <= ~(layer5_out[845] | layer5_out[846]);
     layer6_out[592] <= ~layer5_out[1365];
     layer6_out[593] <= layer5_out[935];
     layer6_out[594] <= layer5_out[358] ^ layer5_out[359];
     layer6_out[595] <= layer5_out[1046];
     layer6_out[596] <= layer5_out[1320];
     layer6_out[597] <= ~layer5_out[1132] | layer5_out[1131];
     layer6_out[598] <= ~(layer5_out[1095] & layer5_out[1096]);
     layer6_out[599] <= ~layer5_out[1236] | layer5_out[1235];
     layer6_out[600] <= layer5_out[1425];
     layer6_out[601] <= ~(layer5_out[732] & layer5_out[733]);
     layer6_out[602] <= layer5_out[1081];
     layer6_out[603] <= layer5_out[924];
     layer6_out[604] <= layer5_out[39] | layer5_out[40];
     layer6_out[605] <= layer5_out[54];
     layer6_out[606] <= ~(layer5_out[1130] | layer5_out[1131]);
     layer6_out[607] <= layer5_out[704] ^ layer5_out[705];
     layer6_out[608] <= layer5_out[337];
     layer6_out[609] <= ~(layer5_out[316] | layer5_out[317]);
     layer6_out[610] <= layer5_out[1288] & ~layer5_out[1287];
     layer6_out[611] <= 1'b0;
     layer6_out[612] <= layer5_out[398];
     layer6_out[613] <= layer5_out[518];
     layer6_out[614] <= ~layer5_out[1306];
     layer6_out[615] <= layer5_out[334];
     layer6_out[616] <= layer5_out[1337] & ~layer5_out[1338];
     layer6_out[617] <= ~layer5_out[1088] | layer5_out[1089];
     layer6_out[618] <= layer5_out[244];
     layer6_out[619] <= ~layer5_out[323] | layer5_out[322];
     layer6_out[620] <= layer5_out[860] & layer5_out[861];
     layer6_out[621] <= layer5_out[653];
     layer6_out[622] <= ~(layer5_out[497] | layer5_out[498]);
     layer6_out[623] <= ~layer5_out[879];
     layer6_out[624] <= layer5_out[1245] ^ layer5_out[1246];
     layer6_out[625] <= ~layer5_out[1274];
     layer6_out[626] <= layer5_out[677] | layer5_out[678];
     layer6_out[627] <= ~layer5_out[355];
     layer6_out[628] <= layer5_out[423] & ~layer5_out[424];
     layer6_out[629] <= ~layer5_out[964];
     layer6_out[630] <= layer5_out[1301] | layer5_out[1302];
     layer6_out[631] <= ~(layer5_out[676] | layer5_out[677]);
     layer6_out[632] <= layer5_out[1318] & ~layer5_out[1317];
     layer6_out[633] <= ~layer5_out[361];
     layer6_out[634] <= ~layer5_out[544];
     layer6_out[635] <= ~layer5_out[925];
     layer6_out[636] <= ~layer5_out[549];
     layer6_out[637] <= ~layer5_out[588];
     layer6_out[638] <= ~layer5_out[1027];
     layer6_out[639] <= ~layer5_out[709];
     layer6_out[640] <= ~(layer5_out[1252] ^ layer5_out[1253]);
     layer6_out[641] <= layer5_out[1279];
     layer6_out[642] <= layer5_out[686] & layer5_out[687];
     layer6_out[643] <= ~(layer5_out[456] | layer5_out[457]);
     layer6_out[644] <= ~layer5_out[1483];
     layer6_out[645] <= layer5_out[886] & layer5_out[887];
     layer6_out[646] <= layer5_out[185];
     layer6_out[647] <= ~layer5_out[66];
     layer6_out[648] <= layer5_out[522] & ~layer5_out[523];
     layer6_out[649] <= ~layer5_out[1449];
     layer6_out[650] <= ~layer5_out[10] | layer5_out[11];
     layer6_out[651] <= layer5_out[934] & ~layer5_out[933];
     layer6_out[652] <= ~layer5_out[864];
     layer6_out[653] <= layer5_out[800] | layer5_out[801];
     layer6_out[654] <= ~layer5_out[1123] | layer5_out[1124];
     layer6_out[655] <= layer5_out[679] & layer5_out[680];
     layer6_out[656] <= layer5_out[755] | layer5_out[756];
     layer6_out[657] <= ~layer5_out[1039] | layer5_out[1038];
     layer6_out[658] <= ~layer5_out[273] | layer5_out[274];
     layer6_out[659] <= ~(layer5_out[931] ^ layer5_out[932]);
     layer6_out[660] <= ~layer5_out[195] | layer5_out[194];
     layer6_out[661] <= ~layer5_out[512];
     layer6_out[662] <= layer5_out[1398] ^ layer5_out[1399];
     layer6_out[663] <= ~layer5_out[88];
     layer6_out[664] <= layer5_out[1345];
     layer6_out[665] <= ~layer5_out[1185] | layer5_out[1186];
     layer6_out[666] <= layer5_out[1321];
     layer6_out[667] <= layer5_out[770] | layer5_out[771];
     layer6_out[668] <= ~(layer5_out[117] ^ layer5_out[118]);
     layer6_out[669] <= layer5_out[21] & ~layer5_out[20];
     layer6_out[670] <= ~(layer5_out[470] ^ layer5_out[471]);
     layer6_out[671] <= ~layer5_out[241];
     layer6_out[672] <= layer5_out[528];
     layer6_out[673] <= ~layer5_out[350];
     layer6_out[674] <= ~layer5_out[936];
     layer6_out[675] <= ~layer5_out[907];
     layer6_out[676] <= layer5_out[469] ^ layer5_out[470];
     layer6_out[677] <= layer5_out[596] & ~layer5_out[595];
     layer6_out[678] <= ~layer5_out[49];
     layer6_out[679] <= ~layer5_out[965] | layer5_out[966];
     layer6_out[680] <= ~layer5_out[265] | layer5_out[264];
     layer6_out[681] <= layer5_out[209];
     layer6_out[682] <= ~layer5_out[838];
     layer6_out[683] <= layer5_out[86] & ~layer5_out[85];
     layer6_out[684] <= layer5_out[1267];
     layer6_out[685] <= ~(layer5_out[1234] & layer5_out[1235]);
     layer6_out[686] <= layer5_out[446] ^ layer5_out[447];
     layer6_out[687] <= 1'b1;
     layer6_out[688] <= ~(layer5_out[1472] & layer5_out[1473]);
     layer6_out[689] <= ~(layer5_out[1003] ^ layer5_out[1004]);
     layer6_out[690] <= ~layer5_out[1269];
     layer6_out[691] <= ~layer5_out[635] | layer5_out[636];
     layer6_out[692] <= ~layer5_out[540];
     layer6_out[693] <= layer5_out[448] & ~layer5_out[449];
     layer6_out[694] <= ~layer5_out[201];
     layer6_out[695] <= ~layer5_out[266] | layer5_out[267];
     layer6_out[696] <= layer5_out[764] ^ layer5_out[765];
     layer6_out[697] <= ~layer5_out[49];
     layer6_out[698] <= layer5_out[175] & ~layer5_out[176];
     layer6_out[699] <= ~layer5_out[459];
     layer6_out[700] <= ~layer5_out[495] | layer5_out[494];
     layer6_out[701] <= ~layer5_out[676];
     layer6_out[702] <= 1'b0;
     layer6_out[703] <= layer5_out[21] & ~layer5_out[22];
     layer6_out[704] <= layer5_out[1071] ^ layer5_out[1072];
     layer6_out[705] <= ~layer5_out[902];
     layer6_out[706] <= layer5_out[1164];
     layer6_out[707] <= layer5_out[229];
     layer6_out[708] <= ~layer5_out[439];
     layer6_out[709] <= layer5_out[120] ^ layer5_out[121];
     layer6_out[710] <= ~(layer5_out[1158] & layer5_out[1159]);
     layer6_out[711] <= layer5_out[1297] | layer5_out[1298];
     layer6_out[712] <= layer5_out[990];
     layer6_out[713] <= 1'b0;
     layer6_out[714] <= layer5_out[1370] ^ layer5_out[1371];
     layer6_out[715] <= layer5_out[762];
     layer6_out[716] <= ~(layer5_out[1453] ^ layer5_out[1454]);
     layer6_out[717] <= layer5_out[1044] | layer5_out[1045];
     layer6_out[718] <= ~layer5_out[675];
     layer6_out[719] <= layer5_out[861] ^ layer5_out[862];
     layer6_out[720] <= ~(layer5_out[479] | layer5_out[480]);
     layer6_out[721] <= ~layer5_out[725] | layer5_out[726];
     layer6_out[722] <= ~layer5_out[83];
     layer6_out[723] <= layer5_out[956] & ~layer5_out[957];
     layer6_out[724] <= ~layer5_out[1058];
     layer6_out[725] <= ~(layer5_out[102] ^ layer5_out[103]);
     layer6_out[726] <= layer5_out[852] & layer5_out[853];
     layer6_out[727] <= ~(layer5_out[607] & layer5_out[608]);
     layer6_out[728] <= layer5_out[665];
     layer6_out[729] <= layer5_out[938] & layer5_out[939];
     layer6_out[730] <= ~layer5_out[1049];
     layer6_out[731] <= layer5_out[123];
     layer6_out[732] <= layer5_out[283];
     layer6_out[733] <= ~layer5_out[309] | layer5_out[308];
     layer6_out[734] <= ~layer5_out[106];
     layer6_out[735] <= ~(layer5_out[105] & layer5_out[106]);
     layer6_out[736] <= layer5_out[890];
     layer6_out[737] <= ~layer5_out[962] | layer5_out[961];
     layer6_out[738] <= ~layer5_out[1272];
     layer6_out[739] <= layer5_out[350] | layer5_out[351];
     layer6_out[740] <= ~layer5_out[866];
     layer6_out[741] <= ~layer5_out[811];
     layer6_out[742] <= layer5_out[170];
     layer6_out[743] <= ~(layer5_out[57] | layer5_out[58]);
     layer6_out[744] <= ~(layer5_out[561] ^ layer5_out[562]);
     layer6_out[745] <= layer5_out[283] & ~layer5_out[284];
     layer6_out[746] <= ~layer5_out[1042];
     layer6_out[747] <= ~layer5_out[179];
     layer6_out[748] <= ~layer5_out[1426];
     layer6_out[749] <= ~layer5_out[1048];
     layer6_out[750] <= layer5_out[1035] & ~layer5_out[1034];
     layer6_out[751] <= ~layer5_out[905] | layer5_out[906];
     layer6_out[752] <= ~layer5_out[1101];
     layer6_out[753] <= layer5_out[157] & ~layer5_out[156];
     layer6_out[754] <= layer5_out[501];
     layer6_out[755] <= ~(layer5_out[292] ^ layer5_out[293]);
     layer6_out[756] <= layer5_out[1099];
     layer6_out[757] <= ~layer5_out[1151];
     layer6_out[758] <= layer5_out[123] ^ layer5_out[124];
     layer6_out[759] <= layer5_out[600];
     layer6_out[760] <= ~layer5_out[268];
     layer6_out[761] <= layer5_out[1212];
     layer6_out[762] <= layer5_out[143];
     layer6_out[763] <= layer5_out[959] | layer5_out[960];
     layer6_out[764] <= layer5_out[502] ^ layer5_out[503];
     layer6_out[765] <= layer5_out[726];
     layer6_out[766] <= layer5_out[448];
     layer6_out[767] <= layer5_out[536];
     layer6_out[768] <= ~layer5_out[1421];
     layer6_out[769] <= layer5_out[274] | layer5_out[275];
     layer6_out[770] <= layer5_out[356] & ~layer5_out[357];
     layer6_out[771] <= ~layer5_out[1005];
     layer6_out[772] <= ~layer5_out[998];
     layer6_out[773] <= ~layer5_out[388];
     layer6_out[774] <= layer5_out[1391];
     layer6_out[775] <= layer5_out[1032];
     layer6_out[776] <= ~layer5_out[1001] | layer5_out[1000];
     layer6_out[777] <= ~(layer5_out[1355] & layer5_out[1356]);
     layer6_out[778] <= ~layer5_out[405];
     layer6_out[779] <= ~(layer5_out[162] ^ layer5_out[163]);
     layer6_out[780] <= layer5_out[1161];
     layer6_out[781] <= ~(layer5_out[636] | layer5_out[637]);
     layer6_out[782] <= ~(layer5_out[242] & layer5_out[243]);
     layer6_out[783] <= ~layer5_out[1356];
     layer6_out[784] <= ~layer5_out[36];
     layer6_out[785] <= ~layer5_out[373];
     layer6_out[786] <= ~(layer5_out[432] ^ layer5_out[433]);
     layer6_out[787] <= ~layer5_out[112];
     layer6_out[788] <= ~layer5_out[1339];
     layer6_out[789] <= layer5_out[1020];
     layer6_out[790] <= layer5_out[1494];
     layer6_out[791] <= ~layer5_out[164];
     layer6_out[792] <= ~layer5_out[1465];
     layer6_out[793] <= layer5_out[1014];
     layer6_out[794] <= layer5_out[1013];
     layer6_out[795] <= ~(layer5_out[1105] | layer5_out[1106]);
     layer6_out[796] <= ~(layer5_out[627] & layer5_out[628]);
     layer6_out[797] <= layer5_out[1321] & ~layer5_out[1322];
     layer6_out[798] <= ~(layer5_out[637] ^ layer5_out[638]);
     layer6_out[799] <= layer5_out[959];
     layer6_out[800] <= layer5_out[594];
     layer6_out[801] <= layer5_out[1291];
     layer6_out[802] <= ~layer5_out[471];
     layer6_out[803] <= layer5_out[729] | layer5_out[730];
     layer6_out[804] <= layer5_out[473] ^ layer5_out[474];
     layer6_out[805] <= ~layer5_out[904] | layer5_out[903];
     layer6_out[806] <= layer5_out[1143];
     layer6_out[807] <= layer5_out[597] & layer5_out[598];
     layer6_out[808] <= ~layer5_out[1108];
     layer6_out[809] <= layer5_out[562];
     layer6_out[810] <= layer5_out[1462];
     layer6_out[811] <= layer5_out[426];
     layer6_out[812] <= layer5_out[1057] | layer5_out[1058];
     layer6_out[813] <= ~(layer5_out[977] ^ layer5_out[978]);
     layer6_out[814] <= layer5_out[137] | layer5_out[138];
     layer6_out[815] <= 1'b0;
     layer6_out[816] <= layer5_out[323] & layer5_out[324];
     layer6_out[817] <= ~(layer5_out[1141] ^ layer5_out[1142]);
     layer6_out[818] <= layer5_out[51];
     layer6_out[819] <= ~layer5_out[1302];
     layer6_out[820] <= ~layer5_out[1077];
     layer6_out[821] <= ~layer5_out[610];
     layer6_out[822] <= ~(layer5_out[124] | layer5_out[125]);
     layer6_out[823] <= ~layer5_out[816];
     layer6_out[824] <= layer5_out[616];
     layer6_out[825] <= ~layer5_out[1159];
     layer6_out[826] <= ~layer5_out[1490] | layer5_out[1491];
     layer6_out[827] <= layer5_out[454] ^ layer5_out[455];
     layer6_out[828] <= layer5_out[1432];
     layer6_out[829] <= layer5_out[1458];
     layer6_out[830] <= layer5_out[579] & ~layer5_out[578];
     layer6_out[831] <= ~layer5_out[344] | layer5_out[345];
     layer6_out[832] <= ~layer5_out[302] | layer5_out[303];
     layer6_out[833] <= layer5_out[689];
     layer6_out[834] <= ~layer5_out[172];
     layer6_out[835] <= layer5_out[595];
     layer6_out[836] <= layer5_out[1404];
     layer6_out[837] <= layer5_out[165];
     layer6_out[838] <= ~(layer5_out[1354] & layer5_out[1355]);
     layer6_out[839] <= ~(layer5_out[15] & layer5_out[16]);
     layer6_out[840] <= ~layer5_out[922];
     layer6_out[841] <= layer5_out[876] & layer5_out[877];
     layer6_out[842] <= ~layer5_out[981];
     layer6_out[843] <= ~(layer5_out[1448] ^ layer5_out[1449]);
     layer6_out[844] <= layer5_out[257] & ~layer5_out[258];
     layer6_out[845] <= ~(layer5_out[696] | layer5_out[697]);
     layer6_out[846] <= ~(layer5_out[284] ^ layer5_out[285]);
     layer6_out[847] <= layer5_out[1191] & layer5_out[1192];
     layer6_out[848] <= layer5_out[1111];
     layer6_out[849] <= ~(layer5_out[281] | layer5_out[282]);
     layer6_out[850] <= ~layer5_out[1082] | layer5_out[1083];
     layer6_out[851] <= layer5_out[1222];
     layer6_out[852] <= layer5_out[62];
     layer6_out[853] <= ~(layer5_out[1056] ^ layer5_out[1057]);
     layer6_out[854] <= layer5_out[798];
     layer6_out[855] <= layer5_out[1218] | layer5_out[1219];
     layer6_out[856] <= ~layer5_out[573];
     layer6_out[857] <= ~(layer5_out[1438] | layer5_out[1439]);
     layer6_out[858] <= layer5_out[871] & ~layer5_out[872];
     layer6_out[859] <= layer5_out[570] & ~layer5_out[571];
     layer6_out[860] <= ~(layer5_out[368] | layer5_out[369]);
     layer6_out[861] <= layer5_out[380] | layer5_out[381];
     layer6_out[862] <= layer5_out[560];
     layer6_out[863] <= layer5_out[682] & ~layer5_out[681];
     layer6_out[864] <= layer5_out[1097];
     layer6_out[865] <= ~(layer5_out[139] | layer5_out[140]);
     layer6_out[866] <= layer5_out[721];
     layer6_out[867] <= ~layer5_out[660] | layer5_out[661];
     layer6_out[868] <= ~(layer5_out[1327] & layer5_out[1328]);
     layer6_out[869] <= layer5_out[141];
     layer6_out[870] <= layer5_out[840] ^ layer5_out[841];
     layer6_out[871] <= ~layer5_out[203] | layer5_out[202];
     layer6_out[872] <= layer5_out[1418] | layer5_out[1419];
     layer6_out[873] <= layer5_out[387] & ~layer5_out[386];
     layer6_out[874] <= layer5_out[1103];
     layer6_out[875] <= ~layer5_out[1332];
     layer6_out[876] <= layer5_out[1228] | layer5_out[1229];
     layer6_out[877] <= layer5_out[357];
     layer6_out[878] <= layer5_out[1443] & ~layer5_out[1442];
     layer6_out[879] <= layer5_out[484] | layer5_out[485];
     layer6_out[880] <= ~(layer5_out[1178] & layer5_out[1179]);
     layer6_out[881] <= layer5_out[19] | layer5_out[20];
     layer6_out[882] <= ~layer5_out[615];
     layer6_out[883] <= layer5_out[220];
     layer6_out[884] <= ~layer5_out[543];
     layer6_out[885] <= ~layer5_out[1262];
     layer6_out[886] <= ~(layer5_out[1362] & layer5_out[1363]);
     layer6_out[887] <= ~layer5_out[808] | layer5_out[809];
     layer6_out[888] <= ~layer5_out[1411];
     layer6_out[889] <= ~(layer5_out[1145] | layer5_out[1146]);
     layer6_out[890] <= ~(layer5_out[480] ^ layer5_out[481]);
     layer6_out[891] <= ~(layer5_out[1104] & layer5_out[1105]);
     layer6_out[892] <= ~(layer5_out[654] | layer5_out[655]);
     layer6_out[893] <= layer5_out[1471];
     layer6_out[894] <= layer5_out[393] & ~layer5_out[392];
     layer6_out[895] <= layer5_out[59] & layer5_out[60];
     layer6_out[896] <= layer5_out[348] & ~layer5_out[349];
     layer6_out[897] <= layer5_out[1293] & ~layer5_out[1294];
     layer6_out[898] <= ~layer5_out[413];
     layer6_out[899] <= ~(layer5_out[1126] & layer5_out[1127]);
     layer6_out[900] <= layer5_out[4];
     layer6_out[901] <= ~layer5_out[576];
     layer6_out[902] <= ~layer5_out[1239];
     layer6_out[903] <= ~layer5_out[747];
     layer6_out[904] <= layer5_out[736] ^ layer5_out[737];
     layer6_out[905] <= layer5_out[706];
     layer6_out[906] <= layer5_out[651];
     layer6_out[907] <= ~(layer5_out[1009] | layer5_out[1010]);
     layer6_out[908] <= layer5_out[812] & layer5_out[813];
     layer6_out[909] <= layer5_out[1113];
     layer6_out[910] <= layer5_out[61] & ~layer5_out[60];
     layer6_out[911] <= ~(layer5_out[1209] | layer5_out[1210]);
     layer6_out[912] <= ~layer5_out[539];
     layer6_out[913] <= layer5_out[694] & layer5_out[695];
     layer6_out[914] <= layer5_out[63] & ~layer5_out[64];
     layer6_out[915] <= ~(layer5_out[144] ^ layer5_out[145]);
     layer6_out[916] <= layer5_out[500] | layer5_out[501];
     layer6_out[917] <= ~layer5_out[1208] | layer5_out[1209];
     layer6_out[918] <= layer5_out[340];
     layer6_out[919] <= ~(layer5_out[546] & layer5_out[547]);
     layer6_out[920] <= ~(layer5_out[495] ^ layer5_out[496]);
     layer6_out[921] <= layer5_out[371];
     layer6_out[922] <= ~(layer5_out[1187] ^ layer5_out[1188]);
     layer6_out[923] <= ~layer5_out[216];
     layer6_out[924] <= layer5_out[0] ^ layer5_out[1];
     layer6_out[925] <= layer5_out[1172] & ~layer5_out[1173];
     layer6_out[926] <= layer5_out[1361] | layer5_out[1362];
     layer6_out[927] <= layer5_out[1094];
     layer6_out[928] <= ~layer5_out[414];
     layer6_out[929] <= ~(layer5_out[1407] | layer5_out[1408]);
     layer6_out[930] <= ~(layer5_out[1289] | layer5_out[1290]);
     layer6_out[931] <= layer5_out[276] ^ layer5_out[277];
     layer6_out[932] <= layer5_out[73] ^ layer5_out[74];
     layer6_out[933] <= ~(layer5_out[84] & layer5_out[85]);
     layer6_out[934] <= ~layer5_out[1052];
     layer6_out[935] <= ~layer5_out[1249];
     layer6_out[936] <= ~layer5_out[745];
     layer6_out[937] <= layer5_out[533] ^ layer5_out[534];
     layer6_out[938] <= ~layer5_out[1381];
     layer6_out[939] <= layer5_out[115];
     layer6_out[940] <= ~(layer5_out[482] | layer5_out[483]);
     layer6_out[941] <= layer5_out[1482];
     layer6_out[942] <= ~(layer5_out[515] ^ layer5_out[516]);
     layer6_out[943] <= ~layer5_out[361];
     layer6_out[944] <= ~(layer5_out[222] | layer5_out[223]);
     layer6_out[945] <= layer5_out[55] & layer5_out[56];
     layer6_out[946] <= layer5_out[1256];
     layer6_out[947] <= layer5_out[1491];
     layer6_out[948] <= layer5_out[433] | layer5_out[434];
     layer6_out[949] <= layer5_out[442] & layer5_out[443];
     layer6_out[950] <= ~(layer5_out[1254] ^ layer5_out[1255]);
     layer6_out[951] <= ~layer5_out[1477];
     layer6_out[952] <= ~layer5_out[68] | layer5_out[67];
     layer6_out[953] <= ~(layer5_out[34] ^ layer5_out[35]);
     layer6_out[954] <= layer5_out[642] & ~layer5_out[641];
     layer6_out[955] <= ~layer5_out[989] | layer5_out[988];
     layer6_out[956] <= ~(layer5_out[1377] | layer5_out[1378]);
     layer6_out[957] <= ~layer5_out[331];
     layer6_out[958] <= layer5_out[1050];
     layer6_out[959] <= ~(layer5_out[1153] | layer5_out[1154]);
     layer6_out[960] <= ~layer5_out[119] | layer5_out[118];
     layer6_out[961] <= ~layer5_out[1070];
     layer6_out[962] <= layer5_out[1002];
     layer6_out[963] <= layer5_out[1414] & ~layer5_out[1415];
     layer6_out[964] <= ~layer5_out[1219] | layer5_out[1220];
     layer6_out[965] <= ~layer5_out[121];
     layer6_out[966] <= ~layer5_out[588];
     layer6_out[967] <= layer5_out[23] & layer5_out[24];
     layer6_out[968] <= layer5_out[80] | layer5_out[81];
     layer6_out[969] <= ~layer5_out[383];
     layer6_out[970] <= layer5_out[1404];
     layer6_out[971] <= ~(layer5_out[1275] ^ layer5_out[1276]);
     layer6_out[972] <= ~(layer5_out[307] ^ layer5_out[308]);
     layer6_out[973] <= layer5_out[376];
     layer6_out[974] <= ~layer5_out[304];
     layer6_out[975] <= layer5_out[540];
     layer6_out[976] <= ~(layer5_out[474] ^ layer5_out[475]);
     layer6_out[977] <= layer5_out[771] ^ layer5_out[772];
     layer6_out[978] <= layer5_out[1090] & layer5_out[1091];
     layer6_out[979] <= ~(layer5_out[287] & layer5_out[288]);
     layer6_out[980] <= ~(layer5_out[901] & layer5_out[902]);
     layer6_out[981] <= ~(layer5_out[250] ^ layer5_out[251]);
     layer6_out[982] <= layer5_out[252];
     layer6_out[983] <= ~layer5_out[1193];
     layer6_out[984] <= ~layer5_out[1393];
     layer6_out[985] <= ~layer5_out[1019];
     layer6_out[986] <= ~(layer5_out[50] | layer5_out[51]);
     layer6_out[987] <= layer5_out[616] & ~layer5_out[617];
     layer6_out[988] <= layer5_out[1144] | layer5_out[1145];
     layer6_out[989] <= ~layer5_out[271];
     layer6_out[990] <= ~layer5_out[599];
     layer6_out[991] <= layer5_out[1054];
     layer6_out[992] <= ~layer5_out[159];
     layer6_out[993] <= ~layer5_out[885] | layer5_out[884];
     layer6_out[994] <= layer5_out[606];
     layer6_out[995] <= layer5_out[630];
     layer6_out[996] <= ~(layer5_out[338] ^ layer5_out[339]);
     layer6_out[997] <= layer5_out[138] ^ layer5_out[139];
     layer6_out[998] <= ~layer5_out[1440] | layer5_out[1439];
     layer6_out[999] <= layer5_out[1424];
     layer6_out[1000] <= ~layer5_out[457];
     layer6_out[1001] <= ~layer5_out[542];
     layer6_out[1002] <= ~layer5_out[618] | layer5_out[619];
     layer6_out[1003] <= ~layer5_out[29];
     layer6_out[1004] <= ~(layer5_out[822] ^ layer5_out[823]);
     layer6_out[1005] <= ~layer5_out[1396];
     layer6_out[1006] <= layer5_out[30];
     layer6_out[1007] <= layer5_out[182] & layer5_out[183];
     layer6_out[1008] <= layer5_out[913] & ~layer5_out[914];
     layer6_out[1009] <= layer5_out[1211] & ~layer5_out[1210];
     layer6_out[1010] <= ~layer5_out[551];
     layer6_out[1011] <= ~layer5_out[662] | layer5_out[663];
     layer6_out[1012] <= layer5_out[190];
     layer6_out[1013] <= layer5_out[153] & ~layer5_out[154];
     layer6_out[1014] <= ~(layer5_out[190] & layer5_out[191]);
     layer6_out[1015] <= layer5_out[146] & ~layer5_out[147];
     layer6_out[1016] <= ~(layer5_out[405] | layer5_out[406]);
     layer6_out[1017] <= ~(layer5_out[1367] ^ layer5_out[1368]);
     layer6_out[1018] <= ~(layer5_out[167] | layer5_out[168]);
     layer6_out[1019] <= layer5_out[336] ^ layer5_out[337];
     layer6_out[1020] <= ~layer5_out[1375];
     layer6_out[1021] <= ~layer5_out[543] | layer5_out[542];
     layer6_out[1022] <= 1'b0;
     layer6_out[1023] <= ~(layer5_out[1399] & layer5_out[1400]);
     layer6_out[1024] <= layer5_out[100] & ~layer5_out[99];
     layer6_out[1025] <= ~layer5_out[295];
     layer6_out[1026] <= ~(layer5_out[2] & layer5_out[3]);
     layer6_out[1027] <= ~layer5_out[343];
     layer6_out[1028] <= ~layer5_out[569];
     layer6_out[1029] <= ~layer5_out[1423];
     layer6_out[1030] <= layer5_out[213] & ~layer5_out[212];
     layer6_out[1031] <= layer5_out[1039] & ~layer5_out[1040];
     layer6_out[1032] <= layer5_out[489];
     layer6_out[1033] <= ~(layer5_out[272] ^ layer5_out[273]);
     layer6_out[1034] <= layer5_out[481] & layer5_out[482];
     layer6_out[1035] <= layer5_out[1022] & ~layer5_out[1021];
     layer6_out[1036] <= layer5_out[94];
     layer6_out[1037] <= layer5_out[1214];
     layer6_out[1038] <= layer5_out[1028];
     layer6_out[1039] <= layer5_out[567] & ~layer5_out[568];
     layer6_out[1040] <= layer5_out[727];
     layer6_out[1041] <= layer5_out[755];
     layer6_out[1042] <= ~layer5_out[253];
     layer6_out[1043] <= layer5_out[874] ^ layer5_out[875];
     layer6_out[1044] <= ~layer5_out[1134];
     layer6_out[1045] <= layer5_out[577] | layer5_out[578];
     layer6_out[1046] <= ~layer5_out[788];
     layer6_out[1047] <= layer5_out[823];
     layer6_out[1048] <= layer5_out[995] | layer5_out[996];
     layer6_out[1049] <= ~(layer5_out[912] & layer5_out[913]);
     layer6_out[1050] <= ~(layer5_out[767] & layer5_out[768]);
     layer6_out[1051] <= layer5_out[78];
     layer6_out[1052] <= ~layer5_out[93];
     layer6_out[1053] <= layer5_out[6] & ~layer5_out[7];
     layer6_out[1054] <= layer5_out[1373];
     layer6_out[1055] <= ~layer5_out[174] | layer5_out[175];
     layer6_out[1056] <= ~layer5_out[1187];
     layer6_out[1057] <= layer5_out[704] & ~layer5_out[703];
     layer6_out[1058] <= ~layer5_out[192] | layer5_out[191];
     layer6_out[1059] <= ~layer5_out[884];
     layer6_out[1060] <= layer5_out[960];
     layer6_out[1061] <= layer5_out[24] | layer5_out[25];
     layer6_out[1062] <= layer5_out[646] & ~layer5_out[647];
     layer6_out[1063] <= ~layer5_out[1398];
     layer6_out[1064] <= ~layer5_out[649];
     layer6_out[1065] <= ~(layer5_out[893] ^ layer5_out[894]);
     layer6_out[1066] <= ~(layer5_out[489] & layer5_out[490]);
     layer6_out[1067] <= ~(layer5_out[839] ^ layer5_out[840]);
     layer6_out[1068] <= ~(layer5_out[127] & layer5_out[128]);
     layer6_out[1069] <= layer5_out[1217] & ~layer5_out[1216];
     layer6_out[1070] <= ~layer5_out[1156];
     layer6_out[1071] <= ~layer5_out[1087];
     layer6_out[1072] <= ~layer5_out[1118];
     layer6_out[1073] <= ~layer5_out[152];
     layer6_out[1074] <= layer5_out[215] | layer5_out[216];
     layer6_out[1075] <= ~layer5_out[204];
     layer6_out[1076] <= ~layer5_out[1137];
     layer6_out[1077] <= ~layer5_out[181];
     layer6_out[1078] <= ~(layer5_out[559] | layer5_out[560]);
     layer6_out[1079] <= layer5_out[1148];
     layer6_out[1080] <= layer5_out[206] & layer5_out[207];
     layer6_out[1081] <= layer5_out[898] ^ layer5_out[899];
     layer6_out[1082] <= layer5_out[558];
     layer6_out[1083] <= ~layer5_out[1470];
     layer6_out[1084] <= layer5_out[1103] ^ layer5_out[1104];
     layer6_out[1085] <= ~(layer5_out[1415] & layer5_out[1416]);
     layer6_out[1086] <= ~layer5_out[1310];
     layer6_out[1087] <= ~layer5_out[935];
     layer6_out[1088] <= ~(layer5_out[201] & layer5_out[202]);
     layer6_out[1089] <= layer5_out[628] & layer5_out[629];
     layer6_out[1090] <= layer5_out[1476] & ~layer5_out[1475];
     layer6_out[1091] <= layer5_out[1372];
     layer6_out[1092] <= ~layer5_out[313];
     layer6_out[1093] <= ~layer5_out[421];
     layer6_out[1094] <= layer5_out[667] & ~layer5_out[668];
     layer6_out[1095] <= ~layer5_out[1110] | layer5_out[1109];
     layer6_out[1096] <= ~layer5_out[1334] | layer5_out[1335];
     layer6_out[1097] <= layer5_out[774];
     layer6_out[1098] <= ~layer5_out[280] | layer5_out[281];
     layer6_out[1099] <= ~layer5_out[911];
     layer6_out[1100] <= ~layer5_out[1329];
     layer6_out[1101] <= 1'b1;
     layer6_out[1102] <= ~(layer5_out[1366] ^ layer5_out[1367]);
     layer6_out[1103] <= layer5_out[1033];
     layer6_out[1104] <= layer5_out[1316];
     layer6_out[1105] <= layer5_out[768];
     layer6_out[1106] <= layer5_out[366];
     layer6_out[1107] <= layer5_out[9];
     layer6_out[1108] <= ~layer5_out[672];
     layer6_out[1109] <= layer5_out[581];
     layer6_out[1110] <= layer5_out[509];
     layer6_out[1111] <= layer5_out[453] & layer5_out[454];
     layer6_out[1112] <= ~layer5_out[919];
     layer6_out[1113] <= layer5_out[772] ^ layer5_out[773];
     layer6_out[1114] <= layer5_out[72] & ~layer5_out[71];
     layer6_out[1115] <= ~layer5_out[156] | layer5_out[155];
     layer6_out[1116] <= layer5_out[866];
     layer6_out[1117] <= layer5_out[937] | layer5_out[938];
     layer6_out[1118] <= layer5_out[55];
     layer6_out[1119] <= layer5_out[1170] & ~layer5_out[1171];
     layer6_out[1120] <= ~layer5_out[1264];
     layer6_out[1121] <= layer5_out[1107];
     layer6_out[1122] <= ~layer5_out[343];
     layer6_out[1123] <= layer5_out[1036] & layer5_out[1037];
     layer6_out[1124] <= layer5_out[1198];
     layer6_out[1125] <= layer5_out[1279];
     layer6_out[1126] <= layer5_out[1127] | layer5_out[1128];
     layer6_out[1127] <= ~(layer5_out[926] ^ layer5_out[927]);
     layer6_out[1128] <= layer5_out[585];
     layer6_out[1129] <= ~layer5_out[496];
     layer6_out[1130] <= layer5_out[79] & ~layer5_out[80];
     layer6_out[1131] <= ~(layer5_out[126] | layer5_out[127]);
     layer6_out[1132] <= layer5_out[437];
     layer6_out[1133] <= layer5_out[525];
     layer6_out[1134] <= ~layer5_out[291];
     layer6_out[1135] <= ~layer5_out[1342] | layer5_out[1343];
     layer6_out[1136] <= ~layer5_out[618];
     layer6_out[1137] <= ~layer5_out[345];
     layer6_out[1138] <= layer5_out[929] & ~layer5_out[928];
     layer6_out[1139] <= ~layer5_out[1204] | layer5_out[1205];
     layer6_out[1140] <= ~layer5_out[1174];
     layer6_out[1141] <= layer5_out[1395];
     layer6_out[1142] <= layer5_out[983];
     layer6_out[1143] <= ~layer5_out[1351];
     layer6_out[1144] <= ~layer5_out[90] | layer5_out[91];
     layer6_out[1145] <= layer5_out[821];
     layer6_out[1146] <= layer5_out[1455] ^ layer5_out[1456];
     layer6_out[1147] <= 1'b1;
     layer6_out[1148] <= layer5_out[892] & ~layer5_out[891];
     layer6_out[1149] <= ~layer5_out[818];
     layer6_out[1150] <= layer5_out[1468] ^ layer5_out[1469];
     layer6_out[1151] <= ~(layer5_out[98] | layer5_out[99]);
     layer6_out[1152] <= layer5_out[42] & ~layer5_out[41];
     layer6_out[1153] <= layer5_out[693];
     layer6_out[1154] <= layer5_out[37];
     layer6_out[1155] <= layer5_out[1467];
     layer6_out[1156] <= ~layer5_out[624];
     layer6_out[1157] <= ~layer5_out[778] | layer5_out[779];
     layer6_out[1158] <= layer5_out[261] & layer5_out[262];
     layer6_out[1159] <= layer5_out[858];
     layer6_out[1160] <= ~layer5_out[409];
     layer6_out[1161] <= layer5_out[1495] & layer5_out[1496];
     layer6_out[1162] <= ~(layer5_out[683] | layer5_out[684]);
     layer6_out[1163] <= 1'b1;
     layer6_out[1164] <= layer5_out[443] ^ layer5_out[444];
     layer6_out[1165] <= ~(layer5_out[633] ^ layer5_out[634]);
     layer6_out[1166] <= layer5_out[869] & ~layer5_out[868];
     layer6_out[1167] <= ~(layer5_out[13] | layer5_out[14]);
     layer6_out[1168] <= ~layer5_out[724];
     layer6_out[1169] <= ~(layer5_out[673] & layer5_out[674]);
     layer6_out[1170] <= layer5_out[806];
     layer6_out[1171] <= layer5_out[1238] & ~layer5_out[1237];
     layer6_out[1172] <= ~layer5_out[853] | layer5_out[854];
     layer6_out[1173] <= ~layer5_out[780];
     layer6_out[1174] <= ~(layer5_out[104] & layer5_out[105]);
     layer6_out[1175] <= ~(layer5_out[289] ^ layer5_out[290]);
     layer6_out[1176] <= ~layer5_out[872] | layer5_out[873];
     layer6_out[1177] <= layer5_out[854] ^ layer5_out[855];
     layer6_out[1178] <= ~layer5_out[389];
     layer6_out[1179] <= layer5_out[587];
     layer6_out[1180] <= layer5_out[1285] | layer5_out[1286];
     layer6_out[1181] <= ~(layer5_out[1401] ^ layer5_out[1402]);
     layer6_out[1182] <= ~layer5_out[668];
     layer6_out[1183] <= ~layer5_out[1173];
     layer6_out[1184] <= ~layer5_out[1409];
     layer6_out[1185] <= layer5_out[680];
     layer6_out[1186] <= layer5_out[757];
     layer6_out[1187] <= ~layer5_out[1380];
     layer6_out[1188] <= ~layer5_out[197];
     layer6_out[1189] <= ~layer5_out[979];
     layer6_out[1190] <= ~layer5_out[603];
     layer6_out[1191] <= ~layer5_out[1191];
     layer6_out[1192] <= layer5_out[915];
     layer6_out[1193] <= layer5_out[1284];
     layer6_out[1194] <= ~layer5_out[797];
     layer6_out[1195] <= layer5_out[1230] & ~layer5_out[1229];
     layer6_out[1196] <= layer5_out[493];
     layer6_out[1197] <= ~layer5_out[1115];
     layer6_out[1198] <= layer5_out[718] & ~layer5_out[717];
     layer6_out[1199] <= layer5_out[1471] | layer5_out[1472];
     layer6_out[1200] <= ~(layer5_out[452] & layer5_out[453]);
     layer6_out[1201] <= ~(layer5_out[619] & layer5_out[620]);
     layer6_out[1202] <= ~layer5_out[687];
     layer6_out[1203] <= ~(layer5_out[327] ^ layer5_out[328]);
     layer6_out[1204] <= layer5_out[224];
     layer6_out[1205] <= ~layer5_out[1363];
     layer6_out[1206] <= layer5_out[1447] & ~layer5_out[1446];
     layer6_out[1207] <= layer5_out[223];
     layer6_out[1208] <= ~(layer5_out[855] | layer5_out[856]);
     layer6_out[1209] <= layer5_out[1436] ^ layer5_out[1437];
     layer6_out[1210] <= ~layer5_out[581] | layer5_out[580];
     layer6_out[1211] <= ~(layer5_out[1040] ^ layer5_out[1041]);
     layer6_out[1212] <= layer5_out[40];
     layer6_out[1213] <= layer5_out[625];
     layer6_out[1214] <= ~layer5_out[1114];
     layer6_out[1215] <= layer5_out[741];
     layer6_out[1216] <= layer5_out[1189];
     layer6_out[1217] <= ~(layer5_out[896] ^ layer5_out[897]);
     layer6_out[1218] <= ~(layer5_out[1345] & layer5_out[1346]);
     layer6_out[1219] <= layer5_out[547];
     layer6_out[1220] <= ~layer5_out[1291] | layer5_out[1292];
     layer6_out[1221] <= layer5_out[1108] & ~layer5_out[1109];
     layer6_out[1222] <= ~layer5_out[1243];
     layer6_out[1223] <= ~layer5_out[639];
     layer6_out[1224] <= ~layer5_out[386];
     layer6_out[1225] <= ~(layer5_out[1309] ^ layer5_out[1310]);
     layer6_out[1226] <= ~layer5_out[149] | layer5_out[150];
     layer6_out[1227] <= ~layer5_out[110];
     layer6_out[1228] <= ~(layer5_out[656] ^ layer5_out[657]);
     layer6_out[1229] <= ~layer5_out[889];
     layer6_out[1230] <= layer5_out[460] & layer5_out[461];
     layer6_out[1231] <= layer5_out[1076];
     layer6_out[1232] <= ~(layer5_out[376] & layer5_out[377]);
     layer6_out[1233] <= ~layer5_out[876] | layer5_out[875];
     layer6_out[1234] <= ~layer5_out[1361] | layer5_out[1360];
     layer6_out[1235] <= ~layer5_out[753] | layer5_out[754];
     layer6_out[1236] <= layer5_out[788] & ~layer5_out[789];
     layer6_out[1237] <= ~(layer5_out[1132] ^ layer5_out[1133]);
     layer6_out[1238] <= layer5_out[1233] & ~layer5_out[1232];
     layer6_out[1239] <= layer5_out[634];
     layer6_out[1240] <= layer5_out[1443];
     layer6_out[1241] <= ~layer5_out[975];
     layer6_out[1242] <= layer5_out[1257];
     layer6_out[1243] <= layer5_out[469];
     layer6_out[1244] <= ~(layer5_out[862] ^ layer5_out[863]);
     layer6_out[1245] <= ~(layer5_out[400] | layer5_out[401]);
     layer6_out[1246] <= layer5_out[844] & ~layer5_out[845];
     layer6_out[1247] <= ~(layer5_out[1244] ^ layer5_out[1245]);
     layer6_out[1248] <= ~layer5_out[1484] | layer5_out[1485];
     layer6_out[1249] <= ~(layer5_out[1053] ^ layer5_out[1054]);
     layer6_out[1250] <= layer5_out[510] & layer5_out[511];
     layer6_out[1251] <= layer5_out[34];
     layer6_out[1252] <= ~layer5_out[1252];
     layer6_out[1253] <= layer5_out[176] ^ layer5_out[177];
     layer6_out[1254] <= ~layer5_out[39];
     layer6_out[1255] <= layer5_out[1265] & ~layer5_out[1266];
     layer6_out[1256] <= layer5_out[1015] & layer5_out[1016];
     layer6_out[1257] <= ~(layer5_out[513] | layer5_out[514]);
     layer6_out[1258] <= layer5_out[916] | layer5_out[917];
     layer6_out[1259] <= ~layer5_out[1263];
     layer6_out[1260] <= ~(layer5_out[1282] ^ layer5_out[1283]);
     layer6_out[1261] <= layer5_out[1369] & layer5_out[1370];
     layer6_out[1262] <= ~(layer5_out[821] | layer5_out[822]);
     layer6_out[1263] <= layer5_out[234];
     layer6_out[1264] <= layer5_out[566] | layer5_out[567];
     layer6_out[1265] <= ~layer5_out[832] | layer5_out[833];
     layer6_out[1266] <= layer5_out[1431];
     layer6_out[1267] <= layer5_out[112] ^ layer5_out[113];
     layer6_out[1268] <= layer5_out[515] & ~layer5_out[514];
     layer6_out[1269] <= layer5_out[414];
     layer6_out[1270] <= layer5_out[827];
     layer6_out[1271] <= ~layer5_out[811];
     layer6_out[1272] <= ~(layer5_out[254] ^ layer5_out[255]);
     layer6_out[1273] <= ~(layer5_out[831] ^ layer5_out[832]);
     layer6_out[1274] <= layer5_out[504] & ~layer5_out[503];
     layer6_out[1275] <= ~layer5_out[1178];
     layer6_out[1276] <= layer5_out[1214] & ~layer5_out[1215];
     layer6_out[1277] <= ~layer5_out[6] | layer5_out[5];
     layer6_out[1278] <= ~layer5_out[1118];
     layer6_out[1279] <= layer5_out[1486] & ~layer5_out[1487];
     layer6_out[1280] <= layer5_out[1091];
     layer6_out[1281] <= ~layer5_out[981] | layer5_out[980];
     layer6_out[1282] <= ~layer5_out[927];
     layer6_out[1283] <= ~layer5_out[13];
     layer6_out[1284] <= layer5_out[390] ^ layer5_out[391];
     layer6_out[1285] <= layer5_out[963];
     layer6_out[1286] <= ~(layer5_out[1169] | layer5_out[1170]);
     layer6_out[1287] <= layer5_out[871];
     layer6_out[1288] <= ~layer5_out[132] | layer5_out[133];
     layer6_out[1289] <= ~layer5_out[912];
     layer6_out[1290] <= layer5_out[556];
     layer6_out[1291] <= ~(layer5_out[942] & layer5_out[943]);
     layer6_out[1292] <= layer5_out[537] & layer5_out[538];
     layer6_out[1293] <= ~(layer5_out[152] | layer5_out[153]);
     layer6_out[1294] <= layer5_out[850] & ~layer5_out[851];
     layer6_out[1295] <= ~layer5_out[1473];
     layer6_out[1296] <= layer5_out[953] | layer5_out[954];
     layer6_out[1297] <= layer5_out[506];
     layer6_out[1298] <= layer5_out[662];
     layer6_out[1299] <= layer5_out[999];
     layer6_out[1300] <= ~(layer5_out[1157] | layer5_out[1158]);
     layer6_out[1301] <= layer5_out[100] ^ layer5_out[101];
     layer6_out[1302] <= layer5_out[608] | layer5_out[609];
     layer6_out[1303] <= layer5_out[650] & ~layer5_out[651];
     layer6_out[1304] <= ~layer5_out[858];
     layer6_out[1305] <= layer5_out[1359];
     layer6_out[1306] <= layer5_out[1466];
     layer6_out[1307] <= ~layer5_out[970];
     layer6_out[1308] <= ~layer5_out[340];
     layer6_out[1309] <= layer5_out[815] & ~layer5_out[814];
     layer6_out[1310] <= ~layer5_out[870];
     layer6_out[1311] <= ~(layer5_out[897] | layer5_out[898]);
     layer6_out[1312] <= ~(layer5_out[147] & layer5_out[148]);
     layer6_out[1313] <= ~layer5_out[1288] | layer5_out[1289];
     layer6_out[1314] <= layer5_out[949] ^ layer5_out[950];
     layer6_out[1315] <= layer5_out[701];
     layer6_out[1316] <= layer5_out[669];
     layer6_out[1317] <= ~layer5_out[189];
     layer6_out[1318] <= ~layer5_out[1406] | layer5_out[1405];
     layer6_out[1319] <= ~layer5_out[1420];
     layer6_out[1320] <= layer5_out[218] & layer5_out[219];
     layer6_out[1321] <= layer5_out[973] ^ layer5_out[974];
     layer6_out[1322] <= ~(layer5_out[829] ^ layer5_out[830]);
     layer6_out[1323] <= ~layer5_out[484] | layer5_out[483];
     layer6_out[1324] <= ~layer5_out[1217];
     layer6_out[1325] <= ~(layer5_out[1242] ^ layer5_out[1243]);
     layer6_out[1326] <= layer5_out[279];
     layer6_out[1327] <= ~(layer5_out[130] | layer5_out[131]);
     layer6_out[1328] <= ~layer5_out[1431];
     layer6_out[1329] <= layer5_out[130];
     layer6_out[1330] <= layer5_out[763] & ~layer5_out[764];
     layer6_out[1331] <= 1'b1;
     layer6_out[1332] <= ~(layer5_out[1068] & layer5_out[1069]);
     layer6_out[1333] <= ~layer5_out[330];
     layer6_out[1334] <= ~layer5_out[246];
     layer6_out[1335] <= ~layer5_out[398];
     layer6_out[1336] <= layer5_out[735];
     layer6_out[1337] <= layer5_out[348] & ~layer5_out[347];
     layer6_out[1338] <= layer5_out[1081] | layer5_out[1082];
     layer6_out[1339] <= layer5_out[1385] & ~layer5_out[1386];
     layer6_out[1340] <= ~(layer5_out[1061] ^ layer5_out[1062]);
     layer6_out[1341] <= layer5_out[885] ^ layer5_out[886];
     layer6_out[1342] <= layer5_out[353];
     layer6_out[1343] <= ~layer5_out[1046];
     layer6_out[1344] <= layer5_out[364] & ~layer5_out[363];
     layer6_out[1345] <= ~layer5_out[1143];
     layer6_out[1346] <= layer5_out[1196];
     layer6_out[1347] <= ~layer5_out[1497] | layer5_out[1498];
     layer6_out[1348] <= layer5_out[579] ^ layer5_out[580];
     layer6_out[1349] <= layer5_out[575];
     layer6_out[1350] <= ~layer5_out[1396] | layer5_out[1395];
     layer6_out[1351] <= ~layer5_out[209];
     layer6_out[1352] <= ~layer5_out[739];
     layer6_out[1353] <= ~(layer5_out[1148] & layer5_out[1149]);
     layer6_out[1354] <= layer5_out[604];
     layer6_out[1355] <= layer5_out[607] & ~layer5_out[606];
     layer6_out[1356] <= ~(layer5_out[296] | layer5_out[297]);
     layer6_out[1357] <= ~layer5_out[1038];
     layer6_out[1358] <= layer5_out[795] & layer5_out[796];
     layer6_out[1359] <= layer5_out[1140] & ~layer5_out[1139];
     layer6_out[1360] <= ~(layer5_out[294] | layer5_out[295]);
     layer6_out[1361] <= ~layer5_out[1452];
     layer6_out[1362] <= ~layer5_out[1117];
     layer6_out[1363] <= layer5_out[8];
     layer6_out[1364] <= layer5_out[731];
     layer6_out[1365] <= ~layer5_out[1308];
     layer6_out[1366] <= ~layer5_out[888];
     layer6_out[1367] <= ~layer5_out[181];
     layer6_out[1368] <= layer5_out[1323];
     layer6_out[1369] <= ~layer5_out[228] | layer5_out[227];
     layer6_out[1370] <= layer5_out[276];
     layer6_out[1371] <= ~(layer5_out[205] | layer5_out[206]);
     layer6_out[1372] <= 1'b1;
     layer6_out[1373] <= layer5_out[665] & layer5_out[666];
     layer6_out[1374] <= layer5_out[873];
     layer6_out[1375] <= layer5_out[737];
     layer6_out[1376] <= layer5_out[1079] & ~layer5_out[1080];
     layer6_out[1377] <= ~layer5_out[1390] | layer5_out[1389];
     layer6_out[1378] <= ~layer5_out[708];
     layer6_out[1379] <= layer5_out[1333] | layer5_out[1334];
     layer6_out[1380] <= ~layer5_out[452];
     layer6_out[1381] <= ~(layer5_out[297] ^ layer5_out[298]);
     layer6_out[1382] <= ~layer5_out[318];
     layer6_out[1383] <= layer5_out[795];
     layer6_out[1384] <= ~layer5_out[597];
     layer6_out[1385] <= layer5_out[799] | layer5_out[800];
     layer6_out[1386] <= ~layer5_out[1112];
     layer6_out[1387] <= layer5_out[658];
     layer6_out[1388] <= layer5_out[334];
     layer6_out[1389] <= layer5_out[411] ^ layer5_out[412];
     layer6_out[1390] <= layer5_out[1434] & layer5_out[1435];
     layer6_out[1391] <= ~layer5_out[246];
     layer6_out[1392] <= layer5_out[880];
     layer6_out[1393] <= ~(layer5_out[1498] | layer5_out[1499]);
     layer6_out[1394] <= ~layer5_out[226];
     layer6_out[1395] <= layer5_out[25];
     layer6_out[1396] <= layer5_out[572];
     layer6_out[1397] <= ~layer5_out[1434];
     layer6_out[1398] <= ~(layer5_out[702] ^ layer5_out[703]);
     layer6_out[1399] <= layer5_out[15] & ~layer5_out[14];
     layer6_out[1400] <= ~layer5_out[1325] | layer5_out[1326];
     layer6_out[1401] <= ~(layer5_out[373] | layer5_out[374]);
     layer6_out[1402] <= ~layer5_out[1311];
     layer6_out[1403] <= layer5_out[992];
     layer6_out[1404] <= ~layer5_out[1220] | layer5_out[1221];
     layer6_out[1405] <= ~layer5_out[2] | layer5_out[1];
     layer6_out[1406] <= ~layer5_out[125] | layer5_out[126];
     layer6_out[1407] <= ~(layer5_out[715] ^ layer5_out[716]);
     layer6_out[1408] <= layer5_out[849];
     layer6_out[1409] <= ~(layer5_out[1182] | layer5_out[1183]);
     layer6_out[1410] <= ~layer5_out[787];
     layer6_out[1411] <= layer5_out[288] ^ layer5_out[289];
     layer6_out[1412] <= ~(layer5_out[248] & layer5_out[249]);
     layer6_out[1413] <= layer5_out[255] | layer5_out[256];
     layer6_out[1414] <= 1'b0;
     layer6_out[1415] <= layer5_out[1125] & layer5_out[1126];
     layer6_out[1416] <= layer5_out[389];
     layer6_out[1417] <= ~layer5_out[445];
     layer6_out[1418] <= layer5_out[1326];
     layer6_out[1419] <= ~layer5_out[193];
     layer6_out[1420] <= layer5_out[74];
     layer6_out[1421] <= 1'b0;
     layer6_out[1422] <= ~(layer5_out[1066] | layer5_out[1067]);
     layer6_out[1423] <= layer5_out[1203] | layer5_out[1204];
     layer6_out[1424] <= ~layer5_out[27] | layer5_out[28];
     layer6_out[1425] <= ~(layer5_out[1099] | layer5_out[1100]);
     layer6_out[1426] <= layer5_out[1025];
     layer6_out[1427] <= ~layer5_out[158];
     layer6_out[1428] <= layer5_out[486] & ~layer5_out[485];
     layer6_out[1429] <= layer5_out[776];
     layer6_out[1430] <= ~layer5_out[1215] | layer5_out[1216];
     layer6_out[1431] <= layer5_out[760] | layer5_out[761];
     layer6_out[1432] <= ~layer5_out[396];
     layer6_out[1433] <= layer5_out[785] & layer5_out[786];
     layer6_out[1434] <= ~layer5_out[19];
     layer6_out[1435] <= layer5_out[450] & ~layer5_out[449];
     layer6_out[1436] <= layer5_out[748] | layer5_out[749];
     layer6_out[1437] <= layer5_out[260] & ~layer5_out[261];
     layer6_out[1438] <= layer5_out[365] & ~layer5_out[366];
     layer6_out[1439] <= ~layer5_out[440];
     layer6_out[1440] <= layer5_out[895];
     layer6_out[1441] <= ~layer5_out[943];
     layer6_out[1442] <= ~layer5_out[403];
     layer6_out[1443] <= ~(layer5_out[1476] & layer5_out[1477]);
     layer6_out[1444] <= layer5_out[1030];
     layer6_out[1445] <= ~layer5_out[569];
     layer6_out[1446] <= layer5_out[1006];
     layer6_out[1447] <= layer5_out[1368];
     layer6_out[1448] <= layer5_out[1258];
     layer6_out[1449] <= layer5_out[957] & ~layer5_out[958];
     layer6_out[1450] <= layer5_out[309];
     layer6_out[1451] <= layer5_out[545];
     layer6_out[1452] <= layer5_out[692] & ~layer5_out[693];
     layer6_out[1453] <= ~layer5_out[564] | layer5_out[563];
     layer6_out[1454] <= ~(layer5_out[1292] | layer5_out[1293]);
     layer6_out[1455] <= ~layer5_out[214];
     layer6_out[1456] <= ~layer5_out[1384];
     layer6_out[1457] <= ~layer5_out[643];
     layer6_out[1458] <= layer5_out[301] & ~layer5_out[302];
     layer6_out[1459] <= ~layer5_out[1018];
     layer6_out[1460] <= ~layer5_out[43];
     layer6_out[1461] <= ~layer5_out[1299];
     layer6_out[1462] <= ~(layer5_out[1205] | layer5_out[1206]);
     layer6_out[1463] <= ~layer5_out[1222] | layer5_out[1221];
     layer6_out[1464] <= layer5_out[756] & layer5_out[757];
     layer6_out[1465] <= ~layer5_out[1444];
     layer6_out[1466] <= 1'b1;
     layer6_out[1467] <= ~layer5_out[792];
     layer6_out[1468] <= layer5_out[791];
     layer6_out[1469] <= ~layer5_out[1339];
     layer6_out[1470] <= layer5_out[534] & ~layer5_out[535];
     layer6_out[1471] <= ~(layer5_out[700] | layer5_out[701]);
     layer6_out[1472] <= layer5_out[442] & ~layer5_out[441];
     layer6_out[1473] <= layer5_out[1224] & ~layer5_out[1223];
     layer6_out[1474] <= ~layer5_out[748] | layer5_out[747];
     layer6_out[1475] <= ~layer5_out[947] | layer5_out[948];
     layer6_out[1476] <= ~layer5_out[1247];
     layer6_out[1477] <= layer5_out[621];
     layer6_out[1478] <= layer5_out[744];
     layer6_out[1479] <= ~layer5_out[752];
     layer6_out[1480] <= layer5_out[479] & ~layer5_out[478];
     layer6_out[1481] <= layer5_out[882];
     layer6_out[1482] <= layer5_out[1005];
     layer6_out[1483] <= layer5_out[1352] & layer5_out[1353];
     layer6_out[1484] <= ~(layer5_out[335] ^ layer5_out[336]);
     layer6_out[1485] <= ~(layer5_out[925] | layer5_out[926]);
     layer6_out[1486] <= layer5_out[624];
     layer6_out[1487] <= ~layer5_out[815];
     layer6_out[1488] <= layer5_out[564];
     layer6_out[1489] <= ~layer5_out[649] | layer5_out[650];
     layer6_out[1490] <= layer5_out[66] ^ layer5_out[67];
     layer6_out[1491] <= ~layer5_out[773] | layer5_out[774];
     layer6_out[1492] <= layer5_out[826] & layer5_out[827];
     layer6_out[1493] <= ~layer5_out[1281];
     layer6_out[1494] <= ~layer5_out[445] | layer5_out[446];
     layer6_out[1495] <= ~layer5_out[65] | layer5_out[64];
     layer6_out[1496] <= layer5_out[264];
     layer6_out[1497] <= ~(layer5_out[1042] & layer5_out[1043]);
     layer6_out[1498] <= layer5_out[313] | layer5_out[314];
     layer6_out[1499] <= 1'b0;
     layer7_out[0] <= layer6_out[892] & layer6_out[893];
     layer7_out[1] <= layer6_out[501];
     layer7_out[2] <= layer6_out[1237] & layer6_out[1238];
     layer7_out[3] <= ~layer6_out[80];
     layer7_out[4] <= ~layer6_out[1325];
     layer7_out[5] <= ~(layer6_out[308] | layer6_out[309]);
     layer7_out[6] <= layer6_out[675] & layer6_out[676];
     layer7_out[7] <= layer6_out[685] & ~layer6_out[686];
     layer7_out[8] <= layer6_out[600] & ~layer6_out[601];
     layer7_out[9] <= layer6_out[1383];
     layer7_out[10] <= ~layer6_out[1002];
     layer7_out[11] <= layer6_out[662];
     layer7_out[12] <= ~(layer6_out[136] & layer6_out[137]);
     layer7_out[13] <= ~(layer6_out[373] | layer6_out[374]);
     layer7_out[14] <= layer6_out[723] & ~layer6_out[724];
     layer7_out[15] <= layer6_out[57] & ~layer6_out[56];
     layer7_out[16] <= ~(layer6_out[399] ^ layer6_out[400]);
     layer7_out[17] <= layer6_out[805] & layer6_out[806];
     layer7_out[18] <= ~(layer6_out[1428] ^ layer6_out[1429]);
     layer7_out[19] <= ~(layer6_out[1136] ^ layer6_out[1137]);
     layer7_out[20] <= layer6_out[441] & ~layer6_out[440];
     layer7_out[21] <= ~layer6_out[769];
     layer7_out[22] <= layer6_out[1210];
     layer7_out[23] <= ~(layer6_out[371] ^ layer6_out[372]);
     layer7_out[24] <= layer6_out[1396] & ~layer6_out[1395];
     layer7_out[25] <= layer6_out[1214];
     layer7_out[26] <= layer6_out[1118];
     layer7_out[27] <= ~(layer6_out[226] | layer6_out[227]);
     layer7_out[28] <= ~(layer6_out[502] ^ layer6_out[503]);
     layer7_out[29] <= ~(layer6_out[787] | layer6_out[788]);
     layer7_out[30] <= layer6_out[1220] & ~layer6_out[1221];
     layer7_out[31] <= ~layer6_out[318];
     layer7_out[32] <= ~layer6_out[1133];
     layer7_out[33] <= ~layer6_out[509];
     layer7_out[34] <= layer6_out[791] ^ layer6_out[792];
     layer7_out[35] <= ~(layer6_out[663] | layer6_out[664]);
     layer7_out[36] <= layer6_out[568];
     layer7_out[37] <= layer6_out[552];
     layer7_out[38] <= ~(layer6_out[327] | layer6_out[328]);
     layer7_out[39] <= layer6_out[822] & ~layer6_out[821];
     layer7_out[40] <= ~layer6_out[415];
     layer7_out[41] <= layer6_out[525];
     layer7_out[42] <= layer6_out[7] & ~layer6_out[8];
     layer7_out[43] <= layer6_out[203];
     layer7_out[44] <= ~(layer6_out[296] ^ layer6_out[297]);
     layer7_out[45] <= ~(layer6_out[479] ^ layer6_out[480]);
     layer7_out[46] <= ~layer6_out[1275] | layer6_out[1274];
     layer7_out[47] <= ~layer6_out[166];
     layer7_out[48] <= ~(layer6_out[602] ^ layer6_out[603]);
     layer7_out[49] <= layer6_out[526] & ~layer6_out[527];
     layer7_out[50] <= layer6_out[893] & ~layer6_out[894];
     layer7_out[51] <= ~layer6_out[160];
     layer7_out[52] <= layer6_out[538];
     layer7_out[53] <= layer6_out[1328] ^ layer6_out[1329];
     layer7_out[54] <= layer6_out[1405] & layer6_out[1406];
     layer7_out[55] <= layer6_out[235] & ~layer6_out[234];
     layer7_out[56] <= ~(layer6_out[365] ^ layer6_out[366]);
     layer7_out[57] <= ~layer6_out[1399];
     layer7_out[58] <= layer6_out[1366];
     layer7_out[59] <= ~(layer6_out[1044] | layer6_out[1045]);
     layer7_out[60] <= layer6_out[717] & ~layer6_out[718];
     layer7_out[61] <= layer6_out[1211];
     layer7_out[62] <= ~layer6_out[208];
     layer7_out[63] <= layer6_out[1197] & ~layer6_out[1196];
     layer7_out[64] <= ~layer6_out[1270];
     layer7_out[65] <= layer6_out[456];
     layer7_out[66] <= layer6_out[1425];
     layer7_out[67] <= layer6_out[1268];
     layer7_out[68] <= ~layer6_out[701];
     layer7_out[69] <= ~(layer6_out[1449] | layer6_out[1450]);
     layer7_out[70] <= ~layer6_out[594];
     layer7_out[71] <= layer6_out[905] & ~layer6_out[906];
     layer7_out[72] <= ~layer6_out[780] | layer6_out[781];
     layer7_out[73] <= layer6_out[1451] & ~layer6_out[1450];
     layer7_out[74] <= ~(layer6_out[1192] | layer6_out[1193]);
     layer7_out[75] <= ~(layer6_out[1042] | layer6_out[1043]);
     layer7_out[76] <= layer6_out[395] & layer6_out[396];
     layer7_out[77] <= layer6_out[710];
     layer7_out[78] <= layer6_out[409] | layer6_out[410];
     layer7_out[79] <= layer6_out[1336];
     layer7_out[80] <= layer6_out[1419];
     layer7_out[81] <= layer6_out[604];
     layer7_out[82] <= ~layer6_out[1277];
     layer7_out[83] <= layer6_out[910];
     layer7_out[84] <= ~(layer6_out[156] | layer6_out[157]);
     layer7_out[85] <= layer6_out[659];
     layer7_out[86] <= ~layer6_out[758];
     layer7_out[87] <= layer6_out[1257];
     layer7_out[88] <= layer6_out[1436] & ~layer6_out[1435];
     layer7_out[89] <= layer6_out[1238] & layer6_out[1239];
     layer7_out[90] <= ~(layer6_out[499] ^ layer6_out[500]);
     layer7_out[91] <= ~layer6_out[100];
     layer7_out[92] <= ~layer6_out[711] | layer6_out[712];
     layer7_out[93] <= layer6_out[800] & ~layer6_out[801];
     layer7_out[94] <= ~(layer6_out[898] | layer6_out[899]);
     layer7_out[95] <= ~layer6_out[530];
     layer7_out[96] <= ~(layer6_out[534] ^ layer6_out[535]);
     layer7_out[97] <= ~layer6_out[612];
     layer7_out[98] <= layer6_out[387];
     layer7_out[99] <= layer6_out[88] & ~layer6_out[87];
     layer7_out[100] <= ~(layer6_out[1041] | layer6_out[1042]);
     layer7_out[101] <= layer6_out[106] & ~layer6_out[105];
     layer7_out[102] <= ~layer6_out[766];
     layer7_out[103] <= ~layer6_out[1323];
     layer7_out[104] <= layer6_out[197] & layer6_out[198];
     layer7_out[105] <= ~layer6_out[1409] | layer6_out[1408];
     layer7_out[106] <= layer6_out[670] & layer6_out[671];
     layer7_out[107] <= layer6_out[857] & ~layer6_out[858];
     layer7_out[108] <= layer6_out[299] ^ layer6_out[300];
     layer7_out[109] <= layer6_out[442] & ~layer6_out[443];
     layer7_out[110] <= ~layer6_out[1301];
     layer7_out[111] <= layer6_out[1017] & layer6_out[1018];
     layer7_out[112] <= ~layer6_out[922];
     layer7_out[113] <= ~(layer6_out[689] | layer6_out[690]);
     layer7_out[114] <= layer6_out[1295] & layer6_out[1296];
     layer7_out[115] <= layer6_out[878];
     layer7_out[116] <= ~layer6_out[631] | layer6_out[632];
     layer7_out[117] <= layer6_out[568] & ~layer6_out[569];
     layer7_out[118] <= ~(layer6_out[745] ^ layer6_out[746]);
     layer7_out[119] <= ~(layer6_out[907] | layer6_out[908]);
     layer7_out[120] <= layer6_out[57];
     layer7_out[121] <= ~layer6_out[913];
     layer7_out[122] <= layer6_out[735];
     layer7_out[123] <= ~(layer6_out[1314] ^ layer6_out[1315]);
     layer7_out[124] <= layer6_out[375] & layer6_out[376];
     layer7_out[125] <= ~layer6_out[1246];
     layer7_out[126] <= layer6_out[1143];
     layer7_out[127] <= ~layer6_out[1002];
     layer7_out[128] <= ~(layer6_out[520] | layer6_out[521]);
     layer7_out[129] <= layer6_out[29];
     layer7_out[130] <= layer6_out[329] & layer6_out[330];
     layer7_out[131] <= layer6_out[423] ^ layer6_out[424];
     layer7_out[132] <= layer6_out[283];
     layer7_out[133] <= layer6_out[1451] & layer6_out[1452];
     layer7_out[134] <= layer6_out[250] & layer6_out[251];
     layer7_out[135] <= ~(layer6_out[1058] ^ layer6_out[1059]);
     layer7_out[136] <= layer6_out[514] ^ layer6_out[515];
     layer7_out[137] <= layer6_out[1103];
     layer7_out[138] <= ~(layer6_out[127] ^ layer6_out[128]);
     layer7_out[139] <= layer6_out[314] & ~layer6_out[315];
     layer7_out[140] <= ~layer6_out[861];
     layer7_out[141] <= ~layer6_out[1410] | layer6_out[1411];
     layer7_out[142] <= layer6_out[649] ^ layer6_out[650];
     layer7_out[143] <= layer6_out[881] & ~layer6_out[880];
     layer7_out[144] <= ~layer6_out[740];
     layer7_out[145] <= ~layer6_out[520];
     layer7_out[146] <= ~layer6_out[1146];
     layer7_out[147] <= ~layer6_out[1379];
     layer7_out[148] <= ~(layer6_out[783] | layer6_out[784]);
     layer7_out[149] <= layer6_out[822];
     layer7_out[150] <= ~(layer6_out[792] | layer6_out[793]);
     layer7_out[151] <= ~(layer6_out[763] | layer6_out[764]);
     layer7_out[152] <= layer6_out[1183] & ~layer6_out[1184];
     layer7_out[153] <= layer6_out[954] ^ layer6_out[955];
     layer7_out[154] <= layer6_out[875];
     layer7_out[155] <= layer6_out[678] & ~layer6_out[679];
     layer7_out[156] <= ~(layer6_out[1344] | layer6_out[1345]);
     layer7_out[157] <= layer6_out[50] & layer6_out[51];
     layer7_out[158] <= ~layer6_out[1011];
     layer7_out[159] <= layer6_out[307];
     layer7_out[160] <= layer6_out[289];
     layer7_out[161] <= layer6_out[643] & ~layer6_out[644];
     layer7_out[162] <= ~(layer6_out[1482] | layer6_out[1483]);
     layer7_out[163] <= ~(layer6_out[458] | layer6_out[459]);
     layer7_out[164] <= layer6_out[181] & layer6_out[182];
     layer7_out[165] <= layer6_out[608] & layer6_out[609];
     layer7_out[166] <= ~(layer6_out[263] | layer6_out[264]);
     layer7_out[167] <= layer6_out[272];
     layer7_out[168] <= layer6_out[915] & ~layer6_out[916];
     layer7_out[169] <= layer6_out[1108] & layer6_out[1109];
     layer7_out[170] <= ~layer6_out[267];
     layer7_out[171] <= layer6_out[1389] & ~layer6_out[1390];
     layer7_out[172] <= layer6_out[289];
     layer7_out[173] <= layer6_out[782] & layer6_out[783];
     layer7_out[174] <= layer6_out[1493];
     layer7_out[175] <= ~layer6_out[180];
     layer7_out[176] <= layer6_out[916] ^ layer6_out[917];
     layer7_out[177] <= layer6_out[1245] & ~layer6_out[1244];
     layer7_out[178] <= layer6_out[1177] & ~layer6_out[1178];
     layer7_out[179] <= layer6_out[443];
     layer7_out[180] <= ~layer6_out[543];
     layer7_out[181] <= ~(layer6_out[1063] | layer6_out[1064]);
     layer7_out[182] <= layer6_out[1142] & ~layer6_out[1143];
     layer7_out[183] <= layer6_out[352];
     layer7_out[184] <= ~(layer6_out[344] | layer6_out[345]);
     layer7_out[185] <= ~layer6_out[379];
     layer7_out[186] <= layer6_out[1037] & layer6_out[1038];
     layer7_out[187] <= ~layer6_out[1377];
     layer7_out[188] <= ~(layer6_out[91] | layer6_out[92]);
     layer7_out[189] <= layer6_out[1161] & ~layer6_out[1162];
     layer7_out[190] <= layer6_out[176];
     layer7_out[191] <= layer6_out[164];
     layer7_out[192] <= layer6_out[324];
     layer7_out[193] <= layer6_out[248] & ~layer6_out[249];
     layer7_out[194] <= ~layer6_out[251];
     layer7_out[195] <= ~(layer6_out[1168] & layer6_out[1169]);
     layer7_out[196] <= layer6_out[1264];
     layer7_out[197] <= layer6_out[336] & layer6_out[337];
     layer7_out[198] <= layer6_out[614] & ~layer6_out[613];
     layer7_out[199] <= ~(layer6_out[958] ^ layer6_out[959]);
     layer7_out[200] <= ~layer6_out[966];
     layer7_out[201] <= layer6_out[842] & ~layer6_out[843];
     layer7_out[202] <= ~(layer6_out[1049] | layer6_out[1050]);
     layer7_out[203] <= layer6_out[1250] ^ layer6_out[1251];
     layer7_out[204] <= ~layer6_out[854];
     layer7_out[205] <= layer6_out[797] & layer6_out[798];
     layer7_out[206] <= ~layer6_out[1094];
     layer7_out[207] <= ~layer6_out[988];
     layer7_out[208] <= layer6_out[1411] ^ layer6_out[1412];
     layer7_out[209] <= layer6_out[804] & ~layer6_out[805];
     layer7_out[210] <= layer6_out[715] & layer6_out[716];
     layer7_out[211] <= layer6_out[1139] & ~layer6_out[1138];
     layer7_out[212] <= layer6_out[34] & layer6_out[35];
     layer7_out[213] <= layer6_out[668] & ~layer6_out[667];
     layer7_out[214] <= layer6_out[1034];
     layer7_out[215] <= layer6_out[772];
     layer7_out[216] <= layer6_out[1167] & ~layer6_out[1166];
     layer7_out[217] <= layer6_out[192] & layer6_out[193];
     layer7_out[218] <= ~layer6_out[1498] | layer6_out[1499];
     layer7_out[219] <= layer6_out[268] & layer6_out[269];
     layer7_out[220] <= ~layer6_out[123];
     layer7_out[221] <= ~(layer6_out[1418] | layer6_out[1419]);
     layer7_out[222] <= layer6_out[533] & layer6_out[534];
     layer7_out[223] <= layer6_out[894];
     layer7_out[224] <= ~layer6_out[210];
     layer7_out[225] <= ~layer6_out[483];
     layer7_out[226] <= layer6_out[1199] & ~layer6_out[1200];
     layer7_out[227] <= ~layer6_out[776] | layer6_out[777];
     layer7_out[228] <= layer6_out[1273] ^ layer6_out[1274];
     layer7_out[229] <= ~layer6_out[618];
     layer7_out[230] <= ~(layer6_out[935] | layer6_out[936]);
     layer7_out[231] <= layer6_out[553];
     layer7_out[232] <= layer6_out[908] & ~layer6_out[909];
     layer7_out[233] <= layer6_out[282] & ~layer6_out[283];
     layer7_out[234] <= layer6_out[563] & ~layer6_out[564];
     layer7_out[235] <= layer6_out[906] ^ layer6_out[907];
     layer7_out[236] <= ~(layer6_out[1467] ^ layer6_out[1468]);
     layer7_out[237] <= layer6_out[1349] & ~layer6_out[1350];
     layer7_out[238] <= ~layer6_out[30];
     layer7_out[239] <= layer6_out[1092] & ~layer6_out[1091];
     layer7_out[240] <= ~(layer6_out[1208] | layer6_out[1209]);
     layer7_out[241] <= layer6_out[719] & ~layer6_out[718];
     layer7_out[242] <= layer6_out[268] & ~layer6_out[267];
     layer7_out[243] <= layer6_out[95] & ~layer6_out[94];
     layer7_out[244] <= layer6_out[983] & ~layer6_out[982];
     layer7_out[245] <= ~(layer6_out[262] | layer6_out[263]);
     layer7_out[246] <= ~(layer6_out[1025] | layer6_out[1026]);
     layer7_out[247] <= layer6_out[781] & layer6_out[782];
     layer7_out[248] <= layer6_out[1248] & ~layer6_out[1249];
     layer7_out[249] <= layer6_out[1333] & ~layer6_out[1334];
     layer7_out[250] <= ~layer6_out[743];
     layer7_out[251] <= layer6_out[625] & ~layer6_out[624];
     layer7_out[252] <= ~(layer6_out[510] ^ layer6_out[511]);
     layer7_out[253] <= ~layer6_out[518];
     layer7_out[254] <= layer6_out[214] & layer6_out[215];
     layer7_out[255] <= layer6_out[244] & layer6_out[245];
     layer7_out[256] <= ~layer6_out[86];
     layer7_out[257] <= layer6_out[1135];
     layer7_out[258] <= layer6_out[247] & layer6_out[248];
     layer7_out[259] <= ~(layer6_out[660] ^ layer6_out[661]);
     layer7_out[260] <= ~(layer6_out[93] | layer6_out[94]);
     layer7_out[261] <= layer6_out[309];
     layer7_out[262] <= layer6_out[1401] & layer6_out[1402];
     layer7_out[263] <= ~(layer6_out[1086] | layer6_out[1087]);
     layer7_out[264] <= layer6_out[1426] & ~layer6_out[1425];
     layer7_out[265] <= layer6_out[1279] & ~layer6_out[1280];
     layer7_out[266] <= ~(layer6_out[417] | layer6_out[418]);
     layer7_out[267] <= ~(layer6_out[716] ^ layer6_out[717]);
     layer7_out[268] <= layer6_out[924] & layer6_out[925];
     layer7_out[269] <= layer6_out[170] & layer6_out[171];
     layer7_out[270] <= layer6_out[575] & ~layer6_out[574];
     layer7_out[271] <= layer6_out[1393];
     layer7_out[272] <= layer6_out[564] ^ layer6_out[565];
     layer7_out[273] <= layer6_out[1361] & ~layer6_out[1360];
     layer7_out[274] <= ~(layer6_out[546] ^ layer6_out[547]);
     layer7_out[275] <= layer6_out[1404] & ~layer6_out[1405];
     layer7_out[276] <= layer6_out[882] & layer6_out[883];
     layer7_out[277] <= ~layer6_out[151];
     layer7_out[278] <= ~(layer6_out[817] | layer6_out[818]);
     layer7_out[279] <= layer6_out[384] ^ layer6_out[385];
     layer7_out[280] <= layer6_out[680] & ~layer6_out[681];
     layer7_out[281] <= layer6_out[383];
     layer7_out[282] <= layer6_out[1340] & layer6_out[1341];
     layer7_out[283] <= ~layer6_out[471];
     layer7_out[284] <= layer6_out[610] & ~layer6_out[611];
     layer7_out[285] <= layer6_out[1089] ^ layer6_out[1090];
     layer7_out[286] <= layer6_out[1222] & ~layer6_out[1223];
     layer7_out[287] <= layer6_out[77] ^ layer6_out[78];
     layer7_out[288] <= layer6_out[362];
     layer7_out[289] <= ~layer6_out[988];
     layer7_out[290] <= layer6_out[1045] & layer6_out[1046];
     layer7_out[291] <= ~layer6_out[1005];
     layer7_out[292] <= ~(layer6_out[1310] ^ layer6_out[1311]);
     layer7_out[293] <= layer6_out[32] & ~layer6_out[33];
     layer7_out[294] <= layer6_out[1181];
     layer7_out[295] <= layer6_out[1490] & layer6_out[1491];
     layer7_out[296] <= ~layer6_out[1096];
     layer7_out[297] <= ~layer6_out[449] | layer6_out[450];
     layer7_out[298] <= layer6_out[1131] & ~layer6_out[1132];
     layer7_out[299] <= ~layer6_out[1061];
     layer7_out[300] <= ~layer6_out[28] | layer6_out[27];
     layer7_out[301] <= layer6_out[722];
     layer7_out[302] <= ~layer6_out[590];
     layer7_out[303] <= ~layer6_out[1269];
     layer7_out[304] <= layer6_out[1185] & layer6_out[1186];
     layer7_out[305] <= ~layer6_out[170];
     layer7_out[306] <= layer6_out[1172] & ~layer6_out[1171];
     layer7_out[307] <= ~layer6_out[871];
     layer7_out[308] <= ~layer6_out[937];
     layer7_out[309] <= ~layer6_out[659];
     layer7_out[310] <= ~layer6_out[1243];
     layer7_out[311] <= ~(layer6_out[996] & layer6_out[997]);
     layer7_out[312] <= layer6_out[1389];
     layer7_out[313] <= ~layer6_out[814];
     layer7_out[314] <= layer6_out[1080] & layer6_out[1081];
     layer7_out[315] <= ~(layer6_out[666] ^ layer6_out[667]);
     layer7_out[316] <= layer6_out[1038];
     layer7_out[317] <= ~(layer6_out[272] | layer6_out[273]);
     layer7_out[318] <= ~(layer6_out[311] ^ layer6_out[312]);
     layer7_out[319] <= ~layer6_out[1265];
     layer7_out[320] <= layer6_out[612] ^ layer6_out[613];
     layer7_out[321] <= ~layer6_out[918];
     layer7_out[322] <= layer6_out[1358];
     layer7_out[323] <= layer6_out[1447] | layer6_out[1448];
     layer7_out[324] <= ~layer6_out[843];
     layer7_out[325] <= layer6_out[831] & ~layer6_out[830];
     layer7_out[326] <= ~layer6_out[575];
     layer7_out[327] <= ~layer6_out[1222];
     layer7_out[328] <= ~(layer6_out[187] | layer6_out[188]);
     layer7_out[329] <= ~layer6_out[279] | layer6_out[278];
     layer7_out[330] <= layer6_out[1444];
     layer7_out[331] <= layer6_out[886] & layer6_out[887];
     layer7_out[332] <= layer6_out[940];
     layer7_out[333] <= ~(layer6_out[531] ^ layer6_out[532]);
     layer7_out[334] <= layer6_out[13];
     layer7_out[335] <= ~layer6_out[673];
     layer7_out[336] <= layer6_out[621] & layer6_out[622];
     layer7_out[337] <= ~(layer6_out[96] ^ layer6_out[97]);
     layer7_out[338] <= layer6_out[232] ^ layer6_out[233];
     layer7_out[339] <= ~layer6_out[865];
     layer7_out[340] <= ~layer6_out[1234];
     layer7_out[341] <= ~layer6_out[310] | layer6_out[311];
     layer7_out[342] <= ~layer6_out[1054];
     layer7_out[343] <= layer6_out[1397] | layer6_out[1398];
     layer7_out[344] <= layer6_out[334] | layer6_out[335];
     layer7_out[345] <= ~(layer6_out[657] ^ layer6_out[658]);
     layer7_out[346] <= layer6_out[584] | layer6_out[585];
     layer7_out[347] <= ~layer6_out[112];
     layer7_out[348] <= layer6_out[900];
     layer7_out[349] <= ~layer6_out[630];
     layer7_out[350] <= layer6_out[10];
     layer7_out[351] <= ~(layer6_out[671] | layer6_out[672]);
     layer7_out[352] <= layer6_out[461];
     layer7_out[353] <= layer6_out[72] & layer6_out[73];
     layer7_out[354] <= layer6_out[1040] ^ layer6_out[1041];
     layer7_out[355] <= ~layer6_out[409];
     layer7_out[356] <= layer6_out[1262];
     layer7_out[357] <= ~layer6_out[616];
     layer7_out[358] <= layer6_out[1420] | layer6_out[1421];
     layer7_out[359] <= ~layer6_out[1332];
     layer7_out[360] <= ~layer6_out[47] | layer6_out[48];
     layer7_out[361] <= ~layer6_out[1354];
     layer7_out[362] <= layer6_out[1035];
     layer7_out[363] <= ~layer6_out[1351];
     layer7_out[364] <= ~(layer6_out[697] | layer6_out[698]);
     layer7_out[365] <= layer6_out[1267] & ~layer6_out[1266];
     layer7_out[366] <= layer6_out[655];
     layer7_out[367] <= layer6_out[1200];
     layer7_out[368] <= ~(layer6_out[1109] | layer6_out[1110]);
     layer7_out[369] <= layer6_out[479] & ~layer6_out[478];
     layer7_out[370] <= ~layer6_out[1202];
     layer7_out[371] <= ~(layer6_out[1306] ^ layer6_out[1307]);
     layer7_out[372] <= ~layer6_out[64];
     layer7_out[373] <= ~(layer6_out[1062] ^ layer6_out[1063]);
     layer7_out[374] <= ~layer6_out[1297];
     layer7_out[375] <= layer6_out[432] & ~layer6_out[433];
     layer7_out[376] <= ~layer6_out[1208];
     layer7_out[377] <= ~(layer6_out[412] & layer6_out[413]);
     layer7_out[378] <= ~(layer6_out[1057] ^ layer6_out[1058]);
     layer7_out[379] <= layer6_out[149];
     layer7_out[380] <= layer6_out[1261] ^ layer6_out[1262];
     layer7_out[381] <= layer6_out[970] & ~layer6_out[971];
     layer7_out[382] <= ~layer6_out[1257];
     layer7_out[383] <= layer6_out[262];
     layer7_out[384] <= ~layer6_out[952];
     layer7_out[385] <= ~(layer6_out[279] ^ layer6_out[280]);
     layer7_out[386] <= ~(layer6_out[1390] | layer6_out[1391]);
     layer7_out[387] <= layer6_out[1053];
     layer7_out[388] <= layer6_out[464] & ~layer6_out[463];
     layer7_out[389] <= layer6_out[427] & ~layer6_out[426];
     layer7_out[390] <= layer6_out[640];
     layer7_out[391] <= layer6_out[58] & ~layer6_out[59];
     layer7_out[392] <= layer6_out[570] & ~layer6_out[569];
     layer7_out[393] <= layer6_out[25] ^ layer6_out[26];
     layer7_out[394] <= layer6_out[950];
     layer7_out[395] <= layer6_out[1289];
     layer7_out[396] <= layer6_out[110] ^ layer6_out[111];
     layer7_out[397] <= ~layer6_out[932] | layer6_out[931];
     layer7_out[398] <= ~layer6_out[937];
     layer7_out[399] <= layer6_out[616] ^ layer6_out[617];
     layer7_out[400] <= layer6_out[1102];
     layer7_out[401] <= ~layer6_out[509] | layer6_out[510];
     layer7_out[402] <= ~layer6_out[475];
     layer7_out[403] <= ~(layer6_out[748] ^ layer6_out[749]);
     layer7_out[404] <= layer6_out[1088] ^ layer6_out[1089];
     layer7_out[405] <= layer6_out[8];
     layer7_out[406] <= ~(layer6_out[784] | layer6_out[785]);
     layer7_out[407] <= ~layer6_out[1287];
     layer7_out[408] <= ~layer6_out[434];
     layer7_out[409] <= layer6_out[1469];
     layer7_out[410] <= ~(layer6_out[1068] ^ layer6_out[1069]);
     layer7_out[411] <= layer6_out[1061] & ~layer6_out[1060];
     layer7_out[412] <= ~layer6_out[687] | layer6_out[686];
     layer7_out[413] <= ~layer6_out[969];
     layer7_out[414] <= layer6_out[915] & ~layer6_out[914];
     layer7_out[415] <= ~(layer6_out[1197] | layer6_out[1198]);
     layer7_out[416] <= ~layer6_out[678];
     layer7_out[417] <= layer6_out[884] ^ layer6_out[885];
     layer7_out[418] <= ~layer6_out[785];
     layer7_out[419] <= layer6_out[1033];
     layer7_out[420] <= ~layer6_out[977];
     layer7_out[421] <= ~(layer6_out[302] & layer6_out[303]);
     layer7_out[422] <= layer6_out[298] & ~layer6_out[297];
     layer7_out[423] <= ~layer6_out[1392];
     layer7_out[424] <= layer6_out[1242] & ~layer6_out[1241];
     layer7_out[425] <= ~layer6_out[495] | layer6_out[496];
     layer7_out[426] <= ~(layer6_out[1366] ^ layer6_out[1367]);
     layer7_out[427] <= ~(layer6_out[1169] ^ layer6_out[1170]);
     layer7_out[428] <= ~layer6_out[825];
     layer7_out[429] <= layer6_out[452] ^ layer6_out[453];
     layer7_out[430] <= ~layer6_out[249];
     layer7_out[431] <= ~layer6_out[354] | layer6_out[355];
     layer7_out[432] <= layer6_out[240];
     layer7_out[433] <= ~layer6_out[99];
     layer7_out[434] <= ~layer6_out[264];
     layer7_out[435] <= ~(layer6_out[1251] | layer6_out[1252]);
     layer7_out[436] <= ~(layer6_out[1440] ^ layer6_out[1441]);
     layer7_out[437] <= layer6_out[930];
     layer7_out[438] <= ~(layer6_out[1317] ^ layer6_out[1318]);
     layer7_out[439] <= ~(layer6_out[544] | layer6_out[545]);
     layer7_out[440] <= layer6_out[1494];
     layer7_out[441] <= layer6_out[920] & layer6_out[921];
     layer7_out[442] <= layer6_out[1226] ^ layer6_out[1227];
     layer7_out[443] <= layer6_out[594];
     layer7_out[444] <= ~layer6_out[1313];
     layer7_out[445] <= ~(layer6_out[1364] ^ layer6_out[1365]);
     layer7_out[446] <= ~(layer6_out[0] ^ layer6_out[2]);
     layer7_out[447] <= ~layer6_out[975];
     layer7_out[448] <= layer6_out[210];
     layer7_out[449] <= ~layer6_out[378];
     layer7_out[450] <= ~layer6_out[1329];
     layer7_out[451] <= ~(layer6_out[1014] | layer6_out[1015]);
     layer7_out[452] <= ~layer6_out[162];
     layer7_out[453] <= ~layer6_out[992];
     layer7_out[454] <= layer6_out[59];
     layer7_out[455] <= layer6_out[1464];
     layer7_out[456] <= layer6_out[693];
     layer7_out[457] <= ~(layer6_out[82] ^ layer6_out[83]);
     layer7_out[458] <= ~layer6_out[1431];
     layer7_out[459] <= layer6_out[935];
     layer7_out[460] <= layer6_out[14];
     layer7_out[461] <= ~layer6_out[1131] | layer6_out[1130];
     layer7_out[462] <= layer6_out[191] ^ layer6_out[192];
     layer7_out[463] <= layer6_out[1338];
     layer7_out[464] <= layer6_out[1402] & ~layer6_out[1403];
     layer7_out[465] <= ~layer6_out[593];
     layer7_out[466] <= layer6_out[986] & ~layer6_out[987];
     layer7_out[467] <= layer6_out[1120] ^ layer6_out[1121];
     layer7_out[468] <= ~layer6_out[255];
     layer7_out[469] <= layer6_out[345] | layer6_out[346];
     layer7_out[470] <= layer6_out[714];
     layer7_out[471] <= ~layer6_out[18];
     layer7_out[472] <= layer6_out[741];
     layer7_out[473] <= layer6_out[225] & layer6_out[226];
     layer7_out[474] <= layer6_out[546];
     layer7_out[475] <= layer6_out[451] & layer6_out[452];
     layer7_out[476] <= layer6_out[1338] & layer6_out[1339];
     layer7_out[477] <= ~(layer6_out[241] & layer6_out[242]);
     layer7_out[478] <= layer6_out[1124] & ~layer6_out[1123];
     layer7_out[479] <= layer6_out[560] | layer6_out[561];
     layer7_out[480] <= ~layer6_out[625];
     layer7_out[481] <= layer6_out[563];
     layer7_out[482] <= ~layer6_out[1454];
     layer7_out[483] <= ~(layer6_out[1145] ^ layer6_out[1146]);
     layer7_out[484] <= layer6_out[1211] | layer6_out[1212];
     layer7_out[485] <= layer6_out[1080];
     layer7_out[486] <= ~layer6_out[307];
     layer7_out[487] <= ~layer6_out[50] | layer6_out[49];
     layer7_out[488] <= layer6_out[142];
     layer7_out[489] <= ~layer6_out[475];
     layer7_out[490] <= layer6_out[647] & ~layer6_out[648];
     layer7_out[491] <= layer6_out[419] & ~layer6_out[420];
     layer7_out[492] <= ~layer6_out[699] | layer6_out[698];
     layer7_out[493] <= ~(layer6_out[1471] | layer6_out[1472]);
     layer7_out[494] <= ~layer6_out[1093];
     layer7_out[495] <= ~layer6_out[835];
     layer7_out[496] <= ~(layer6_out[472] ^ layer6_out[473]);
     layer7_out[497] <= ~layer6_out[127];
     layer7_out[498] <= layer6_out[855] & ~layer6_out[856];
     layer7_out[499] <= layer6_out[125] & ~layer6_out[124];
     layer7_out[500] <= layer6_out[854] & layer6_out[855];
     layer7_out[501] <= ~layer6_out[1189] | layer6_out[1190];
     layer7_out[502] <= layer6_out[1386] ^ layer6_out[1387];
     layer7_out[503] <= ~layer6_out[19];
     layer7_out[504] <= layer6_out[1232];
     layer7_out[505] <= ~(layer6_out[182] | layer6_out[183]);
     layer7_out[506] <= layer6_out[333] | layer6_out[334];
     layer7_out[507] <= ~layer6_out[543];
     layer7_out[508] <= ~layer6_out[888];
     layer7_out[509] <= ~layer6_out[139];
     layer7_out[510] <= ~(layer6_out[1214] | layer6_out[1215]);
     layer7_out[511] <= ~layer6_out[352];
     layer7_out[512] <= layer6_out[446] & ~layer6_out[447];
     layer7_out[513] <= ~(layer6_out[1110] | layer6_out[1111]);
     layer7_out[514] <= layer6_out[1008] & ~layer6_out[1009];
     layer7_out[515] <= layer6_out[1193] & ~layer6_out[1194];
     layer7_out[516] <= layer6_out[219] & layer6_out[220];
     layer7_out[517] <= layer6_out[380];
     layer7_out[518] <= ~layer6_out[1369];
     layer7_out[519] <= layer6_out[157] & layer6_out[158];
     layer7_out[520] <= layer6_out[393] & ~layer6_out[392];
     layer7_out[521] <= ~layer6_out[84];
     layer7_out[522] <= layer6_out[1464];
     layer7_out[523] <= layer6_out[316] & layer6_out[317];
     layer7_out[524] <= layer6_out[998] | layer6_out[999];
     layer7_out[525] <= ~(layer6_out[1235] ^ layer6_out[1236]);
     layer7_out[526] <= ~layer6_out[7];
     layer7_out[527] <= layer6_out[1176] & ~layer6_out[1177];
     layer7_out[528] <= layer6_out[385];
     layer7_out[529] <= ~layer6_out[107];
     layer7_out[530] <= ~layer6_out[1478];
     layer7_out[531] <= layer6_out[601];
     layer7_out[532] <= layer6_out[883] | layer6_out[884];
     layer7_out[533] <= ~(layer6_out[41] ^ layer6_out[42]);
     layer7_out[534] <= layer6_out[867] & ~layer6_out[866];
     layer7_out[535] <= layer6_out[969] & layer6_out[970];
     layer7_out[536] <= ~layer6_out[507] | layer6_out[508];
     layer7_out[537] <= layer6_out[1309] & ~layer6_out[1308];
     layer7_out[538] <= layer6_out[901];
     layer7_out[539] <= layer6_out[366];
     layer7_out[540] <= ~(layer6_out[83] ^ layer6_out[84]);
     layer7_out[541] <= ~layer6_out[504];
     layer7_out[542] <= ~layer6_out[1408];
     layer7_out[543] <= layer6_out[844];
     layer7_out[544] <= layer6_out[67];
     layer7_out[545] <= layer6_out[1171];
     layer7_out[546] <= layer6_out[1289];
     layer7_out[547] <= ~layer6_out[1095];
     layer7_out[548] <= ~layer6_out[846];
     layer7_out[549] <= layer6_out[756] ^ layer6_out[757];
     layer7_out[550] <= layer6_out[1360];
     layer7_out[551] <= layer6_out[769] & ~layer6_out[768];
     layer7_out[552] <= ~(layer6_out[387] ^ layer6_out[388]);
     layer7_out[553] <= ~layer6_out[752];
     layer7_out[554] <= layer6_out[416] ^ layer6_out[417];
     layer7_out[555] <= layer6_out[572] ^ layer6_out[573];
     layer7_out[556] <= layer6_out[738] & layer6_out[739];
     layer7_out[557] <= layer6_out[356];
     layer7_out[558] <= layer6_out[153];
     layer7_out[559] <= ~layer6_out[856];
     layer7_out[560] <= ~layer6_out[590];
     layer7_out[561] <= layer6_out[1299] ^ layer6_out[1300];
     layer7_out[562] <= layer6_out[878];
     layer7_out[563] <= ~layer6_out[786] | layer6_out[787];
     layer7_out[564] <= layer6_out[690];
     layer7_out[565] <= ~layer6_out[498];
     layer7_out[566] <= layer6_out[775] & layer6_out[776];
     layer7_out[567] <= ~layer6_out[40] | layer6_out[41];
     layer7_out[568] <= ~layer6_out[260];
     layer7_out[569] <= layer6_out[46] & layer6_out[47];
     layer7_out[570] <= ~(layer6_out[679] ^ layer6_out[680]);
     layer7_out[571] <= layer6_out[125];
     layer7_out[572] <= layer6_out[1443] & ~layer6_out[1442];
     layer7_out[573] <= layer6_out[104] & ~layer6_out[105];
     layer7_out[574] <= ~(layer6_out[456] | layer6_out[457]);
     layer7_out[575] <= layer6_out[505];
     layer7_out[576] <= layer6_out[1342];
     layer7_out[577] <= layer6_out[1356] & ~layer6_out[1355];
     layer7_out[578] <= ~layer6_out[995];
     layer7_out[579] <= layer6_out[577];
     layer7_out[580] <= ~layer6_out[1301];
     layer7_out[581] <= ~layer6_out[242] | layer6_out[243];
     layer7_out[582] <= layer6_out[1069];
     layer7_out[583] <= ~(layer6_out[21] ^ layer6_out[22]);
     layer7_out[584] <= layer6_out[1182] & ~layer6_out[1181];
     layer7_out[585] <= layer6_out[1150] & layer6_out[1151];
     layer7_out[586] <= ~(layer6_out[403] | layer6_out[404]);
     layer7_out[587] <= ~layer6_out[558];
     layer7_out[588] <= layer6_out[103] & layer6_out[104];
     layer7_out[589] <= ~(layer6_out[38] ^ layer6_out[39]);
     layer7_out[590] <= ~layer6_out[12];
     layer7_out[591] <= layer6_out[305] ^ layer6_out[306];
     layer7_out[592] <= ~layer6_out[255];
     layer7_out[593] <= ~layer6_out[719];
     layer7_out[594] <= layer6_out[153] & ~layer6_out[152];
     layer7_out[595] <= layer6_out[454];
     layer7_out[596] <= layer6_out[282];
     layer7_out[597] <= layer6_out[1335] & ~layer6_out[1334];
     layer7_out[598] <= ~layer6_out[1373];
     layer7_out[599] <= ~layer6_out[529] | layer6_out[528];
     layer7_out[600] <= layer6_out[322];
     layer7_out[601] <= layer6_out[393] & ~layer6_out[394];
     layer7_out[602] <= layer6_out[1249] ^ layer6_out[1250];
     layer7_out[603] <= ~(layer6_out[203] | layer6_out[204]);
     layer7_out[604] <= layer6_out[193] & ~layer6_out[194];
     layer7_out[605] <= layer6_out[71];
     layer7_out[606] <= ~layer6_out[1048] | layer6_out[1047];
     layer7_out[607] <= layer6_out[872] & layer6_out[873];
     layer7_out[608] <= ~layer6_out[1482];
     layer7_out[609] <= layer6_out[260];
     layer7_out[610] <= ~layer6_out[623] | layer6_out[624];
     layer7_out[611] <= layer6_out[1324];
     layer7_out[612] <= ~layer6_out[891];
     layer7_out[613] <= layer6_out[60] & layer6_out[61];
     layer7_out[614] <= layer6_out[155];
     layer7_out[615] <= layer6_out[961] | layer6_out[962];
     layer7_out[616] <= layer6_out[411] | layer6_out[412];
     layer7_out[617] <= layer6_out[246];
     layer7_out[618] <= layer6_out[558];
     layer7_out[619] <= ~layer6_out[429];
     layer7_out[620] <= ~(layer6_out[1172] | layer6_out[1173]);
     layer7_out[621] <= layer6_out[1487] | layer6_out[1488];
     layer7_out[622] <= layer6_out[398] ^ layer6_out[399];
     layer7_out[623] <= layer6_out[462] & layer6_out[463];
     layer7_out[624] <= layer6_out[1093] & ~layer6_out[1094];
     layer7_out[625] <= layer6_out[115];
     layer7_out[626] <= layer6_out[704] ^ layer6_out[705];
     layer7_out[627] <= layer6_out[1441];
     layer7_out[628] <= layer6_out[552];
     layer7_out[629] <= ~layer6_out[1048];
     layer7_out[630] <= ~(layer6_out[945] ^ layer6_out[946]);
     layer7_out[631] <= layer6_out[218] & layer6_out[219];
     layer7_out[632] <= ~layer6_out[1285];
     layer7_out[633] <= ~layer6_out[1106];
     layer7_out[634] <= ~layer6_out[620];
     layer7_out[635] <= layer6_out[199];
     layer7_out[636] <= ~(layer6_out[980] & layer6_out[981]);
     layer7_out[637] <= ~layer6_out[565];
     layer7_out[638] <= layer6_out[1246];
     layer7_out[639] <= ~(layer6_out[851] ^ layer6_out[852]);
     layer7_out[640] <= ~(layer6_out[1055] & layer6_out[1056]);
     layer7_out[641] <= layer6_out[1194];
     layer7_out[642] <= layer6_out[827] & layer6_out[828];
     layer7_out[643] <= ~layer6_out[766];
     layer7_out[644] <= layer6_out[246] & ~layer6_out[245];
     layer7_out[645] <= layer6_out[637];
     layer7_out[646] <= ~layer6_out[1406];
     layer7_out[647] <= layer6_out[839] & layer6_out[840];
     layer7_out[648] <= ~(layer6_out[1371] ^ layer6_out[1372]);
     layer7_out[649] <= ~(layer6_out[835] | layer6_out[836]);
     layer7_out[650] <= layer6_out[1076];
     layer7_out[651] <= layer6_out[1448] | layer6_out[1449];
     layer7_out[652] <= layer6_out[839] & ~layer6_out[838];
     layer7_out[653] <= ~(layer6_out[859] ^ layer6_out[860]);
     layer7_out[654] <= ~layer6_out[795];
     layer7_out[655] <= layer6_out[75] & ~layer6_out[74];
     layer7_out[656] <= ~layer6_out[853];
     layer7_out[657] <= ~(layer6_out[1056] ^ layer6_out[1057]);
     layer7_out[658] <= layer6_out[450];
     layer7_out[659] <= ~layer6_out[1240];
     layer7_out[660] <= ~layer6_out[1456];
     layer7_out[661] <= layer6_out[436] & ~layer6_out[437];
     layer7_out[662] <= layer6_out[978] | layer6_out[979];
     layer7_out[663] <= layer6_out[828];
     layer7_out[664] <= ~layer6_out[54] | layer6_out[53];
     layer7_out[665] <= layer6_out[1371];
     layer7_out[666] <= layer6_out[774];
     layer7_out[667] <= layer6_out[1255] & ~layer6_out[1254];
     layer7_out[668] <= ~layer6_out[957];
     layer7_out[669] <= ~(layer6_out[471] & layer6_out[472]);
     layer7_out[670] <= layer6_out[369];
     layer7_out[671] <= ~(layer6_out[881] ^ layer6_out[882]);
     layer7_out[672] <= layer6_out[1480] ^ layer6_out[1481];
     layer7_out[673] <= ~layer6_out[1167];
     layer7_out[674] <= ~layer6_out[34];
     layer7_out[675] <= layer6_out[1467];
     layer7_out[676] <= layer6_out[1312] & ~layer6_out[1311];
     layer7_out[677] <= layer6_out[292];
     layer7_out[678] <= ~(layer6_out[1293] | layer6_out[1294]);
     layer7_out[679] <= layer6_out[62];
     layer7_out[680] <= layer6_out[1470] ^ layer6_out[1471];
     layer7_out[681] <= ~layer6_out[128];
     layer7_out[682] <= ~layer6_out[131];
     layer7_out[683] <= ~layer6_out[693];
     layer7_out[684] <= ~layer6_out[1014];
     layer7_out[685] <= ~layer6_out[1083];
     layer7_out[686] <= layer6_out[1114];
     layer7_out[687] <= ~(layer6_out[1375] ^ layer6_out[1376]);
     layer7_out[688] <= ~(layer6_out[492] | layer6_out[493]);
     layer7_out[689] <= layer6_out[1428] & ~layer6_out[1427];
     layer7_out[690] <= layer6_out[771];
     layer7_out[691] <= ~layer6_out[488];
     layer7_out[692] <= layer6_out[1047];
     layer7_out[693] <= ~layer6_out[421];
     layer7_out[694] <= ~(layer6_out[874] & layer6_out[875]);
     layer7_out[695] <= layer6_out[995];
     layer7_out[696] <= ~(layer6_out[913] | layer6_out[914]);
     layer7_out[697] <= layer6_out[691] ^ layer6_out[692];
     layer7_out[698] <= layer6_out[389];
     layer7_out[699] <= layer6_out[1153];
     layer7_out[700] <= ~layer6_out[579] | layer6_out[578];
     layer7_out[701] <= ~layer6_out[340] | layer6_out[339];
     layer7_out[702] <= layer6_out[591];
     layer7_out[703] <= layer6_out[619];
     layer7_out[704] <= ~(layer6_out[1260] | layer6_out[1261]);
     layer7_out[705] <= ~layer6_out[133];
     layer7_out[706] <= layer6_out[644] ^ layer6_out[645];
     layer7_out[707] <= layer6_out[115];
     layer7_out[708] <= layer6_out[943] & ~layer6_out[942];
     layer7_out[709] <= ~layer6_out[113];
     layer7_out[710] <= layer6_out[406];
     layer7_out[711] <= ~(layer6_out[863] ^ layer6_out[864]);
     layer7_out[712] <= ~layer6_out[570];
     layer7_out[713] <= layer6_out[847];
     layer7_out[714] <= layer6_out[771] & ~layer6_out[772];
     layer7_out[715] <= ~layer6_out[79];
     layer7_out[716] <= ~layer6_out[823];
     layer7_out[717] <= layer6_out[1019] & layer6_out[1020];
     layer7_out[718] <= layer6_out[137] & ~layer6_out[138];
     layer7_out[719] <= layer6_out[175] | layer6_out[176];
     layer7_out[720] <= ~(layer6_out[909] | layer6_out[910]);
     layer7_out[721] <= layer6_out[24];
     layer7_out[722] <= ~layer6_out[806];
     layer7_out[723] <= ~layer6_out[1159];
     layer7_out[724] <= layer6_out[39] & layer6_out[40];
     layer7_out[725] <= layer6_out[1295] & ~layer6_out[1294];
     layer7_out[726] <= ~layer6_out[440];
     layer7_out[727] <= ~layer6_out[891];
     layer7_out[728] <= layer6_out[16] | layer6_out[17];
     layer7_out[729] <= layer6_out[1015];
     layer7_out[730] <= ~layer6_out[238];
     layer7_out[731] <= ~(layer6_out[276] | layer6_out[277]);
     layer7_out[732] <= layer6_out[75];
     layer7_out[733] <= ~layer6_out[1088];
     layer7_out[734] <= ~layer6_out[3];
     layer7_out[735] <= layer6_out[1439] & ~layer6_out[1440];
     layer7_out[736] <= ~(layer6_out[1271] & layer6_out[1272]);
     layer7_out[737] <= layer6_out[212] ^ layer6_out[213];
     layer7_out[738] <= layer6_out[979];
     layer7_out[739] <= ~(layer6_out[460] | layer6_out[461]);
     layer7_out[740] <= ~layer6_out[1435];
     layer7_out[741] <= ~layer6_out[286];
     layer7_out[742] <= layer6_out[418];
     layer7_out[743] <= layer6_out[162];
     layer7_out[744] <= layer6_out[867] & ~layer6_out[868];
     layer7_out[745] <= layer6_out[581];
     layer7_out[746] <= ~layer6_out[1386];
     layer7_out[747] <= layer6_out[990] & ~layer6_out[991];
     layer7_out[748] <= layer6_out[423] & ~layer6_out[422];
     layer7_out[749] <= layer6_out[150];
     layer7_out[750] <= layer6_out[360] ^ layer6_out[361];
     layer7_out[751] <= ~layer6_out[365] | layer6_out[364];
     layer7_out[752] <= layer6_out[940] & ~layer6_out[939];
     layer7_out[753] <= ~layer6_out[1459] | layer6_out[1458];
     layer7_out[754] <= ~(layer6_out[1187] & layer6_out[1188]);
     layer7_out[755] <= layer6_out[807];
     layer7_out[756] <= layer6_out[36] | layer6_out[37];
     layer7_out[757] <= ~(layer6_out[118] | layer6_out[119]);
     layer7_out[758] <= layer6_out[1287];
     layer7_out[759] <= layer6_out[1004];
     layer7_out[760] <= layer6_out[425];
     layer7_out[761] <= layer6_out[223] & ~layer6_out[222];
     layer7_out[762] <= ~layer6_out[982];
     layer7_out[763] <= ~layer6_out[318];
     layer7_out[764] <= ~layer6_out[1077];
     layer7_out[765] <= layer6_out[1309] & layer6_out[1310];
     layer7_out[766] <= ~layer6_out[1291] | layer6_out[1292];
     layer7_out[767] <= ~(layer6_out[758] ^ layer6_out[759]);
     layer7_out[768] <= layer6_out[583] & ~layer6_out[582];
     layer7_out[769] <= layer6_out[469];
     layer7_out[770] <= layer6_out[1141];
     layer7_out[771] <= ~layer6_out[301];
     layer7_out[772] <= ~layer6_out[498];
     layer7_out[773] <= layer6_out[1160] ^ layer6_out[1161];
     layer7_out[774] <= layer6_out[1474];
     layer7_out[775] <= ~(layer6_out[720] ^ layer6_out[721]);
     layer7_out[776] <= layer6_out[561] ^ layer6_out[562];
     layer7_out[777] <= ~(layer6_out[500] | layer6_out[501]);
     layer7_out[778] <= layer6_out[469];
     layer7_out[779] <= ~layer6_out[964];
     layer7_out[780] <= ~(layer6_out[831] ^ layer6_out[832]);
     layer7_out[781] <= ~layer6_out[747];
     layer7_out[782] <= layer6_out[871] & layer6_out[872];
     layer7_out[783] <= ~layer6_out[1104];
     layer7_out[784] <= ~layer6_out[596];
     layer7_out[785] <= ~layer6_out[826] | layer6_out[825];
     layer7_out[786] <= ~layer6_out[1145];
     layer7_out[787] <= layer6_out[467];
     layer7_out[788] <= layer6_out[833] ^ layer6_out[834];
     layer7_out[789] <= layer6_out[89] ^ layer6_out[90];
     layer7_out[790] <= ~(layer6_out[1387] ^ layer6_out[1388]);
     layer7_out[791] <= ~layer6_out[332];
     layer7_out[792] <= ~layer6_out[506];
     layer7_out[793] <= layer6_out[1276] & ~layer6_out[1275];
     layer7_out[794] <= ~layer6_out[411];
     layer7_out[795] <= layer6_out[1433];
     layer7_out[796] <= layer6_out[1037] & ~layer6_out[1036];
     layer7_out[797] <= layer6_out[700] & layer6_out[701];
     layer7_out[798] <= ~layer6_out[477] | layer6_out[478];
     layer7_out[799] <= layer6_out[133];
     layer7_out[800] <= layer6_out[608] & ~layer6_out[607];
     layer7_out[801] <= layer6_out[1065];
     layer7_out[802] <= layer6_out[1000] ^ layer6_out[1001];
     layer7_out[803] <= layer6_out[1098];
     layer7_out[804] <= ~layer6_out[747];
     layer7_out[805] <= layer6_out[92];
     layer7_out[806] <= layer6_out[1016] ^ layer6_out[1017];
     layer7_out[807] <= layer6_out[1456] & ~layer6_out[1457];
     layer7_out[808] <= ~layer6_out[1302] | layer6_out[1303];
     layer7_out[809] <= layer6_out[1462] & layer6_out[1463];
     layer7_out[810] <= ~layer6_out[1362];
     layer7_out[811] <= ~layer6_out[755];
     layer7_out[812] <= ~layer6_out[862];
     layer7_out[813] <= layer6_out[295] ^ layer6_out[296];
     layer7_out[814] <= ~(layer6_out[1362] | layer6_out[1363]);
     layer7_out[815] <= ~layer6_out[1322];
     layer7_out[816] <= layer6_out[1296] ^ layer6_out[1297];
     layer7_out[817] <= layer6_out[80] & ~layer6_out[79];
     layer7_out[818] <= layer6_out[504] & ~layer6_out[505];
     layer7_out[819] <= layer6_out[918] ^ layer6_out[919];
     layer7_out[820] <= layer6_out[325];
     layer7_out[821] <= layer6_out[155] & layer6_out[156];
     layer7_out[822] <= ~layer6_out[448];
     layer7_out[823] <= layer6_out[391];
     layer7_out[824] <= ~(layer6_out[252] & layer6_out[253]);
     layer7_out[825] <= ~layer6_out[123];
     layer7_out[826] <= layer6_out[1176];
     layer7_out[827] <= ~layer6_out[491];
     layer7_out[828] <= ~layer6_out[1];
     layer7_out[829] <= layer6_out[1140] & layer6_out[1141];
     layer7_out[830] <= layer6_out[228] & ~layer6_out[227];
     layer7_out[831] <= layer6_out[1313] & ~layer6_out[1312];
     layer7_out[832] <= layer6_out[1483];
     layer7_out[833] <= layer6_out[270] & ~layer6_out[271];
     layer7_out[834] <= layer6_out[1422];
     layer7_out[835] <= ~layer6_out[284];
     layer7_out[836] <= layer6_out[513] ^ layer6_out[514];
     layer7_out[837] <= ~(layer6_out[636] ^ layer6_out[637]);
     layer7_out[838] <= ~layer6_out[497];
     layer7_out[839] <= ~layer6_out[696];
     layer7_out[840] <= layer6_out[932] ^ layer6_out[933];
     layer7_out[841] <= ~layer6_out[1348];
     layer7_out[842] <= ~layer6_out[86];
     layer7_out[843] <= layer6_out[556];
     layer7_out[844] <= ~(layer6_out[239] ^ layer6_out[240]);
     layer7_out[845] <= layer6_out[346] | layer6_out[347];
     layer7_out[846] <= ~layer6_out[1205];
     layer7_out[847] <= ~layer6_out[641];
     layer7_out[848] <= layer6_out[67] & ~layer6_out[66];
     layer7_out[849] <= ~layer6_out[989];
     layer7_out[850] <= layer6_out[343] ^ layer6_out[344];
     layer7_out[851] <= ~layer6_out[1267];
     layer7_out[852] <= ~(layer6_out[635] ^ layer6_out[636]);
     layer7_out[853] <= ~(layer6_out[1070] | layer6_out[1071]);
     layer7_out[854] <= ~(layer6_out[1326] | layer6_out[1327]);
     layer7_out[855] <= ~layer6_out[1];
     layer7_out[856] <= layer6_out[542];
     layer7_out[857] <= ~layer6_out[1139];
     layer7_out[858] <= ~layer6_out[1125];
     layer7_out[859] <= ~(layer6_out[465] | layer6_out[466]);
     layer7_out[860] <= layer6_out[1292] | layer6_out[1293];
     layer7_out[861] <= layer6_out[1347] & ~layer6_out[1346];
     layer7_out[862] <= layer6_out[376];
     layer7_out[863] <= layer6_out[1179] & ~layer6_out[1180];
     layer7_out[864] <= layer6_out[483];
     layer7_out[865] <= layer6_out[635];
     layer7_out[866] <= ~layer6_out[186];
     layer7_out[867] <= ~(layer6_out[547] ^ layer6_out[548]);
     layer7_out[868] <= ~layer6_out[813] | layer6_out[814];
     layer7_out[869] <= ~layer6_out[874] | layer6_out[873];
     layer7_out[870] <= layer6_out[62] ^ layer6_out[63];
     layer7_out[871] <= layer6_out[167] ^ layer6_out[168];
     layer7_out[872] <= layer6_out[434];
     layer7_out[873] <= layer6_out[1422];
     layer7_out[874] <= layer6_out[208] & layer6_out[209];
     layer7_out[875] <= layer6_out[1066];
     layer7_out[876] <= layer6_out[556];
     layer7_out[877] <= layer6_out[1284] & layer6_out[1285];
     layer7_out[878] <= layer6_out[1320];
     layer7_out[879] <= layer6_out[754] & ~layer6_out[755];
     layer7_out[880] <= layer6_out[583] | layer6_out[584];
     layer7_out[881] <= ~(layer6_out[911] | layer6_out[912]);
     layer7_out[882] <= layer6_out[1461];
     layer7_out[883] <= layer6_out[1115] ^ layer6_out[1116];
     layer7_out[884] <= ~layer6_out[615];
     layer7_out[885] <= ~layer6_out[1339];
     layer7_out[886] <= ~layer6_out[1379] | layer6_out[1380];
     layer7_out[887] <= ~layer6_out[1203];
     layer7_out[888] <= layer6_out[714] & layer6_out[715];
     layer7_out[889] <= ~(layer6_out[1012] | layer6_out[1013]);
     layer7_out[890] <= ~(layer6_out[63] ^ layer6_out[64]);
     layer7_out[891] <= layer6_out[1491] ^ layer6_out[1492];
     layer7_out[892] <= ~layer6_out[626];
     layer7_out[893] <= ~(layer6_out[448] | layer6_out[449]);
     layer7_out[894] <= ~layer6_out[531] | layer6_out[530];
     layer7_out[895] <= layer6_out[1392];
     layer7_out[896] <= layer6_out[1343] | layer6_out[1344];
     layer7_out[897] <= layer6_out[391];
     layer7_out[898] <= layer6_out[429] & ~layer6_out[430];
     layer7_out[899] <= layer6_out[1306];
     layer7_out[900] <= ~layer6_out[1349];
     layer7_out[901] <= layer6_out[523] & ~layer6_out[524];
     layer7_out[902] <= layer6_out[291];
     layer7_out[903] <= layer6_out[438];
     layer7_out[904] <= ~layer6_out[1216];
     layer7_out[905] <= layer6_out[73] & ~layer6_out[74];
     layer7_out[906] <= layer6_out[445];
     layer7_out[907] <= ~(layer6_out[1219] & layer6_out[1220]);
     layer7_out[908] <= layer6_out[1303];
     layer7_out[909] <= layer6_out[1460] & ~layer6_out[1459];
     layer7_out[910] <= ~layer6_out[436];
     layer7_out[911] <= ~(layer6_out[1316] ^ layer6_out[1317]);
     layer7_out[912] <= layer6_out[796] & ~layer6_out[795];
     layer7_out[913] <= ~layer6_out[148];
     layer7_out[914] <= layer6_out[682];
     layer7_out[915] <= ~(layer6_out[1350] & layer6_out[1351]);
     layer7_out[916] <= layer6_out[274] | layer6_out[275];
     layer7_out[917] <= layer6_out[1010];
     layer7_out[918] <= ~layer6_out[425];
     layer7_out[919] <= ~(layer6_out[1121] ^ layer6_out[1122]);
     layer7_out[920] <= ~(layer6_out[1479] ^ layer6_out[1480]);
     layer7_out[921] <= layer6_out[11] & ~layer6_out[10];
     layer7_out[922] <= layer6_out[742] & layer6_out[743];
     layer7_out[923] <= ~(layer6_out[1429] ^ layer6_out[1430]);
     layer7_out[924] <= ~(layer6_out[638] ^ layer6_out[639]);
     layer7_out[925] <= ~layer6_out[1468];
     layer7_out[926] <= layer6_out[1315] ^ layer6_out[1316];
     layer7_out[927] <= ~(layer6_out[189] ^ layer6_out[190]);
     layer7_out[928] <= ~(layer6_out[363] ^ layer6_out[364]);
     layer7_out[929] <= ~(layer6_out[1067] & layer6_out[1068]);
     layer7_out[930] <= layer6_out[1098];
     layer7_out[931] <= ~(layer6_out[326] | layer6_out[327]);
     layer7_out[932] <= layer6_out[991] & layer6_out[992];
     layer7_out[933] <= ~layer6_out[711];
     layer7_out[934] <= ~layer6_out[1282];
     layer7_out[935] <= layer6_out[331];
     layer7_out[936] <= layer6_out[1437];
     layer7_out[937] <= layer6_out[1413];
     layer7_out[938] <= ~(layer6_out[1373] | layer6_out[1374]);
     layer7_out[939] <= layer6_out[135] & ~layer6_out[134];
     layer7_out[940] <= layer6_out[702] ^ layer6_out[703];
     layer7_out[941] <= layer6_out[342] & ~layer6_out[343];
     layer7_out[942] <= layer6_out[865];
     layer7_out[943] <= layer6_out[605];
     layer7_out[944] <= layer6_out[274] & ~layer6_out[273];
     layer7_out[945] <= ~layer6_out[1367];
     layer7_out[946] <= ~layer6_out[1060] | layer6_out[1059];
     layer7_out[947] <= layer6_out[759] & ~layer6_out[760];
     layer7_out[948] <= ~layer6_out[221];
     layer7_out[949] <= layer6_out[819] & layer6_out[820];
     layer7_out[950] <= layer6_out[1184];
     layer7_out[951] <= ~layer6_out[348];
     layer7_out[952] <= ~(layer6_out[370] & layer6_out[371]);
     layer7_out[953] <= layer6_out[1147] ^ layer6_out[1148];
     layer7_out[954] <= ~(layer6_out[517] | layer6_out[518]);
     layer7_out[955] <= layer6_out[1021];
     layer7_out[956] <= layer6_out[628];
     layer7_out[957] <= layer6_out[1010] & layer6_out[1011];
     layer7_out[958] <= layer6_out[523] & ~layer6_out[522];
     layer7_out[959] <= layer6_out[457] & layer6_out[458];
     layer7_out[960] <= layer6_out[402] & layer6_out[403];
     layer7_out[961] <= layer6_out[90] & ~layer6_out[91];
     layer7_out[962] <= ~(layer6_out[897] ^ layer6_out[898]);
     layer7_out[963] <= ~layer6_out[677];
     layer7_out[964] <= layer6_out[325];
     layer7_out[965] <= layer6_out[244] & ~layer6_out[243];
     layer7_out[966] <= layer6_out[1280] ^ layer6_out[1281];
     layer7_out[967] <= layer6_out[1028] ^ layer6_out[1029];
     layer7_out[968] <= ~(layer6_out[1218] & layer6_out[1219]);
     layer7_out[969] <= layer6_out[293];
     layer7_out[970] <= ~(layer6_out[221] | layer6_out[222]);
     layer7_out[971] <= layer6_out[761] | layer6_out[762];
     layer7_out[972] <= ~layer6_out[231];
     layer7_out[973] <= layer6_out[1132];
     layer7_out[974] <= ~layer6_out[328];
     layer7_out[975] <= layer6_out[548];
     layer7_out[976] <= layer6_out[213] & ~layer6_out[214];
     layer7_out[977] <= ~layer6_out[276] | layer6_out[275];
     layer7_out[978] <= layer6_out[721] & layer6_out[722];
     layer7_out[979] <= layer6_out[465];
     layer7_out[980] <= layer6_out[359] & ~layer6_out[360];
     layer7_out[981] <= layer6_out[1085] & ~layer6_out[1086];
     layer7_out[982] <= layer6_out[427];
     layer7_out[983] <= layer6_out[947];
     layer7_out[984] <= ~(layer6_out[848] ^ layer6_out[849]);
     layer7_out[985] <= ~layer6_out[512];
     layer7_out[986] <= layer6_out[1478];
     layer7_out[987] <= layer6_out[180];
     layer7_out[988] <= layer6_out[1233] & ~layer6_out[1232];
     layer7_out[989] <= ~layer6_out[233];
     layer7_out[990] <= layer6_out[574];
     layer7_out[991] <= ~layer6_out[481];
     layer7_out[992] <= layer6_out[224] & ~layer6_out[223];
     layer7_out[993] <= layer6_out[1345] ^ layer6_out[1346];
     layer7_out[994] <= ~layer6_out[237];
     layer7_out[995] <= ~layer6_out[1307];
     layer7_out[996] <= layer6_out[372] | layer6_out[373];
     layer7_out[997] <= ~layer6_out[190];
     layer7_out[998] <= layer6_out[1476] & ~layer6_out[1477];
     layer7_out[999] <= layer6_out[312];
     layer7_out[1000] <= layer6_out[406];
     layer7_out[1001] <= ~(layer6_out[257] | layer6_out[258]);
     layer7_out[1002] <= layer6_out[631];
     layer7_out[1003] <= layer6_out[1240] & ~layer6_out[1241];
     layer7_out[1004] <= ~layer6_out[533];
     layer7_out[1005] <= ~(layer6_out[211] ^ layer6_out[212]);
     layer7_out[1006] <= layer6_out[1260];
     layer7_out[1007] <= layer6_out[42] ^ layer6_out[43];
     layer7_out[1008] <= ~layer6_out[1054];
     layer7_out[1009] <= layer6_out[931];
     layer7_out[1010] <= layer6_out[1081];
     layer7_out[1011] <= layer6_out[1160] & ~layer6_out[1159];
     layer7_out[1012] <= layer6_out[337] ^ layer6_out[338];
     layer7_out[1013] <= ~layer6_out[733];
     layer7_out[1014] <= layer6_out[798] & ~layer6_out[799];
     layer7_out[1015] <= layer6_out[525] & layer6_out[526];
     layer7_out[1016] <= ~layer6_out[81];
     layer7_out[1017] <= ~(layer6_out[217] | layer6_out[218]);
     layer7_out[1018] <= ~layer6_out[1182] | layer6_out[1183];
     layer7_out[1019] <= layer6_out[97];
     layer7_out[1020] <= ~(layer6_out[973] ^ layer6_out[974]);
     layer7_out[1021] <= layer6_out[682];
     layer7_out[1022] <= ~layer6_out[1074];
     layer7_out[1023] <= layer6_out[6];
     layer7_out[1024] <= layer6_out[395] & ~layer6_out[394];
     layer7_out[1025] <= layer6_out[1130];
     layer7_out[1026] <= ~layer6_out[708];
     layer7_out[1027] <= layer6_out[774];
     layer7_out[1028] <= layer6_out[1281] ^ layer6_out[1282];
     layer7_out[1029] <= layer6_out[1253] & ~layer6_out[1254];
     layer7_out[1030] <= layer6_out[1032] & ~layer6_out[1031];
     layer7_out[1031] <= ~layer6_out[225];
     layer7_out[1032] <= layer6_out[820] & ~layer6_out[821];
     layer7_out[1033] <= ~(layer6_out[340] ^ layer6_out[341]);
     layer7_out[1034] <= layer6_out[1410] & ~layer6_out[1409];
     layer7_out[1035] <= layer6_out[662] & ~layer6_out[663];
     layer7_out[1036] <= layer6_out[581];
     layer7_out[1037] <= layer6_out[972];
     layer7_out[1038] <= layer6_out[1021];
     layer7_out[1039] <= layer6_out[174] & layer6_out[175];
     layer7_out[1040] <= ~layer6_out[733];
     layer7_out[1041] <= layer6_out[869];
     layer7_out[1042] <= ~layer6_out[699];
     layer7_out[1043] <= layer6_out[490];
     layer7_out[1044] <= ~(layer6_out[1127] & layer6_out[1128]);
     layer7_out[1045] <= ~layer6_out[1298];
     layer7_out[1046] <= ~(layer6_out[172] | layer6_out[173]);
     layer7_out[1047] <= ~layer6_out[708];
     layer7_out[1048] <= ~layer6_out[486];
     layer7_out[1049] <= layer6_out[788];
     layer7_out[1050] <= ~layer6_out[653];
     layer7_out[1051] <= ~(layer6_out[1460] & layer6_out[1461]);
     layer7_out[1052] <= ~layer6_out[70];
     layer7_out[1053] <= layer6_out[397] | layer6_out[398];
     layer7_out[1054] <= layer6_out[512] & layer6_out[513];
     layer7_out[1055] <= layer6_out[955];
     layer7_out[1056] <= layer6_out[431] & layer6_out[432];
     layer7_out[1057] <= layer6_out[760] & ~layer6_out[761];
     layer7_out[1058] <= ~layer6_out[1119];
     layer7_out[1059] <= ~layer6_out[304];
     layer7_out[1060] <= ~layer6_out[933] | layer6_out[934];
     layer7_out[1061] <= ~layer6_out[477];
     layer7_out[1062] <= layer6_out[1149] & layer6_out[1150];
     layer7_out[1063] <= layer6_out[1465];
     layer7_out[1064] <= ~layer6_out[974] | layer6_out[975];
     layer7_out[1065] <= ~(layer6_out[1154] ^ layer6_out[1155]);
     layer7_out[1066] <= layer6_out[749];
     layer7_out[1067] <= layer6_out[315] ^ layer6_out[316];
     layer7_out[1068] <= ~layer6_out[354];
     layer7_out[1069] <= layer6_out[1137] ^ layer6_out[1138];
     layer7_out[1070] <= layer6_out[1066];
     layer7_out[1071] <= layer6_out[780];
     layer7_out[1072] <= ~layer6_out[587];
     layer7_out[1073] <= layer6_out[656] & ~layer6_out[657];
     layer7_out[1074] <= layer6_out[253];
     layer7_out[1075] <= ~layer6_out[620];
     layer7_out[1076] <= ~layer6_out[1189];
     layer7_out[1077] <= layer6_out[651] & ~layer6_out[650];
     layer7_out[1078] <= layer6_out[229] & ~layer6_out[228];
     layer7_out[1079] <= layer6_out[815] ^ layer6_out[816];
     layer7_out[1080] <= ~layer6_out[21];
     layer7_out[1081] <= layer6_out[1116] | layer6_out[1117];
     layer7_out[1082] <= layer6_out[1050] & layer6_out[1051];
     layer7_out[1083] <= layer6_out[809];
     layer7_out[1084] <= layer6_out[764] ^ layer6_out[765];
     layer7_out[1085] <= ~layer6_out[727];
     layer7_out[1086] <= ~layer6_out[819];
     layer7_out[1087] <= ~(layer6_out[1099] ^ layer6_out[1100]);
     layer7_out[1088] <= ~layer6_out[742];
     layer7_out[1089] <= ~layer6_out[920];
     layer7_out[1090] <= ~layer6_out[730] | layer6_out[729];
     layer7_out[1091] <= layer6_out[1400];
     layer7_out[1092] <= ~layer6_out[540];
     layer7_out[1093] <= layer6_out[288];
     layer7_out[1094] <= layer6_out[1205] & ~layer6_out[1206];
     layer7_out[1095] <= layer6_out[1357] & layer6_out[1358];
     layer7_out[1096] <= layer6_out[803] & ~layer6_out[802];
     layer7_out[1097] <= ~layer6_out[16];
     layer7_out[1098] <= ~layer6_out[1255];
     layer7_out[1099] <= ~(layer6_out[14] & layer6_out[15]);
     layer7_out[1100] <= layer6_out[1198] ^ layer6_out[1199];
     layer7_out[1101] <= ~layer6_out[572] | layer6_out[571];
     layer7_out[1102] <= ~layer6_out[235];
     layer7_out[1103] <= layer6_out[183] | layer6_out[184];
     layer7_out[1104] <= layer6_out[381];
     layer7_out[1105] <= ~(layer6_out[645] | layer6_out[646]);
     layer7_out[1106] <= layer6_out[977];
     layer7_out[1107] <= layer6_out[200];
     layer7_out[1108] <= ~layer6_out[604];
     layer7_out[1109] <= layer6_out[1273];
     layer7_out[1110] <= ~(layer6_out[338] ^ layer6_out[339]);
     layer7_out[1111] <= layer6_out[358];
     layer7_out[1112] <= ~(layer6_out[999] ^ layer6_out[1000]);
     layer7_out[1113] <= layer6_out[1424] & ~layer6_out[1423];
     layer7_out[1114] <= layer6_out[549] ^ layer6_out[550];
     layer7_out[1115] <= layer6_out[1165] & ~layer6_out[1164];
     layer7_out[1116] <= layer6_out[230] & ~layer6_out[231];
     layer7_out[1117] <= layer6_out[1376] & layer6_out[1377];
     layer7_out[1118] <= ~layer6_out[675];
     layer7_out[1119] <= layer6_out[1231];
     layer7_out[1120] <= layer6_out[1071] & layer6_out[1072];
     layer7_out[1121] <= layer6_out[1414] | layer6_out[1415];
     layer7_out[1122] <= layer6_out[44] & layer6_out[45];
     layer7_out[1123] <= ~layer6_out[1229];
     layer7_out[1124] <= layer6_out[1247] & ~layer6_out[1248];
     layer7_out[1125] <= layer6_out[941] & layer6_out[942];
     layer7_out[1126] <= layer6_out[1030] & layer6_out[1031];
     layer7_out[1127] <= layer6_out[229] & layer6_out[230];
     layer7_out[1128] <= ~layer6_out[402];
     layer7_out[1129] <= layer6_out[793];
     layer7_out[1130] <= layer6_out[217];
     layer7_out[1131] <= ~(layer6_out[31] ^ layer6_out[32]);
     layer7_out[1132] <= layer6_out[382];
     layer7_out[1133] <= ~(layer6_out[688] & layer6_out[689]);
     layer7_out[1134] <= ~layer6_out[342];
     layer7_out[1135] <= ~(layer6_out[1190] ^ layer6_out[1191]);
     layer7_out[1136] <= ~layer6_out[1191];
     layer7_out[1137] <= ~layer6_out[336];
     layer7_out[1138] <= ~layer6_out[688];
     layer7_out[1139] <= ~layer6_out[670];
     layer7_out[1140] <= ~layer6_out[1258];
     layer7_out[1141] <= ~layer6_out[727];
     layer7_out[1142] <= ~layer6_out[37];
     layer7_out[1143] <= layer6_out[68];
     layer7_out[1144] <= ~(layer6_out[1233] | layer6_out[1234]);
     layer7_out[1145] <= layer6_out[320] | layer6_out[321];
     layer7_out[1146] <= ~layer6_out[1320] | layer6_out[1319];
     layer7_out[1147] <= ~(layer6_out[71] & layer6_out[72]);
     layer7_out[1148] <= layer6_out[538] & ~layer6_out[539];
     layer7_out[1149] <= layer6_out[1100];
     layer7_out[1150] <= ~layer6_out[494];
     layer7_out[1151] <= layer6_out[683];
     layer7_out[1152] <= ~layer6_out[752] | layer6_out[753];
     layer7_out[1153] <= layer6_out[173] & layer6_out[174];
     layer7_out[1154] <= layer6_out[131] & layer6_out[132];
     layer7_out[1155] <= layer6_out[320];
     layer7_out[1156] <= layer6_out[488];
     layer7_out[1157] <= ~layer6_out[1229];
     layer7_out[1158] <= ~(layer6_out[101] & layer6_out[102]);
     layer7_out[1159] <= ~layer6_out[947];
     layer7_out[1160] <= layer6_out[767] ^ layer6_out[768];
     layer7_out[1161] <= layer6_out[1252] & ~layer6_out[1253];
     layer7_out[1162] <= layer6_out[117] | layer6_out[118];
     layer7_out[1163] <= layer6_out[1035];
     layer7_out[1164] <= ~(layer6_out[1242] & layer6_out[1243]);
     layer7_out[1165] <= layer6_out[1447];
     layer7_out[1166] <= ~layer6_out[1135];
     layer7_out[1167] <= ~(layer6_out[437] ^ layer6_out[438]);
     layer7_out[1168] <= layer6_out[1290] ^ layer6_out[1291];
     layer7_out[1169] <= ~layer6_out[536];
     layer7_out[1170] <= layer6_out[790];
     layer7_out[1171] <= layer6_out[1433];
     layer7_out[1172] <= ~layer6_out[1104];
     layer7_out[1173] <= ~layer6_out[171] | layer6_out[172];
     layer7_out[1174] <= layer6_out[1153] & layer6_out[1154];
     layer7_out[1175] <= layer6_out[896] ^ layer6_out[897];
     layer7_out[1176] <= ~(layer6_out[694] ^ layer6_out[695]);
     layer7_out[1177] <= layer6_out[1174] & ~layer6_out[1173];
     layer7_out[1178] <= ~(layer6_out[76] ^ layer6_out[77]);
     layer7_out[1179] <= layer6_out[195] & ~layer6_out[196];
     layer7_out[1180] <= ~(layer6_out[1084] ^ layer6_out[1085]);
     layer7_out[1181] <= ~layer6_out[1472];
     layer7_out[1182] <= layer6_out[803] ^ layer6_out[804];
     layer7_out[1183] <= layer6_out[56] & ~layer6_out[55];
     layer7_out[1184] <= layer6_out[1174] & layer6_out[1175];
     layer7_out[1185] <= ~layer6_out[551];
     layer7_out[1186] <= ~(layer6_out[559] | layer6_out[560]);
     layer7_out[1187] <= ~layer6_out[357] | layer6_out[358];
     layer7_out[1188] <= layer6_out[184];
     layer7_out[1189] <= layer6_out[44] & ~layer6_out[43];
     layer7_out[1190] <= ~(layer6_out[1128] ^ layer6_out[1129]);
     layer7_out[1191] <= layer6_out[404] ^ layer6_out[405];
     layer7_out[1192] <= layer6_out[1025];
     layer7_out[1193] <= ~layer6_out[1385];
     layer7_out[1194] <= layer6_out[960];
     layer7_out[1195] <= layer6_out[51];
     layer7_out[1196] <= ~layer6_out[966];
     layer7_out[1197] <= ~layer6_out[704];
     layer7_out[1198] <= layer6_out[301] & layer6_out[302];
     layer7_out[1199] <= ~(layer6_out[887] | layer6_out[888]);
     layer7_out[1200] <= ~layer6_out[1304];
     layer7_out[1201] <= ~layer6_out[1383];
     layer7_out[1202] <= ~(layer6_out[1488] ^ layer6_out[1489]);
     layer7_out[1203] <= ~(layer6_out[1494] & layer6_out[1495]);
     layer7_out[1204] <= layer6_out[1395];
     layer7_out[1205] <= ~layer6_out[355];
     layer7_out[1206] <= layer6_out[515];
     layer7_out[1207] <= layer6_out[1122] & ~layer6_out[1123];
     layer7_out[1208] <= ~layer6_out[904];
     layer7_out[1209] <= ~layer6_out[1415];
     layer7_out[1210] <= layer6_out[862];
     layer7_out[1211] <= ~layer6_out[1156];
     layer7_out[1212] <= ~layer6_out[1330];
     layer7_out[1213] <= ~(layer6_out[135] ^ layer6_out[136]);
     layer7_out[1214] <= ~layer6_out[652];
     layer7_out[1215] <= layer6_out[1106];
     layer7_out[1216] <= ~layer6_out[1040];
     layer7_out[1217] <= ~layer6_out[753];
     layer7_out[1218] <= layer6_out[1399];
     layer7_out[1219] <= layer6_out[1283] & ~layer6_out[1284];
     layer7_out[1220] <= ~layer6_out[1078];
     layer7_out[1221] <= ~layer6_out[1126];
     layer7_out[1222] <= layer6_out[849] ^ layer6_out[850];
     layer7_out[1223] <= ~layer6_out[642] | layer6_out[643];
     layer7_out[1224] <= ~layer6_out[1201];
     layer7_out[1225] <= layer6_out[535] ^ layer6_out[536];
     layer7_out[1226] <= layer6_out[35] & layer6_out[36];
     layer7_out[1227] <= layer6_out[368] & ~layer6_out[367];
     layer7_out[1228] <= layer6_out[1216] & layer6_out[1217];
     layer7_out[1229] <= ~layer6_out[1277];
     layer7_out[1230] <= layer6_out[1444] ^ layer6_out[1445];
     layer7_out[1231] <= ~layer6_out[266];
     layer7_out[1232] <= ~(layer6_out[972] & layer6_out[973]);
     layer7_out[1233] <= ~layer6_out[726];
     layer7_out[1234] <= layer6_out[730] ^ layer6_out[731];
     layer7_out[1235] <= ~layer6_out[927];
     layer7_out[1236] <= layer6_out[832];
     layer7_out[1237] <= ~(layer6_out[597] & layer6_out[598]);
     layer7_out[1238] <= ~(layer6_out[368] ^ layer6_out[369]);
     layer7_out[1239] <= layer6_out[841];
     layer7_out[1240] <= layer6_out[178] & layer6_out[179];
     layer7_out[1241] <= ~layer6_out[486] | layer6_out[487];
     layer7_out[1242] <= layer6_out[801] & layer6_out[802];
     layer7_out[1243] <= ~layer6_out[269] | layer6_out[270];
     layer7_out[1244] <= ~(layer6_out[1023] ^ layer6_out[1024]);
     layer7_out[1245] <= layer6_out[5] & ~layer6_out[4];
     layer7_out[1246] <= ~layer6_out[925];
     layer7_out[1247] <= layer6_out[817];
     layer7_out[1248] <= layer6_out[541];
     layer7_out[1249] <= ~(layer6_out[1227] | layer6_out[1228]);
     layer7_out[1250] <= ~layer6_out[195] | layer6_out[194];
     layer7_out[1251] <= ~(layer6_out[799] & layer6_out[800]);
     layer7_out[1252] <= ~(layer6_out[113] ^ layer6_out[114]);
     layer7_out[1253] <= ~(layer6_out[796] & layer6_out[797]);
     layer7_out[1254] <= layer6_out[54] ^ layer6_out[55];
     layer7_out[1255] <= layer6_out[491] & ~layer6_out[490];
     layer7_out[1256] <= layer6_out[45] & ~layer6_out[46];
     layer7_out[1257] <= layer6_out[587];
     layer7_out[1258] <= ~layer6_out[168];
     layer7_out[1259] <= ~layer6_out[944];
     layer7_out[1260] <= layer6_out[579] ^ layer6_out[580];
     layer7_out[1261] <= layer6_out[408] & ~layer6_out[407];
     layer7_out[1262] <= layer6_out[144] & layer6_out[145];
     layer7_out[1263] <= layer6_out[964] & ~layer6_out[963];
     layer7_out[1264] <= ~layer6_out[1353];
     layer7_out[1265] <= layer6_out[348];
     layer7_out[1266] <= layer6_out[522] & ~layer6_out[521];
     layer7_out[1267] <= ~layer6_out[633] | layer6_out[632];
     layer7_out[1268] <= layer6_out[160] & layer6_out[161];
     layer7_out[1269] <= ~layer6_out[1023];
     layer7_out[1270] <= layer6_out[1381];
     layer7_out[1271] <= layer6_out[381] ^ layer6_out[382];
     layer7_out[1272] <= layer6_out[596] & ~layer6_out[595];
     layer7_out[1273] <= ~layer6_out[838];
     layer7_out[1274] <= ~layer6_out[287];
     layer7_out[1275] <= layer6_out[712];
     layer7_out[1276] <= ~layer6_out[1454];
     layer7_out[1277] <= ~layer6_out[1078];
     layer7_out[1278] <= layer6_out[985];
     layer7_out[1279] <= ~(layer6_out[331] | layer6_out[332]);
     layer7_out[1280] <= ~layer6_out[322];
     layer7_out[1281] <= ~layer6_out[779];
     layer7_out[1282] <= ~(layer6_out[1497] ^ layer6_out[1498]);
     layer7_out[1283] <= ~layer6_out[1369];
     layer7_out[1284] <= layer6_out[1007] ^ layer6_out[1008];
     layer7_out[1285] <= ~layer6_out[1090] | layer6_out[1091];
     layer7_out[1286] <= ~layer6_out[886] | layer6_out[885];
     layer7_out[1287] <= ~layer6_out[1446] | layer6_out[1445];
     layer7_out[1288] <= layer6_out[1164];
     layer7_out[1289] <= ~layer6_out[1124] | layer6_out[1125];
     layer7_out[1290] <= ~(layer6_out[576] ^ layer6_out[577]);
     layer7_out[1291] <= ~layer6_out[728];
     layer7_out[1292] <= layer6_out[585] ^ layer6_out[586];
     layer7_out[1293] <= layer6_out[566] & ~layer6_out[567];
     layer7_out[1294] <= layer6_out[1486];
     layer7_out[1295] <= layer6_out[889];
     layer7_out[1296] <= ~layer6_out[777];
     layer7_out[1297] <= layer6_out[1374] ^ layer6_out[1375];
     layer7_out[1298] <= layer6_out[847] ^ layer6_out[848];
     layer7_out[1299] <= ~(layer6_out[1111] | layer6_out[1112]);
     layer7_out[1300] <= ~layer6_out[414];
     layer7_out[1301] <= layer6_out[100] & layer6_out[101];
     layer7_out[1302] <= layer6_out[1458];
     layer7_out[1303] <= layer6_out[697];
     layer7_out[1304] <= layer6_out[280];
     layer7_out[1305] <= ~(layer6_out[628] ^ layer6_out[629]);
     layer7_out[1306] <= layer6_out[1224];
     layer7_out[1307] <= layer6_out[1412] ^ layer6_out[1413];
     layer7_out[1308] <= layer6_out[52] & ~layer6_out[53];
     layer7_out[1309] <= ~layer6_out[901];
     layer7_out[1310] <= layer6_out[493] & layer6_out[494];
     layer7_out[1311] <= ~layer6_out[121];
     layer7_out[1312] <= ~layer6_out[130];
     layer7_out[1313] <= layer6_out[967];
     layer7_out[1314] <= layer6_out[350] & ~layer6_out[351];
     layer7_out[1315] <= layer6_out[1381];
     layer7_out[1316] <= ~(layer6_out[119] ^ layer6_out[120]);
     layer7_out[1317] <= ~layer6_out[1417];
     layer7_out[1318] <= ~layer6_out[983] | layer6_out[984];
     layer7_out[1319] <= layer6_out[1436] ^ layer6_out[1437];
     layer7_out[1320] <= ~layer6_out[445];
     layer7_out[1321] <= layer6_out[201] | layer6_out[202];
     layer7_out[1322] <= layer6_out[641] & ~layer6_out[642];
     layer7_out[1323] <= layer6_out[441] & layer6_out[442];
     layer7_out[1324] <= layer6_out[144] & ~layer6_out[143];
     layer7_out[1325] <= ~(layer6_out[858] | layer6_out[859]);
     layer7_out[1326] <= layer6_out[151] & ~layer6_out[150];
     layer7_out[1327] <= ~(layer6_out[1324] & layer6_out[1325]);
     layer7_out[1328] <= ~layer6_out[960] | layer6_out[961];
     layer7_out[1329] <= layer6_out[623] & ~layer6_out[622];
     layer7_out[1330] <= ~layer6_out[238] | layer6_out[239];
     layer7_out[1331] <= layer6_out[850] ^ layer6_out[851];
     layer7_out[1332] <= ~layer6_out[106];
     layer7_out[1333] <= layer6_out[1217] & layer6_out[1218];
     layer7_out[1334] <= layer6_out[205] & ~layer6_out[204];
     layer7_out[1335] <= ~layer6_out[65] | layer6_out[66];
     layer7_out[1336] <= ~(layer6_out[158] ^ layer6_out[159]);
     layer7_out[1337] <= layer6_out[1328];
     layer7_out[1338] <= ~layer6_out[648];
     layer7_out[1339] <= layer6_out[1162] ^ layer6_out[1163];
     layer7_out[1340] <= ~(layer6_out[186] | layer6_out[187]);
     layer7_out[1341] <= layer6_out[1356] ^ layer6_out[1357];
     layer7_out[1342] <= layer6_out[1237];
     layer7_out[1343] <= layer6_out[188];
     layer7_out[1344] <= ~layer6_out[108];
     layer7_out[1345] <= layer6_out[705];
     layer7_out[1346] <= ~(layer6_out[48] ^ layer6_out[49]);
     layer7_out[1347] <= ~layer6_out[1364];
     layer7_out[1348] <= ~(layer6_out[166] ^ layer6_out[167]);
     layer7_out[1349] <= ~layer6_out[652];
     layer7_out[1350] <= ~layer6_out[950];
     layer7_out[1351] <= ~(layer6_out[1403] | layer6_out[1404]);
     layer7_out[1352] <= layer6_out[790];
     layer7_out[1353] <= ~layer6_out[948] | layer6_out[949];
     layer7_out[1354] <= ~(layer6_out[921] ^ layer6_out[922]);
     layer7_out[1355] <= ~layer6_out[647] | layer6_out[646];
     layer7_out[1356] <= layer6_out[1072] & ~layer6_out[1073];
     layer7_out[1357] <= layer6_out[1186] & ~layer6_out[1187];
     layer7_out[1358] <= ~(layer6_out[1018] | layer6_out[1019]);
     layer7_out[1359] <= ~(layer6_out[812] & layer6_out[813]);
     layer7_out[1360] <= ~layer6_out[633];
     layer7_out[1361] <= ~(layer6_out[879] | layer6_out[880]);
     layer7_out[1362] <= ~layer6_out[1157];
     layer7_out[1363] <= ~layer6_out[206];
     layer7_out[1364] <= ~layer6_out[928];
     layer7_out[1365] <= layer6_out[259];
     layer7_out[1366] <= layer6_out[673];
     layer7_out[1367] <= layer6_out[1224];
     layer7_out[1368] <= ~(layer6_out[1452] ^ layer6_out[1453]);
     layer7_out[1369] <= ~(layer6_out[997] | layer6_out[998]);
     layer7_out[1370] <= layer6_out[763] & ~layer6_out[762];
     layer7_out[1371] <= layer6_out[28] & ~layer6_out[29];
     layer7_out[1372] <= ~layer6_out[164];
     layer7_out[1373] <= ~(layer6_out[1117] ^ layer6_out[1118]);
     layer7_out[1374] <= ~(layer6_out[1212] ^ layer6_out[1213]);
     layer7_out[1375] <= ~layer6_out[294];
     layer7_out[1376] <= layer6_out[1004];
     layer7_out[1377] <= layer6_out[145] ^ layer6_out[146];
     layer7_out[1378] <= ~layer6_out[414];
     layer7_out[1379] <= layer6_out[1474] & ~layer6_out[1473];
     layer7_out[1380] <= layer6_out[808] ^ layer6_out[809];
     layer7_out[1381] <= layer6_out[1426] & layer6_out[1427];
     layer7_out[1382] <= layer6_out[1075];
     layer7_out[1383] <= ~layer6_out[1178];
     layer7_out[1384] <= layer6_out[24];
     layer7_out[1385] <= ~layer6_out[459];
     layer7_out[1386] <= ~(layer6_out[836] & layer6_out[837]);
     layer7_out[1387] <= layer6_out[23] & ~layer6_out[22];
     layer7_out[1388] <= layer6_out[389];
     layer7_out[1389] <= layer6_out[952];
     layer7_out[1390] <= layer6_out[1113] & ~layer6_out[1112];
     layer7_out[1391] <= layer6_out[102];
     layer7_out[1392] <= layer6_out[607];
     layer7_out[1393] <= ~(layer6_out[1083] | layer6_out[1084]);
     layer7_out[1394] <= ~(layer6_out[598] ^ layer6_out[599]);
     layer7_out[1395] <= layer6_out[927] & ~layer6_out[928];
     layer7_out[1396] <= ~(layer6_out[1318] | layer6_out[1319]);
     layer7_out[1397] <= ~layer6_out[923];
     layer7_out[1398] <= ~layer6_out[1152];
     layer7_out[1399] <= layer6_out[1052];
     layer7_out[1400] <= layer6_out[397];
     layer7_out[1401] <= layer6_out[1355];
     layer7_out[1402] <= layer6_out[298] & layer6_out[299];
     layer7_out[1403] <= ~(layer6_out[1396] | layer6_out[1397]);
     layer7_out[1404] <= layer6_out[178];
     layer7_out[1405] <= layer6_out[1149] & ~layer6_out[1148];
     layer7_out[1406] <= ~layer6_out[811];
     layer7_out[1407] <= layer6_out[870];
     layer7_out[1408] <= ~(layer6_out[744] ^ layer6_out[745]);
     layer7_out[1409] <= layer6_out[1027];
     layer7_out[1410] <= ~layer6_out[811];
     layer7_out[1411] <= ~(layer6_out[215] ^ layer6_out[216]);
     layer7_out[1412] <= layer6_out[1113] | layer6_out[1114];
     layer7_out[1413] <= layer6_out[1484] ^ layer6_out[1485];
     layer7_out[1414] <= layer6_out[666] & ~layer6_out[665];
     layer7_out[1415] <= layer6_out[993] ^ layer6_out[994];
     layer7_out[1416] <= ~(layer6_out[1156] | layer6_out[1157]);
     layer7_out[1417] <= ~layer6_out[1207];
     layer7_out[1418] <= layer6_out[954];
     layer7_out[1419] <= layer6_out[481];
     layer7_out[1420] <= ~(layer6_out[903] | layer6_out[904]);
     layer7_out[1421] <= layer6_out[292] & ~layer6_out[293];
     layer7_out[1422] <= ~layer6_out[706];
     layer7_out[1423] <= layer6_out[599];
     layer7_out[1424] <= ~layer6_out[473];
     layer7_out[1425] <= ~(layer6_out[484] | layer6_out[485]);
     layer7_out[1426] <= layer6_out[669] & ~layer6_out[668];
     layer7_out[1427] <= layer6_out[1343];
     layer7_out[1428] <= layer6_out[750];
     layer7_out[1429] <= layer6_out[143] & ~layer6_out[142];
     layer7_out[1430] <= layer6_out[528];
     layer7_out[1431] <= layer6_out[1475];
     layer7_out[1432] <= layer6_out[1332] & ~layer6_out[1333];
     layer7_out[1433] <= ~layer6_out[199];
     layer7_out[1434] <= ~layer6_out[1006];
     layer7_out[1435] <= ~layer6_out[304];
     layer7_out[1436] <= layer6_out[147];
     layer7_out[1437] <= ~(layer6_out[277] | layer6_out[278]);
     layer7_out[1438] <= layer6_out[140] & ~layer6_out[141];
     layer7_out[1439] <= layer6_out[1278];
     layer7_out[1440] <= layer6_out[26];
     layer7_out[1441] <= layer6_out[88];
     layer7_out[1442] <= layer6_out[1044];
     layer7_out[1443] <= layer6_out[827];
     layer7_out[1444] <= ~(layer6_out[453] | layer6_out[454]);
     layer7_out[1445] <= layer6_out[313] ^ layer6_out[314];
     layer7_out[1446] <= layer6_out[256];
     layer7_out[1447] <= ~(layer6_out[609] | layer6_out[610]);
     layer7_out[1448] <= layer6_out[840] & layer6_out[841];
     layer7_out[1449] <= ~layer6_out[736];
     layer7_out[1450] <= layer6_out[1265];
     layer7_out[1451] <= layer6_out[1490] & ~layer6_out[1489];
     layer7_out[1452] <= layer6_out[1438];
     layer7_out[1453] <= layer6_out[724] & layer6_out[725];
     layer7_out[1454] <= layer6_out[1497] & ~layer6_out[1496];
     layer7_out[1455] <= layer6_out[422];
     layer7_out[1456] <= layer6_out[962];
     layer7_out[1457] <= layer6_out[656] & ~layer6_out[655];
     layer7_out[1458] <= layer6_out[737] & ~layer6_out[736];
     layer7_out[1459] <= layer6_out[362] ^ layer6_out[363];
     layer7_out[1460] <= layer6_out[985];
     layer7_out[1461] <= ~layer6_out[943];
     layer7_out[1462] <= layer6_out[374] & layer6_out[375];
     layer7_out[1463] <= layer6_out[116] ^ layer6_out[117];
     layer7_out[1464] <= ~(layer6_out[1195] | layer6_out[1196]);
     layer7_out[1465] <= layer6_out[466] & layer6_out[467];
     layer7_out[1466] <= ~layer6_out[206];
     layer7_out[1467] <= ~layer6_out[829];
     layer7_out[1468] <= ~(layer6_out[876] & layer6_out[877]);
     layer7_out[1469] <= ~layer6_out[4];
     layer7_out[1470] <= layer6_out[1431] & ~layer6_out[1432];
     layer7_out[1471] <= layer6_out[401];
     layer7_out[1472] <= ~(layer6_out[902] ^ layer6_out[903]);
     layer7_out[1473] <= layer6_out[896];
     layer7_out[1474] <= layer6_out[197] & ~layer6_out[196];
     layer7_out[1475] <= layer6_out[1416] & ~layer6_out[1417];
     layer7_out[1476] <= layer6_out[1165] | layer6_out[1166];
     layer7_out[1477] <= layer6_out[1225] ^ layer6_out[1226];
     layer7_out[1478] <= layer6_out[350];
     layer7_out[1479] <= ~(layer6_out[684] & layer6_out[685]);
     layer7_out[1480] <= ~layer6_out[18];
     layer7_out[1481] <= layer6_out[1108] & ~layer6_out[1107];
     layer7_out[1482] <= layer6_out[939];
     layer7_out[1483] <= layer6_out[1486] ^ layer6_out[1487];
     layer7_out[1484] <= layer6_out[121] | layer6_out[122];
     layer7_out[1485] <= layer6_out[737] & ~layer6_out[738];
     layer7_out[1486] <= ~layer6_out[732];
     layer7_out[1487] <= ~layer6_out[589];
     layer7_out[1488] <= layer6_out[96] & ~layer6_out[95];
     layer7_out[1489] <= layer6_out[1030] & ~layer6_out[1029];
     layer7_out[1490] <= ~layer6_out[109];
     layer7_out[1491] <= ~(layer6_out[664] | layer6_out[665]);
     layer7_out[1492] <= layer6_out[554];
     layer7_out[1493] <= layer6_out[1336];
     layer7_out[1494] <= layer6_out[517];
     layer7_out[1495] <= ~(layer6_out[957] & layer6_out[958]);
     layer7_out[1496] <= layer6_out[140];
     layer7_out[1497] <= layer6_out[1027];
     layer7_out[1498] <= layer6_out[1495] ^ layer6_out[1496];
     layer7_out[1499] <= ~layer6_out[430];
      last_layer_output <= layer7_out;

      result[0] <= last_layer_output[0] + last_layer_output[1] + last_layer_output[2] + last_layer_output[3] + last_layer_output[4] + last_layer_output[5] + last_layer_output[6] + last_layer_output[7] + last_layer_output[8] + last_layer_output[9] + last_layer_output[10] + last_layer_output[11] + last_layer_output[12] + last_layer_output[13] + last_layer_output[14] + last_layer_output[15] + last_layer_output[16] + last_layer_output[17] + last_layer_output[18] + last_layer_output[19] + last_layer_output[20] + last_layer_output[21] + last_layer_output[22] + last_layer_output[23] + last_layer_output[24] + last_layer_output[25] + last_layer_output[26] + last_layer_output[27] + last_layer_output[28] + last_layer_output[29] + last_layer_output[30] + last_layer_output[31] + last_layer_output[32] + last_layer_output[33] + last_layer_output[34] + last_layer_output[35] + last_layer_output[36] + last_layer_output[37] + last_layer_output[38] + last_layer_output[39] + last_layer_output[40] + last_layer_output[41] + last_layer_output[42] + last_layer_output[43] + last_layer_output[44] + last_layer_output[45] + last_layer_output[46] + last_layer_output[47] + last_layer_output[48] + last_layer_output[49] + last_layer_output[50] + last_layer_output[51] + last_layer_output[52] + last_layer_output[53] + last_layer_output[54] + last_layer_output[55] + last_layer_output[56] + last_layer_output[57] + last_layer_output[58] + last_layer_output[59] + last_layer_output[60] + last_layer_output[61] + last_layer_output[62] + last_layer_output[63] + last_layer_output[64] + last_layer_output[65] + last_layer_output[66] + last_layer_output[67] + last_layer_output[68] + last_layer_output[69] + last_layer_output[70] + last_layer_output[71] + last_layer_output[72] + last_layer_output[73] + last_layer_output[74] + last_layer_output[75] + last_layer_output[76] + last_layer_output[77] + last_layer_output[78] + last_layer_output[79] + last_layer_output[80] + last_layer_output[81] + last_layer_output[82] + last_layer_output[83] + last_layer_output[84] + last_layer_output[85] + last_layer_output[86] + last_layer_output[87] + last_layer_output[88] + last_layer_output[89] + last_layer_output[90] + last_layer_output[91] + last_layer_output[92] + last_layer_output[93] + last_layer_output[94] + last_layer_output[95] + last_layer_output[96] + last_layer_output[97] + last_layer_output[98] + last_layer_output[99] + last_layer_output[100] + last_layer_output[101] + last_layer_output[102] + last_layer_output[103] + last_layer_output[104] + last_layer_output[105] + last_layer_output[106] + last_layer_output[107] + last_layer_output[108] + last_layer_output[109] + last_layer_output[110] + last_layer_output[111] + last_layer_output[112] + last_layer_output[113] + last_layer_output[114] + last_layer_output[115] + last_layer_output[116] + last_layer_output[117] + last_layer_output[118] + last_layer_output[119] + last_layer_output[120] + last_layer_output[121] + last_layer_output[122] + last_layer_output[123] + last_layer_output[124] + last_layer_output[125] + last_layer_output[126] + last_layer_output[127] + last_layer_output[128] + last_layer_output[129] + last_layer_output[130] + last_layer_output[131] + last_layer_output[132] + last_layer_output[133] + last_layer_output[134] + last_layer_output[135] + last_layer_output[136] + last_layer_output[137] + last_layer_output[138] + last_layer_output[139] + last_layer_output[140] + last_layer_output[141] + last_layer_output[142] + last_layer_output[143] + last_layer_output[144] + last_layer_output[145] + last_layer_output[146] + last_layer_output[147] + last_layer_output[148] + last_layer_output[149];
      result[1] <= last_layer_output[150] + last_layer_output[151] + last_layer_output[152] + last_layer_output[153] + last_layer_output[154] + last_layer_output[155] + last_layer_output[156] + last_layer_output[157] + last_layer_output[158] + last_layer_output[159] + last_layer_output[160] + last_layer_output[161] + last_layer_output[162] + last_layer_output[163] + last_layer_output[164] + last_layer_output[165] + last_layer_output[166] + last_layer_output[167] + last_layer_output[168] + last_layer_output[169] + last_layer_output[170] + last_layer_output[171] + last_layer_output[172] + last_layer_output[173] + last_layer_output[174] + last_layer_output[175] + last_layer_output[176] + last_layer_output[177] + last_layer_output[178] + last_layer_output[179] + last_layer_output[180] + last_layer_output[181] + last_layer_output[182] + last_layer_output[183] + last_layer_output[184] + last_layer_output[185] + last_layer_output[186] + last_layer_output[187] + last_layer_output[188] + last_layer_output[189] + last_layer_output[190] + last_layer_output[191] + last_layer_output[192] + last_layer_output[193] + last_layer_output[194] + last_layer_output[195] + last_layer_output[196] + last_layer_output[197] + last_layer_output[198] + last_layer_output[199] + last_layer_output[200] + last_layer_output[201] + last_layer_output[202] + last_layer_output[203] + last_layer_output[204] + last_layer_output[205] + last_layer_output[206] + last_layer_output[207] + last_layer_output[208] + last_layer_output[209] + last_layer_output[210] + last_layer_output[211] + last_layer_output[212] + last_layer_output[213] + last_layer_output[214] + last_layer_output[215] + last_layer_output[216] + last_layer_output[217] + last_layer_output[218] + last_layer_output[219] + last_layer_output[220] + last_layer_output[221] + last_layer_output[222] + last_layer_output[223] + last_layer_output[224] + last_layer_output[225] + last_layer_output[226] + last_layer_output[227] + last_layer_output[228] + last_layer_output[229] + last_layer_output[230] + last_layer_output[231] + last_layer_output[232] + last_layer_output[233] + last_layer_output[234] + last_layer_output[235] + last_layer_output[236] + last_layer_output[237] + last_layer_output[238] + last_layer_output[239] + last_layer_output[240] + last_layer_output[241] + last_layer_output[242] + last_layer_output[243] + last_layer_output[244] + last_layer_output[245] + last_layer_output[246] + last_layer_output[247] + last_layer_output[248] + last_layer_output[249] + last_layer_output[250] + last_layer_output[251] + last_layer_output[252] + last_layer_output[253] + last_layer_output[254] + last_layer_output[255] + last_layer_output[256] + last_layer_output[257] + last_layer_output[258] + last_layer_output[259] + last_layer_output[260] + last_layer_output[261] + last_layer_output[262] + last_layer_output[263] + last_layer_output[264] + last_layer_output[265] + last_layer_output[266] + last_layer_output[267] + last_layer_output[268] + last_layer_output[269] + last_layer_output[270] + last_layer_output[271] + last_layer_output[272] + last_layer_output[273] + last_layer_output[274] + last_layer_output[275] + last_layer_output[276] + last_layer_output[277] + last_layer_output[278] + last_layer_output[279] + last_layer_output[280] + last_layer_output[281] + last_layer_output[282] + last_layer_output[283] + last_layer_output[284] + last_layer_output[285] + last_layer_output[286] + last_layer_output[287] + last_layer_output[288] + last_layer_output[289] + last_layer_output[290] + last_layer_output[291] + last_layer_output[292] + last_layer_output[293] + last_layer_output[294] + last_layer_output[295] + last_layer_output[296] + last_layer_output[297] + last_layer_output[298] + last_layer_output[299];
      result[2] <= last_layer_output[300] + last_layer_output[301] + last_layer_output[302] + last_layer_output[303] + last_layer_output[304] + last_layer_output[305] + last_layer_output[306] + last_layer_output[307] + last_layer_output[308] + last_layer_output[309] + last_layer_output[310] + last_layer_output[311] + last_layer_output[312] + last_layer_output[313] + last_layer_output[314] + last_layer_output[315] + last_layer_output[316] + last_layer_output[317] + last_layer_output[318] + last_layer_output[319] + last_layer_output[320] + last_layer_output[321] + last_layer_output[322] + last_layer_output[323] + last_layer_output[324] + last_layer_output[325] + last_layer_output[326] + last_layer_output[327] + last_layer_output[328] + last_layer_output[329] + last_layer_output[330] + last_layer_output[331] + last_layer_output[332] + last_layer_output[333] + last_layer_output[334] + last_layer_output[335] + last_layer_output[336] + last_layer_output[337] + last_layer_output[338] + last_layer_output[339] + last_layer_output[340] + last_layer_output[341] + last_layer_output[342] + last_layer_output[343] + last_layer_output[344] + last_layer_output[345] + last_layer_output[346] + last_layer_output[347] + last_layer_output[348] + last_layer_output[349] + last_layer_output[350] + last_layer_output[351] + last_layer_output[352] + last_layer_output[353] + last_layer_output[354] + last_layer_output[355] + last_layer_output[356] + last_layer_output[357] + last_layer_output[358] + last_layer_output[359] + last_layer_output[360] + last_layer_output[361] + last_layer_output[362] + last_layer_output[363] + last_layer_output[364] + last_layer_output[365] + last_layer_output[366] + last_layer_output[367] + last_layer_output[368] + last_layer_output[369] + last_layer_output[370] + last_layer_output[371] + last_layer_output[372] + last_layer_output[373] + last_layer_output[374] + last_layer_output[375] + last_layer_output[376] + last_layer_output[377] + last_layer_output[378] + last_layer_output[379] + last_layer_output[380] + last_layer_output[381] + last_layer_output[382] + last_layer_output[383] + last_layer_output[384] + last_layer_output[385] + last_layer_output[386] + last_layer_output[387] + last_layer_output[388] + last_layer_output[389] + last_layer_output[390] + last_layer_output[391] + last_layer_output[392] + last_layer_output[393] + last_layer_output[394] + last_layer_output[395] + last_layer_output[396] + last_layer_output[397] + last_layer_output[398] + last_layer_output[399] + last_layer_output[400] + last_layer_output[401] + last_layer_output[402] + last_layer_output[403] + last_layer_output[404] + last_layer_output[405] + last_layer_output[406] + last_layer_output[407] + last_layer_output[408] + last_layer_output[409] + last_layer_output[410] + last_layer_output[411] + last_layer_output[412] + last_layer_output[413] + last_layer_output[414] + last_layer_output[415] + last_layer_output[416] + last_layer_output[417] + last_layer_output[418] + last_layer_output[419] + last_layer_output[420] + last_layer_output[421] + last_layer_output[422] + last_layer_output[423] + last_layer_output[424] + last_layer_output[425] + last_layer_output[426] + last_layer_output[427] + last_layer_output[428] + last_layer_output[429] + last_layer_output[430] + last_layer_output[431] + last_layer_output[432] + last_layer_output[433] + last_layer_output[434] + last_layer_output[435] + last_layer_output[436] + last_layer_output[437] + last_layer_output[438] + last_layer_output[439] + last_layer_output[440] + last_layer_output[441] + last_layer_output[442] + last_layer_output[443] + last_layer_output[444] + last_layer_output[445] + last_layer_output[446] + last_layer_output[447] + last_layer_output[448] + last_layer_output[449];
      result[3] <= last_layer_output[450] + last_layer_output[451] + last_layer_output[452] + last_layer_output[453] + last_layer_output[454] + last_layer_output[455] + last_layer_output[456] + last_layer_output[457] + last_layer_output[458] + last_layer_output[459] + last_layer_output[460] + last_layer_output[461] + last_layer_output[462] + last_layer_output[463] + last_layer_output[464] + last_layer_output[465] + last_layer_output[466] + last_layer_output[467] + last_layer_output[468] + last_layer_output[469] + last_layer_output[470] + last_layer_output[471] + last_layer_output[472] + last_layer_output[473] + last_layer_output[474] + last_layer_output[475] + last_layer_output[476] + last_layer_output[477] + last_layer_output[478] + last_layer_output[479] + last_layer_output[480] + last_layer_output[481] + last_layer_output[482] + last_layer_output[483] + last_layer_output[484] + last_layer_output[485] + last_layer_output[486] + last_layer_output[487] + last_layer_output[488] + last_layer_output[489] + last_layer_output[490] + last_layer_output[491] + last_layer_output[492] + last_layer_output[493] + last_layer_output[494] + last_layer_output[495] + last_layer_output[496] + last_layer_output[497] + last_layer_output[498] + last_layer_output[499] + last_layer_output[500] + last_layer_output[501] + last_layer_output[502] + last_layer_output[503] + last_layer_output[504] + last_layer_output[505] + last_layer_output[506] + last_layer_output[507] + last_layer_output[508] + last_layer_output[509] + last_layer_output[510] + last_layer_output[511] + last_layer_output[512] + last_layer_output[513] + last_layer_output[514] + last_layer_output[515] + last_layer_output[516] + last_layer_output[517] + last_layer_output[518] + last_layer_output[519] + last_layer_output[520] + last_layer_output[521] + last_layer_output[522] + last_layer_output[523] + last_layer_output[524] + last_layer_output[525] + last_layer_output[526] + last_layer_output[527] + last_layer_output[528] + last_layer_output[529] + last_layer_output[530] + last_layer_output[531] + last_layer_output[532] + last_layer_output[533] + last_layer_output[534] + last_layer_output[535] + last_layer_output[536] + last_layer_output[537] + last_layer_output[538] + last_layer_output[539] + last_layer_output[540] + last_layer_output[541] + last_layer_output[542] + last_layer_output[543] + last_layer_output[544] + last_layer_output[545] + last_layer_output[546] + last_layer_output[547] + last_layer_output[548] + last_layer_output[549] + last_layer_output[550] + last_layer_output[551] + last_layer_output[552] + last_layer_output[553] + last_layer_output[554] + last_layer_output[555] + last_layer_output[556] + last_layer_output[557] + last_layer_output[558] + last_layer_output[559] + last_layer_output[560] + last_layer_output[561] + last_layer_output[562] + last_layer_output[563] + last_layer_output[564] + last_layer_output[565] + last_layer_output[566] + last_layer_output[567] + last_layer_output[568] + last_layer_output[569] + last_layer_output[570] + last_layer_output[571] + last_layer_output[572] + last_layer_output[573] + last_layer_output[574] + last_layer_output[575] + last_layer_output[576] + last_layer_output[577] + last_layer_output[578] + last_layer_output[579] + last_layer_output[580] + last_layer_output[581] + last_layer_output[582] + last_layer_output[583] + last_layer_output[584] + last_layer_output[585] + last_layer_output[586] + last_layer_output[587] + last_layer_output[588] + last_layer_output[589] + last_layer_output[590] + last_layer_output[591] + last_layer_output[592] + last_layer_output[593] + last_layer_output[594] + last_layer_output[595] + last_layer_output[596] + last_layer_output[597] + last_layer_output[598] + last_layer_output[599];
      result[4] <= last_layer_output[600] + last_layer_output[601] + last_layer_output[602] + last_layer_output[603] + last_layer_output[604] + last_layer_output[605] + last_layer_output[606] + last_layer_output[607] + last_layer_output[608] + last_layer_output[609] + last_layer_output[610] + last_layer_output[611] + last_layer_output[612] + last_layer_output[613] + last_layer_output[614] + last_layer_output[615] + last_layer_output[616] + last_layer_output[617] + last_layer_output[618] + last_layer_output[619] + last_layer_output[620] + last_layer_output[621] + last_layer_output[622] + last_layer_output[623] + last_layer_output[624] + last_layer_output[625] + last_layer_output[626] + last_layer_output[627] + last_layer_output[628] + last_layer_output[629] + last_layer_output[630] + last_layer_output[631] + last_layer_output[632] + last_layer_output[633] + last_layer_output[634] + last_layer_output[635] + last_layer_output[636] + last_layer_output[637] + last_layer_output[638] + last_layer_output[639] + last_layer_output[640] + last_layer_output[641] + last_layer_output[642] + last_layer_output[643] + last_layer_output[644] + last_layer_output[645] + last_layer_output[646] + last_layer_output[647] + last_layer_output[648] + last_layer_output[649] + last_layer_output[650] + last_layer_output[651] + last_layer_output[652] + last_layer_output[653] + last_layer_output[654] + last_layer_output[655] + last_layer_output[656] + last_layer_output[657] + last_layer_output[658] + last_layer_output[659] + last_layer_output[660] + last_layer_output[661] + last_layer_output[662] + last_layer_output[663] + last_layer_output[664] + last_layer_output[665] + last_layer_output[666] + last_layer_output[667] + last_layer_output[668] + last_layer_output[669] + last_layer_output[670] + last_layer_output[671] + last_layer_output[672] + last_layer_output[673] + last_layer_output[674] + last_layer_output[675] + last_layer_output[676] + last_layer_output[677] + last_layer_output[678] + last_layer_output[679] + last_layer_output[680] + last_layer_output[681] + last_layer_output[682] + last_layer_output[683] + last_layer_output[684] + last_layer_output[685] + last_layer_output[686] + last_layer_output[687] + last_layer_output[688] + last_layer_output[689] + last_layer_output[690] + last_layer_output[691] + last_layer_output[692] + last_layer_output[693] + last_layer_output[694] + last_layer_output[695] + last_layer_output[696] + last_layer_output[697] + last_layer_output[698] + last_layer_output[699] + last_layer_output[700] + last_layer_output[701] + last_layer_output[702] + last_layer_output[703] + last_layer_output[704] + last_layer_output[705] + last_layer_output[706] + last_layer_output[707] + last_layer_output[708] + last_layer_output[709] + last_layer_output[710] + last_layer_output[711] + last_layer_output[712] + last_layer_output[713] + last_layer_output[714] + last_layer_output[715] + last_layer_output[716] + last_layer_output[717] + last_layer_output[718] + last_layer_output[719] + last_layer_output[720] + last_layer_output[721] + last_layer_output[722] + last_layer_output[723] + last_layer_output[724] + last_layer_output[725] + last_layer_output[726] + last_layer_output[727] + last_layer_output[728] + last_layer_output[729] + last_layer_output[730] + last_layer_output[731] + last_layer_output[732] + last_layer_output[733] + last_layer_output[734] + last_layer_output[735] + last_layer_output[736] + last_layer_output[737] + last_layer_output[738] + last_layer_output[739] + last_layer_output[740] + last_layer_output[741] + last_layer_output[742] + last_layer_output[743] + last_layer_output[744] + last_layer_output[745] + last_layer_output[746] + last_layer_output[747] + last_layer_output[748] + last_layer_output[749];
      result[5] <= last_layer_output[750] + last_layer_output[751] + last_layer_output[752] + last_layer_output[753] + last_layer_output[754] + last_layer_output[755] + last_layer_output[756] + last_layer_output[757] + last_layer_output[758] + last_layer_output[759] + last_layer_output[760] + last_layer_output[761] + last_layer_output[762] + last_layer_output[763] + last_layer_output[764] + last_layer_output[765] + last_layer_output[766] + last_layer_output[767] + last_layer_output[768] + last_layer_output[769] + last_layer_output[770] + last_layer_output[771] + last_layer_output[772] + last_layer_output[773] + last_layer_output[774] + last_layer_output[775] + last_layer_output[776] + last_layer_output[777] + last_layer_output[778] + last_layer_output[779] + last_layer_output[780] + last_layer_output[781] + last_layer_output[782] + last_layer_output[783] + last_layer_output[784] + last_layer_output[785] + last_layer_output[786] + last_layer_output[787] + last_layer_output[788] + last_layer_output[789] + last_layer_output[790] + last_layer_output[791] + last_layer_output[792] + last_layer_output[793] + last_layer_output[794] + last_layer_output[795] + last_layer_output[796] + last_layer_output[797] + last_layer_output[798] + last_layer_output[799] + last_layer_output[800] + last_layer_output[801] + last_layer_output[802] + last_layer_output[803] + last_layer_output[804] + last_layer_output[805] + last_layer_output[806] + last_layer_output[807] + last_layer_output[808] + last_layer_output[809] + last_layer_output[810] + last_layer_output[811] + last_layer_output[812] + last_layer_output[813] + last_layer_output[814] + last_layer_output[815] + last_layer_output[816] + last_layer_output[817] + last_layer_output[818] + last_layer_output[819] + last_layer_output[820] + last_layer_output[821] + last_layer_output[822] + last_layer_output[823] + last_layer_output[824] + last_layer_output[825] + last_layer_output[826] + last_layer_output[827] + last_layer_output[828] + last_layer_output[829] + last_layer_output[830] + last_layer_output[831] + last_layer_output[832] + last_layer_output[833] + last_layer_output[834] + last_layer_output[835] + last_layer_output[836] + last_layer_output[837] + last_layer_output[838] + last_layer_output[839] + last_layer_output[840] + last_layer_output[841] + last_layer_output[842] + last_layer_output[843] + last_layer_output[844] + last_layer_output[845] + last_layer_output[846] + last_layer_output[847] + last_layer_output[848] + last_layer_output[849] + last_layer_output[850] + last_layer_output[851] + last_layer_output[852] + last_layer_output[853] + last_layer_output[854] + last_layer_output[855] + last_layer_output[856] + last_layer_output[857] + last_layer_output[858] + last_layer_output[859] + last_layer_output[860] + last_layer_output[861] + last_layer_output[862] + last_layer_output[863] + last_layer_output[864] + last_layer_output[865] + last_layer_output[866] + last_layer_output[867] + last_layer_output[868] + last_layer_output[869] + last_layer_output[870] + last_layer_output[871] + last_layer_output[872] + last_layer_output[873] + last_layer_output[874] + last_layer_output[875] + last_layer_output[876] + last_layer_output[877] + last_layer_output[878] + last_layer_output[879] + last_layer_output[880] + last_layer_output[881] + last_layer_output[882] + last_layer_output[883] + last_layer_output[884] + last_layer_output[885] + last_layer_output[886] + last_layer_output[887] + last_layer_output[888] + last_layer_output[889] + last_layer_output[890] + last_layer_output[891] + last_layer_output[892] + last_layer_output[893] + last_layer_output[894] + last_layer_output[895] + last_layer_output[896] + last_layer_output[897] + last_layer_output[898] + last_layer_output[899];
      result[6] <= last_layer_output[900] + last_layer_output[901] + last_layer_output[902] + last_layer_output[903] + last_layer_output[904] + last_layer_output[905] + last_layer_output[906] + last_layer_output[907] + last_layer_output[908] + last_layer_output[909] + last_layer_output[910] + last_layer_output[911] + last_layer_output[912] + last_layer_output[913] + last_layer_output[914] + last_layer_output[915] + last_layer_output[916] + last_layer_output[917] + last_layer_output[918] + last_layer_output[919] + last_layer_output[920] + last_layer_output[921] + last_layer_output[922] + last_layer_output[923] + last_layer_output[924] + last_layer_output[925] + last_layer_output[926] + last_layer_output[927] + last_layer_output[928] + last_layer_output[929] + last_layer_output[930] + last_layer_output[931] + last_layer_output[932] + last_layer_output[933] + last_layer_output[934] + last_layer_output[935] + last_layer_output[936] + last_layer_output[937] + last_layer_output[938] + last_layer_output[939] + last_layer_output[940] + last_layer_output[941] + last_layer_output[942] + last_layer_output[943] + last_layer_output[944] + last_layer_output[945] + last_layer_output[946] + last_layer_output[947] + last_layer_output[948] + last_layer_output[949] + last_layer_output[950] + last_layer_output[951] + last_layer_output[952] + last_layer_output[953] + last_layer_output[954] + last_layer_output[955] + last_layer_output[956] + last_layer_output[957] + last_layer_output[958] + last_layer_output[959] + last_layer_output[960] + last_layer_output[961] + last_layer_output[962] + last_layer_output[963] + last_layer_output[964] + last_layer_output[965] + last_layer_output[966] + last_layer_output[967] + last_layer_output[968] + last_layer_output[969] + last_layer_output[970] + last_layer_output[971] + last_layer_output[972] + last_layer_output[973] + last_layer_output[974] + last_layer_output[975] + last_layer_output[976] + last_layer_output[977] + last_layer_output[978] + last_layer_output[979] + last_layer_output[980] + last_layer_output[981] + last_layer_output[982] + last_layer_output[983] + last_layer_output[984] + last_layer_output[985] + last_layer_output[986] + last_layer_output[987] + last_layer_output[988] + last_layer_output[989] + last_layer_output[990] + last_layer_output[991] + last_layer_output[992] + last_layer_output[993] + last_layer_output[994] + last_layer_output[995] + last_layer_output[996] + last_layer_output[997] + last_layer_output[998] + last_layer_output[999] + last_layer_output[1000] + last_layer_output[1001] + last_layer_output[1002] + last_layer_output[1003] + last_layer_output[1004] + last_layer_output[1005] + last_layer_output[1006] + last_layer_output[1007] + last_layer_output[1008] + last_layer_output[1009] + last_layer_output[1010] + last_layer_output[1011] + last_layer_output[1012] + last_layer_output[1013] + last_layer_output[1014] + last_layer_output[1015] + last_layer_output[1016] + last_layer_output[1017] + last_layer_output[1018] + last_layer_output[1019] + last_layer_output[1020] + last_layer_output[1021] + last_layer_output[1022] + last_layer_output[1023] + last_layer_output[1024] + last_layer_output[1025] + last_layer_output[1026] + last_layer_output[1027] + last_layer_output[1028] + last_layer_output[1029] + last_layer_output[1030] + last_layer_output[1031] + last_layer_output[1032] + last_layer_output[1033] + last_layer_output[1034] + last_layer_output[1035] + last_layer_output[1036] + last_layer_output[1037] + last_layer_output[1038] + last_layer_output[1039] + last_layer_output[1040] + last_layer_output[1041] + last_layer_output[1042] + last_layer_output[1043] + last_layer_output[1044] + last_layer_output[1045] + last_layer_output[1046] + last_layer_output[1047] + last_layer_output[1048] + last_layer_output[1049];
      result[7] <= last_layer_output[1050] + last_layer_output[1051] + last_layer_output[1052] + last_layer_output[1053] + last_layer_output[1054] + last_layer_output[1055] + last_layer_output[1056] + last_layer_output[1057] + last_layer_output[1058] + last_layer_output[1059] + last_layer_output[1060] + last_layer_output[1061] + last_layer_output[1062] + last_layer_output[1063] + last_layer_output[1064] + last_layer_output[1065] + last_layer_output[1066] + last_layer_output[1067] + last_layer_output[1068] + last_layer_output[1069] + last_layer_output[1070] + last_layer_output[1071] + last_layer_output[1072] + last_layer_output[1073] + last_layer_output[1074] + last_layer_output[1075] + last_layer_output[1076] + last_layer_output[1077] + last_layer_output[1078] + last_layer_output[1079] + last_layer_output[1080] + last_layer_output[1081] + last_layer_output[1082] + last_layer_output[1083] + last_layer_output[1084] + last_layer_output[1085] + last_layer_output[1086] + last_layer_output[1087] + last_layer_output[1088] + last_layer_output[1089] + last_layer_output[1090] + last_layer_output[1091] + last_layer_output[1092] + last_layer_output[1093] + last_layer_output[1094] + last_layer_output[1095] + last_layer_output[1096] + last_layer_output[1097] + last_layer_output[1098] + last_layer_output[1099] + last_layer_output[1100] + last_layer_output[1101] + last_layer_output[1102] + last_layer_output[1103] + last_layer_output[1104] + last_layer_output[1105] + last_layer_output[1106] + last_layer_output[1107] + last_layer_output[1108] + last_layer_output[1109] + last_layer_output[1110] + last_layer_output[1111] + last_layer_output[1112] + last_layer_output[1113] + last_layer_output[1114] + last_layer_output[1115] + last_layer_output[1116] + last_layer_output[1117] + last_layer_output[1118] + last_layer_output[1119] + last_layer_output[1120] + last_layer_output[1121] + last_layer_output[1122] + last_layer_output[1123] + last_layer_output[1124] + last_layer_output[1125] + last_layer_output[1126] + last_layer_output[1127] + last_layer_output[1128] + last_layer_output[1129] + last_layer_output[1130] + last_layer_output[1131] + last_layer_output[1132] + last_layer_output[1133] + last_layer_output[1134] + last_layer_output[1135] + last_layer_output[1136] + last_layer_output[1137] + last_layer_output[1138] + last_layer_output[1139] + last_layer_output[1140] + last_layer_output[1141] + last_layer_output[1142] + last_layer_output[1143] + last_layer_output[1144] + last_layer_output[1145] + last_layer_output[1146] + last_layer_output[1147] + last_layer_output[1148] + last_layer_output[1149] + last_layer_output[1150] + last_layer_output[1151] + last_layer_output[1152] + last_layer_output[1153] + last_layer_output[1154] + last_layer_output[1155] + last_layer_output[1156] + last_layer_output[1157] + last_layer_output[1158] + last_layer_output[1159] + last_layer_output[1160] + last_layer_output[1161] + last_layer_output[1162] + last_layer_output[1163] + last_layer_output[1164] + last_layer_output[1165] + last_layer_output[1166] + last_layer_output[1167] + last_layer_output[1168] + last_layer_output[1169] + last_layer_output[1170] + last_layer_output[1171] + last_layer_output[1172] + last_layer_output[1173] + last_layer_output[1174] + last_layer_output[1175] + last_layer_output[1176] + last_layer_output[1177] + last_layer_output[1178] + last_layer_output[1179] + last_layer_output[1180] + last_layer_output[1181] + last_layer_output[1182] + last_layer_output[1183] + last_layer_output[1184] + last_layer_output[1185] + last_layer_output[1186] + last_layer_output[1187] + last_layer_output[1188] + last_layer_output[1189] + last_layer_output[1190] + last_layer_output[1191] + last_layer_output[1192] + last_layer_output[1193] + last_layer_output[1194] + last_layer_output[1195] + last_layer_output[1196] + last_layer_output[1197] + last_layer_output[1198] + last_layer_output[1199];
      result[8] <= last_layer_output[1200] + last_layer_output[1201] + last_layer_output[1202] + last_layer_output[1203] + last_layer_output[1204] + last_layer_output[1205] + last_layer_output[1206] + last_layer_output[1207] + last_layer_output[1208] + last_layer_output[1209] + last_layer_output[1210] + last_layer_output[1211] + last_layer_output[1212] + last_layer_output[1213] + last_layer_output[1214] + last_layer_output[1215] + last_layer_output[1216] + last_layer_output[1217] + last_layer_output[1218] + last_layer_output[1219] + last_layer_output[1220] + last_layer_output[1221] + last_layer_output[1222] + last_layer_output[1223] + last_layer_output[1224] + last_layer_output[1225] + last_layer_output[1226] + last_layer_output[1227] + last_layer_output[1228] + last_layer_output[1229] + last_layer_output[1230] + last_layer_output[1231] + last_layer_output[1232] + last_layer_output[1233] + last_layer_output[1234] + last_layer_output[1235] + last_layer_output[1236] + last_layer_output[1237] + last_layer_output[1238] + last_layer_output[1239] + last_layer_output[1240] + last_layer_output[1241] + last_layer_output[1242] + last_layer_output[1243] + last_layer_output[1244] + last_layer_output[1245] + last_layer_output[1246] + last_layer_output[1247] + last_layer_output[1248] + last_layer_output[1249] + last_layer_output[1250] + last_layer_output[1251] + last_layer_output[1252] + last_layer_output[1253] + last_layer_output[1254] + last_layer_output[1255] + last_layer_output[1256] + last_layer_output[1257] + last_layer_output[1258] + last_layer_output[1259] + last_layer_output[1260] + last_layer_output[1261] + last_layer_output[1262] + last_layer_output[1263] + last_layer_output[1264] + last_layer_output[1265] + last_layer_output[1266] + last_layer_output[1267] + last_layer_output[1268] + last_layer_output[1269] + last_layer_output[1270] + last_layer_output[1271] + last_layer_output[1272] + last_layer_output[1273] + last_layer_output[1274] + last_layer_output[1275] + last_layer_output[1276] + last_layer_output[1277] + last_layer_output[1278] + last_layer_output[1279] + last_layer_output[1280] + last_layer_output[1281] + last_layer_output[1282] + last_layer_output[1283] + last_layer_output[1284] + last_layer_output[1285] + last_layer_output[1286] + last_layer_output[1287] + last_layer_output[1288] + last_layer_output[1289] + last_layer_output[1290] + last_layer_output[1291] + last_layer_output[1292] + last_layer_output[1293] + last_layer_output[1294] + last_layer_output[1295] + last_layer_output[1296] + last_layer_output[1297] + last_layer_output[1298] + last_layer_output[1299] + last_layer_output[1300] + last_layer_output[1301] + last_layer_output[1302] + last_layer_output[1303] + last_layer_output[1304] + last_layer_output[1305] + last_layer_output[1306] + last_layer_output[1307] + last_layer_output[1308] + last_layer_output[1309] + last_layer_output[1310] + last_layer_output[1311] + last_layer_output[1312] + last_layer_output[1313] + last_layer_output[1314] + last_layer_output[1315] + last_layer_output[1316] + last_layer_output[1317] + last_layer_output[1318] + last_layer_output[1319] + last_layer_output[1320] + last_layer_output[1321] + last_layer_output[1322] + last_layer_output[1323] + last_layer_output[1324] + last_layer_output[1325] + last_layer_output[1326] + last_layer_output[1327] + last_layer_output[1328] + last_layer_output[1329] + last_layer_output[1330] + last_layer_output[1331] + last_layer_output[1332] + last_layer_output[1333] + last_layer_output[1334] + last_layer_output[1335] + last_layer_output[1336] + last_layer_output[1337] + last_layer_output[1338] + last_layer_output[1339] + last_layer_output[1340] + last_layer_output[1341] + last_layer_output[1342] + last_layer_output[1343] + last_layer_output[1344] + last_layer_output[1345] + last_layer_output[1346] + last_layer_output[1347] + last_layer_output[1348] + last_layer_output[1349];
      result[9] <= last_layer_output[1350] + last_layer_output[1351] + last_layer_output[1352] + last_layer_output[1353] + last_layer_output[1354] + last_layer_output[1355] + last_layer_output[1356] + last_layer_output[1357] + last_layer_output[1358] + last_layer_output[1359] + last_layer_output[1360] + last_layer_output[1361] + last_layer_output[1362] + last_layer_output[1363] + last_layer_output[1364] + last_layer_output[1365] + last_layer_output[1366] + last_layer_output[1367] + last_layer_output[1368] + last_layer_output[1369] + last_layer_output[1370] + last_layer_output[1371] + last_layer_output[1372] + last_layer_output[1373] + last_layer_output[1374] + last_layer_output[1375] + last_layer_output[1376] + last_layer_output[1377] + last_layer_output[1378] + last_layer_output[1379] + last_layer_output[1380] + last_layer_output[1381] + last_layer_output[1382] + last_layer_output[1383] + last_layer_output[1384] + last_layer_output[1385] + last_layer_output[1386] + last_layer_output[1387] + last_layer_output[1388] + last_layer_output[1389] + last_layer_output[1390] + last_layer_output[1391] + last_layer_output[1392] + last_layer_output[1393] + last_layer_output[1394] + last_layer_output[1395] + last_layer_output[1396] + last_layer_output[1397] + last_layer_output[1398] + last_layer_output[1399] + last_layer_output[1400] + last_layer_output[1401] + last_layer_output[1402] + last_layer_output[1403] + last_layer_output[1404] + last_layer_output[1405] + last_layer_output[1406] + last_layer_output[1407] + last_layer_output[1408] + last_layer_output[1409] + last_layer_output[1410] + last_layer_output[1411] + last_layer_output[1412] + last_layer_output[1413] + last_layer_output[1414] + last_layer_output[1415] + last_layer_output[1416] + last_layer_output[1417] + last_layer_output[1418] + last_layer_output[1419] + last_layer_output[1420] + last_layer_output[1421] + last_layer_output[1422] + last_layer_output[1423] + last_layer_output[1424] + last_layer_output[1425] + last_layer_output[1426] + last_layer_output[1427] + last_layer_output[1428] + last_layer_output[1429] + last_layer_output[1430] + last_layer_output[1431] + last_layer_output[1432] + last_layer_output[1433] + last_layer_output[1434] + last_layer_output[1435] + last_layer_output[1436] + last_layer_output[1437] + last_layer_output[1438] + last_layer_output[1439] + last_layer_output[1440] + last_layer_output[1441] + last_layer_output[1442] + last_layer_output[1443] + last_layer_output[1444] + last_layer_output[1445] + last_layer_output[1446] + last_layer_output[1447] + last_layer_output[1448] + last_layer_output[1449] + last_layer_output[1450] + last_layer_output[1451] + last_layer_output[1452] + last_layer_output[1453] + last_layer_output[1454] + last_layer_output[1455] + last_layer_output[1456] + last_layer_output[1457] + last_layer_output[1458] + last_layer_output[1459] + last_layer_output[1460] + last_layer_output[1461] + last_layer_output[1462] + last_layer_output[1463] + last_layer_output[1464] + last_layer_output[1465] + last_layer_output[1466] + last_layer_output[1467] + last_layer_output[1468] + last_layer_output[1469] + last_layer_output[1470] + last_layer_output[1471] + last_layer_output[1472] + last_layer_output[1473] + last_layer_output[1474] + last_layer_output[1475] + last_layer_output[1476] + last_layer_output[1477] + last_layer_output[1478] + last_layer_output[1479] + last_layer_output[1480] + last_layer_output[1481] + last_layer_output[1482] + last_layer_output[1483] + last_layer_output[1484] + last_layer_output[1485] + last_layer_output[1486] + last_layer_output[1487] + last_layer_output[1488] + last_layer_output[1489] + last_layer_output[1490] + last_layer_output[1491] + last_layer_output[1492] + last_layer_output[1493] + last_layer_output[1494] + last_layer_output[1495] + last_layer_output[1496] + last_layer_output[1497] + last_layer_output[1498] + last_layer_output[1499];
end
      assign y[79:72]=result[0];
      assign y[71:64]=result[1];
      assign y[63:56]=result[2];
      assign y[55:48]=result[3];
      assign y[47:40]=result[4];
      assign y[39:32]=result[5];
      assign y[31:24]=result[6];
      assign y[23:16]=result[7];
      assign y[15:8]=result[8];
      assign y[7:0]=result[9];
endmodule