module logic_network (    input clk,
    input wire [399:0] x,
    output wire [69:0] y
);
      reg [799:0] layer0_out = 0;
      reg [799:0] layer1_out = 0;
      reg [799:0] layer2_out = 0;
      reg [799:0] layer3_out = 0;
      reg [799:0] layer4_out = 0;
      reg [799:0] layer5_out = 0;
      reg [799:0] last_layer_output = 0;
      reg [6:0] result [9:0];
      always @(posedge clk) begin
     layer0_out[0] <= ~(x[29] | x[31]);
     layer0_out[1] <= ~(x[157] & x[159]);
     layer0_out[2] <= x[59] | x[61];
     layer0_out[3] <= 1'b1;
     layer0_out[4] <= 1'b1;
     layer0_out[5] <= ~x[163];
     layer0_out[6] <= ~x[27] | x[29];
     layer0_out[7] <= x[106] & x[107];
     layer0_out[8] <= x[324] | x[325];
     layer0_out[9] <= ~(x[215] & x[216]);
     layer0_out[10] <= ~x[225];
     layer0_out[11] <= ~(x[90] | x[91]);
     layer0_out[12] <= x[74];
     layer0_out[13] <= 1'b1;
     layer0_out[14] <= x[369] | x[371];
     layer0_out[15] <= ~(x[16] | x[17]);
     layer0_out[16] <= 1'b0;
     layer0_out[17] <= 1'b0;
     layer0_out[18] <= 1'b1;
     layer0_out[19] <= x[382] | x[383];
     layer0_out[20] <= x[255] | x[257];
     layer0_out[21] <= ~(x[42] | x[44]);
     layer0_out[22] <= 1'b0;
     layer0_out[23] <= x[179] | x[180];
     layer0_out[24] <= 1'b0;
     layer0_out[25] <= x[302] | x[303];
     layer0_out[26] <= x[69] | x[70];
     layer0_out[27] <= ~x[367];
     layer0_out[28] <= ~x[332];
     layer0_out[29] <= x[362] | x[364];
     layer0_out[30] <= x[267];
     layer0_out[31] <= ~(x[330] | x[331]);
     layer0_out[32] <= x[9] | x[10];
     layer0_out[33] <= ~(x[48] | x[49]);
     layer0_out[34] <= x[308] | x[309];
     layer0_out[35] <= x[210] | x[211];
     layer0_out[36] <= ~x[94];
     layer0_out[37] <= ~(x[284] | x[286]);
     layer0_out[38] <= x[308];
     layer0_out[39] <= ~(x[212] | x[214]);
     layer0_out[40] <= ~(x[173] | x[175]);
     layer0_out[41] <= ~(x[96] | x[98]);
     layer0_out[42] <= ~x[132];
     layer0_out[43] <= 1'b0;
     layer0_out[44] <= x[372] | x[374];
     layer0_out[45] <= x[110] | x[112];
     layer0_out[46] <= x[250] | x[252];
     layer0_out[47] <= x[196];
     layer0_out[48] <= x[142];
     layer0_out[49] <= 1'b0;
     layer0_out[50] <= ~(x[161] | x[162]);
     layer0_out[51] <= x[207] | x[208];
     layer0_out[52] <= ~(x[209] | x[211]);
     layer0_out[53] <= x[149] | x[151];
     layer0_out[54] <= ~(x[67] | x[68]);
     layer0_out[55] <= ~(x[83] | x[84]);
     layer0_out[56] <= ~x[108] | x[106];
     layer0_out[57] <= x[139];
     layer0_out[58] <= x[73] | x[74];
     layer0_out[59] <= x[95] & ~x[93];
     layer0_out[60] <= 1'b1;
     layer0_out[61] <= x[307] | x[309];
     layer0_out[62] <= x[370] & x[372];
     layer0_out[63] <= ~(x[38] | x[39]);
     layer0_out[64] <= ~x[281];
     layer0_out[65] <= ~x[208] | x[206];
     layer0_out[66] <= x[340] | x[342];
     layer0_out[67] <= x[109];
     layer0_out[68] <= 1'b1;
     layer0_out[69] <= x[197];
     layer0_out[70] <= x[225] | x[227];
     layer0_out[71] <= ~x[342];
     layer0_out[72] <= ~(x[20] & x[21]);
     layer0_out[73] <= x[236] | x[238];
     layer0_out[74] <= ~(x[185] | x[187]);
     layer0_out[75] <= ~(x[282] | x[283]);
     layer0_out[76] <= x[262] | x[263];
     layer0_out[77] <= ~x[77] | x[76];
     layer0_out[78] <= x[139] | x[140];
     layer0_out[79] <= ~(x[239] | x[240]);
     layer0_out[80] <= x[44] | x[46];
     layer0_out[81] <= 1'b1;
     layer0_out[82] <= 1'b0;
     layer0_out[83] <= ~(x[255] | x[256]);
     layer0_out[84] <= ~x[343];
     layer0_out[85] <= ~(x[163] | x[165]);
     layer0_out[86] <= x[14] | x[15];
     layer0_out[87] <= ~x[190];
     layer0_out[88] <= x[211];
     layer0_out[89] <= 1'b1;
     layer0_out[90] <= x[328] | x[330];
     layer0_out[91] <= ~x[268];
     layer0_out[92] <= x[386];
     layer0_out[93] <= ~x[50];
     layer0_out[94] <= ~(x[88] | x[89]);
     layer0_out[95] <= x[158] | x[159];
     layer0_out[96] <= x[200] | x[202];
     layer0_out[97] <= x[166] | x[167];
     layer0_out[98] <= 1'b1;
     layer0_out[99] <= x[358] | x[359];
     layer0_out[100] <= ~(x[351] | x[352]);
     layer0_out[101] <= ~(x[355] | x[357]);
     layer0_out[102] <= x[78] | x[79];
     layer0_out[103] <= x[243] | x[244];
     layer0_out[104] <= 1'b0;
     layer0_out[105] <= x[325];
     layer0_out[106] <= ~(x[278] | x[280]);
     layer0_out[107] <= ~(x[6] & x[8]);
     layer0_out[108] <= ~(x[2] | x[4]);
     layer0_out[109] <= 1'b1;
     layer0_out[110] <= ~x[220];
     layer0_out[111] <= x[168] & ~x[166];
     layer0_out[112] <= ~(x[58] | x[59]);
     layer0_out[113] <= x[41] | x[42];
     layer0_out[114] <= x[130] & ~x[128];
     layer0_out[115] <= x[40] | x[41];
     layer0_out[116] <= x[59];
     layer0_out[117] <= ~(x[129] | x[130]);
     layer0_out[118] <= x[296] | x[298];
     layer0_out[119] <= x[394] | x[396];
     layer0_out[120] <= 1'b1;
     layer0_out[121] <= 1'b0;
     layer0_out[122] <= 1'b1;
     layer0_out[123] <= ~(x[182] | x[183]);
     layer0_out[124] <= ~(x[195] | x[197]);
     layer0_out[125] <= x[295] & ~x[293];
     layer0_out[126] <= x[213];
     layer0_out[127] <= ~(x[270] ^ x[271]);
     layer0_out[128] <= ~(x[334] | x[335]);
     layer0_out[129] <= x[338] & x[340];
     layer0_out[130] <= x[246] | x[248];
     layer0_out[131] <= x[159];
     layer0_out[132] <= ~(x[125] | x[127]);
     layer0_out[133] <= ~x[18] | x[19];
     layer0_out[134] <= ~(x[14] | x[16]);
     layer0_out[135] <= ~(x[378] | x[379]);
     layer0_out[136] <= 1'b1;
     layer0_out[137] <= x[396] & x[397];
     layer0_out[138] <= x[84] | x[85];
     layer0_out[139] <= 1'b0;
     layer0_out[140] <= x[35];
     layer0_out[141] <= ~(x[336] | x[337]);
     layer0_out[142] <= ~x[375];
     layer0_out[143] <= ~x[209];
     layer0_out[144] <= 1'b0;
     layer0_out[145] <= ~(x[68] | x[70]);
     layer0_out[146] <= ~x[387];
     layer0_out[147] <= ~(x[344] | x[345]);
     layer0_out[148] <= x[45];
     layer0_out[149] <= ~x[57] | x[56];
     layer0_out[150] <= x[225] & x[226];
     layer0_out[151] <= ~(x[199] | x[200]);
     layer0_out[152] <= ~x[395] | x[393];
     layer0_out[153] <= x[112] & x[114];
     layer0_out[154] <= 1'b0;
     layer0_out[155] <= ~(x[354] | x[355]);
     layer0_out[156] <= ~x[265] | x[267];
     layer0_out[157] <= ~(x[311] | x[312]);
     layer0_out[158] <= ~x[159];
     layer0_out[159] <= 1'b0;
     layer0_out[160] <= ~x[10];
     layer0_out[161] <= ~(x[165] & x[167]);
     layer0_out[162] <= ~x[350];
     layer0_out[163] <= x[275] | x[277];
     layer0_out[164] <= ~(x[109] & x[111]);
     layer0_out[165] <= ~(x[391] | x[392]);
     layer0_out[166] <= ~x[73];
     layer0_out[167] <= 1'b0;
     layer0_out[168] <= ~(x[30] ^ x[32]);
     layer0_out[169] <= x[63] | x[65];
     layer0_out[170] <= x[7] | x[8];
     layer0_out[171] <= x[152] | x[153];
     layer0_out[172] <= x[160] | x[162];
     layer0_out[173] <= x[253];
     layer0_out[174] <= ~x[345];
     layer0_out[175] <= 1'b1;
     layer0_out[176] <= x[250];
     layer0_out[177] <= 1'b0;
     layer0_out[178] <= x[69] | x[71];
     layer0_out[179] <= 1'b1;
     layer0_out[180] <= x[155] | x[157];
     layer0_out[181] <= ~(x[104] ^ x[105]);
     layer0_out[182] <= ~x[308];
     layer0_out[183] <= x[82] | x[83];
     layer0_out[184] <= ~(x[247] | x[248]);
     layer0_out[185] <= 1'b1;
     layer0_out[186] <= x[295] | x[296];
     layer0_out[187] <= ~x[264];
     layer0_out[188] <= x[204] | x[205];
     layer0_out[189] <= x[201];
     layer0_out[190] <= ~(x[156] | x[158]);
     layer0_out[191] <= 1'b1;
     layer0_out[192] <= x[97] | x[99];
     layer0_out[193] <= ~(x[316] | x[318]);
     layer0_out[194] <= 1'b0;
     layer0_out[195] <= x[158] | x[160];
     layer0_out[196] <= ~(x[374] | x[376]);
     layer0_out[197] <= x[46];
     layer0_out[198] <= x[386] | x[388];
     layer0_out[199] <= x[254] | x[256];
     layer0_out[200] <= x[330] | x[332];
     layer0_out[201] <= 1'b0;
     layer0_out[202] <= 1'b0;
     layer0_out[203] <= 1'b0;
     layer0_out[204] <= 1'b1;
     layer0_out[205] <= 1'b0;
     layer0_out[206] <= x[173] & ~x[171];
     layer0_out[207] <= x[341] | x[343];
     layer0_out[208] <= ~(x[365] | x[367]);
     layer0_out[209] <= x[123] & ~x[121];
     layer0_out[210] <= x[64];
     layer0_out[211] <= ~(x[391] | x[393]);
     layer0_out[212] <= x[15] | x[16];
     layer0_out[213] <= x[277] | x[278];
     layer0_out[214] <= x[319] | x[321];
     layer0_out[215] <= 1'b1;
     layer0_out[216] <= ~x[280] | x[279];
     layer0_out[217] <= ~(x[136] & x[137]);
     layer0_out[218] <= ~x[145] | x[147];
     layer0_out[219] <= x[115] | x[117];
     layer0_out[220] <= x[234];
     layer0_out[221] <= ~(x[2] | x[5]);
     layer0_out[222] <= x[339];
     layer0_out[223] <= 1'b1;
     layer0_out[224] <= ~x[28];
     layer0_out[225] <= ~x[150];
     layer0_out[226] <= ~x[397] | x[398];
     layer0_out[227] <= ~(x[68] | x[69]);
     layer0_out[228] <= x[120];
     layer0_out[229] <= x[77] | x[78];
     layer0_out[230] <= x[320] & ~x[321];
     layer0_out[231] <= x[355];
     layer0_out[232] <= x[313] & ~x[315];
     layer0_out[233] <= 1'b0;
     layer0_out[234] <= x[357] | x[358];
     layer0_out[235] <= ~(x[39] | x[41]);
     layer0_out[236] <= ~x[276];
     layer0_out[237] <= x[135] | x[136];
     layer0_out[238] <= ~x[129] | x[127];
     layer0_out[239] <= ~(x[181] | x[183]);
     layer0_out[240] <= ~(x[30] | x[31]);
     layer0_out[241] <= ~(x[382] | x[384]);
     layer0_out[242] <= x[51];
     layer0_out[243] <= ~(x[18] | x[20]);
     layer0_out[244] <= ~x[137] | x[139];
     layer0_out[245] <= x[186] | x[188];
     layer0_out[246] <= 1'b0;
     layer0_out[247] <= 1'b1;
     layer0_out[248] <= x[377];
     layer0_out[249] <= ~(x[174] | x[175]);
     layer0_out[250] <= ~(x[257] | x[259]);
     layer0_out[251] <= x[140] | x[141];
     layer0_out[252] <= ~x[249] | x[251];
     layer0_out[253] <= ~(x[194] | x[196]);
     layer0_out[254] <= ~(x[55] & x[57]);
     layer0_out[255] <= x[328] & x[329];
     layer0_out[256] <= 1'b1;
     layer0_out[257] <= ~(x[0] | x[3]);
     layer0_out[258] <= ~(x[108] | x[110]);
     layer0_out[259] <= x[150] | x[152];
     layer0_out[260] <= 1'b1;
     layer0_out[261] <= ~(x[243] | x[245]);
     layer0_out[262] <= ~(x[244] & x[246]);
     layer0_out[263] <= x[50] | x[51];
     layer0_out[264] <= ~(x[368] | x[370]);
     layer0_out[265] <= x[93] | x[94];
     layer0_out[266] <= x[229] | x[231];
     layer0_out[267] <= x[68];
     layer0_out[268] <= 1'b0;
     layer0_out[269] <= ~(x[381] & x[382]);
     layer0_out[270] <= ~(x[3] | x[4]);
     layer0_out[271] <= 1'b0;
     layer0_out[272] <= 1'b1;
     layer0_out[273] <= x[273] | x[275];
     layer0_out[274] <= ~(x[302] | x[304]);
     layer0_out[275] <= 1'b0;
     layer0_out[276] <= ~(x[179] | x[181]);
     layer0_out[277] <= x[363];
     layer0_out[278] <= ~(x[205] | x[206]);
     layer0_out[279] <= x[10] | x[11];
     layer0_out[280] <= x[133] ^ x[134];
     layer0_out[281] <= ~(x[267] | x[268]);
     layer0_out[282] <= ~x[54];
     layer0_out[283] <= x[219];
     layer0_out[284] <= ~(x[56] | x[58]);
     layer0_out[285] <= x[24] | x[26];
     layer0_out[286] <= ~x[171];
     layer0_out[287] <= x[188] ^ x[189];
     layer0_out[288] <= x[29] | x[30];
     layer0_out[289] <= x[352] & ~x[353];
     layer0_out[290] <= x[172] | x[174];
     layer0_out[291] <= 1'b1;
     layer0_out[292] <= 1'b0;
     layer0_out[293] <= x[333];
     layer0_out[294] <= x[208] | x[209];
     layer0_out[295] <= x[28] | x[30];
     layer0_out[296] <= x[388] | x[390];
     layer0_out[297] <= x[164];
     layer0_out[298] <= ~(x[252] | x[254]);
     layer0_out[299] <= x[194] | x[195];
     layer0_out[300] <= ~(x[189] & x[191]);
     layer0_out[301] <= ~x[198];
     layer0_out[302] <= x[233];
     layer0_out[303] <= x[222] | x[223];
     layer0_out[304] <= ~(x[79] | x[81]);
     layer0_out[305] <= ~x[385] | x[384];
     layer0_out[306] <= ~(x[276] | x[278]);
     layer0_out[307] <= 1'b0;
     layer0_out[308] <= ~x[19];
     layer0_out[309] <= x[13];
     layer0_out[310] <= x[126] ^ x[127];
     layer0_out[311] <= 1'b0;
     layer0_out[312] <= ~x[313];
     layer0_out[313] <= x[246] ^ x[247];
     layer0_out[314] <= ~(x[182] & x[184]);
     layer0_out[315] <= ~x[275] | x[274];
     layer0_out[316] <= ~x[116];
     layer0_out[317] <= x[341] | x[342];
     layer0_out[318] <= ~x[283] | x[284];
     layer0_out[319] <= ~x[38];
     layer0_out[320] <= x[349] | x[351];
     layer0_out[321] <= ~x[189];
     layer0_out[322] <= 1'b0;
     layer0_out[323] <= ~x[265];
     layer0_out[324] <= ~(x[116] | x[118]);
     layer0_out[325] <= ~x[206];
     layer0_out[326] <= ~x[310];
     layer0_out[327] <= ~x[76];
     layer0_out[328] <= x[88] | x[90];
     layer0_out[329] <= x[45] | x[47];
     layer0_out[330] <= x[13];
     layer0_out[331] <= 1'b1;
     layer0_out[332] <= x[269] | x[271];
     layer0_out[333] <= x[285];
     layer0_out[334] <= ~x[82];
     layer0_out[335] <= x[164] | x[166];
     layer0_out[336] <= ~(x[115] | x[116]);
     layer0_out[337] <= x[121] & x[122];
     layer0_out[338] <= x[355] | x[356];
     layer0_out[339] <= ~(x[248] | x[250]);
     layer0_out[340] <= x[261] | x[263];
     layer0_out[341] <= ~x[135];
     layer0_out[342] <= ~x[287];
     layer0_out[343] <= x[213] ^ x[214];
     layer0_out[344] <= 1'b1;
     layer0_out[345] <= 1'b0;
     layer0_out[346] <= 1'b0;
     layer0_out[347] <= x[300] | x[301];
     layer0_out[348] <= x[1] | x[4];
     layer0_out[349] <= ~(x[362] | x[363]);
     layer0_out[350] <= ~(x[379] | x[380]);
     layer0_out[351] <= ~x[194];
     layer0_out[352] <= x[147] & x[148];
     layer0_out[353] <= 1'b1;
     layer0_out[354] <= ~(x[198] | x[200]);
     layer0_out[355] <= ~(x[89] | x[90]);
     layer0_out[356] <= ~(x[364] | x[365]);
     layer0_out[357] <= 1'b0;
     layer0_out[358] <= 1'b0;
     layer0_out[359] <= x[234] | x[236];
     layer0_out[360] <= x[245] & ~x[246];
     layer0_out[361] <= ~(x[137] | x[138]);
     layer0_out[362] <= x[157] | x[158];
     layer0_out[363] <= x[238] | x[239];
     layer0_out[364] <= x[12] | x[13];
     layer0_out[365] <= x[44] & ~x[43];
     layer0_out[366] <= 1'b1;
     layer0_out[367] <= x[231] | x[232];
     layer0_out[368] <= ~(x[262] | x[264]);
     layer0_out[369] <= x[368] & ~x[369];
     layer0_out[370] <= ~(x[95] | x[96]);
     layer0_out[371] <= 1'b1;
     layer0_out[372] <= 1'b0;
     layer0_out[373] <= ~x[148] | x[149];
     layer0_out[374] <= x[109] | x[110];
     layer0_out[375] <= x[23] & ~x[21];
     layer0_out[376] <= x[299] | x[300];
     layer0_out[377] <= ~(x[367] | x[368]);
     layer0_out[378] <= x[119] | x[120];
     layer0_out[379] <= x[50] & ~x[52];
     layer0_out[380] <= ~(x[32] | x[34]);
     layer0_out[381] <= x[226] & ~x[224];
     layer0_out[382] <= x[232] | x[233];
     layer0_out[383] <= ~(x[80] | x[81]);
     layer0_out[384] <= x[49] | x[51];
     layer0_out[385] <= ~(x[72] | x[74]);
     layer0_out[386] <= ~(x[398] | x[399]);
     layer0_out[387] <= 1'b1;
     layer0_out[388] <= 1'b1;
     layer0_out[389] <= 1'b0;
     layer0_out[390] <= 1'b0;
     layer0_out[391] <= 1'b1;
     layer0_out[392] <= x[336] | x[338];
     layer0_out[393] <= 1'b0;
     layer0_out[394] <= ~x[253] | x[255];
     layer0_out[395] <= ~(x[62] | x[64]);
     layer0_out[396] <= 1'b0;
     layer0_out[397] <= x[111] | x[113];
     layer0_out[398] <= x[288];
     layer0_out[399] <= ~(x[164] | x[165]);
     layer0_out[400] <= 1'b1;
     layer0_out[401] <= ~x[398];
     layer0_out[402] <= ~(x[301] | x[302]);
     layer0_out[403] <= x[81] | x[82];
     layer0_out[404] <= ~(x[378] | x[380]);
     layer0_out[405] <= 1'b0;
     layer0_out[406] <= ~(x[323] | x[324]);
     layer0_out[407] <= x[54];
     layer0_out[408] <= ~(x[5] | x[6]);
     layer0_out[409] <= x[26];
     layer0_out[410] <= ~(x[47] & x[48]);
     layer0_out[411] <= x[33] | x[35];
     layer0_out[412] <= 1'b0;
     layer0_out[413] <= ~(x[42] | x[43]);
     layer0_out[414] <= 1'b0;
     layer0_out[415] <= x[74] | x[75];
     layer0_out[416] <= ~(x[123] | x[124]);
     layer0_out[417] <= 1'b1;
     layer0_out[418] <= ~x[397] | x[395];
     layer0_out[419] <= ~(x[350] | x[351]);
     layer0_out[420] <= 1'b1;
     layer0_out[421] <= x[131] | x[132];
     layer0_out[422] <= ~x[119];
     layer0_out[423] <= ~(x[184] | x[185]);
     layer0_out[424] <= ~x[372];
     layer0_out[425] <= 1'b0;
     layer0_out[426] <= x[208] | x[210];
     layer0_out[427] <= ~(x[79] | x[80]);
     layer0_out[428] <= 1'b1;
     layer0_out[429] <= 1'b1;
     layer0_out[430] <= ~(x[248] | x[249]);
     layer0_out[431] <= ~(x[290] | x[292]);
     layer0_out[432] <= x[65];
     layer0_out[433] <= 1'b0;
     layer0_out[434] <= x[315] | x[317];
     layer0_out[435] <= x[171] | x[172];
     layer0_out[436] <= 1'b0;
     layer0_out[437] <= ~(x[184] & x[186]);
     layer0_out[438] <= x[371] | x[373];
     layer0_out[439] <= x[153] | x[155];
     layer0_out[440] <= ~(x[291] | x[292]);
     layer0_out[441] <= x[181] | x[182];
     layer0_out[442] <= x[188] | x[190];
     layer0_out[443] <= ~x[327];
     layer0_out[444] <= ~(x[326] | x[327]);
     layer0_out[445] <= ~(x[124] | x[126]);
     layer0_out[446] <= ~(x[332] | x[334]);
     layer0_out[447] <= x[252] | x[253];
     layer0_out[448] <= x[259] | x[261];
     layer0_out[449] <= x[228] | x[230];
     layer0_out[450] <= x[254] | x[255];
     layer0_out[451] <= ~(x[200] | x[201]);
     layer0_out[452] <= ~(x[263] | x[264]);
     layer0_out[453] <= x[203] | x[205];
     layer0_out[454] <= 1'b0;
     layer0_out[455] <= ~(x[122] | x[123]);
     layer0_out[456] <= 1'b0;
     layer0_out[457] <= ~(x[9] & x[11]);
     layer0_out[458] <= x[53] | x[55];
     layer0_out[459] <= 1'b1;
     layer0_out[460] <= 1'b0;
     layer0_out[461] <= x[113] | x[115];
     layer0_out[462] <= x[370] & ~x[369];
     layer0_out[463] <= 1'b0;
     layer0_out[464] <= x[221] | x[222];
     layer0_out[465] <= ~x[201];
     layer0_out[466] <= 1'b0;
     layer0_out[467] <= x[126] | x[128];
     layer0_out[468] <= 1'b0;
     layer0_out[469] <= x[226] | x[227];
     layer0_out[470] <= ~(x[250] ^ x[251]);
     layer0_out[471] <= ~(x[289] & x[291]);
     layer0_out[472] <= x[277] | x[279];
     layer0_out[473] <= ~(x[367] | x[369]);
     layer0_out[474] <= x[59] | x[60];
     layer0_out[475] <= ~x[302] | x[300];
     layer0_out[476] <= 1'b0;
     layer0_out[477] <= 1'b1;
     layer0_out[478] <= 1'b1;
     layer0_out[479] <= x[37];
     layer0_out[480] <= ~x[63];
     layer0_out[481] <= ~x[176] | x[175];
     layer0_out[482] <= 1'b1;
     layer0_out[483] <= ~x[27] | x[26];
     layer0_out[484] <= x[103];
     layer0_out[485] <= 1'b0;
     layer0_out[486] <= x[122] | x[124];
     layer0_out[487] <= x[104] & ~x[103];
     layer0_out[488] <= ~x[278] | x[279];
     layer0_out[489] <= x[35];
     layer0_out[490] <= x[244] & ~x[242];
     layer0_out[491] <= ~(x[395] | x[396]);
     layer0_out[492] <= ~(x[22] | x[23]);
     layer0_out[493] <= x[256] | x[257];
     layer0_out[494] <= x[345] | x[347];
     layer0_out[495] <= x[348] | x[349];
     layer0_out[496] <= x[293];
     layer0_out[497] <= 1'b1;
     layer0_out[498] <= 1'b1;
     layer0_out[499] <= ~(x[156] | x[157]);
     layer0_out[500] <= x[114] | x[116];
     layer0_out[501] <= ~(x[169] | x[170]);
     layer0_out[502] <= ~x[284];
     layer0_out[503] <= ~(x[1] | x[3]);
     layer0_out[504] <= ~(x[125] | x[126]);
     layer0_out[505] <= x[73];
     layer0_out[506] <= ~(x[87] | x[88]);
     layer0_out[507] <= ~(x[236] | x[237]);
     layer0_out[508] <= x[147] | x[149];
     layer0_out[509] <= x[258];
     layer0_out[510] <= x[385];
     layer0_out[511] <= x[91] | x[93];
     layer0_out[512] <= x[316];
     layer0_out[513] <= ~(x[284] | x[285]);
     layer0_out[514] <= 1'b0;
     layer0_out[515] <= ~(x[100] | x[101]);
     layer0_out[516] <= x[223] | x[224];
     layer0_out[517] <= ~(x[365] | x[366]);
     layer0_out[518] <= ~(x[383] | x[384]);
     layer0_out[519] <= ~x[124];
     layer0_out[520] <= ~x[207];
     layer0_out[521] <= ~(x[110] | x[111]);
     layer0_out[522] <= 1'b0;
     layer0_out[523] <= ~x[193];
     layer0_out[524] <= 1'b0;
     layer0_out[525] <= x[60] | x[61];
     layer0_out[526] <= ~(x[129] & x[131]);
     layer0_out[527] <= ~(x[97] & x[98]);
     layer0_out[528] <= 1'b0;
     layer0_out[529] <= ~x[113] | x[112];
     layer0_out[530] <= ~(x[190] | x[191]);
     layer0_out[531] <= x[281] & x[283];
     layer0_out[532] <= x[134] & x[136];
     layer0_out[533] <= x[37] | x[38];
     layer0_out[534] <= x[170] & x[172];
     layer0_out[535] <= x[292] & x[294];
     layer0_out[536] <= x[121] & ~x[120];
     layer0_out[537] <= ~x[117];
     layer0_out[538] <= x[12];
     layer0_out[539] <= ~(x[364] & x[366]);
     layer0_out[540] <= x[239] | x[241];
     layer0_out[541] <= 1'b0;
     layer0_out[542] <= ~x[301];
     layer0_out[543] <= ~(x[31] & x[32]);
     layer0_out[544] <= 1'b1;
     layer0_out[545] <= x[226];
     layer0_out[546] <= ~(x[134] | x[135]);
     layer0_out[547] <= ~(x[325] | x[327]);
     layer0_out[548] <= x[288] | x[289];
     layer0_out[549] <= x[390] | x[392];
     layer0_out[550] <= ~(x[96] | x[97]);
     layer0_out[551] <= ~(x[23] ^ x[25]);
     layer0_out[552] <= x[392] | x[393];
     layer0_out[553] <= ~(x[350] | x[352]);
     layer0_out[554] <= x[380] & x[382];
     layer0_out[555] <= 1'b0;
     layer0_out[556] <= x[78] | x[80];
     layer0_out[557] <= x[130];
     layer0_out[558] <= x[107] | x[109];
     layer0_out[559] <= 1'b1;
     layer0_out[560] <= x[138] | x[140];
     layer0_out[561] <= ~x[128] | x[129];
     layer0_out[562] <= x[271] | x[272];
     layer0_out[563] <= 1'b1;
     layer0_out[564] <= 1'b1;
     layer0_out[565] <= 1'b1;
     layer0_out[566] <= ~(x[283] | x[285]);
     layer0_out[567] <= ~(x[120] | x[122]);
     layer0_out[568] <= x[67];
     layer0_out[569] <= 1'b1;
     layer0_out[570] <= ~x[234];
     layer0_out[571] <= x[84] & x[86];
     layer0_out[572] <= x[304] & ~x[305];
     layer0_out[573] <= x[376] | x[378];
     layer0_out[574] <= ~(x[292] | x[293]);
     layer0_out[575] <= ~(x[373] | x[375]);
     layer0_out[576] <= x[25];
     layer0_out[577] <= x[313] | x[314];
     layer0_out[578] <= ~(x[220] | x[222]);
     layer0_out[579] <= ~(x[363] | x[365]);
     layer0_out[580] <= x[397];
     layer0_out[581] <= 1'b1;
     layer0_out[582] <= ~x[60] | x[58];
     layer0_out[583] <= ~(x[345] | x[346]);
     layer0_out[584] <= ~x[326] | x[328];
     layer0_out[585] <= ~(x[389] | x[390]);
     layer0_out[586] <= x[289] | x[290];
     layer0_out[587] <= 1'b0;
     layer0_out[588] <= 1'b0;
     layer0_out[589] <= x[65] | x[66];
     layer0_out[590] <= ~x[24];
     layer0_out[591] <= ~(x[52] | x[53]);
     layer0_out[592] <= ~x[89];
     layer0_out[593] <= x[201] & x[203];
     layer0_out[594] <= ~(x[19] | x[21]);
     layer0_out[595] <= 1'b1;
     layer0_out[596] <= ~(x[215] | x[217]);
     layer0_out[597] <= x[168] | x[169];
     layer0_out[598] <= ~(x[270] | x[272]);
     layer0_out[599] <= x[339];
     layer0_out[600] <= ~x[335];
     layer0_out[601] <= x[55] ^ x[56];
     layer0_out[602] <= x[133] & ~x[135];
     layer0_out[603] <= ~(x[102] | x[103]);
     layer0_out[604] <= x[258] | x[260];
     layer0_out[605] <= x[99] | x[100];
     layer0_out[606] <= ~(x[388] & x[389]);
     layer0_out[607] <= x[354] | x[356];
     layer0_out[608] <= ~x[298];
     layer0_out[609] <= x[180];
     layer0_out[610] <= 1'b0;
     layer0_out[611] <= ~x[88];
     layer0_out[612] <= x[101];
     layer0_out[613] <= x[314];
     layer0_out[614] <= x[145] ^ x[146];
     layer0_out[615] <= x[290] | x[291];
     layer0_out[616] <= x[243] & ~x[242];
     layer0_out[617] <= x[195] | x[196];
     layer0_out[618] <= x[346];
     layer0_out[619] <= x[167] | x[168];
     layer0_out[620] <= x[83] | x[85];
     layer0_out[621] <= 1'b0;
     layer0_out[622] <= ~(x[17] | x[18]);
     layer0_out[623] <= ~(x[356] | x[357]);
     layer0_out[624] <= x[107] | x[108];
     layer0_out[625] <= ~(x[39] & x[40]);
     layer0_out[626] <= 1'b0;
     layer0_out[627] <= x[63] | x[64];
     layer0_out[628] <= ~x[394] | x[395];
     layer0_out[629] <= ~(x[347] | x[349]);
     layer0_out[630] <= 1'b0;
     layer0_out[631] <= 1'b1;
     layer0_out[632] <= ~(x[196] | x[197]);
     layer0_out[633] <= ~(x[360] ^ x[361]);
     layer0_out[634] <= x[46] | x[47];
     layer0_out[635] <= ~(x[377] | x[379]);
     layer0_out[636] <= ~(x[324] | x[326]);
     layer0_out[637] <= ~x[107];
     layer0_out[638] <= ~(x[392] | x[394]);
     layer0_out[639] <= x[214] | x[215];
     layer0_out[640] <= 1'b0;
     layer0_out[641] <= ~x[162] | x[163];
     layer0_out[642] <= x[7] | x[9];
     layer0_out[643] <= 1'b0;
     layer0_out[644] <= x[260] & ~x[261];
     layer0_out[645] <= x[342] | x[344];
     layer0_out[646] <= x[85] | x[87];
     layer0_out[647] <= ~(x[318] | x[320]);
     layer0_out[648] <= ~(x[377] | x[378]);
     layer0_out[649] <= ~(x[216] | x[218]);
     layer0_out[650] <= x[94] & x[96];
     layer0_out[651] <= 1'b1;
     layer0_out[652] <= x[316];
     layer0_out[653] <= ~(x[316] | x[317]);
     layer0_out[654] <= x[80] | x[82];
     layer0_out[655] <= x[67] | x[69];
     layer0_out[656] <= ~(x[294] | x[296]);
     layer0_out[657] <= ~x[336];
     layer0_out[658] <= ~x[143];
     layer0_out[659] <= ~(x[303] | x[304]);
     layer0_out[660] <= x[177] | x[179];
     layer0_out[661] <= ~(x[98] & x[100]);
     layer0_out[662] <= ~x[37];
     layer0_out[663] <= 1'b0;
     layer0_out[664] <= x[384] | x[386];
     layer0_out[665] <= x[136] | x[138];
     layer0_out[666] <= 1'b1;
     layer0_out[667] <= x[178] | x[179];
     layer0_out[668] <= x[286] | x[287];
     layer0_out[669] <= ~x[47];
     layer0_out[670] <= x[216] | x[217];
     layer0_out[671] <= x[325] | x[326];
     layer0_out[672] <= 1'b0;
     layer0_out[673] <= x[22] & ~x[21];
     layer0_out[674] <= x[173] | x[174];
     layer0_out[675] <= ~x[138];
     layer0_out[676] <= ~(x[309] | x[311]);
     layer0_out[677] <= 1'b0;
     layer0_out[678] <= x[238] | x[240];
     layer0_out[679] <= x[321] | x[323];
     layer0_out[680] <= x[141] | x[143];
     layer0_out[681] <= x[247] & ~x[249];
     layer0_out[682] <= x[23] | x[24];
     layer0_out[683] <= x[161];
     layer0_out[684] <= ~(x[155] & x[156]);
     layer0_out[685] <= x[176] & ~x[178];
     layer0_out[686] <= ~(x[337] | x[338]);
     layer0_out[687] <= x[217] | x[218];
     layer0_out[688] <= ~(x[390] | x[391]);
     layer0_out[689] <= 1'b0;
     layer0_out[690] <= x[12] & ~x[14];
     layer0_out[691] <= ~(x[130] | x[132]);
     layer0_out[692] <= x[148];
     layer0_out[693] <= 1'b0;
     layer0_out[694] <= x[366] | x[368];
     layer0_out[695] <= x[144] | x[145];
     layer0_out[696] <= x[17] & ~x[15];
     layer0_out[697] <= x[321] | x[322];
     layer0_out[698] <= ~(x[32] | x[33]);
     layer0_out[699] <= ~(x[322] & x[323]);
     layer0_out[700] <= ~(x[329] | x[330]);
     layer0_out[701] <= 1'b1;
     layer0_out[702] <= ~(x[4] | x[6]);
     layer0_out[703] <= 1'b1;
     layer0_out[704] <= x[25] | x[27];
     layer0_out[705] <= x[240] | x[241];
     layer0_out[706] <= x[189] & ~x[190];
     layer0_out[707] <= ~(x[57] | x[58]);
     layer0_out[708] <= ~x[376];
     layer0_out[709] <= ~(x[140] | x[142]);
     layer0_out[710] <= x[153] | x[154];
     layer0_out[711] <= ~(x[176] | x[177]);
     layer0_out[712] <= ~(x[46] | x[48]);
     layer0_out[713] <= ~(x[288] | x[290]);
     layer0_out[714] <= 1'b0;
     layer0_out[715] <= x[86] | x[87];
     layer0_out[716] <= 1'b0;
     layer0_out[717] <= ~x[268] | x[270];
     layer0_out[718] <= x[228] | x[229];
     layer0_out[719] <= 1'b0;
     layer0_out[720] <= x[178] & ~x[177];
     layer0_out[721] <= x[295];
     layer0_out[722] <= ~(x[168] | x[170]);
     layer0_out[723] <= x[117] & ~x[119];
     layer0_out[724] <= ~x[358] | x[360];
     layer0_out[725] <= x[114] | x[115];
     layer0_out[726] <= x[241] | x[243];
     layer0_out[727] <= ~(x[6] | x[7]);
     layer0_out[728] <= ~x[317];
     layer0_out[729] <= ~x[299] | x[298];
     layer0_out[730] <= ~x[235];
     layer0_out[731] <= 1'b1;
     layer0_out[732] <= 1'b1;
     layer0_out[733] <= ~(x[71] & x[73]);
     layer0_out[734] <= ~(x[193] | x[195]);
     layer0_out[735] <= x[211] | x[212];
     layer0_out[736] <= x[346] | x[347];
     layer0_out[737] <= x[285];
     layer0_out[738] <= x[3];
     layer0_out[739] <= x[186] & ~x[187];
     layer0_out[740] <= ~(x[65] | x[67]);
     layer0_out[741] <= ~(x[227] | x[229]);
     layer0_out[742] <= x[346];
     layer0_out[743] <= ~(x[94] | x[95]);
     layer0_out[744] <= x[180] | x[181];
     layer0_out[745] <= x[282];
     layer0_out[746] <= 1'b1;
     layer0_out[747] <= 1'b0;
     layer0_out[748] <= x[151] | x[152];
     layer0_out[749] <= x[320];
     layer0_out[750] <= ~(x[34] | x[36]);
     layer0_out[751] <= x[362];
     layer0_out[752] <= ~(x[202] | x[204]);
     layer0_out[753] <= ~(x[359] | x[360]);
     layer0_out[754] <= 1'b0;
     layer0_out[755] <= ~(x[230] | x[232]);
     layer0_out[756] <= x[13];
     layer0_out[757] <= 1'b0;
     layer0_out[758] <= 1'b0;
     layer0_out[759] <= ~x[185];
     layer0_out[760] <= ~(x[127] | x[128]);
     layer0_out[761] <= 1'b1;
     layer0_out[762] <= ~x[146];
     layer0_out[763] <= ~x[175];
     layer0_out[764] <= 1'b0;
     layer0_out[765] <= x[1] | x[2];
     layer0_out[766] <= ~x[101] | x[99];
     layer0_out[767] <= 1'b1;
     layer0_out[768] <= 1'b0;
     layer0_out[769] <= 1'b1;
     layer0_out[770] <= 1'b1;
     layer0_out[771] <= 1'b0;
     layer0_out[772] <= 1'b0;
     layer0_out[773] <= ~(x[356] | x[358]);
     layer0_out[774] <= ~(x[317] | x[318]);
     layer0_out[775] <= ~x[221] | x[220];
     layer0_out[776] <= x[370] | x[371];
     layer0_out[777] <= x[203];
     layer0_out[778] <= ~(x[219] | x[221]);
     layer0_out[779] <= x[349] | x[350];
     layer0_out[780] <= ~(x[191] | x[193]);
     layer0_out[781] <= x[28];
     layer0_out[782] <= x[351] | x[353];
     layer0_out[783] <= 1'b0;
     layer0_out[784] <= ~(x[231] | x[233]);
     layer0_out[785] <= ~x[322] | x[320];
     layer0_out[786] <= x[305] ^ x[307];
     layer0_out[787] <= ~(x[240] & x[242]);
     layer0_out[788] <= ~(x[87] | x[89]);
     layer0_out[789] <= x[332];
     layer0_out[790] <= ~(x[305] & x[306]);
     layer0_out[791] <= x[192] | x[193];
     layer0_out[792] <= x[256] | x[258];
     layer0_out[793] <= x[31] ^ x[33];
     layer0_out[794] <= ~(x[383] ^ x[385]);
     layer0_out[795] <= x[43];
     layer0_out[796] <= x[304] ^ x[306];
     layer0_out[797] <= x[393];
     layer0_out[798] <= 1'b0;
     layer0_out[799] <= 1'b1;
     layer1_out[0] <= ~layer0_out[270];
     layer1_out[1] <= layer0_out[325];
     layer1_out[2] <= layer0_out[760];
     layer1_out[3] <= layer0_out[150];
     layer1_out[4] <= ~layer0_out[674];
     layer1_out[5] <= layer0_out[199];
     layer1_out[6] <= ~(layer0_out[206] | layer0_out[207]);
     layer1_out[7] <= ~layer0_out[32] | layer0_out[31];
     layer1_out[8] <= ~layer0_out[366];
     layer1_out[9] <= ~(layer0_out[639] & layer0_out[640]);
     layer1_out[10] <= ~layer0_out[467] | layer0_out[466];
     layer1_out[11] <= layer0_out[198] | layer0_out[199];
     layer1_out[12] <= ~(layer0_out[482] | layer0_out[483]);
     layer1_out[13] <= ~(layer0_out[65] | layer0_out[66]);
     layer1_out[14] <= ~layer0_out[712] | layer0_out[713];
     layer1_out[15] <= layer0_out[275] & layer0_out[276];
     layer1_out[16] <= ~layer0_out[450];
     layer1_out[17] <= ~layer0_out[708] | layer0_out[709];
     layer1_out[18] <= layer0_out[762] & ~layer0_out[761];
     layer1_out[19] <= layer0_out[768] | layer0_out[769];
     layer1_out[20] <= layer0_out[522] & ~layer0_out[521];
     layer1_out[21] <= ~(layer0_out[164] | layer0_out[165]);
     layer1_out[22] <= layer0_out[0] & ~layer0_out[1];
     layer1_out[23] <= ~layer0_out[691] | layer0_out[692];
     layer1_out[24] <= ~layer0_out[110];
     layer1_out[25] <= layer0_out[692] & ~layer0_out[693];
     layer1_out[26] <= layer0_out[330] & layer0_out[331];
     layer1_out[27] <= 1'b0;
     layer1_out[28] <= 1'b0;
     layer1_out[29] <= ~layer0_out[282] | layer0_out[283];
     layer1_out[30] <= ~(layer0_out[655] | layer0_out[656]);
     layer1_out[31] <= 1'b1;
     layer1_out[32] <= ~layer0_out[95] | layer0_out[96];
     layer1_out[33] <= layer0_out[327] | layer0_out[328];
     layer1_out[34] <= 1'b1;
     layer1_out[35] <= ~layer0_out[454];
     layer1_out[36] <= layer0_out[244];
     layer1_out[37] <= ~layer0_out[612] | layer0_out[613];
     layer1_out[38] <= 1'b1;
     layer1_out[39] <= 1'b0;
     layer1_out[40] <= layer0_out[334] & ~layer0_out[335];
     layer1_out[41] <= ~layer0_out[603];
     layer1_out[42] <= layer0_out[208];
     layer1_out[43] <= layer0_out[323];
     layer1_out[44] <= 1'b0;
     layer1_out[45] <= layer0_out[656];
     layer1_out[46] <= layer0_out[34] & ~layer0_out[33];
     layer1_out[47] <= 1'b0;
     layer1_out[48] <= layer0_out[271] | layer0_out[272];
     layer1_out[49] <= layer0_out[528] & ~layer0_out[527];
     layer1_out[50] <= ~(layer0_out[389] ^ layer0_out[390]);
     layer1_out[51] <= ~layer0_out[8];
     layer1_out[52] <= ~layer0_out[661] | layer0_out[662];
     layer1_out[53] <= 1'b0;
     layer1_out[54] <= layer0_out[232];
     layer1_out[55] <= ~(layer0_out[416] & layer0_out[417]);
     layer1_out[56] <= ~layer0_out[641] | layer0_out[642];
     layer1_out[57] <= layer0_out[4];
     layer1_out[58] <= layer0_out[317];
     layer1_out[59] <= 1'b1;
     layer1_out[60] <= 1'b1;
     layer1_out[61] <= ~(layer0_out[126] & layer0_out[127]);
     layer1_out[62] <= ~layer0_out[556] | layer0_out[557];
     layer1_out[63] <= layer0_out[152];
     layer1_out[64] <= 1'b0;
     layer1_out[65] <= ~layer0_out[743];
     layer1_out[66] <= ~layer0_out[461] | layer0_out[462];
     layer1_out[67] <= layer0_out[606] & ~layer0_out[605];
     layer1_out[68] <= 1'b1;
     layer1_out[69] <= ~(layer0_out[56] ^ layer0_out[57]);
     layer1_out[70] <= ~layer0_out[347];
     layer1_out[71] <= ~(layer0_out[599] & layer0_out[600]);
     layer1_out[72] <= ~layer0_out[35] | layer0_out[36];
     layer1_out[73] <= layer0_out[513];
     layer1_out[74] <= layer0_out[391];
     layer1_out[75] <= layer0_out[681];
     layer1_out[76] <= layer0_out[284] | layer0_out[285];
     layer1_out[77] <= layer0_out[81];
     layer1_out[78] <= layer0_out[161] & ~layer0_out[162];
     layer1_out[79] <= layer0_out[298];
     layer1_out[80] <= 1'b0;
     layer1_out[81] <= ~layer0_out[502] | layer0_out[503];
     layer1_out[82] <= layer0_out[168];
     layer1_out[83] <= layer0_out[91] & ~layer0_out[90];
     layer1_out[84] <= ~(layer0_out[695] | layer0_out[696]);
     layer1_out[85] <= ~(layer0_out[499] | layer0_out[500]);
     layer1_out[86] <= ~layer0_out[223];
     layer1_out[87] <= layer0_out[664];
     layer1_out[88] <= layer0_out[402];
     layer1_out[89] <= layer0_out[400];
     layer1_out[90] <= layer0_out[173] & ~layer0_out[174];
     layer1_out[91] <= ~(layer0_out[105] & layer0_out[106]);
     layer1_out[92] <= ~layer0_out[358] | layer0_out[357];
     layer1_out[93] <= ~layer0_out[181];
     layer1_out[94] <= ~layer0_out[638];
     layer1_out[95] <= 1'b0;
     layer1_out[96] <= 1'b0;
     layer1_out[97] <= 1'b0;
     layer1_out[98] <= layer0_out[134];
     layer1_out[99] <= layer0_out[439] & layer0_out[440];
     layer1_out[100] <= layer0_out[754] & ~layer0_out[755];
     layer1_out[101] <= ~layer0_out[118] | layer0_out[119];
     layer1_out[102] <= layer0_out[20] | layer0_out[21];
     layer1_out[103] <= layer0_out[781];
     layer1_out[104] <= layer0_out[497] & layer0_out[498];
     layer1_out[105] <= layer0_out[566] | layer0_out[567];
     layer1_out[106] <= ~layer0_out[724] | layer0_out[725];
     layer1_out[107] <= layer0_out[786] | layer0_out[787];
     layer1_out[108] <= layer0_out[417];
     layer1_out[109] <= layer0_out[505] | layer0_out[506];
     layer1_out[110] <= layer0_out[292];
     layer1_out[111] <= 1'b0;
     layer1_out[112] <= 1'b1;
     layer1_out[113] <= 1'b0;
     layer1_out[114] <= layer0_out[418] | layer0_out[419];
     layer1_out[115] <= layer0_out[677] | layer0_out[678];
     layer1_out[116] <= ~(layer0_out[476] & layer0_out[477]);
     layer1_out[117] <= ~layer0_out[165];
     layer1_out[118] <= layer0_out[35] & ~layer0_out[34];
     layer1_out[119] <= 1'b1;
     layer1_out[120] <= layer0_out[534] & ~layer0_out[535];
     layer1_out[121] <= layer0_out[632] & layer0_out[633];
     layer1_out[122] <= ~(layer0_out[340] & layer0_out[341]);
     layer1_out[123] <= ~layer0_out[172] | layer0_out[173];
     layer1_out[124] <= 1'b1;
     layer1_out[125] <= layer0_out[264] | layer0_out[265];
     layer1_out[126] <= ~layer0_out[243];
     layer1_out[127] <= ~layer0_out[437];
     layer1_out[128] <= layer0_out[397] | layer0_out[398];
     layer1_out[129] <= 1'b0;
     layer1_out[130] <= ~layer0_out[541];
     layer1_out[131] <= ~layer0_out[84];
     layer1_out[132] <= layer0_out[10] & ~layer0_out[9];
     layer1_out[133] <= ~(layer0_out[696] | layer0_out[697]);
     layer1_out[134] <= ~layer0_out[311] | layer0_out[310];
     layer1_out[135] <= ~layer0_out[303];
     layer1_out[136] <= ~(layer0_out[39] & layer0_out[40]);
     layer1_out[137] <= layer0_out[430];
     layer1_out[138] <= 1'b1;
     layer1_out[139] <= layer0_out[629] & layer0_out[630];
     layer1_out[140] <= ~layer0_out[333];
     layer1_out[141] <= layer0_out[396] & layer0_out[397];
     layer1_out[142] <= 1'b1;
     layer1_out[143] <= layer0_out[472] & ~layer0_out[471];
     layer1_out[144] <= 1'b1;
     layer1_out[145] <= layer0_out[639];
     layer1_out[146] <= 1'b1;
     layer1_out[147] <= ~layer0_out[355] | layer0_out[356];
     layer1_out[148] <= layer0_out[644] & layer0_out[645];
     layer1_out[149] <= ~(layer0_out[789] | layer0_out[790]);
     layer1_out[150] <= ~layer0_out[564] | layer0_out[563];
     layer1_out[151] <= layer0_out[654];
     layer1_out[152] <= 1'b0;
     layer1_out[153] <= layer0_out[771];
     layer1_out[154] <= ~layer0_out[327];
     layer1_out[155] <= layer0_out[248];
     layer1_out[156] <= ~(layer0_out[259] | layer0_out[260]);
     layer1_out[157] <= layer0_out[253];
     layer1_out[158] <= ~layer0_out[263];
     layer1_out[159] <= 1'b1;
     layer1_out[160] <= ~layer0_out[478];
     layer1_out[161] <= ~layer0_out[70];
     layer1_out[162] <= ~layer0_out[730] | layer0_out[731];
     layer1_out[163] <= layer0_out[336] & layer0_out[337];
     layer1_out[164] <= layer0_out[544];
     layer1_out[165] <= layer0_out[214];
     layer1_out[166] <= ~(layer0_out[584] & layer0_out[585]);
     layer1_out[167] <= layer0_out[354];
     layer1_out[168] <= ~layer0_out[595];
     layer1_out[169] <= ~layer0_out[713] | layer0_out[714];
     layer1_out[170] <= layer0_out[329] | layer0_out[330];
     layer1_out[171] <= layer0_out[539];
     layer1_out[172] <= ~(layer0_out[434] | layer0_out[435]);
     layer1_out[173] <= layer0_out[633];
     layer1_out[174] <= layer0_out[450] & ~layer0_out[451];
     layer1_out[175] <= layer0_out[764] & layer0_out[765];
     layer1_out[176] <= ~(layer0_out[710] | layer0_out[711]);
     layer1_out[177] <= layer0_out[352];
     layer1_out[178] <= ~(layer0_out[438] & layer0_out[439]);
     layer1_out[179] <= layer0_out[494] & layer0_out[495];
     layer1_out[180] <= ~(layer0_out[548] & layer0_out[549]);
     layer1_out[181] <= ~layer0_out[99];
     layer1_out[182] <= layer0_out[177] | layer0_out[178];
     layer1_out[183] <= ~(layer0_out[788] | layer0_out[789]);
     layer1_out[184] <= 1'b0;
     layer1_out[185] <= layer0_out[79] | layer0_out[80];
     layer1_out[186] <= ~layer0_out[266] | layer0_out[267];
     layer1_out[187] <= 1'b1;
     layer1_out[188] <= ~layer0_out[374] | layer0_out[373];
     layer1_out[189] <= layer0_out[370] | layer0_out[371];
     layer1_out[190] <= ~layer0_out[560];
     layer1_out[191] <= layer0_out[606] & layer0_out[607];
     layer1_out[192] <= ~(layer0_out[117] & layer0_out[118]);
     layer1_out[193] <= ~layer0_out[381];
     layer1_out[194] <= ~layer0_out[675];
     layer1_out[195] <= ~(layer0_out[659] | layer0_out[660]);
     layer1_out[196] <= ~layer0_out[716];
     layer1_out[197] <= ~layer0_out[16] | layer0_out[15];
     layer1_out[198] <= layer0_out[667];
     layer1_out[199] <= ~(layer0_out[580] | layer0_out[581]);
     layer1_out[200] <= ~layer0_out[773];
     layer1_out[201] <= layer0_out[643];
     layer1_out[202] <= ~(layer0_out[487] | layer0_out[488]);
     layer1_out[203] <= layer0_out[104];
     layer1_out[204] <= ~layer0_out[185] | layer0_out[186];
     layer1_out[205] <= layer0_out[627] | layer0_out[628];
     layer1_out[206] <= ~layer0_out[779] | layer0_out[778];
     layer1_out[207] <= layer0_out[211] | layer0_out[212];
     layer1_out[208] <= layer0_out[658] & ~layer0_out[659];
     layer1_out[209] <= layer0_out[532] & layer0_out[533];
     layer1_out[210] <= layer0_out[279] & ~layer0_out[280];
     layer1_out[211] <= ~layer0_out[8] | layer0_out[9];
     layer1_out[212] <= 1'b1;
     layer1_out[213] <= ~(layer0_out[578] & layer0_out[579]);
     layer1_out[214] <= ~layer0_out[72];
     layer1_out[215] <= ~(layer0_out[210] & layer0_out[211]);
     layer1_out[216] <= ~(layer0_out[70] & layer0_out[71]);
     layer1_out[217] <= layer0_out[115] | layer0_out[116];
     layer1_out[218] <= 1'b1;
     layer1_out[219] <= layer0_out[568];
     layer1_out[220] <= layer0_out[720];
     layer1_out[221] <= ~(layer0_out[619] | layer0_out[620]);
     layer1_out[222] <= 1'b0;
     layer1_out[223] <= 1'b0;
     layer1_out[224] <= ~(layer0_out[733] & layer0_out[734]);
     layer1_out[225] <= layer0_out[44] | layer0_out[45];
     layer1_out[226] <= layer0_out[209];
     layer1_out[227] <= layer0_out[234];
     layer1_out[228] <= layer0_out[495] | layer0_out[496];
     layer1_out[229] <= ~(layer0_out[672] & layer0_out[673]);
     layer1_out[230] <= layer0_out[125];
     layer1_out[231] <= ~(layer0_out[26] & layer0_out[27]);
     layer1_out[232] <= ~layer0_out[458] | layer0_out[457];
     layer1_out[233] <= layer0_out[102] | layer0_out[103];
     layer1_out[234] <= layer0_out[519];
     layer1_out[235] <= ~layer0_out[0] | layer0_out[2];
     layer1_out[236] <= 1'b1;
     layer1_out[237] <= layer0_out[279] & ~layer0_out[278];
     layer1_out[238] <= layer0_out[343] & ~layer0_out[344];
     layer1_out[239] <= ~(layer0_out[709] & layer0_out[710]);
     layer1_out[240] <= layer0_out[166];
     layer1_out[241] <= 1'b1;
     layer1_out[242] <= layer0_out[722];
     layer1_out[243] <= layer0_out[729];
     layer1_out[244] <= layer0_out[323] & ~layer0_out[322];
     layer1_out[245] <= layer0_out[223];
     layer1_out[246] <= ~layer0_out[704] | layer0_out[703];
     layer1_out[247] <= layer0_out[59] & ~layer0_out[60];
     layer1_out[248] <= 1'b0;
     layer1_out[249] <= ~layer0_out[701];
     layer1_out[250] <= 1'b1;
     layer1_out[251] <= layer0_out[396];
     layer1_out[252] <= layer0_out[16] & ~layer0_out[17];
     layer1_out[253] <= layer0_out[562];
     layer1_out[254] <= ~layer0_out[106];
     layer1_out[255] <= ~(layer0_out[759] & layer0_out[760]);
     layer1_out[256] <= 1'b0;
     layer1_out[257] <= ~layer0_out[405] | layer0_out[404];
     layer1_out[258] <= layer0_out[777] & layer0_out[778];
     layer1_out[259] <= layer0_out[740] & layer0_out[741];
     layer1_out[260] <= layer0_out[545];
     layer1_out[261] <= layer0_out[414] & ~layer0_out[413];
     layer1_out[262] <= layer0_out[60] & ~layer0_out[61];
     layer1_out[263] <= ~layer0_out[456];
     layer1_out[264] <= ~(layer0_out[514] | layer0_out[515]);
     layer1_out[265] <= ~layer0_out[232];
     layer1_out[266] <= ~layer0_out[348];
     layer1_out[267] <= ~layer0_out[309];
     layer1_out[268] <= ~(layer0_out[419] & layer0_out[420]);
     layer1_out[269] <= 1'b0;
     layer1_out[270] <= layer0_out[345] & layer0_out[346];
     layer1_out[271] <= 1'b1;
     layer1_out[272] <= 1'b1;
     layer1_out[273] <= layer0_out[160] | layer0_out[161];
     layer1_out[274] <= layer0_out[737] & layer0_out[738];
     layer1_out[275] <= layer0_out[770] & ~layer0_out[769];
     layer1_out[276] <= 1'b1;
     layer1_out[277] <= ~layer0_out[685] | layer0_out[684];
     layer1_out[278] <= layer0_out[339];
     layer1_out[279] <= ~layer0_out[537] | layer0_out[536];
     layer1_out[280] <= ~layer0_out[83] | layer0_out[82];
     layer1_out[281] <= ~(layer0_out[762] ^ layer0_out[763]);
     layer1_out[282] <= ~(layer0_out[375] | layer0_out[376]);
     layer1_out[283] <= layer0_out[256] & ~layer0_out[255];
     layer1_out[284] <= ~layer0_out[717] | layer0_out[718];
     layer1_out[285] <= layer0_out[422] & ~layer0_out[423];
     layer1_out[286] <= layer0_out[580];
     layer1_out[287] <= ~layer0_out[490];
     layer1_out[288] <= ~layer0_out[183];
     layer1_out[289] <= ~layer0_out[50];
     layer1_out[290] <= ~layer0_out[485];
     layer1_out[291] <= ~(layer0_out[321] & layer0_out[322]);
     layer1_out[292] <= 1'b1;
     layer1_out[293] <= 1'b0;
     layer1_out[294] <= layer0_out[28];
     layer1_out[295] <= 1'b0;
     layer1_out[296] <= layer0_out[435] | layer0_out[436];
     layer1_out[297] <= 1'b0;
     layer1_out[298] <= 1'b1;
     layer1_out[299] <= layer0_out[275] & ~layer0_out[274];
     layer1_out[300] <= 1'b1;
     layer1_out[301] <= ~layer0_out[184];
     layer1_out[302] <= ~layer0_out[281];
     layer1_out[303] <= 1'b1;
     layer1_out[304] <= ~layer0_out[766];
     layer1_out[305] <= ~layer0_out[52];
     layer1_out[306] <= ~layer0_out[241];
     layer1_out[307] <= 1'b0;
     layer1_out[308] <= ~layer0_out[129] | layer0_out[128];
     layer1_out[309] <= ~(layer0_out[673] & layer0_out[674]);
     layer1_out[310] <= ~layer0_out[324] | layer0_out[325];
     layer1_out[311] <= layer0_out[602] & ~layer0_out[603];
     layer1_out[312] <= 1'b1;
     layer1_out[313] <= ~layer0_out[188];
     layer1_out[314] <= layer0_out[178] & layer0_out[179];
     layer1_out[315] <= 1'b0;
     layer1_out[316] <= ~layer0_out[575] | layer0_out[576];
     layer1_out[317] <= ~layer0_out[87];
     layer1_out[318] <= 1'b0;
     layer1_out[319] <= layer0_out[624] & ~layer0_out[625];
     layer1_out[320] <= layer0_out[748] | layer0_out[749];
     layer1_out[321] <= ~(layer0_out[205] & layer0_out[206]);
     layer1_out[322] <= 1'b1;
     layer1_out[323] <= ~layer0_out[794] | layer0_out[795];
     layer1_out[324] <= ~layer0_out[284] | layer0_out[283];
     layer1_out[325] <= layer0_out[18] & ~layer0_out[17];
     layer1_out[326] <= layer0_out[644];
     layer1_out[327] <= layer0_out[380] ^ layer0_out[381];
     layer1_out[328] <= 1'b0;
     layer1_out[329] <= layer0_out[785] & ~layer0_out[784];
     layer1_out[330] <= layer0_out[682] ^ layer0_out[683];
     layer1_out[331] <= layer0_out[635] & ~layer0_out[636];
     layer1_out[332] <= ~layer0_out[461];
     layer1_out[333] <= layer0_out[409] & ~layer0_out[410];
     layer1_out[334] <= 1'b1;
     layer1_out[335] <= layer0_out[66];
     layer1_out[336] <= ~layer0_out[226];
     layer1_out[337] <= layer0_out[705] & layer0_out[706];
     layer1_out[338] <= layer0_out[386];
     layer1_out[339] <= ~layer0_out[651] | layer0_out[652];
     layer1_out[340] <= 1'b0;
     layer1_out[341] <= 1'b1;
     layer1_out[342] <= ~layer0_out[272];
     layer1_out[343] <= layer0_out[615];
     layer1_out[344] <= 1'b1;
     layer1_out[345] <= ~layer0_out[156] | layer0_out[157];
     layer1_out[346] <= ~layer0_out[246] | layer0_out[245];
     layer1_out[347] <= 1'b1;
     layer1_out[348] <= layer0_out[94] & ~layer0_out[95];
     layer1_out[349] <= ~layer0_out[443] | layer0_out[444];
     layer1_out[350] <= 1'b0;
     layer1_out[351] <= layer0_out[715] | layer0_out[716];
     layer1_out[352] <= ~layer0_out[695];
     layer1_out[353] <= 1'b1;
     layer1_out[354] <= layer0_out[492] & ~layer0_out[491];
     layer1_out[355] <= layer0_out[133] & ~layer0_out[134];
     layer1_out[356] <= ~(layer0_out[468] | layer0_out[469]);
     layer1_out[357] <= 1'b1;
     layer1_out[358] <= ~layer0_out[702];
     layer1_out[359] <= ~(layer0_out[191] | layer0_out[192]);
     layer1_out[360] <= layer0_out[136] & ~layer0_out[135];
     layer1_out[361] <= 1'b1;
     layer1_out[362] <= 1'b1;
     layer1_out[363] <= layer0_out[197] | layer0_out[198];
     layer1_out[364] <= layer0_out[295];
     layer1_out[365] <= ~(layer0_out[242] | layer0_out[243]);
     layer1_out[366] <= 1'b0;
     layer1_out[367] <= layer0_out[497];
     layer1_out[368] <= 1'b0;
     layer1_out[369] <= ~layer0_out[566];
     layer1_out[370] <= ~layer0_out[679] | layer0_out[680];
     layer1_out[371] <= layer0_out[507];
     layer1_out[372] <= layer0_out[154] & layer0_out[155];
     layer1_out[373] <= layer0_out[41] | layer0_out[42];
     layer1_out[374] <= layer0_out[101] & layer0_out[102];
     layer1_out[375] <= layer0_out[315];
     layer1_out[376] <= layer0_out[293];
     layer1_out[377] <= layer0_out[45] | layer0_out[46];
     layer1_out[378] <= layer0_out[763];
     layer1_out[379] <= 1'b1;
     layer1_out[380] <= ~layer0_out[203];
     layer1_out[381] <= ~layer0_out[792] | layer0_out[791];
     layer1_out[382] <= layer0_out[507] & ~layer0_out[508];
     layer1_out[383] <= ~(layer0_out[475] ^ layer0_out[476]);
     layer1_out[384] <= 1'b1;
     layer1_out[385] <= 1'b0;
     layer1_out[386] <= ~(layer0_out[503] | layer0_out[504]);
     layer1_out[387] <= layer0_out[446];
     layer1_out[388] <= 1'b0;
     layer1_out[389] <= ~layer0_out[597] | layer0_out[596];
     layer1_out[390] <= ~(layer0_out[174] | layer0_out[175]);
     layer1_out[391] <= layer0_out[312] | layer0_out[313];
     layer1_out[392] <= 1'b1;
     layer1_out[393] <= ~layer0_out[408] | layer0_out[407];
     layer1_out[394] <= ~(layer0_out[465] | layer0_out[466]);
     layer1_out[395] <= layer0_out[235] | layer0_out[236];
     layer1_out[396] <= 1'b1;
     layer1_out[397] <= ~layer0_out[239] | layer0_out[240];
     layer1_out[398] <= layer0_out[23];
     layer1_out[399] <= 1'b0;
     layer1_out[400] <= ~layer0_out[69] | layer0_out[68];
     layer1_out[401] <= ~(layer0_out[570] & layer0_out[571]);
     layer1_out[402] <= ~layer0_out[303];
     layer1_out[403] <= layer0_out[316] & layer0_out[317];
     layer1_out[404] <= layer0_out[201];
     layer1_out[405] <= ~layer0_out[753];
     layer1_out[406] <= ~(layer0_out[749] ^ layer0_out[750]);
     layer1_out[407] <= ~layer0_out[736];
     layer1_out[408] <= layer0_out[94] & ~layer0_out[93];
     layer1_out[409] <= layer0_out[572];
     layer1_out[410] <= 1'b1;
     layer1_out[411] <= 1'b1;
     layer1_out[412] <= ~(layer0_out[351] & layer0_out[352]);
     layer1_out[413] <= layer0_out[448] & layer0_out[449];
     layer1_out[414] <= layer0_out[547] & layer0_out[548];
     layer1_out[415] <= layer0_out[220] & ~layer0_out[221];
     layer1_out[416] <= layer0_out[732];
     layer1_out[417] <= ~layer0_out[61];
     layer1_out[418] <= layer0_out[651] & ~layer0_out[650];
     layer1_out[419] <= ~layer0_out[338];
     layer1_out[420] <= ~layer0_out[137] | layer0_out[136];
     layer1_out[421] <= layer0_out[540];
     layer1_out[422] <= ~layer0_out[573];
     layer1_out[423] <= ~layer0_out[292];
     layer1_out[424] <= 1'b0;
     layer1_out[425] <= ~layer0_out[658];
     layer1_out[426] <= layer0_out[116] & layer0_out[117];
     layer1_out[427] <= ~layer0_out[28];
     layer1_out[428] <= ~layer0_out[170] | layer0_out[171];
     layer1_out[429] <= layer0_out[687] | layer0_out[688];
     layer1_out[430] <= ~layer0_out[200];
     layer1_out[431] <= layer0_out[158] ^ layer0_out[159];
     layer1_out[432] <= layer0_out[702] | layer0_out[703];
     layer1_out[433] <= 1'b1;
     layer1_out[434] <= ~layer0_out[163] | layer0_out[164];
     layer1_out[435] <= ~layer0_out[65];
     layer1_out[436] <= layer0_out[23] & ~layer0_out[24];
     layer1_out[437] <= 1'b1;
     layer1_out[438] <= 1'b0;
     layer1_out[439] <= layer0_out[678] & layer0_out[679];
     layer1_out[440] <= layer0_out[464];
     layer1_out[441] <= ~layer0_out[186] | layer0_out[187];
     layer1_out[442] <= ~(layer0_out[287] & layer0_out[288]);
     layer1_out[443] <= layer0_out[287];
     layer1_out[444] <= layer0_out[551];
     layer1_out[445] <= layer0_out[747];
     layer1_out[446] <= layer0_out[712];
     layer1_out[447] <= layer0_out[574] & layer0_out[575];
     layer1_out[448] <= layer0_out[234];
     layer1_out[449] <= layer0_out[72] & layer0_out[73];
     layer1_out[450] <= ~layer0_out[547] | layer0_out[546];
     layer1_out[451] <= layer0_out[786] & ~layer0_out[785];
     layer1_out[452] <= ~(layer0_out[256] & layer0_out[257]);
     layer1_out[453] <= 1'b1;
     layer1_out[454] <= layer0_out[641] & ~layer0_out[640];
     layer1_out[455] <= ~layer0_out[649];
     layer1_out[456] <= ~layer0_out[502];
     layer1_out[457] <= ~layer0_out[226] | layer0_out[227];
     layer1_out[458] <= layer0_out[141] & ~layer0_out[140];
     layer1_out[459] <= ~(layer0_out[263] & layer0_out[264]);
     layer1_out[460] <= layer0_out[157] & layer0_out[158];
     layer1_out[461] <= layer0_out[366] & ~layer0_out[367];
     layer1_out[462] <= ~layer0_out[669];
     layer1_out[463] <= layer0_out[793] | layer0_out[794];
     layer1_out[464] <= ~layer0_out[597] | layer0_out[598];
     layer1_out[465] <= ~layer0_out[780];
     layer1_out[466] <= layer0_out[441];
     layer1_out[467] <= layer0_out[425];
     layer1_out[468] <= layer0_out[471];
     layer1_out[469] <= layer0_out[137];
     layer1_out[470] <= ~layer0_out[483] | layer0_out[484];
     layer1_out[471] <= 1'b0;
     layer1_out[472] <= 1'b0;
     layer1_out[473] <= layer0_out[662] & layer0_out[663];
     layer1_out[474] <= ~layer0_out[357];
     layer1_out[475] <= layer0_out[646];
     layer1_out[476] <= ~layer0_out[590] | layer0_out[589];
     layer1_out[477] <= ~layer0_out[395] | layer0_out[394];
     layer1_out[478] <= ~layer0_out[475];
     layer1_out[479] <= ~layer0_out[494];
     layer1_out[480] <= ~layer0_out[453] | layer0_out[452];
     layer1_out[481] <= ~(layer0_out[62] | layer0_out[63]);
     layer1_out[482] <= 1'b1;
     layer1_out[483] <= layer0_out[53] & layer0_out[54];
     layer1_out[484] <= ~layer0_out[759];
     layer1_out[485] <= ~layer0_out[472] | layer0_out[473];
     layer1_out[486] <= layer0_out[260];
     layer1_out[487] <= ~layer0_out[683];
     layer1_out[488] <= ~layer0_out[349] | layer0_out[350];
     layer1_out[489] <= ~layer0_out[195];
     layer1_out[490] <= layer0_out[790];
     layer1_out[491] <= layer0_out[490];
     layer1_out[492] <= ~layer0_out[554];
     layer1_out[493] <= ~layer0_out[528];
     layer1_out[494] <= ~layer0_out[270];
     layer1_out[495] <= layer0_out[114];
     layer1_out[496] <= ~(layer0_out[522] & layer0_out[523]);
     layer1_out[497] <= layer0_out[1];
     layer1_out[498] <= ~(layer0_out[688] & layer0_out[689]);
     layer1_out[499] <= layer0_out[228] | layer0_out[229];
     layer1_out[500] <= 1'b0;
     layer1_out[501] <= ~layer0_out[715];
     layer1_out[502] <= layer0_out[721] & ~layer0_out[722];
     layer1_out[503] <= layer0_out[19] & ~layer0_out[20];
     layer1_out[504] <= layer0_out[305] | layer0_out[306];
     layer1_out[505] <= ~layer0_out[570];
     layer1_out[506] <= ~layer0_out[742];
     layer1_out[507] <= ~layer0_out[43];
     layer1_out[508] <= layer0_out[149];
     layer1_out[509] <= ~layer0_out[757];
     layer1_out[510] <= ~(layer0_out[169] | layer0_out[170]);
     layer1_out[511] <= layer0_out[482];
     layer1_out[512] <= layer0_out[511];
     layer1_out[513] <= layer0_out[589];
     layer1_out[514] <= ~layer0_out[289];
     layer1_out[515] <= ~layer0_out[130];
     layer1_out[516] <= layer0_out[328] | layer0_out[329];
     layer1_out[517] <= layer0_out[389] & ~layer0_out[388];
     layer1_out[518] <= ~layer0_out[780];
     layer1_out[519] <= ~layer0_out[797];
     layer1_out[520] <= ~layer0_out[408] | layer0_out[409];
     layer1_out[521] <= layer0_out[159] | layer0_out[160];
     layer1_out[522] <= ~layer0_out[616];
     layer1_out[523] <= layer0_out[276] | layer0_out[277];
     layer1_out[524] <= layer0_out[216];
     layer1_out[525] <= ~layer0_out[552] | layer0_out[551];
     layer1_out[526] <= ~(layer0_out[442] | layer0_out[443]);
     layer1_out[527] <= ~layer0_out[41] | layer0_out[40];
     layer1_out[528] <= layer0_out[751];
     layer1_out[529] <= ~layer0_out[250];
     layer1_out[530] <= 1'b1;
     layer1_out[531] <= layer0_out[212];
     layer1_out[532] <= ~(layer0_out[308] & layer0_out[309]);
     layer1_out[533] <= layer0_out[610] & ~layer0_out[609];
     layer1_out[534] <= ~(layer0_out[143] & layer0_out[144]);
     layer1_out[535] <= 1'b0;
     layer1_out[536] <= layer0_out[720] | layer0_out[721];
     layer1_out[537] <= ~layer0_out[636];
     layer1_out[538] <= layer0_out[480] | layer0_out[481];
     layer1_out[539] <= layer0_out[376] & ~layer0_out[377];
     layer1_out[540] <= ~layer0_out[247] | layer0_out[246];
     layer1_out[541] <= layer0_out[776];
     layer1_out[542] <= layer0_out[519] | layer0_out[520];
     layer1_out[543] <= ~layer0_out[121] | layer0_out[122];
     layer1_out[544] <= layer0_out[424] & layer0_out[425];
     layer1_out[545] <= ~(layer0_out[458] & layer0_out[459]);
     layer1_out[546] <= ~layer0_out[399] | layer0_out[400];
     layer1_out[547] <= 1'b1;
     layer1_out[548] <= ~layer0_out[214] | layer0_out[213];
     layer1_out[549] <= ~layer0_out[36];
     layer1_out[550] <= ~layer0_out[259] | layer0_out[258];
     layer1_out[551] <= layer0_out[108];
     layer1_out[552] <= layer0_out[576] & ~layer0_out[577];
     layer1_out[553] <= layer0_out[163];
     layer1_out[554] <= ~layer0_out[426] | layer0_out[427];
     layer1_out[555] <= layer0_out[76] & ~layer0_out[77];
     layer1_out[556] <= layer0_out[222] & ~layer0_out[221];
     layer1_out[557] <= ~layer0_out[402] | layer0_out[401];
     layer1_out[558] <= layer0_out[153] & ~layer0_out[152];
     layer1_out[559] <= ~layer0_out[120];
     layer1_out[560] <= ~layer0_out[153];
     layer1_out[561] <= layer0_out[433];
     layer1_out[562] <= ~(layer0_out[192] & layer0_out[193]);
     layer1_out[563] <= 1'b0;
     layer1_out[564] <= layer0_out[768] & ~layer0_out[767];
     layer1_out[565] <= 1'b0;
     layer1_out[566] <= layer0_out[87];
     layer1_out[567] <= layer0_out[342];
     layer1_out[568] <= ~layer0_out[730];
     layer1_out[569] <= layer0_out[51] & layer0_out[52];
     layer1_out[570] <= ~layer0_out[647];
     layer1_out[571] <= 1'b1;
     layer1_out[572] <= layer0_out[427] & layer0_out[428];
     layer1_out[573] <= ~layer0_out[132] | layer0_out[131];
     layer1_out[574] <= ~layer0_out[792];
     layer1_out[575] <= layer0_out[447];
     layer1_out[576] <= ~(layer0_out[251] & layer0_out[252]);
     layer1_out[577] <= 1'b1;
     layer1_out[578] <= ~layer0_out[277];
     layer1_out[579] <= layer0_out[141];
     layer1_out[580] <= layer0_out[771];
     layer1_out[581] <= 1'b1;
     layer1_out[582] <= layer0_out[796] | layer0_out[797];
     layer1_out[583] <= layer0_out[583] & ~layer0_out[584];
     layer1_out[584] <= layer0_out[653] & ~layer0_out[652];
     layer1_out[585] <= ~layer0_out[677];
     layer1_out[586] <= 1'b0;
     layer1_out[587] <= layer0_out[249];
     layer1_out[588] <= ~layer0_out[92];
     layer1_out[589] <= layer0_out[505] & ~layer0_out[504];
     layer1_out[590] <= ~layer0_out[474] | layer0_out[473];
     layer1_out[591] <= layer0_out[689];
     layer1_out[592] <= 1'b0;
     layer1_out[593] <= layer0_out[123] & layer0_out[124];
     layer1_out[594] <= layer0_out[442];
     layer1_out[595] <= 1'b0;
     layer1_out[596] <= 1'b1;
     layer1_out[597] <= ~(layer0_out[139] | layer0_out[140]);
     layer1_out[598] <= ~layer0_out[220];
     layer1_out[599] <= 1'b0;
     layer1_out[600] <= layer0_out[57];
     layer1_out[601] <= layer0_out[197];
     layer1_out[602] <= 1'b1;
     layer1_out[603] <= ~layer0_out[195];
     layer1_out[604] <= layer0_out[795] & ~layer0_out[796];
     layer1_out[605] <= ~layer0_out[588];
     layer1_out[606] <= ~(layer0_out[333] & layer0_out[334]);
     layer1_out[607] <= 1'b1;
     layer1_out[608] <= ~(layer0_out[451] & layer0_out[452]);
     layer1_out[609] <= 1'b0;
     layer1_out[610] <= 1'b0;
     layer1_out[611] <= ~layer0_out[268] | layer0_out[267];
     layer1_out[612] <= layer0_out[10] & ~layer0_out[11];
     layer1_out[613] <= ~layer0_out[444] | layer0_out[445];
     layer1_out[614] <= ~layer0_out[735] | layer0_out[734];
     layer1_out[615] <= ~layer0_out[257] | layer0_out[258];
     layer1_out[616] <= layer0_out[182];
     layer1_out[617] <= ~layer0_out[299];
     layer1_out[618] <= layer0_out[236];
     layer1_out[619] <= layer0_out[587];
     layer1_out[620] <= ~(layer0_out[187] | layer0_out[188]);
     layer1_out[621] <= 1'b0;
     layer1_out[622] <= layer0_out[516] & ~layer0_out[517];
     layer1_out[623] <= 1'b0;
     layer1_out[624] <= 1'b1;
     layer1_out[625] <= layer0_out[765];
     layer1_out[626] <= ~layer0_out[544];
     layer1_out[627] <= layer0_out[727] & ~layer0_out[726];
     layer1_out[628] <= ~layer0_out[530] | layer0_out[531];
     layer1_out[629] <= layer0_out[369] & layer0_out[370];
     layer1_out[630] <= ~layer0_out[708];
     layer1_out[631] <= layer0_out[145];
     layer1_out[632] <= 1'b1;
     layer1_out[633] <= 1'b1;
     layer1_out[634] <= ~layer0_out[609] | layer0_out[608];
     layer1_out[635] <= ~layer0_out[388] | layer0_out[387];
     layer1_out[636] <= layer0_out[299];
     layer1_out[637] <= ~layer0_out[30] | layer0_out[29];
     layer1_out[638] <= ~layer0_out[237] | layer0_out[238];
     layer1_out[639] <= ~layer0_out[177];
     layer1_out[640] <= layer0_out[313];
     layer1_out[641] <= ~layer0_out[15] | layer0_out[14];
     layer1_out[642] <= 1'b0;
     layer1_out[643] <= ~layer0_out[339];
     layer1_out[644] <= ~(layer0_out[549] | layer0_out[550]);
     layer1_out[645] <= ~(layer0_out[364] & layer0_out[365]);
     layer1_out[646] <= ~layer0_out[582] | layer0_out[583];
     layer1_out[647] <= ~(layer0_out[552] & layer0_out[553]);
     layer1_out[648] <= layer0_out[594] & layer0_out[595];
     layer1_out[649] <= layer0_out[312];
     layer1_out[650] <= ~layer0_out[301];
     layer1_out[651] <= layer0_out[559] & ~layer0_out[558];
     layer1_out[652] <= layer0_out[109] & ~layer0_out[108];
     layer1_out[653] <= layer0_out[217] & layer0_out[218];
     layer1_out[654] <= layer0_out[755] & ~layer0_out[756];
     layer1_out[655] <= layer0_out[752];
     layer1_out[656] <= layer0_out[619];
     layer1_out[657] <= ~layer0_out[648] | layer0_out[647];
     layer1_out[658] <= ~layer0_out[306] | layer0_out[307];
     layer1_out[659] <= ~layer0_out[290];
     layer1_out[660] <= 1'b0;
     layer1_out[661] <= 1'b0;
     layer1_out[662] <= ~layer0_out[269];
     layer1_out[663] <= 1'b1;
     layer1_out[664] <= 1'b0;
     layer1_out[665] <= 1'b0;
     layer1_out[666] <= ~layer0_out[556];
     layer1_out[667] <= ~layer0_out[705] | layer0_out[704];
     layer1_out[668] <= ~layer0_out[104];
     layer1_out[669] <= layer0_out[605];
     layer1_out[670] <= 1'b1;
     layer1_out[671] <= ~(layer0_out[621] & layer0_out[622]);
     layer1_out[672] <= ~layer0_out[290] | layer0_out[289];
     layer1_out[673] <= ~layer0_out[694];
     layer1_out[674] <= 1'b1;
     layer1_out[675] <= 1'b0;
     layer1_out[676] <= ~layer0_out[98];
     layer1_out[677] <= ~(layer0_out[138] | layer0_out[139]);
     layer1_out[678] <= layer0_out[412];
     layer1_out[679] <= ~layer0_out[85] | layer0_out[86];
     layer1_out[680] <= ~layer0_out[433] | layer0_out[434];
     layer1_out[681] <= layer0_out[774] | layer0_out[775];
     layer1_out[682] <= layer0_out[375];
     layer1_out[683] <= ~layer0_out[430];
     layer1_out[684] <= 1'b0;
     layer1_out[685] <= ~layer0_out[274] | layer0_out[273];
     layer1_out[686] <= ~layer0_out[88] | layer0_out[89];
     layer1_out[687] <= layer0_out[634] & layer0_out[635];
     layer1_out[688] <= ~(layer0_out[611] & layer0_out[612]);
     layer1_out[689] <= ~layer0_out[687];
     layer1_out[690] <= ~layer0_out[410];
     layer1_out[691] <= layer0_out[132] | layer0_out[133];
     layer1_out[692] <= layer0_out[33] & ~layer0_out[32];
     layer1_out[693] <= ~layer0_out[592];
     layer1_out[694] <= 1'b0;
     layer1_out[695] <= 1'b0;
     layer1_out[696] <= 1'b0;
     layer1_out[697] <= ~layer0_out[593];
     layer1_out[698] <= ~layer0_out[96] | layer0_out[97];
     layer1_out[699] <= layer0_out[773];
     layer1_out[700] <= layer0_out[536];
     layer1_out[701] <= layer0_out[742];
     layer1_out[702] <= 1'b1;
     layer1_out[703] <= layer0_out[685] & layer0_out[686];
     layer1_out[704] <= 1'b0;
     layer1_out[705] <= ~layer0_out[345] | layer0_out[344];
     layer1_out[706] <= 1'b1;
     layer1_out[707] <= 1'b0;
     layer1_out[708] <= ~layer0_out[698];
     layer1_out[709] <= layer0_out[586] & ~layer0_out[585];
     layer1_out[710] <= layer0_out[732] & ~layer0_out[731];
     layer1_out[711] <= layer0_out[367] & ~layer0_out[368];
     layer1_out[712] <= layer0_out[666] & ~layer0_out[667];
     layer1_out[713] <= 1'b1;
     layer1_out[714] <= layer0_out[512];
     layer1_out[715] <= ~layer0_out[631] | layer0_out[630];
     layer1_out[716] <= layer0_out[404];
     layer1_out[717] <= ~layer0_out[204];
     layer1_out[718] <= ~(layer0_out[669] & layer0_out[670]);
     layer1_out[719] <= layer0_out[127] & layer0_out[128];
     layer1_out[720] <= ~layer0_out[301];
     layer1_out[721] <= layer0_out[384];
     layer1_out[722] <= ~layer0_out[361] | layer0_out[360];
     layer1_out[723] <= 1'b1;
     layer1_out[724] <= layer0_out[567] & layer0_out[568];
     layer1_out[725] <= ~(layer0_out[539] ^ layer0_out[540]);
     layer1_out[726] <= ~(layer0_out[577] & layer0_out[578]);
     layer1_out[727] <= ~layer0_out[241] | layer0_out[242];
     layer1_out[728] <= ~layer0_out[378] | layer0_out[377];
     layer1_out[729] <= ~layer0_out[464] | layer0_out[463];
     layer1_out[730] <= ~layer0_out[227] | layer0_out[228];
     layer1_out[731] <= layer0_out[406] | layer0_out[407];
     layer1_out[732] <= layer0_out[530] & ~layer0_out[529];
     layer1_out[733] <= ~(layer0_out[613] & layer0_out[614]);
     layer1_out[734] <= layer0_out[351];
     layer1_out[735] <= ~layer0_out[307] | layer0_out[308];
     layer1_out[736] <= 1'b1;
     layer1_out[737] <= 1'b1;
     layer1_out[738] <= 1'b0;
     layer1_out[739] <= ~(layer0_out[238] | layer0_out[239]);
     layer1_out[740] <= layer0_out[113] & ~layer0_out[112];
     layer1_out[741] <= 1'b1;
     layer1_out[742] <= ~(layer0_out[146] & layer0_out[147]);
     layer1_out[743] <= layer0_out[510];
     layer1_out[744] <= layer0_out[745];
     layer1_out[745] <= ~(layer0_out[486] | layer0_out[487]);
     layer1_out[746] <= layer0_out[363];
     layer1_out[747] <= layer0_out[631] & layer0_out[632];
     layer1_out[748] <= ~layer0_out[43];
     layer1_out[749] <= ~(layer0_out[38] & layer0_out[39]);
     layer1_out[750] <= layer0_out[392];
     layer1_out[751] <= layer0_out[740];
     layer1_out[752] <= layer0_out[379];
     layer1_out[753] <= ~(layer0_out[229] | layer0_out[230]);
     layer1_out[754] <= layer0_out[318] | layer0_out[319];
     layer1_out[755] <= layer0_out[670] | layer0_out[671];
     layer1_out[756] <= ~layer0_out[532];
     layer1_out[757] <= layer0_out[752];
     layer1_out[758] <= ~layer0_out[725];
     layer1_out[759] <= layer0_out[437] | layer0_out[438];
     layer1_out[760] <= 1'b0;
     layer1_out[761] <= 1'b0;
     layer1_out[762] <= layer0_out[254] & ~layer0_out[255];
     layer1_out[763] <= ~layer0_out[315];
     layer1_out[764] <= ~layer0_out[294];
     layer1_out[765] <= ~layer0_out[460] | layer0_out[459];
     layer1_out[766] <= ~layer0_out[520];
     layer1_out[767] <= ~(layer0_out[462] & layer0_out[463]);
     layer1_out[768] <= layer0_out[347];
     layer1_out[769] <= 1'b0;
     layer1_out[770] <= 1'b0;
     layer1_out[771] <= ~(layer0_out[167] & layer0_out[168]);
     layer1_out[772] <= 1'b1;
     layer1_out[773] <= 1'b1;
     layer1_out[774] <= layer0_out[783];
     layer1_out[775] <= 1'b0;
     layer1_out[776] <= layer0_out[304] & layer0_out[305];
     layer1_out[777] <= layer0_out[265];
     layer1_out[778] <= ~layer0_out[2];
     layer1_out[779] <= layer0_out[493];
     layer1_out[780] <= ~layer0_out[543] | layer0_out[542];
     layer1_out[781] <= layer0_out[147];
     layer1_out[782] <= 1'b1;
     layer1_out[783] <= 1'b0;
     layer1_out[784] <= 1'b0;
     layer1_out[785] <= 1'b1;
     layer1_out[786] <= ~(layer0_out[411] & layer0_out[412]);
     layer1_out[787] <= layer0_out[64];
     layer1_out[788] <= ~layer0_out[55];
     layer1_out[789] <= layer0_out[554];
     layer1_out[790] <= ~layer0_out[372];
     layer1_out[791] <= layer0_out[736] | layer0_out[737];
     layer1_out[792] <= ~(layer0_out[99] | layer0_out[100]);
     layer1_out[793] <= ~layer0_out[90];
     layer1_out[794] <= ~layer0_out[372] | layer0_out[371];
     layer1_out[795] <= ~layer0_out[468] | layer0_out[467];
     layer1_out[796] <= layer0_out[224] | layer0_out[225];
     layer1_out[797] <= ~layer0_out[126];
     layer1_out[798] <= layer0_out[598];
     layer1_out[799] <= layer0_out[691] & ~layer0_out[690];
     layer2_out[0] <= ~layer1_out[663] | layer1_out[662];
     layer2_out[1] <= layer1_out[93] & ~layer1_out[92];
     layer2_out[2] <= ~layer1_out[629] | layer1_out[628];
     layer2_out[3] <= layer1_out[186];
     layer2_out[4] <= ~layer1_out[378];
     layer2_out[5] <= 1'b0;
     layer2_out[6] <= ~layer1_out[501];
     layer2_out[7] <= ~layer1_out[494];
     layer2_out[8] <= ~layer1_out[613];
     layer2_out[9] <= layer1_out[408] & ~layer1_out[407];
     layer2_out[10] <= layer1_out[186];
     layer2_out[11] <= layer1_out[359] & layer1_out[360];
     layer2_out[12] <= 1'b1;
     layer2_out[13] <= ~layer1_out[219] | layer1_out[220];
     layer2_out[14] <= layer1_out[671] & ~layer1_out[670];
     layer2_out[15] <= ~layer1_out[224];
     layer2_out[16] <= layer1_out[8] & ~layer1_out[7];
     layer2_out[17] <= layer1_out[199];
     layer2_out[18] <= layer1_out[33] & layer1_out[34];
     layer2_out[19] <= layer1_out[165] & layer1_out[166];
     layer2_out[20] <= 1'b1;
     layer2_out[21] <= layer1_out[617] | layer1_out[618];
     layer2_out[22] <= layer1_out[195] | layer1_out[196];
     layer2_out[23] <= layer1_out[758] & ~layer1_out[757];
     layer2_out[24] <= layer1_out[792];
     layer2_out[25] <= layer1_out[532] | layer1_out[533];
     layer2_out[26] <= ~layer1_out[733];
     layer2_out[27] <= layer1_out[353] & ~layer1_out[354];
     layer2_out[28] <= 1'b1;
     layer2_out[29] <= layer1_out[489];
     layer2_out[30] <= layer1_out[707] & ~layer1_out[708];
     layer2_out[31] <= ~layer1_out[173];
     layer2_out[32] <= layer1_out[690];
     layer2_out[33] <= layer1_out[318];
     layer2_out[34] <= 1'b0;
     layer2_out[35] <= ~layer1_out[328];
     layer2_out[36] <= layer1_out[73];
     layer2_out[37] <= 1'b1;
     layer2_out[38] <= ~layer1_out[216];
     layer2_out[39] <= ~layer1_out[196];
     layer2_out[40] <= layer1_out[753];
     layer2_out[41] <= ~layer1_out[799];
     layer2_out[42] <= layer1_out[546] & ~layer1_out[545];
     layer2_out[43] <= layer1_out[40] & layer1_out[41];
     layer2_out[44] <= layer1_out[449] & layer1_out[450];
     layer2_out[45] <= layer1_out[439] & ~layer1_out[440];
     layer2_out[46] <= 1'b0;
     layer2_out[47] <= layer1_out[534] & layer1_out[535];
     layer2_out[48] <= ~layer1_out[741];
     layer2_out[49] <= layer1_out[430] & ~layer1_out[429];
     layer2_out[50] <= ~(layer1_out[151] & layer1_out[152]);
     layer2_out[51] <= layer1_out[401];
     layer2_out[52] <= layer1_out[518] & layer1_out[519];
     layer2_out[53] <= layer1_out[534];
     layer2_out[54] <= ~layer1_out[202];
     layer2_out[55] <= layer1_out[697];
     layer2_out[56] <= layer1_out[549] & layer1_out[550];
     layer2_out[57] <= ~layer1_out[311] | layer1_out[310];
     layer2_out[58] <= layer1_out[155];
     layer2_out[59] <= layer1_out[529] & ~layer1_out[530];
     layer2_out[60] <= ~layer1_out[789] | layer1_out[788];
     layer2_out[61] <= ~(layer1_out[681] & layer1_out[682]);
     layer2_out[62] <= layer1_out[632] & layer1_out[633];
     layer2_out[63] <= 1'b0;
     layer2_out[64] <= ~layer1_out[175];
     layer2_out[65] <= layer1_out[298] & ~layer1_out[297];
     layer2_out[66] <= ~(layer1_out[648] | layer1_out[649]);
     layer2_out[67] <= ~(layer1_out[777] | layer1_out[778]);
     layer2_out[68] <= layer1_out[120] & layer1_out[121];
     layer2_out[69] <= layer1_out[206] & ~layer1_out[205];
     layer2_out[70] <= ~layer1_out[148];
     layer2_out[71] <= ~layer1_out[500] | layer1_out[499];
     layer2_out[72] <= layer1_out[333] & ~layer1_out[332];
     layer2_out[73] <= layer1_out[1] | layer1_out[2];
     layer2_out[74] <= ~layer1_out[387];
     layer2_out[75] <= ~layer1_out[512];
     layer2_out[76] <= layer1_out[716];
     layer2_out[77] <= layer1_out[414] & ~layer1_out[415];
     layer2_out[78] <= layer1_out[616];
     layer2_out[79] <= layer1_out[123] & ~layer1_out[124];
     layer2_out[80] <= ~layer1_out[598];
     layer2_out[81] <= layer1_out[410];
     layer2_out[82] <= layer1_out[620] & ~layer1_out[619];
     layer2_out[83] <= layer1_out[517];
     layer2_out[84] <= layer1_out[323];
     layer2_out[85] <= ~layer1_out[692];
     layer2_out[86] <= ~layer1_out[270];
     layer2_out[87] <= layer1_out[307] | layer1_out[308];
     layer2_out[88] <= ~layer1_out[285];
     layer2_out[89] <= 1'b0;
     layer2_out[90] <= layer1_out[559] & layer1_out[560];
     layer2_out[91] <= layer1_out[751];
     layer2_out[92] <= layer1_out[261] & layer1_out[262];
     layer2_out[93] <= 1'b0;
     layer2_out[94] <= layer1_out[392] & ~layer1_out[393];
     layer2_out[95] <= layer1_out[791];
     layer2_out[96] <= layer1_out[54] | layer1_out[55];
     layer2_out[97] <= ~layer1_out[80] | layer1_out[81];
     layer2_out[98] <= layer1_out[625];
     layer2_out[99] <= layer1_out[462];
     layer2_out[100] <= layer1_out[421];
     layer2_out[101] <= ~layer1_out[643];
     layer2_out[102] <= ~layer1_out[127];
     layer2_out[103] <= layer1_out[63];
     layer2_out[104] <= layer1_out[581] | layer1_out[582];
     layer2_out[105] <= layer1_out[349];
     layer2_out[106] <= layer1_out[723];
     layer2_out[107] <= 1'b0;
     layer2_out[108] <= layer1_out[37] & ~layer1_out[38];
     layer2_out[109] <= 1'b1;
     layer2_out[110] <= layer1_out[26];
     layer2_out[111] <= layer1_out[319];
     layer2_out[112] <= ~layer1_out[159] | layer1_out[158];
     layer2_out[113] <= ~layer1_out[188] | layer1_out[187];
     layer2_out[114] <= layer1_out[467];
     layer2_out[115] <= ~layer1_out[159];
     layer2_out[116] <= layer1_out[87] & ~layer1_out[86];
     layer2_out[117] <= layer1_out[363] & ~layer1_out[362];
     layer2_out[118] <= layer1_out[106];
     layer2_out[119] <= layer1_out[422] & ~layer1_out[423];
     layer2_out[120] <= ~(layer1_out[345] & layer1_out[346]);
     layer2_out[121] <= layer1_out[646];
     layer2_out[122] <= ~(layer1_out[411] & layer1_out[412]);
     layer2_out[123] <= layer1_out[267] | layer1_out[268];
     layer2_out[124] <= ~layer1_out[70];
     layer2_out[125] <= layer1_out[408];
     layer2_out[126] <= layer1_out[388];
     layer2_out[127] <= layer1_out[695];
     layer2_out[128] <= ~layer1_out[389] | layer1_out[390];
     layer2_out[129] <= layer1_out[436] | layer1_out[437];
     layer2_out[130] <= ~(layer1_out[303] | layer1_out[304]);
     layer2_out[131] <= layer1_out[561] & ~layer1_out[562];
     layer2_out[132] <= layer1_out[413];
     layer2_out[133] <= ~layer1_out[256] | layer1_out[257];
     layer2_out[134] <= layer1_out[90];
     layer2_out[135] <= 1'b0;
     layer2_out[136] <= ~(layer1_out[18] | layer1_out[19]);
     layer2_out[137] <= 1'b1;
     layer2_out[138] <= layer1_out[361];
     layer2_out[139] <= layer1_out[588] & layer1_out[589];
     layer2_out[140] <= layer1_out[660];
     layer2_out[141] <= layer1_out[3];
     layer2_out[142] <= ~layer1_out[554] | layer1_out[553];
     layer2_out[143] <= layer1_out[3] & layer1_out[4];
     layer2_out[144] <= ~layer1_out[685] | layer1_out[686];
     layer2_out[145] <= layer1_out[639];
     layer2_out[146] <= ~layer1_out[4];
     layer2_out[147] <= ~layer1_out[249] | layer1_out[248];
     layer2_out[148] <= layer1_out[255] | layer1_out[256];
     layer2_out[149] <= ~(layer1_out[455] & layer1_out[456]);
     layer2_out[150] <= layer1_out[236] | layer1_out[237];
     layer2_out[151] <= layer1_out[88] & layer1_out[89];
     layer2_out[152] <= layer1_out[360] & layer1_out[361];
     layer2_out[153] <= ~layer1_out[289];
     layer2_out[154] <= layer1_out[688] & layer1_out[689];
     layer2_out[155] <= layer1_out[668];
     layer2_out[156] <= ~layer1_out[571];
     layer2_out[157] <= layer1_out[57] & ~layer1_out[56];
     layer2_out[158] <= layer1_out[467] & ~layer1_out[466];
     layer2_out[159] <= ~layer1_out[679];
     layer2_out[160] <= 1'b1;
     layer2_out[161] <= ~layer1_out[8];
     layer2_out[162] <= 1'b1;
     layer2_out[163] <= ~(layer1_out[721] & layer1_out[722]);
     layer2_out[164] <= 1'b1;
     layer2_out[165] <= ~layer1_out[521] | layer1_out[522];
     layer2_out[166] <= layer1_out[508] & layer1_out[509];
     layer2_out[167] <= ~layer1_out[110];
     layer2_out[168] <= layer1_out[650];
     layer2_out[169] <= layer1_out[104];
     layer2_out[170] <= ~layer1_out[195] | layer1_out[194];
     layer2_out[171] <= layer1_out[507] ^ layer1_out[508];
     layer2_out[172] <= layer1_out[495] | layer1_out[496];
     layer2_out[173] <= 1'b1;
     layer2_out[174] <= ~layer1_out[572] | layer1_out[573];
     layer2_out[175] <= layer1_out[66];
     layer2_out[176] <= ~layer1_out[730];
     layer2_out[177] <= ~(layer1_out[673] | layer1_out[674]);
     layer2_out[178] <= layer1_out[63] & layer1_out[64];
     layer2_out[179] <= layer1_out[755];
     layer2_out[180] <= 1'b0;
     layer2_out[181] <= layer1_out[219] & ~layer1_out[218];
     layer2_out[182] <= ~(layer1_out[376] ^ layer1_out[377]);
     layer2_out[183] <= layer1_out[393];
     layer2_out[184] <= layer1_out[305];
     layer2_out[185] <= ~layer1_out[464];
     layer2_out[186] <= ~layer1_out[306];
     layer2_out[187] <= ~layer1_out[89] | layer1_out[90];
     layer2_out[188] <= layer1_out[580] & layer1_out[581];
     layer2_out[189] <= ~layer1_out[365];
     layer2_out[190] <= layer1_out[333];
     layer2_out[191] <= layer1_out[252] ^ layer1_out[253];
     layer2_out[192] <= ~layer1_out[595] | layer1_out[594];
     layer2_out[193] <= layer1_out[397];
     layer2_out[194] <= ~layer1_out[488] | layer1_out[489];
     layer2_out[195] <= layer1_out[358] & ~layer1_out[357];
     layer2_out[196] <= ~layer1_out[69];
     layer2_out[197] <= 1'b0;
     layer2_out[198] <= ~layer1_out[474] | layer1_out[475];
     layer2_out[199] <= layer1_out[450] & ~layer1_out[451];
     layer2_out[200] <= ~(layer1_out[433] | layer1_out[434]);
     layer2_out[201] <= layer1_out[156] & ~layer1_out[157];
     layer2_out[202] <= layer1_out[276];
     layer2_out[203] <= layer1_out[794] & layer1_out[795];
     layer2_out[204] <= 1'b1;
     layer2_out[205] <= ~(layer1_out[21] | layer1_out[22]);
     layer2_out[206] <= layer1_out[728];
     layer2_out[207] <= ~layer1_out[319];
     layer2_out[208] <= ~layer1_out[106];
     layer2_out[209] <= ~(layer1_out[346] & layer1_out[347]);
     layer2_out[210] <= ~layer1_out[540];
     layer2_out[211] <= ~layer1_out[303] | layer1_out[302];
     layer2_out[212] <= ~layer1_out[781];
     layer2_out[213] <= layer1_out[184];
     layer2_out[214] <= 1'b0;
     layer2_out[215] <= layer1_out[325] & layer1_out[326];
     layer2_out[216] <= ~(layer1_out[391] ^ layer1_out[392]);
     layer2_out[217] <= layer1_out[181] | layer1_out[182];
     layer2_out[218] <= layer1_out[629];
     layer2_out[219] <= ~layer1_out[726] | layer1_out[727];
     layer2_out[220] <= ~layer1_out[21] | layer1_out[20];
     layer2_out[221] <= layer1_out[797];
     layer2_out[222] <= layer1_out[275] | layer1_out[276];
     layer2_out[223] <= ~(layer1_out[459] | layer1_out[460]);
     layer2_out[224] <= ~layer1_out[309];
     layer2_out[225] <= ~(layer1_out[701] | layer1_out[702]);
     layer2_out[226] <= ~layer1_out[515];
     layer2_out[227] <= layer1_out[53];
     layer2_out[228] <= ~layer1_out[10];
     layer2_out[229] <= 1'b1;
     layer2_out[230] <= layer1_out[35];
     layer2_out[231] <= layer1_out[444] & layer1_out[445];
     layer2_out[232] <= layer1_out[511] & ~layer1_out[510];
     layer2_out[233] <= layer1_out[50] & ~layer1_out[51];
     layer2_out[234] <= layer1_out[479];
     layer2_out[235] <= layer1_out[717];
     layer2_out[236] <= layer1_out[300];
     layer2_out[237] <= ~layer1_out[175];
     layer2_out[238] <= ~layer1_out[640];
     layer2_out[239] <= ~layer1_out[226];
     layer2_out[240] <= layer1_out[483] & layer1_out[484];
     layer2_out[241] <= layer1_out[241] & ~layer1_out[240];
     layer2_out[242] <= layer1_out[5];
     layer2_out[243] <= layer1_out[296];
     layer2_out[244] <= ~(layer1_out[273] & layer1_out[274]);
     layer2_out[245] <= 1'b0;
     layer2_out[246] <= layer1_out[455] & ~layer1_out[454];
     layer2_out[247] <= ~layer1_out[752];
     layer2_out[248] <= ~layer1_out[796] | layer1_out[795];
     layer2_out[249] <= layer1_out[121] & layer1_out[122];
     layer2_out[250] <= layer1_out[544] & ~layer1_out[543];
     layer2_out[251] <= layer1_out[564] | layer1_out[565];
     layer2_out[252] <= layer1_out[62] & ~layer1_out[61];
     layer2_out[253] <= layer1_out[316] & ~layer1_out[315];
     layer2_out[254] <= layer1_out[476];
     layer2_out[255] <= 1'b0;
     layer2_out[256] <= layer1_out[745] & ~layer1_out[744];
     layer2_out[257] <= layer1_out[28] & ~layer1_out[29];
     layer2_out[258] <= ~layer1_out[731];
     layer2_out[259] <= ~layer1_out[316] | layer1_out[317];
     layer2_out[260] <= 1'b0;
     layer2_out[261] <= ~layer1_out[536];
     layer2_out[262] <= layer1_out[59] | layer1_out[60];
     layer2_out[263] <= layer1_out[296];
     layer2_out[264] <= layer1_out[458] & layer1_out[459];
     layer2_out[265] <= ~layer1_out[45];
     layer2_out[266] <= layer1_out[779] & ~layer1_out[780];
     layer2_out[267] <= layer1_out[230] & layer1_out[231];
     layer2_out[268] <= ~layer1_out[740];
     layer2_out[269] <= layer1_out[77] | layer1_out[78];
     layer2_out[270] <= ~layer1_out[707];
     layer2_out[271] <= ~(layer1_out[591] | layer1_out[592]);
     layer2_out[272] <= ~layer1_out[52];
     layer2_out[273] <= ~(layer1_out[447] & layer1_out[448]);
     layer2_out[274] <= ~layer1_out[773];
     layer2_out[275] <= ~(layer1_out[456] | layer1_out[457]);
     layer2_out[276] <= ~(layer1_out[75] & layer1_out[76]);
     layer2_out[277] <= ~(layer1_out[271] | layer1_out[272]);
     layer2_out[278] <= layer1_out[525] & layer1_out[526];
     layer2_out[279] <= ~(layer1_out[385] | layer1_out[386]);
     layer2_out[280] <= ~layer1_out[644];
     layer2_out[281] <= ~layer1_out[453] | layer1_out[454];
     layer2_out[282] <= layer1_out[441] & ~layer1_out[440];
     layer2_out[283] <= layer1_out[690] ^ layer1_out[691];
     layer2_out[284] <= layer1_out[473] & layer1_out[474];
     layer2_out[285] <= ~layer1_out[611];
     layer2_out[286] <= layer1_out[426] & ~layer1_out[425];
     layer2_out[287] <= layer1_out[567] & layer1_out[568];
     layer2_out[288] <= layer1_out[118] & layer1_out[119];
     layer2_out[289] <= 1'b1;
     layer2_out[290] <= layer1_out[438];
     layer2_out[291] <= layer1_out[532];
     layer2_out[292] <= layer1_out[284];
     layer2_out[293] <= ~layer1_out[255] | layer1_out[254];
     layer2_out[294] <= 1'b1;
     layer2_out[295] <= ~layer1_out[569];
     layer2_out[296] <= ~layer1_out[213] | layer1_out[212];
     layer2_out[297] <= 1'b1;
     layer2_out[298] <= ~(layer1_out[435] & layer1_out[436]);
     layer2_out[299] <= ~layer1_out[527] | layer1_out[528];
     layer2_out[300] <= ~layer1_out[702];
     layer2_out[301] <= ~layer1_out[403];
     layer2_out[302] <= layer1_out[531] & ~layer1_out[530];
     layer2_out[303] <= ~(layer1_out[550] & layer1_out[551]);
     layer2_out[304] <= layer1_out[133];
     layer2_out[305] <= ~layer1_out[43];
     layer2_out[306] <= layer1_out[374] & ~layer1_out[373];
     layer2_out[307] <= ~layer1_out[478];
     layer2_out[308] <= layer1_out[161] & ~layer1_out[162];
     layer2_out[309] <= ~(layer1_out[584] & layer1_out[585]);
     layer2_out[310] <= ~layer1_out[385];
     layer2_out[311] <= ~(layer1_out[771] & layer1_out[772]);
     layer2_out[312] <= layer1_out[774] | layer1_out[775];
     layer2_out[313] <= layer1_out[188];
     layer2_out[314] <= ~layer1_out[85] | layer1_out[86];
     layer2_out[315] <= 1'b1;
     layer2_out[316] <= ~(layer1_out[700] ^ layer1_out[701]);
     layer2_out[317] <= ~layer1_out[78];
     layer2_out[318] <= ~layer1_out[715] | layer1_out[716];
     layer2_out[319] <= layer1_out[300] ^ layer1_out[301];
     layer2_out[320] <= ~(layer1_out[180] & layer1_out[181]);
     layer2_out[321] <= ~layer1_out[163];
     layer2_out[322] <= 1'b1;
     layer2_out[323] <= layer1_out[586] | layer1_out[587];
     layer2_out[324] <= layer1_out[84];
     layer2_out[325] <= layer1_out[129] ^ layer1_out[130];
     layer2_out[326] <= ~(layer1_out[516] | layer1_out[517]);
     layer2_out[327] <= layer1_out[235];
     layer2_out[328] <= ~layer1_out[492] | layer1_out[491];
     layer2_out[329] <= layer1_out[565] & ~layer1_out[566];
     layer2_out[330] <= ~layer1_out[263];
     layer2_out[331] <= 1'b0;
     layer2_out[332] <= layer1_out[254];
     layer2_out[333] <= ~(layer1_out[352] | layer1_out[353]);
     layer2_out[334] <= ~layer1_out[497] | layer1_out[496];
     layer2_out[335] <= layer1_out[44] & ~layer1_out[45];
     layer2_out[336] <= ~layer1_out[666] | layer1_out[667];
     layer2_out[337] <= ~layer1_out[523] | layer1_out[524];
     layer2_out[338] <= layer1_out[658];
     layer2_out[339] <= layer1_out[555];
     layer2_out[340] <= ~(layer1_out[734] & layer1_out[735]);
     layer2_out[341] <= ~layer1_out[564];
     layer2_out[342] <= ~(layer1_out[645] | layer1_out[646]);
     layer2_out[343] <= layer1_out[179];
     layer2_out[344] <= ~layer1_out[443];
     layer2_out[345] <= layer1_out[222] | layer1_out[223];
     layer2_out[346] <= layer1_out[469] | layer1_out[470];
     layer2_out[347] <= ~layer1_out[430] | layer1_out[431];
     layer2_out[348] <= ~layer1_out[615] | layer1_out[616];
     layer2_out[349] <= ~layer1_out[438] | layer1_out[439];
     layer2_out[350] <= layer1_out[150] ^ layer1_out[151];
     layer2_out[351] <= 1'b0;
     layer2_out[352] <= ~layer1_out[427];
     layer2_out[353] <= layer1_out[481] & layer1_out[482];
     layer2_out[354] <= layer1_out[604] | layer1_out[605];
     layer2_out[355] <= ~layer1_out[312];
     layer2_out[356] <= ~layer1_out[674];
     layer2_out[357] <= ~layer1_out[55] | layer1_out[56];
     layer2_out[358] <= ~(layer1_out[215] | layer1_out[216]);
     layer2_out[359] <= 1'b0;
     layer2_out[360] <= layer1_out[773];
     layer2_out[361] <= layer1_out[761];
     layer2_out[362] <= ~layer1_out[13];
     layer2_out[363] <= layer1_out[0] & layer1_out[2];
     layer2_out[364] <= ~layer1_out[88] | layer1_out[87];
     layer2_out[365] <= 1'b0;
     layer2_out[366] <= layer1_out[73] & ~layer1_out[72];
     layer2_out[367] <= ~layer1_out[279] | layer1_out[280];
     layer2_out[368] <= layer1_out[278];
     layer2_out[369] <= layer1_out[326] | layer1_out[327];
     layer2_out[370] <= layer1_out[283] | layer1_out[284];
     layer2_out[371] <= layer1_out[245] & layer1_out[246];
     layer2_out[372] <= ~layer1_out[720] | layer1_out[719];
     layer2_out[373] <= ~(layer1_out[144] | layer1_out[145]);
     layer2_out[374] <= ~layer1_out[743];
     layer2_out[375] <= ~layer1_out[790];
     layer2_out[376] <= ~layer1_out[135] | layer1_out[134];
     layer2_out[377] <= layer1_out[217];
     layer2_out[378] <= ~(layer1_out[631] | layer1_out[632]);
     layer2_out[379] <= ~layer1_out[260] | layer1_out[261];
     layer2_out[380] <= 1'b1;
     layer2_out[381] <= layer1_out[37];
     layer2_out[382] <= layer1_out[662] & ~layer1_out[661];
     layer2_out[383] <= ~layer1_out[519] | layer1_out[520];
     layer2_out[384] <= ~layer1_out[782] | layer1_out[783];
     layer2_out[385] <= ~(layer1_out[93] & layer1_out[94]);
     layer2_out[386] <= ~layer1_out[759];
     layer2_out[387] <= layer1_out[28];
     layer2_out[388] <= layer1_out[351] & ~layer1_out[350];
     layer2_out[389] <= ~(layer1_out[277] & layer1_out[278]);
     layer2_out[390] <= ~layer1_out[664] | layer1_out[665];
     layer2_out[391] <= ~layer1_out[473] | layer1_out[472];
     layer2_out[392] <= ~layer1_out[101];
     layer2_out[393] <= layer1_out[693];
     layer2_out[394] <= layer1_out[200] & ~layer1_out[201];
     layer2_out[395] <= ~layer1_out[709];
     layer2_out[396] <= layer1_out[291] & layer1_out[292];
     layer2_out[397] <= layer1_out[582] & ~layer1_out[583];
     layer2_out[398] <= layer1_out[67];
     layer2_out[399] <= layer1_out[153];
     layer2_out[400] <= ~layer1_out[566];
     layer2_out[401] <= layer1_out[630];
     layer2_out[402] <= ~layer1_out[15];
     layer2_out[403] <= layer1_out[57];
     layer2_out[404] <= ~layer1_out[482];
     layer2_out[405] <= 1'b0;
     layer2_out[406] <= layer1_out[797];
     layer2_out[407] <= ~layer1_out[258];
     layer2_out[408] <= layer1_out[770] & layer1_out[771];
     layer2_out[409] <= ~layer1_out[341];
     layer2_out[410] <= layer1_out[335];
     layer2_out[411] <= ~layer1_out[676] | layer1_out[675];
     layer2_out[412] <= layer1_out[756] | layer1_out[757];
     layer2_out[413] <= ~layer1_out[681];
     layer2_out[414] <= 1'b1;
     layer2_out[415] <= ~(layer1_out[418] & layer1_out[419]);
     layer2_out[416] <= ~(layer1_out[107] & layer1_out[108]);
     layer2_out[417] <= ~layer1_out[287];
     layer2_out[418] <= 1'b1;
     layer2_out[419] <= layer1_out[226] & layer1_out[227];
     layer2_out[420] <= ~(layer1_out[81] | layer1_out[82]);
     layer2_out[421] <= layer1_out[423];
     layer2_out[422] <= layer1_out[612];
     layer2_out[423] <= layer1_out[612];
     layer2_out[424] <= layer1_out[359];
     layer2_out[425] <= ~layer1_out[497];
     layer2_out[426] <= ~layer1_out[668] | layer1_out[667];
     layer2_out[427] <= ~layer1_out[619] | layer1_out[618];
     layer2_out[428] <= ~(layer1_out[595] | layer1_out[596]);
     layer2_out[429] <= ~layer1_out[99] | layer1_out[100];
     layer2_out[430] <= ~layer1_out[1] | layer1_out[0];
     layer2_out[431] <= layer1_out[113] | layer1_out[114];
     layer2_out[432] <= ~(layer1_out[286] | layer1_out[287]);
     layer2_out[433] <= layer1_out[752];
     layer2_out[434] <= layer1_out[607] & layer1_out[608];
     layer2_out[435] <= layer1_out[575] & ~layer1_out[576];
     layer2_out[436] <= ~(layer1_out[463] & layer1_out[464]);
     layer2_out[437] <= layer1_out[658] & ~layer1_out[657];
     layer2_out[438] <= ~layer1_out[243];
     layer2_out[439] <= layer1_out[549] & ~layer1_out[548];
     layer2_out[440] <= 1'b1;
     layer2_out[441] <= layer1_out[24] & layer1_out[25];
     layer2_out[442] <= ~(layer1_out[602] | layer1_out[603]);
     layer2_out[443] <= layer1_out[683];
     layer2_out[444] <= layer1_out[660] & ~layer1_out[659];
     layer2_out[445] <= ~layer1_out[244];
     layer2_out[446] <= ~(layer1_out[410] & layer1_out[411]);
     layer2_out[447] <= layer1_out[155];
     layer2_out[448] <= ~layer1_out[77];
     layer2_out[449] <= layer1_out[114] & ~layer1_out[115];
     layer2_out[450] <= layer1_out[204] | layer1_out[205];
     layer2_out[451] <= ~(layer1_out[546] | layer1_out[547]);
     layer2_out[452] <= layer1_out[46] & ~layer1_out[47];
     layer2_out[453] <= ~layer1_out[294];
     layer2_out[454] <= ~layer1_out[36];
     layer2_out[455] <= layer1_out[457] & ~layer1_out[458];
     layer2_out[456] <= layer1_out[693] & ~layer1_out[692];
     layer2_out[457] <= 1'b1;
     layer2_out[458] <= 1'b0;
     layer2_out[459] <= layer1_out[640];
     layer2_out[460] <= layer1_out[104];
     layer2_out[461] <= layer1_out[178];
     layer2_out[462] <= layer1_out[418];
     layer2_out[463] <= 1'b1;
     layer2_out[464] <= ~layer1_out[543];
     layer2_out[465] <= ~layer1_out[471];
     layer2_out[466] <= 1'b0;
     layer2_out[467] <= ~layer1_out[451];
     layer2_out[468] <= layer1_out[499] & ~layer1_out[498];
     layer2_out[469] <= ~layer1_out[65] | layer1_out[64];
     layer2_out[470] <= layer1_out[364] & ~layer1_out[363];
     layer2_out[471] <= layer1_out[29] & ~layer1_out[30];
     layer2_out[472] <= ~layer1_out[764] | layer1_out[765];
     layer2_out[473] <= ~layer1_out[340] | layer1_out[339];
     layer2_out[474] <= ~layer1_out[539];
     layer2_out[475] <= ~layer1_out[578];
     layer2_out[476] <= ~(layer1_out[570] & layer1_out[571]);
     layer2_out[477] <= ~layer1_out[420];
     layer2_out[478] <= layer1_out[330] ^ layer1_out[331];
     layer2_out[479] <= layer1_out[335] | layer1_out[336];
     layer2_out[480] <= ~layer1_out[524] | layer1_out[525];
     layer2_out[481] <= layer1_out[491];
     layer2_out[482] <= ~layer1_out[141];
     layer2_out[483] <= ~layer1_out[583];
     layer2_out[484] <= layer1_out[657];
     layer2_out[485] <= layer1_out[762];
     layer2_out[486] <= ~(layer1_out[22] & layer1_out[23]);
     layer2_out[487] <= layer1_out[488] & ~layer1_out[487];
     layer2_out[488] <= ~layer1_out[569];
     layer2_out[489] <= ~layer1_out[369];
     layer2_out[490] <= ~layer1_out[434] | layer1_out[435];
     layer2_out[491] <= 1'b1;
     layer2_out[492] <= 1'b0;
     layer2_out[493] <= layer1_out[465];
     layer2_out[494] <= ~layer1_out[112] | layer1_out[113];
     layer2_out[495] <= ~layer1_out[529] | layer1_out[528];
     layer2_out[496] <= layer1_out[72];
     layer2_out[497] <= 1'b1;
     layer2_out[498] <= layer1_out[190] & ~layer1_out[191];
     layer2_out[499] <= ~layer1_out[313] | layer1_out[314];
     layer2_out[500] <= layer1_out[677];
     layer2_out[501] <= layer1_out[194];
     layer2_out[502] <= layer1_out[349];
     layer2_out[503] <= layer1_out[623];
     layer2_out[504] <= layer1_out[537] | layer1_out[538];
     layer2_out[505] <= layer1_out[540] & layer1_out[541];
     layer2_out[506] <= layer1_out[235] | layer1_out[236];
     layer2_out[507] <= layer1_out[274];
     layer2_out[508] <= layer1_out[593] | layer1_out[594];
     layer2_out[509] <= ~(layer1_out[432] | layer1_out[433]);
     layer2_out[510] <= layer1_out[780];
     layer2_out[511] <= ~layer1_out[97] | layer1_out[96];
     layer2_out[512] <= layer1_out[625] & ~layer1_out[626];
     layer2_out[513] <= ~layer1_out[329];
     layer2_out[514] <= 1'b0;
     layer2_out[515] <= ~layer1_out[371] | layer1_out[370];
     layer2_out[516] <= layer1_out[221] & ~layer1_out[220];
     layer2_out[517] <= layer1_out[327];
     layer2_out[518] <= layer1_out[592];
     layer2_out[519] <= layer1_out[311];
     layer2_out[520] <= 1'b0;
     layer2_out[521] <= layer1_out[281] & ~layer1_out[280];
     layer2_out[522] <= ~(layer1_out[597] | layer1_out[598]);
     layer2_out[523] <= ~(layer1_out[754] & layer1_out[755]);
     layer2_out[524] <= 1'b1;
     layer2_out[525] <= ~layer1_out[24];
     layer2_out[526] <= layer1_out[400];
     layer2_out[527] <= layer1_out[147];
     layer2_out[528] <= 1'b0;
     layer2_out[529] <= ~(layer1_out[207] ^ layer1_out[208]);
     layer2_out[530] <= ~layer1_out[621] | layer1_out[620];
     layer2_out[531] <= layer1_out[506] & layer1_out[507];
     layer2_out[532] <= layer1_out[260];
     layer2_out[533] <= layer1_out[655];
     layer2_out[534] <= ~layer1_out[401];
     layer2_out[535] <= layer1_out[673];
     layer2_out[536] <= ~layer1_out[419] | layer1_out[420];
     layer2_out[537] <= ~layer1_out[41];
     layer2_out[538] <= layer1_out[634] & layer1_out[635];
     layer2_out[539] <= ~(layer1_out[562] | layer1_out[563]);
     layer2_out[540] <= ~layer1_out[19];
     layer2_out[541] <= ~layer1_out[14];
     layer2_out[542] <= ~(layer1_out[342] | layer1_out[343]);
     layer2_out[543] <= ~(layer1_out[127] | layer1_out[128]);
     layer2_out[544] <= ~layer1_out[368] | layer1_out[367];
     layer2_out[545] <= ~layer1_out[264] | layer1_out[265];
     layer2_out[546] <= ~layer1_out[669];
     layer2_out[547] <= layer1_out[230] & ~layer1_out[229];
     layer2_out[548] <= layer1_out[203];
     layer2_out[549] <= ~layer1_out[737];
     layer2_out[550] <= ~layer1_out[714] | layer1_out[715];
     layer2_out[551] <= ~layer1_out[185];
     layer2_out[552] <= ~layer1_out[137];
     layer2_out[553] <= layer1_out[413] | layer1_out[414];
     layer2_out[554] <= ~layer1_out[728];
     layer2_out[555] <= layer1_out[504];
     layer2_out[556] <= layer1_out[602];
     layer2_out[557] <= layer1_out[97] | layer1_out[98];
     layer2_out[558] <= ~layer1_out[137];
     layer2_out[559] <= layer1_out[263] & ~layer1_out[264];
     layer2_out[560] <= layer1_out[242] | layer1_out[243];
     layer2_out[561] <= layer1_out[43] & layer1_out[44];
     layer2_out[562] <= 1'b0;
     layer2_out[563] <= layer1_out[269] & ~layer1_out[268];
     layer2_out[564] <= ~(layer1_out[355] & layer1_out[356]);
     layer2_out[565] <= layer1_out[314] & layer1_out[315];
     layer2_out[566] <= layer1_out[341] & layer1_out[342];
     layer2_out[567] <= ~(layer1_out[266] | layer1_out[267]);
     layer2_out[568] <= layer1_out[677];
     layer2_out[569] <= layer1_out[232];
     layer2_out[570] <= ~layer1_out[448];
     layer2_out[571] <= ~layer1_out[555];
     layer2_out[572] <= ~layer1_out[171] | layer1_out[172];
     layer2_out[573] <= ~layer1_out[609];
     layer2_out[574] <= layer1_out[168];
     layer2_out[575] <= layer1_out[30];
     layer2_out[576] <= ~layer1_out[688];
     layer2_out[577] <= layer1_out[124];
     layer2_out[578] <= layer1_out[66] & layer1_out[67];
     layer2_out[579] <= 1'b1;
     layer2_out[580] <= layer1_out[71];
     layer2_out[581] <= layer1_out[96] & ~layer1_out[95];
     layer2_out[582] <= layer1_out[377];
     layer2_out[583] <= ~(layer1_out[164] | layer1_out[165]);
     layer2_out[584] <= layer1_out[735] & ~layer1_out[736];
     layer2_out[585] <= layer1_out[443] & layer1_out[444];
     layer2_out[586] <= ~layer1_out[560];
     layer2_out[587] <= ~layer1_out[725];
     layer2_out[588] <= layer1_out[38] & layer1_out[39];
     layer2_out[589] <= layer1_out[609] & layer1_out[610];
     layer2_out[590] <= layer1_out[339] & ~layer1_out[338];
     layer2_out[591] <= ~layer1_out[388];
     layer2_out[592] <= ~layer1_out[354];
     layer2_out[593] <= layer1_out[510];
     layer2_out[594] <= ~layer1_out[736];
     layer2_out[595] <= ~layer1_out[724];
     layer2_out[596] <= layer1_out[684];
     layer2_out[597] <= ~layer1_out[504] | layer1_out[503];
     layer2_out[598] <= ~layer1_out[101] | layer1_out[100];
     layer2_out[599] <= ~(layer1_out[119] & layer1_out[120]);
     layer2_out[600] <= ~(layer1_out[192] | layer1_out[193]);
     layer2_out[601] <= ~(layer1_out[709] | layer1_out[710]);
     layer2_out[602] <= 1'b0;
     layer2_out[603] <= layer1_out[495];
     layer2_out[604] <= 1'b0;
     layer2_out[605] <= ~(layer1_out[380] | layer1_out[381]);
     layer2_out[606] <= ~layer1_out[183];
     layer2_out[607] <= ~layer1_out[394];
     layer2_out[608] <= layer1_out[768] & layer1_out[769];
     layer2_out[609] <= layer1_out[99];
     layer2_out[610] <= ~layer1_out[645];
     layer2_out[611] <= layer1_out[642];
     layer2_out[612] <= ~(layer1_out[241] & layer1_out[242]);
     layer2_out[613] <= layer1_out[628];
     layer2_out[614] <= ~layer1_out[373] | layer1_out[372];
     layer2_out[615] <= ~layer1_out[548];
     layer2_out[616] <= layer1_out[767] & layer1_out[768];
     layer2_out[617] <= ~layer1_out[247];
     layer2_out[618] <= 1'b0;
     layer2_out[619] <= layer1_out[229];
     layer2_out[620] <= layer1_out[492];
     layer2_out[621] <= ~(layer1_out[484] & layer1_out[485]);
     layer2_out[622] <= layer1_out[10] & layer1_out[11];
     layer2_out[623] <= ~layer1_out[204];
     layer2_out[624] <= layer1_out[95];
     layer2_out[625] <= layer1_out[777] & ~layer1_out[776];
     layer2_out[626] <= layer1_out[227];
     layer2_out[627] <= ~layer1_out[273];
     layer2_out[628] <= ~layer1_out[678] | layer1_out[679];
     layer2_out[629] <= ~layer1_out[654] | layer1_out[653];
     layer2_out[630] <= ~(layer1_out[786] ^ layer1_out[787]);
     layer2_out[631] <= layer1_out[291];
     layer2_out[632] <= layer1_out[480] & layer1_out[481];
     layer2_out[633] <= ~(layer1_out[710] & layer1_out[711]);
     layer2_out[634] <= ~layer1_out[321];
     layer2_out[635] <= ~layer1_out[247] | layer1_out[246];
     layer2_out[636] <= layer1_out[380];
     layer2_out[637] <= ~layer1_out[221];
     layer2_out[638] <= ~layer1_out[178] | layer1_out[177];
     layer2_out[639] <= layer1_out[168];
     layer2_out[640] <= layer1_out[294] & ~layer1_out[295];
     layer2_out[641] <= ~(layer1_out[308] & layer1_out[309]);
     layer2_out[642] <= ~layer1_out[209];
     layer2_out[643] <= layer1_out[624] & ~layer1_out[623];
     layer2_out[644] <= 1'b0;
     layer2_out[645] <= layer1_out[742] & layer1_out[743];
     layer2_out[646] <= layer1_out[138] | layer1_out[139];
     layer2_out[647] <= layer1_out[102];
     layer2_out[648] <= layer1_out[347] | layer1_out[348];
     layer2_out[649] <= layer1_out[206] & layer1_out[207];
     layer2_out[650] <= layer1_out[502] | layer1_out[503];
     layer2_out[651] <= layer1_out[636];
     layer2_out[652] <= ~layer1_out[7];
     layer2_out[653] <= ~(layer1_out[427] & layer1_out[428]);
     layer2_out[654] <= 1'b0;
     layer2_out[655] <= layer1_out[621] & ~layer1_out[622];
     layer2_out[656] <= 1'b0;
     layer2_out[657] <= layer1_out[672];
     layer2_out[658] <= ~layer1_out[634] | layer1_out[633];
     layer2_out[659] <= ~layer1_out[108] | layer1_out[109];
     layer2_out[660] <= layer1_out[551] & ~layer1_out[552];
     layer2_out[661] <= layer1_out[390];
     layer2_out[662] <= ~(layer1_out[152] & layer1_out[153]);
     layer2_out[663] <= ~layer1_out[14];
     layer2_out[664] <= ~layer1_out[527];
     layer2_out[665] <= layer1_out[405] & layer1_out[406];
     layer2_out[666] <= layer1_out[749] ^ layer1_out[750];
     layer2_out[667] <= ~layer1_out[557];
     layer2_out[668] <= ~layer1_out[699];
     layer2_out[669] <= layer1_out[665] ^ layer1_out[666];
     layer2_out[670] <= layer1_out[761];
     layer2_out[671] <= layer1_out[724] | layer1_out[725];
     layer2_out[672] <= layer1_out[375] ^ layer1_out[376];
     layer2_out[673] <= ~(layer1_out[505] | layer1_out[506]);
     layer2_out[674] <= layer1_out[486] & layer1_out[487];
     layer2_out[675] <= ~layer1_out[574];
     layer2_out[676] <= ~layer1_out[131] | layer1_out[132];
     layer2_out[677] <= layer1_out[270];
     layer2_out[678] <= ~(layer1_out[130] | layer1_out[131]);
     layer2_out[679] <= layer1_out[157];
     layer2_out[680] <= layer1_out[587] & layer1_out[588];
     layer2_out[681] <= ~(layer1_out[416] | layer1_out[417]);
     layer2_out[682] <= ~layer1_out[425];
     layer2_out[683] <= ~layer1_out[537];
     layer2_out[684] <= ~layer1_out[714] | layer1_out[713];
     layer2_out[685] <= layer1_out[60] & ~layer1_out[61];
     layer2_out[686] <= ~layer1_out[197];
     layer2_out[687] <= layer1_out[173];
     layer2_out[688] <= layer1_out[384] & ~layer1_out[383];
     layer2_out[689] <= ~layer1_out[344];
     layer2_out[690] <= 1'b0;
     layer2_out[691] <= ~(layer1_out[322] | layer1_out[323]);
     layer2_out[692] <= ~(layer1_out[398] & layer1_out[399]);
     layer2_out[693] <= ~layer1_out[357];
     layer2_out[694] <= ~layer1_out[237];
     layer2_out[695] <= layer1_out[299];
     layer2_out[696] <= ~layer1_out[332] | layer1_out[331];
     layer2_out[697] <= ~layer1_out[685];
     layer2_out[698] <= layer1_out[626];
     layer2_out[699] <= layer1_out[345] & ~layer1_out[344];
     layer2_out[700] <= layer1_out[596];
     layer2_out[701] <= ~layer1_out[321];
     layer2_out[702] <= layer1_out[416] & ~layer1_out[415];
     layer2_out[703] <= layer1_out[513] ^ layer1_out[514];
     layer2_out[704] <= ~layer1_out[764] | layer1_out[763];
     layer2_out[705] <= ~layer1_out[170] | layer1_out[169];
     layer2_out[706] <= layer1_out[460] | layer1_out[461];
     layer2_out[707] <= layer1_out[699];
     layer2_out[708] <= layer1_out[712];
     layer2_out[709] <= 1'b0;
     layer2_out[710] <= ~layer1_out[591];
     layer2_out[711] <= ~(layer1_out[16] ^ layer1_out[17]);
     layer2_out[712] <= layer1_out[402];
     layer2_out[713] <= ~layer1_out[791];
     layer2_out[714] <= layer1_out[374];
     layer2_out[715] <= layer1_out[110];
     layer2_out[716] <= layer1_out[704] & ~layer1_out[703];
     layer2_out[717] <= ~layer1_out[463];
     layer2_out[718] <= ~layer1_out[606] | layer1_out[605];
     layer2_out[719] <= ~(layer1_out[306] ^ layer1_out[307]);
     layer2_out[720] <= ~layer1_out[606];
     layer2_out[721] <= ~layer1_out[784];
     layer2_out[722] <= layer1_out[364] & ~layer1_out[365];
     layer2_out[723] <= ~(layer1_out[208] & layer1_out[209]);
     layer2_out[724] <= ~layer1_out[778] | layer1_out[779];
     layer2_out[725] <= layer1_out[139] & ~layer1_out[140];
     layer2_out[726] <= layer1_out[367];
     layer2_out[727] <= ~layer1_out[785];
     layer2_out[728] <= layer1_out[83];
     layer2_out[729] <= layer1_out[210] & layer1_out[211];
     layer2_out[730] <= layer1_out[573] | layer1_out[574];
     layer2_out[731] <= ~(layer1_out[117] & layer1_out[118]);
     layer2_out[732] <= ~layer1_out[232] | layer1_out[231];
     layer2_out[733] <= layer1_out[84] & ~layer1_out[83];
     layer2_out[734] <= ~layer1_out[17] | layer1_out[18];
     layer2_out[735] <= ~(layer1_out[552] | layer1_out[553]);
     layer2_out[736] <= layer1_out[211] | layer1_out[212];
     layer2_out[737] <= layer1_out[784];
     layer2_out[738] <= layer1_out[614] ^ layer1_out[615];
     layer2_out[739] <= layer1_out[75];
     layer2_out[740] <= ~layer1_out[650];
     layer2_out[741] <= layer1_out[149] & ~layer1_out[150];
     layer2_out[742] <= layer1_out[164] & ~layer1_out[163];
     layer2_out[743] <= layer1_out[647];
     layer2_out[744] <= layer1_out[190] & ~layer1_out[189];
     layer2_out[745] <= ~(layer1_out[128] & layer1_out[129]);
     layer2_out[746] <= 1'b0;
     layer2_out[747] <= 1'b1;
     layer2_out[748] <= layer1_out[92];
     layer2_out[749] <= layer1_out[705] & ~layer1_out[704];
     layer2_out[750] <= 1'b1;
     layer2_out[751] <= ~layer1_out[170];
     layer2_out[752] <= ~(layer1_out[368] & layer1_out[369]);
     layer2_out[753] <= ~(layer1_out[651] & layer1_out[652]);
     layer2_out[754] <= layer1_out[288] & ~layer1_out[289];
     layer2_out[755] <= ~(layer1_out[511] & layer1_out[512]);
     layer2_out[756] <= ~(layer1_out[281] | layer1_out[282]);
     layer2_out[757] <= layer1_out[213] & ~layer1_out[214];
     layer2_out[758] <= layer1_out[429] & ~layer1_out[428];
     layer2_out[759] <= ~layer1_out[148];
     layer2_out[760] <= ~(layer1_out[214] & layer1_out[215]);
     layer2_out[761] <= ~layer1_out[576];
     layer2_out[762] <= layer1_out[453];
     layer2_out[763] <= ~layer1_out[238];
     layer2_out[764] <= layer1_out[39];
     layer2_out[765] <= ~layer1_out[302];
     layer2_out[766] <= layer1_out[265];
     layer2_out[767] <= ~(layer1_out[396] & layer1_out[397]);
     layer2_out[768] <= layer1_out[26];
     layer2_out[769] <= ~layer1_out[600] | layer1_out[601];
     layer2_out[770] <= ~layer1_out[697] | layer1_out[698];
     layer2_out[771] <= ~layer1_out[233] | layer1_out[234];
     layer2_out[772] <= layer1_out[766] & ~layer1_out[765];
     layer2_out[773] <= layer1_out[446] | layer1_out[447];
     layer2_out[774] <= layer1_out[478] & layer1_out[479];
     layer2_out[775] <= ~layer1_out[663];
     layer2_out[776] <= ~layer1_out[325] | layer1_out[324];
     layer2_out[777] <= layer1_out[337];
     layer2_out[778] <= layer1_out[718] & ~layer1_out[719];
     layer2_out[779] <= layer1_out[395];
     layer2_out[780] <= layer1_out[589] | layer1_out[590];
     layer2_out[781] <= layer1_out[733];
     layer2_out[782] <= 1'b1;
     layer2_out[783] <= layer1_out[176] & ~layer1_out[177];
     layer2_out[784] <= layer1_out[636] ^ layer1_out[637];
     layer2_out[785] <= layer1_out[652];
     layer2_out[786] <= layer1_out[766];
     layer2_out[787] <= layer1_out[441] & ~layer1_out[442];
     layer2_out[788] <= layer1_out[293];
     layer2_out[789] <= ~(layer1_out[544] & layer1_out[545]);
     layer2_out[790] <= layer1_out[143] | layer1_out[144];
     layer2_out[791] <= layer1_out[655] | layer1_out[656];
     layer2_out[792] <= layer1_out[336];
     layer2_out[793] <= ~layer1_out[475];
     layer2_out[794] <= ~(layer1_out[404] | layer1_out[405]);
     layer2_out[795] <= ~(layer1_out[115] & layer1_out[116]);
     layer2_out[796] <= ~(layer1_out[11] & layer1_out[12]);
     layer2_out[797] <= ~layer1_out[117] | layer1_out[116];
     layer2_out[798] <= layer1_out[579] | layer1_out[580];
     layer2_out[799] <= layer1_out[637] & ~layer1_out[638];
     layer3_out[0] <= ~layer2_out[745];
     layer3_out[1] <= layer2_out[219];
     layer3_out[2] <= layer2_out[721] & ~layer2_out[722];
     layer3_out[3] <= ~layer2_out[517] | layer2_out[516];
     layer3_out[4] <= ~layer2_out[156];
     layer3_out[5] <= layer2_out[515] & ~layer2_out[514];
     layer3_out[6] <= layer2_out[639];
     layer3_out[7] <= layer2_out[780];
     layer3_out[8] <= ~layer2_out[418] | layer2_out[417];
     layer3_out[9] <= ~layer2_out[490];
     layer3_out[10] <= layer2_out[280];
     layer3_out[11] <= ~layer2_out[217] | layer2_out[218];
     layer3_out[12] <= ~layer2_out[193];
     layer3_out[13] <= layer2_out[527] & ~layer2_out[526];
     layer3_out[14] <= ~layer2_out[634];
     layer3_out[15] <= layer2_out[0] & layer2_out[2];
     layer3_out[16] <= layer2_out[272] | layer2_out[273];
     layer3_out[17] <= ~layer2_out[761];
     layer3_out[18] <= layer2_out[491] & ~layer2_out[492];
     layer3_out[19] <= ~(layer2_out[594] | layer2_out[595]);
     layer3_out[20] <= ~layer2_out[52];
     layer3_out[21] <= layer2_out[441] ^ layer2_out[442];
     layer3_out[22] <= ~layer2_out[269];
     layer3_out[23] <= layer2_out[636];
     layer3_out[24] <= ~(layer2_out[778] & layer2_out[779]);
     layer3_out[25] <= layer2_out[516];
     layer3_out[26] <= layer2_out[782];
     layer3_out[27] <= ~layer2_out[571];
     layer3_out[28] <= layer2_out[349];
     layer3_out[29] <= ~(layer2_out[590] | layer2_out[591]);
     layer3_out[30] <= layer2_out[795];
     layer3_out[31] <= layer2_out[453] & ~layer2_out[454];
     layer3_out[32] <= ~layer2_out[382];
     layer3_out[33] <= ~layer2_out[657] | layer2_out[656];
     layer3_out[34] <= layer2_out[414];
     layer3_out[35] <= 1'b0;
     layer3_out[36] <= layer2_out[2];
     layer3_out[37] <= ~(layer2_out[757] & layer2_out[758]);
     layer3_out[38] <= ~(layer2_out[445] & layer2_out[446]);
     layer3_out[39] <= ~(layer2_out[783] & layer2_out[784]);
     layer3_out[40] <= layer2_out[548] & layer2_out[549];
     layer3_out[41] <= layer2_out[552] | layer2_out[553];
     layer3_out[42] <= layer2_out[11];
     layer3_out[43] <= ~(layer2_out[677] & layer2_out[678]);
     layer3_out[44] <= ~layer2_out[377];
     layer3_out[45] <= ~layer2_out[187] | layer2_out[188];
     layer3_out[46] <= ~layer2_out[67];
     layer3_out[47] <= layer2_out[786] & ~layer2_out[785];
     layer3_out[48] <= layer2_out[96];
     layer3_out[49] <= ~layer2_out[317];
     layer3_out[50] <= ~layer2_out[71] | layer2_out[72];
     layer3_out[51] <= layer2_out[80];
     layer3_out[52] <= ~layer2_out[694] | layer2_out[695];
     layer3_out[53] <= ~layer2_out[254];
     layer3_out[54] <= layer2_out[35] & layer2_out[36];
     layer3_out[55] <= ~layer2_out[653] | layer2_out[654];
     layer3_out[56] <= layer2_out[681] | layer2_out[682];
     layer3_out[57] <= ~layer2_out[315] | layer2_out[314];
     layer3_out[58] <= ~(layer2_out[378] & layer2_out[379]);
     layer3_out[59] <= ~layer2_out[83];
     layer3_out[60] <= ~layer2_out[274];
     layer3_out[61] <= layer2_out[422];
     layer3_out[62] <= ~layer2_out[82];
     layer3_out[63] <= layer2_out[247];
     layer3_out[64] <= layer2_out[167] | layer2_out[168];
     layer3_out[65] <= ~layer2_out[162];
     layer3_out[66] <= layer2_out[483];
     layer3_out[67] <= layer2_out[623];
     layer3_out[68] <= ~(layer2_out[86] & layer2_out[87]);
     layer3_out[69] <= layer2_out[482];
     layer3_out[70] <= layer2_out[11] & ~layer2_out[10];
     layer3_out[71] <= ~layer2_out[23];
     layer3_out[72] <= ~(layer2_out[254] | layer2_out[255]);
     layer3_out[73] <= ~(layer2_out[746] | layer2_out[747]);
     layer3_out[74] <= layer2_out[73] & layer2_out[74];
     layer3_out[75] <= layer2_out[137] & ~layer2_out[136];
     layer3_out[76] <= layer2_out[191];
     layer3_out[77] <= layer2_out[258] & layer2_out[259];
     layer3_out[78] <= layer2_out[367] | layer2_out[368];
     layer3_out[79] <= ~layer2_out[494];
     layer3_out[80] <= layer2_out[687];
     layer3_out[81] <= layer2_out[721];
     layer3_out[82] <= layer2_out[203];
     layer3_out[83] <= ~layer2_out[734];
     layer3_out[84] <= layer2_out[743] ^ layer2_out[744];
     layer3_out[85] <= layer2_out[268];
     layer3_out[86] <= 1'b1;
     layer3_out[87] <= layer2_out[247] & ~layer2_out[246];
     layer3_out[88] <= layer2_out[336] & ~layer2_out[335];
     layer3_out[89] <= layer2_out[87];
     layer3_out[90] <= ~layer2_out[769] | layer2_out[770];
     layer3_out[91] <= 1'b1;
     layer3_out[92] <= ~(layer2_out[408] | layer2_out[409]);
     layer3_out[93] <= ~layer2_out[207] | layer2_out[206];
     layer3_out[94] <= layer2_out[252];
     layer3_out[95] <= layer2_out[175];
     layer3_out[96] <= layer2_out[325] & layer2_out[326];
     layer3_out[97] <= layer2_out[593] & layer2_out[594];
     layer3_out[98] <= 1'b1;
     layer3_out[99] <= ~layer2_out[517];
     layer3_out[100] <= 1'b1;
     layer3_out[101] <= ~layer2_out[587] | layer2_out[588];
     layer3_out[102] <= layer2_out[110] & layer2_out[111];
     layer3_out[103] <= ~(layer2_out[279] | layer2_out[280]);
     layer3_out[104] <= ~(layer2_out[595] ^ layer2_out[596]);
     layer3_out[105] <= ~(layer2_out[107] & layer2_out[108]);
     layer3_out[106] <= ~layer2_out[700];
     layer3_out[107] <= layer2_out[403] & ~layer2_out[404];
     layer3_out[108] <= ~(layer2_out[100] & layer2_out[101]);
     layer3_out[109] <= ~layer2_out[96] | layer2_out[97];
     layer3_out[110] <= ~(layer2_out[4] & layer2_out[5]);
     layer3_out[111] <= layer2_out[194];
     layer3_out[112] <= layer2_out[78] & ~layer2_out[79];
     layer3_out[113] <= layer2_out[688];
     layer3_out[114] <= layer2_out[633];
     layer3_out[115] <= layer2_out[494] & ~layer2_out[495];
     layer3_out[116] <= layer2_out[303] | layer2_out[304];
     layer3_out[117] <= layer2_out[41] & ~layer2_out[42];
     layer3_out[118] <= ~layer2_out[791];
     layer3_out[119] <= 1'b0;
     layer3_out[120] <= ~layer2_out[514];
     layer3_out[121] <= layer2_out[257] | layer2_out[258];
     layer3_out[122] <= ~layer2_out[2] | layer2_out[3];
     layer3_out[123] <= ~(layer2_out[622] ^ layer2_out[623]);
     layer3_out[124] <= ~(layer2_out[380] | layer2_out[381]);
     layer3_out[125] <= layer2_out[13];
     layer3_out[126] <= ~layer2_out[704];
     layer3_out[127] <= layer2_out[141] & ~layer2_out[142];
     layer3_out[128] <= layer2_out[70] & ~layer2_out[71];
     layer3_out[129] <= ~layer2_out[499];
     layer3_out[130] <= 1'b0;
     layer3_out[131] <= layer2_out[120] | layer2_out[121];
     layer3_out[132] <= layer2_out[172] & ~layer2_out[171];
     layer3_out[133] <= 1'b0;
     layer3_out[134] <= layer2_out[658] & ~layer2_out[659];
     layer3_out[135] <= ~(layer2_out[138] | layer2_out[139]);
     layer3_out[136] <= layer2_out[64] & layer2_out[65];
     layer3_out[137] <= layer2_out[600] & layer2_out[601];
     layer3_out[138] <= layer2_out[465];
     layer3_out[139] <= ~layer2_out[376];
     layer3_out[140] <= ~layer2_out[506];
     layer3_out[141] <= layer2_out[430] & layer2_out[431];
     layer3_out[142] <= ~layer2_out[522] | layer2_out[523];
     layer3_out[143] <= layer2_out[210];
     layer3_out[144] <= layer2_out[304];
     layer3_out[145] <= ~layer2_out[681] | layer2_out[680];
     layer3_out[146] <= ~layer2_out[548];
     layer3_out[147] <= layer2_out[260] & ~layer2_out[259];
     layer3_out[148] <= ~(layer2_out[326] & layer2_out[327]);
     layer3_out[149] <= ~layer2_out[228];
     layer3_out[150] <= ~layer2_out[143];
     layer3_out[151] <= ~layer2_out[121];
     layer3_out[152] <= ~(layer2_out[573] ^ layer2_out[574]);
     layer3_out[153] <= ~layer2_out[567] | layer2_out[566];
     layer3_out[154] <= ~(layer2_out[369] & layer2_out[370]);
     layer3_out[155] <= layer2_out[732] | layer2_out[733];
     layer3_out[156] <= ~(layer2_out[189] | layer2_out[190]);
     layer3_out[157] <= ~layer2_out[461];
     layer3_out[158] <= layer2_out[584] & ~layer2_out[585];
     layer3_out[159] <= ~layer2_out[133];
     layer3_out[160] <= layer2_out[648];
     layer3_out[161] <= ~layer2_out[157];
     layer3_out[162] <= layer2_out[395];
     layer3_out[163] <= layer2_out[47];
     layer3_out[164] <= layer2_out[406] & ~layer2_out[407];
     layer3_out[165] <= layer2_out[191] | layer2_out[192];
     layer3_out[166] <= ~layer2_out[204];
     layer3_out[167] <= layer2_out[282];
     layer3_out[168] <= ~(layer2_out[150] | layer2_out[151]);
     layer3_out[169] <= ~layer2_out[382];
     layer3_out[170] <= layer2_out[324] | layer2_out[325];
     layer3_out[171] <= ~layer2_out[39] | layer2_out[38];
     layer3_out[172] <= layer2_out[231];
     layer3_out[173] <= layer2_out[456];
     layer3_out[174] <= layer2_out[425];
     layer3_out[175] <= ~layer2_out[709] | layer2_out[708];
     layer3_out[176] <= layer2_out[367] & ~layer2_out[366];
     layer3_out[177] <= 1'b0;
     layer3_out[178] <= layer2_out[37] & ~layer2_out[38];
     layer3_out[179] <= ~layer2_out[100];
     layer3_out[180] <= ~layer2_out[184] | layer2_out[185];
     layer3_out[181] <= layer2_out[607];
     layer3_out[182] <= layer2_out[48];
     layer3_out[183] <= layer2_out[129] | layer2_out[130];
     layer3_out[184] <= ~(layer2_out[649] & layer2_out[650]);
     layer3_out[185] <= ~layer2_out[463];
     layer3_out[186] <= ~(layer2_out[296] | layer2_out[297]);
     layer3_out[187] <= 1'b1;
     layer3_out[188] <= layer2_out[217];
     layer3_out[189] <= layer2_out[271] & ~layer2_out[270];
     layer3_out[190] <= layer2_out[624];
     layer3_out[191] <= ~layer2_out[550];
     layer3_out[192] <= ~(layer2_out[521] & layer2_out[522]);
     layer3_out[193] <= ~layer2_out[149];
     layer3_out[194] <= 1'b1;
     layer3_out[195] <= 1'b0;
     layer3_out[196] <= 1'b0;
     layer3_out[197] <= layer2_out[114] & layer2_out[115];
     layer3_out[198] <= ~layer2_out[529];
     layer3_out[199] <= 1'b0;
     layer3_out[200] <= layer2_out[689] ^ layer2_out[690];
     layer3_out[201] <= ~(layer2_out[690] & layer2_out[691]);
     layer3_out[202] <= layer2_out[245] & layer2_out[246];
     layer3_out[203] <= ~(layer2_out[126] | layer2_out[127]);
     layer3_out[204] <= ~(layer2_out[756] | layer2_out[757]);
     layer3_out[205] <= ~(layer2_out[527] ^ layer2_out[528]);
     layer3_out[206] <= ~(layer2_out[84] | layer2_out[85]);
     layer3_out[207] <= layer2_out[135];
     layer3_out[208] <= 1'b1;
     layer3_out[209] <= ~layer2_out[457];
     layer3_out[210] <= layer2_out[166];
     layer3_out[211] <= layer2_out[796];
     layer3_out[212] <= layer2_out[738];
     layer3_out[213] <= ~(layer2_out[766] ^ layer2_out[767]);
     layer3_out[214] <= layer2_out[292] & ~layer2_out[293];
     layer3_out[215] <= layer2_out[255] & layer2_out[256];
     layer3_out[216] <= ~layer2_out[569];
     layer3_out[217] <= layer2_out[670];
     layer3_out[218] <= layer2_out[641];
     layer3_out[219] <= ~(layer2_out[602] & layer2_out[603]);
     layer3_out[220] <= layer2_out[119] | layer2_out[120];
     layer3_out[221] <= ~(layer2_out[358] | layer2_out[359]);
     layer3_out[222] <= layer2_out[211] | layer2_out[212];
     layer3_out[223] <= layer2_out[75] | layer2_out[76];
     layer3_out[224] <= ~(layer2_out[446] | layer2_out[447]);
     layer3_out[225] <= ~layer2_out[778];
     layer3_out[226] <= layer2_out[56];
     layer3_out[227] <= layer2_out[320] ^ layer2_out[321];
     layer3_out[228] <= layer2_out[271] & layer2_out[272];
     layer3_out[229] <= ~layer2_out[712] | layer2_out[713];
     layer3_out[230] <= layer2_out[639] ^ layer2_out[640];
     layer3_out[231] <= ~layer2_out[532] | layer2_out[531];
     layer3_out[232] <= ~layer2_out[234] | layer2_out[233];
     layer3_out[233] <= layer2_out[483];
     layer3_out[234] <= layer2_out[28];
     layer3_out[235] <= ~layer2_out[43];
     layer3_out[236] <= ~layer2_out[620];
     layer3_out[237] <= ~layer2_out[558];
     layer3_out[238] <= layer2_out[294];
     layer3_out[239] <= ~layer2_out[90];
     layer3_out[240] <= layer2_out[348] & ~layer2_out[349];
     layer3_out[241] <= ~(layer2_out[582] & layer2_out[583]);
     layer3_out[242] <= ~(layer2_out[628] | layer2_out[629]);
     layer3_out[243] <= ~layer2_out[507] | layer2_out[508];
     layer3_out[244] <= ~(layer2_out[687] & layer2_out[688]);
     layer3_out[245] <= layer2_out[154] & ~layer2_out[153];
     layer3_out[246] <= ~(layer2_out[754] & layer2_out[755]);
     layer3_out[247] <= layer2_out[459];
     layer3_out[248] <= layer2_out[760];
     layer3_out[249] <= layer2_out[88] & ~layer2_out[89];
     layer3_out[250] <= ~layer2_out[94];
     layer3_out[251] <= layer2_out[64];
     layer3_out[252] <= layer2_out[302];
     layer3_out[253] <= layer2_out[603];
     layer3_out[254] <= ~(layer2_out[509] ^ layer2_out[510]);
     layer3_out[255] <= layer2_out[668] & ~layer2_out[667];
     layer3_out[256] <= ~layer2_out[682];
     layer3_out[257] <= ~layer2_out[147] | layer2_out[148];
     layer3_out[258] <= ~layer2_out[579];
     layer3_out[259] <= layer2_out[467] | layer2_out[468];
     layer3_out[260] <= layer2_out[164];
     layer3_out[261] <= layer2_out[149] & ~layer2_out[150];
     layer3_out[262] <= layer2_out[208];
     layer3_out[263] <= ~layer2_out[431];
     layer3_out[264] <= layer2_out[331] & ~layer2_out[332];
     layer3_out[265] <= ~(layer2_out[30] & layer2_out[31]);
     layer3_out[266] <= 1'b1;
     layer3_out[267] <= layer2_out[402];
     layer3_out[268] <= layer2_out[745] & ~layer2_out[744];
     layer3_out[269] <= ~(layer2_out[659] & layer2_out[660]);
     layer3_out[270] <= ~(layer2_out[267] | layer2_out[268]);
     layer3_out[271] <= layer2_out[596];
     layer3_out[272] <= layer2_out[537] ^ layer2_out[538];
     layer3_out[273] <= layer2_out[25] | layer2_out[26];
     layer3_out[274] <= ~(layer2_out[711] | layer2_out[712]);
     layer3_out[275] <= ~layer2_out[736];
     layer3_out[276] <= ~layer2_out[334] | layer2_out[335];
     layer3_out[277] <= ~layer2_out[587] | layer2_out[586];
     layer3_out[278] <= ~(layer2_out[644] | layer2_out[645]);
     layer3_out[279] <= layer2_out[170] & ~layer2_out[171];
     layer3_out[280] <= layer2_out[538];
     layer3_out[281] <= ~(layer2_out[322] ^ layer2_out[323]);
     layer3_out[282] <= ~layer2_out[443];
     layer3_out[283] <= ~(layer2_out[613] ^ layer2_out[614]);
     layer3_out[284] <= layer2_out[342] | layer2_out[343];
     layer3_out[285] <= ~(layer2_out[31] ^ layer2_out[32]);
     layer3_out[286] <= ~layer2_out[717];
     layer3_out[287] <= ~layer2_out[523];
     layer3_out[288] <= layer2_out[437] & ~layer2_out[436];
     layer3_out[289] <= ~(layer2_out[664] ^ layer2_out[665]);
     layer3_out[290] <= ~layer2_out[93] | layer2_out[92];
     layer3_out[291] <= layer2_out[379] & ~layer2_out[380];
     layer3_out[292] <= layer2_out[432];
     layer3_out[293] <= ~layer2_out[572] | layer2_out[571];
     layer3_out[294] <= ~(layer2_out[543] | layer2_out[544]);
     layer3_out[295] <= ~layer2_out[651] | layer2_out[652];
     layer3_out[296] <= layer2_out[417] & ~layer2_out[416];
     layer3_out[297] <= ~layer2_out[700];
     layer3_out[298] <= layer2_out[410] & ~layer2_out[409];
     layer3_out[299] <= layer2_out[155];
     layer3_out[300] <= ~(layer2_out[140] & layer2_out[141]);
     layer3_out[301] <= ~layer2_out[153];
     layer3_out[302] <= layer2_out[614] & ~layer2_out[615];
     layer3_out[303] <= layer2_out[240] & ~layer2_out[239];
     layer3_out[304] <= layer2_out[180];
     layer3_out[305] <= layer2_out[410] & ~layer2_out[411];
     layer3_out[306] <= ~(layer2_out[278] & layer2_out[279]);
     layer3_out[307] <= ~(layer2_out[212] & layer2_out[213]);
     layer3_out[308] <= layer2_out[484];
     layer3_out[309] <= ~layer2_out[47];
     layer3_out[310] <= 1'b0;
     layer3_out[311] <= layer2_out[54];
     layer3_out[312] <= layer2_out[500] | layer2_out[501];
     layer3_out[313] <= layer2_out[496] & ~layer2_out[495];
     layer3_out[314] <= layer2_out[128] | layer2_out[129];
     layer3_out[315] <= ~layer2_out[124];
     layer3_out[316] <= ~(layer2_out[158] | layer2_out[159]);
     layer3_out[317] <= layer2_out[350];
     layer3_out[318] <= ~layer2_out[14];
     layer3_out[319] <= ~layer2_out[610];
     layer3_out[320] <= ~layer2_out[281];
     layer3_out[321] <= ~layer2_out[525] | layer2_out[524];
     layer3_out[322] <= layer2_out[427] | layer2_out[428];
     layer3_out[323] <= layer2_out[336] | layer2_out[337];
     layer3_out[324] <= layer2_out[230] & ~layer2_out[231];
     layer3_out[325] <= layer2_out[221];
     layer3_out[326] <= layer2_out[377] & ~layer2_out[376];
     layer3_out[327] <= ~(layer2_out[283] & layer2_out[284]);
     layer3_out[328] <= ~layer2_out[771];
     layer3_out[329] <= ~layer2_out[720];
     layer3_out[330] <= layer2_out[503] & ~layer2_out[502];
     layer3_out[331] <= layer2_out[371];
     layer3_out[332] <= ~(layer2_out[792] | layer2_out[793]);
     layer3_out[333] <= 1'b0;
     layer3_out[334] <= layer2_out[361];
     layer3_out[335] <= ~layer2_out[399] | layer2_out[398];
     layer3_out[336] <= ~layer2_out[615];
     layer3_out[337] <= ~layer2_out[202] | layer2_out[203];
     layer3_out[338] <= ~layer2_out[356] | layer2_out[357];
     layer3_out[339] <= ~layer2_out[774];
     layer3_out[340] <= ~layer2_out[529] | layer2_out[530];
     layer3_out[341] <= ~layer2_out[61] | layer2_out[62];
     layer3_out[342] <= layer2_out[274];
     layer3_out[343] <= layer2_out[276] | layer2_out[277];
     layer3_out[344] <= ~(layer2_out[787] & layer2_out[788]);
     layer3_out[345] <= layer2_out[511];
     layer3_out[346] <= ~(layer2_out[591] & layer2_out[592]);
     layer3_out[347] <= ~layer2_out[227] | layer2_out[226];
     layer3_out[348] <= ~layer2_out[116];
     layer3_out[349] <= ~layer2_out[209];
     layer3_out[350] <= layer2_out[661] & ~layer2_out[662];
     layer3_out[351] <= layer2_out[793] & layer2_out[794];
     layer3_out[352] <= ~(layer2_out[532] & layer2_out[533]);
     layer3_out[353] <= ~layer2_out[461] | layer2_out[462];
     layer3_out[354] <= layer2_out[213];
     layer3_out[355] <= ~layer2_out[702];
     layer3_out[356] <= ~layer2_out[759] | layer2_out[758];
     layer3_out[357] <= ~layer2_out[570];
     layer3_out[358] <= 1'b1;
     layer3_out[359] <= layer2_out[630];
     layer3_out[360] <= layer2_out[790] ^ layer2_out[791];
     layer3_out[361] <= ~(layer2_out[776] & layer2_out[777]);
     layer3_out[362] <= ~layer2_out[311] | layer2_out[310];
     layer3_out[363] <= ~(layer2_out[68] ^ layer2_out[69]);
     layer3_out[364] <= layer2_out[487] & ~layer2_out[488];
     layer3_out[365] <= layer2_out[775] & ~layer2_out[774];
     layer3_out[366] <= ~layer2_out[198];
     layer3_out[367] <= ~layer2_out[498] | layer2_out[497];
     layer3_out[368] <= ~(layer2_out[359] | layer2_out[360]);
     layer3_out[369] <= layer2_out[122] & ~layer2_out[123];
     layer3_out[370] <= layer2_out[540] | layer2_out[541];
     layer3_out[371] <= ~layer2_out[452];
     layer3_out[372] <= layer2_out[542] & ~layer2_out[543];
     layer3_out[373] <= layer2_out[276];
     layer3_out[374] <= 1'b1;
     layer3_out[375] <= ~layer2_out[52];
     layer3_out[376] <= layer2_out[340];
     layer3_out[377] <= ~layer2_out[284];
     layer3_out[378] <= layer2_out[90] | layer2_out[91];
     layer3_out[379] <= layer2_out[263];
     layer3_out[380] <= 1'b0;
     layer3_out[381] <= layer2_out[75];
     layer3_out[382] <= ~layer2_out[627];
     layer3_out[383] <= layer2_out[670] ^ layer2_out[671];
     layer3_out[384] <= layer2_out[227] | layer2_out[228];
     layer3_out[385] <= layer2_out[160] | layer2_out[161];
     layer3_out[386] <= layer2_out[104];
     layer3_out[387] <= layer2_out[384] & ~layer2_out[385];
     layer3_out[388] <= ~(layer2_out[166] | layer2_out[167]);
     layer3_out[389] <= layer2_out[238];
     layer3_out[390] <= ~layer2_out[589] | layer2_out[588];
     layer3_out[391] <= layer2_out[9] & ~layer2_out[8];
     layer3_out[392] <= 1'b1;
     layer3_out[393] <= ~(layer2_out[442] | layer2_out[443]);
     layer3_out[394] <= ~layer2_out[225];
     layer3_out[395] <= layer2_out[119];
     layer3_out[396] <= layer2_out[510] & layer2_out[511];
     layer3_out[397] <= 1'b0;
     layer3_out[398] <= ~layer2_out[341] | layer2_out[342];
     layer3_out[399] <= ~layer2_out[696];
     layer3_out[400] <= ~(layer2_out[134] | layer2_out[135]);
     layer3_out[401] <= 1'b0;
     layer3_out[402] <= ~layer2_out[201];
     layer3_out[403] <= ~layer2_out[647];
     layer3_out[404] <= ~layer2_out[222];
     layer3_out[405] <= layer2_out[173] & ~layer2_out[174];
     layer3_out[406] <= layer2_out[565] ^ layer2_out[566];
     layer3_out[407] <= layer2_out[572];
     layer3_out[408] <= layer2_out[605];
     layer3_out[409] <= layer2_out[199];
     layer3_out[410] <= ~layer2_out[474];
     layer3_out[411] <= layer2_out[400] & layer2_out[401];
     layer3_out[412] <= ~(layer2_out[332] & layer2_out[333]);
     layer3_out[413] <= layer2_out[116] & ~layer2_out[115];
     layer3_out[414] <= ~layer2_out[521];
     layer3_out[415] <= ~(layer2_out[668] | layer2_out[669]);
     layer3_out[416] <= ~layer2_out[24];
     layer3_out[417] <= layer2_out[607] & ~layer2_out[608];
     layer3_out[418] <= layer2_out[250];
     layer3_out[419] <= layer2_out[242] & ~layer2_out[243];
     layer3_out[420] <= layer2_out[783];
     layer3_out[421] <= layer2_out[740];
     layer3_out[422] <= layer2_out[319] | layer2_out[320];
     layer3_out[423] <= layer2_out[598] | layer2_out[599];
     layer3_out[424] <= layer2_out[57] & ~layer2_out[56];
     layer3_out[425] <= ~(layer2_out[168] & layer2_out[169]);
     layer3_out[426] <= ~(layer2_out[641] ^ layer2_out[642]);
     layer3_out[427] <= ~layer2_out[450] | layer2_out[449];
     layer3_out[428] <= ~layer2_out[455];
     layer3_out[429] <= layer2_out[646] & ~layer2_out[645];
     layer3_out[430] <= layer2_out[631] & ~layer2_out[632];
     layer3_out[431] <= ~(layer2_out[374] & layer2_out[375]);
     layer3_out[432] <= layer2_out[236];
     layer3_out[433] <= ~(layer2_out[159] | layer2_out[160]);
     layer3_out[434] <= ~(layer2_out[767] & layer2_out[768]);
     layer3_out[435] <= layer2_out[702] & layer2_out[703];
     layer3_out[436] <= 1'b1;
     layer3_out[437] <= layer2_out[294] | layer2_out[295];
     layer3_out[438] <= ~layer2_out[751] | layer2_out[752];
     layer3_out[439] <= layer2_out[423];
     layer3_out[440] <= ~layer2_out[133];
     layer3_out[441] <= layer2_out[740] & ~layer2_out[741];
     layer3_out[442] <= ~layer2_out[501] | layer2_out[502];
     layer3_out[443] <= layer2_out[12] & ~layer2_out[13];
     layer3_out[444] <= layer2_out[724];
     layer3_out[445] <= ~layer2_out[239];
     layer3_out[446] <= layer2_out[161] & layer2_out[162];
     layer3_out[447] <= ~layer2_out[725];
     layer3_out[448] <= layer2_out[124] | layer2_out[125];
     layer3_out[449] <= ~layer2_out[578];
     layer3_out[450] <= layer2_out[146] | layer2_out[147];
     layer3_out[451] <= ~layer2_out[21] | layer2_out[22];
     layer3_out[452] <= layer2_out[399] & layer2_out[400];
     layer3_out[453] <= ~layer2_out[20];
     layer3_out[454] <= layer2_out[333] & layer2_out[334];
     layer3_out[455] <= layer2_out[219] & ~layer2_out[220];
     layer3_out[456] <= ~(layer2_out[475] ^ layer2_out[476]);
     layer3_out[457] <= ~layer2_out[328];
     layer3_out[458] <= ~layer2_out[187] | layer2_out[186];
     layer3_out[459] <= 1'b1;
     layer3_out[460] <= layer2_out[707] & ~layer2_out[708];
     layer3_out[461] <= layer2_out[756] & ~layer2_out[755];
     layer3_out[462] <= layer2_out[439] & ~layer2_out[440];
     layer3_out[463] <= layer2_out[364] & layer2_out[365];
     layer3_out[464] <= layer2_out[288];
     layer3_out[465] <= layer2_out[224];
     layer3_out[466] <= ~layer2_out[27];
     layer3_out[467] <= 1'b1;
     layer3_out[468] <= layer2_out[575];
     layer3_out[469] <= ~layer2_out[222];
     layer3_out[470] <= ~layer2_out[711] | layer2_out[710];
     layer3_out[471] <= layer2_out[210] & layer2_out[211];
     layer3_out[472] <= layer2_out[192] & layer2_out[193];
     layer3_out[473] <= ~layer2_out[16] | layer2_out[15];
     layer3_out[474] <= ~layer2_out[695];
     layer3_out[475] <= layer2_out[631];
     layer3_out[476] <= layer2_out[737] | layer2_out[738];
     layer3_out[477] <= ~layer2_out[60];
     layer3_out[478] <= ~layer2_out[489];
     layer3_out[479] <= layer2_out[340] | layer2_out[341];
     layer3_out[480] <= ~layer2_out[513];
     layer3_out[481] <= ~layer2_out[713];
     layer3_out[482] <= ~(layer2_out[433] & layer2_out[434]);
     layer3_out[483] <= layer2_out[545] ^ layer2_out[546];
     layer3_out[484] <= layer2_out[574];
     layer3_out[485] <= layer2_out[781];
     layer3_out[486] <= ~layer2_out[518];
     layer3_out[487] <= layer2_out[608] & ~layer2_out[609];
     layer3_out[488] <= ~layer2_out[590];
     layer3_out[489] <= layer2_out[45] | layer2_out[46];
     layer3_out[490] <= 1'b0;
     layer3_out[491] <= ~layer2_out[308] | layer2_out[307];
     layer3_out[492] <= layer2_out[264] & layer2_out[265];
     layer3_out[493] <= 1'b0;
     layer3_out[494] <= ~layer2_out[389] | layer2_out[390];
     layer3_out[495] <= layer2_out[583];
     layer3_out[496] <= layer2_out[506] & ~layer2_out[507];
     layer3_out[497] <= layer2_out[585] & ~layer2_out[586];
     layer3_out[498] <= ~layer2_out[112] | layer2_out[111];
     layer3_out[499] <= layer2_out[421];
     layer3_out[500] <= ~layer2_out[555];
     layer3_out[501] <= layer2_out[41] & ~layer2_out[40];
     layer3_out[502] <= ~(layer2_out[243] | layer2_out[244]);
     layer3_out[503] <= ~layer2_out[139];
     layer3_out[504] <= ~(layer2_out[611] | layer2_out[612]);
     layer3_out[505] <= layer2_out[784] & layer2_out[785];
     layer3_out[506] <= layer2_out[61] & ~layer2_out[60];
     layer3_out[507] <= ~layer2_out[343];
     layer3_out[508] <= layer2_out[109];
     layer3_out[509] <= ~layer2_out[266];
     layer3_out[510] <= layer2_out[373];
     layer3_out[511] <= ~layer2_out[562] | layer2_out[563];
     layer3_out[512] <= layer2_out[329] & ~layer2_out[330];
     layer3_out[513] <= ~layer2_out[444] | layer2_out[445];
     layer3_out[514] <= ~(layer2_out[544] | layer2_out[545]);
     layer3_out[515] <= layer2_out[6] | layer2_out[7];
     layer3_out[516] <= layer2_out[285];
     layer3_out[517] <= layer2_out[557] ^ layer2_out[558];
     layer3_out[518] <= layer2_out[296] & ~layer2_out[295];
     layer3_out[519] <= ~layer2_out[613];
     layer3_out[520] <= layer2_out[102];
     layer3_out[521] <= layer2_out[54] ^ layer2_out[55];
     layer3_out[522] <= layer2_out[323] | layer2_out[324];
     layer3_out[523] <= 1'b0;
     layer3_out[524] <= ~layer2_out[679];
     layer3_out[525] <= layer2_out[627];
     layer3_out[526] <= ~layer2_out[547];
     layer3_out[527] <= 1'b0;
     layer3_out[528] <= layer2_out[257];
     layer3_out[529] <= ~(layer2_out[469] | layer2_out[470]);
     layer3_out[530] <= ~(layer2_out[395] ^ layer2_out[396]);
     layer3_out[531] <= ~layer2_out[80];
     layer3_out[532] <= ~layer2_out[787];
     layer3_out[533] <= ~(layer2_out[69] | layer2_out[70]);
     layer3_out[534] <= ~layer2_out[292];
     layer3_out[535] <= ~layer2_out[300];
     layer3_out[536] <= layer2_out[790];
     layer3_out[537] <= layer2_out[10];
     layer3_out[538] <= ~layer2_out[39] | layer2_out[40];
     layer3_out[539] <= ~layer2_out[170] | layer2_out[169];
     layer3_out[540] <= layer2_out[728] & ~layer2_out[729];
     layer3_out[541] <= ~layer2_out[568] | layer2_out[567];
     layer3_out[542] <= layer2_out[202] & ~layer2_out[201];
     layer3_out[543] <= ~(layer2_out[260] & layer2_out[261]);
     layer3_out[544] <= layer2_out[196];
     layer3_out[545] <= ~layer2_out[769];
     layer3_out[546] <= layer2_out[397];
     layer3_out[547] <= layer2_out[653] & ~layer2_out[652];
     layer3_out[548] <= layer2_out[44] & ~layer2_out[45];
     layer3_out[549] <= layer2_out[112] & layer2_out[113];
     layer3_out[550] <= ~layer2_out[519];
     layer3_out[551] <= ~layer2_out[253];
     layer3_out[552] <= 1'b0;
     layer3_out[553] <= ~(layer2_out[318] & layer2_out[319]);
     layer3_out[554] <= layer2_out[478];
     layer3_out[555] <= layer2_out[662] ^ layer2_out[663];
     layer3_out[556] <= ~layer2_out[651];
     layer3_out[557] <= ~layer2_out[59];
     layer3_out[558] <= ~(layer2_out[244] | layer2_out[245]);
     layer3_out[559] <= ~layer2_out[561];
     layer3_out[560] <= ~layer2_out[599];
     layer3_out[561] <= layer2_out[145] ^ layer2_out[146];
     layer3_out[562] <= ~layer2_out[492];
     layer3_out[563] <= layer2_out[91] & layer2_out[92];
     layer3_out[564] <= 1'b0;
     layer3_out[565] <= layer2_out[23] | layer2_out[24];
     layer3_out[566] <= layer2_out[51];
     layer3_out[567] <= layer2_out[72] & layer2_out[73];
     layer3_out[568] <= layer2_out[609] & layer2_out[610];
     layer3_out[569] <= ~layer2_out[354] | layer2_out[353];
     layer3_out[570] <= layer2_out[387];
     layer3_out[571] <= layer2_out[789] & ~layer2_out[788];
     layer3_out[572] <= ~layer2_out[298] | layer2_out[299];
     layer3_out[573] <= ~(layer2_out[592] | layer2_out[593]);
     layer3_out[574] <= layer2_out[535];
     layer3_out[575] <= layer2_out[436] & ~layer2_out[435];
     layer3_out[576] <= ~layer2_out[463] | layer2_out[464];
     layer3_out[577] <= layer2_out[151];
     layer3_out[578] <= ~layer2_out[564];
     layer3_out[579] <= ~layer2_out[33];
     layer3_out[580] <= layer2_out[347];
     layer3_out[581] <= layer2_out[509];
     layer3_out[582] <= ~layer2_out[665];
     layer3_out[583] <= layer2_out[480];
     layer3_out[584] <= layer2_out[534];
     layer3_out[585] <= ~layer2_out[531];
     layer3_out[586] <= layer2_out[130] | layer2_out[131];
     layer3_out[587] <= ~layer2_out[407];
     layer3_out[588] <= layer2_out[318] & ~layer2_out[317];
     layer3_out[589] <= ~layer2_out[581];
     layer3_out[590] <= layer2_out[727] & ~layer2_out[726];
     layer3_out[591] <= layer2_out[391];
     layer3_out[592] <= layer2_out[419];
     layer3_out[593] <= layer2_out[799];
     layer3_out[594] <= ~layer2_out[99];
     layer3_out[595] <= layer2_out[368];
     layer3_out[596] <= ~layer2_out[173];
     layer3_out[597] <= layer2_out[655];
     layer3_out[598] <= ~(layer2_out[49] | layer2_out[50]);
     layer3_out[599] <= layer2_out[344] | layer2_out[345];
     layer3_out[600] <= 1'b1;
     layer3_out[601] <= ~layer2_out[365] | layer2_out[366];
     layer3_out[602] <= ~(layer2_out[362] | layer2_out[363]);
     layer3_out[603] <= layer2_out[229] & ~layer2_out[230];
     layer3_out[604] <= ~layer2_out[302] | layer2_out[303];
     layer3_out[605] <= ~(layer2_out[525] & layer2_out[526]);
     layer3_out[606] <= layer2_out[387];
     layer3_out[607] <= 1'b1;
     layer3_out[608] <= ~layer2_out[616] | layer2_out[617];
     layer3_out[609] <= ~layer2_out[86] | layer2_out[85];
     layer3_out[610] <= layer2_out[126];
     layer3_out[611] <= layer2_out[182] & ~layer2_out[181];
     layer3_out[612] <= layer2_out[411] | layer2_out[412];
     layer3_out[613] <= ~layer2_out[634];
     layer3_out[614] <= 1'b0;
     layer3_out[615] <= ~layer2_out[618];
     layer3_out[616] <= layer2_out[32] ^ layer2_out[33];
     layer3_out[617] <= layer2_out[473];
     layer3_out[618] <= ~layer2_out[315];
     layer3_out[619] <= ~layer2_out[453];
     layer3_out[620] <= layer2_out[312];
     layer3_out[621] <= ~layer2_out[684] | layer2_out[683];
     layer3_out[622] <= layer2_out[684];
     layer3_out[623] <= ~layer2_out[673];
     layer3_out[624] <= ~layer2_out[189] | layer2_out[188];
     layer3_out[625] <= layer2_out[504];
     layer3_out[626] <= ~(layer2_out[706] & layer2_out[707]);
     layer3_out[627] <= layer2_out[102];
     layer3_out[628] <= ~layer2_out[215];
     layer3_out[629] <= layer2_out[234] ^ layer2_out[235];
     layer3_out[630] <= ~(layer2_out[601] & layer2_out[602]);
     layer3_out[631] <= ~layer2_out[371] | layer2_out[370];
     layer3_out[632] <= ~layer2_out[564];
     layer3_out[633] <= layer2_out[250] & layer2_out[251];
     layer3_out[634] <= ~(layer2_out[405] ^ layer2_out[406]);
     layer3_out[635] <= layer2_out[248] | layer2_out[249];
     layer3_out[636] <= ~layer2_out[331];
     layer3_out[637] <= ~layer2_out[470] | layer2_out[471];
     layer3_out[638] <= ~layer2_out[94] | layer2_out[93];
     layer3_out[639] <= layer2_out[131] & ~layer2_out[132];
     layer3_out[640] <= ~layer2_out[180];
     layer3_out[641] <= ~layer2_out[383];
     layer3_out[642] <= ~layer2_out[772];
     layer3_out[643] <= ~layer2_out[224] | layer2_out[225];
     layer3_out[644] <= layer2_out[328] & ~layer2_out[327];
     layer3_out[645] <= ~layer2_out[4] | layer2_out[3];
     layer3_out[646] <= layer2_out[698] ^ layer2_out[699];
     layer3_out[647] <= ~layer2_out[576];
     layer3_out[648] <= ~(layer2_out[795] ^ layer2_out[796]);
     layer3_out[649] <= ~(layer2_out[763] & layer2_out[764]);
     layer3_out[650] <= layer2_out[388] | layer2_out[389];
     layer3_out[651] <= ~layer2_out[459] | layer2_out[460];
     layer3_out[652] <= layer2_out[195];
     layer3_out[653] <= layer2_out[447] & ~layer2_out[448];
     layer3_out[654] <= layer2_out[215];
     layer3_out[655] <= ~layer2_out[287];
     layer3_out[656] <= layer2_out[391];
     layer3_out[657] <= layer2_out[658];
     layer3_out[658] <= ~layer2_out[82];
     layer3_out[659] <= ~(layer2_out[736] | layer2_out[737]);
     layer3_out[660] <= ~(layer2_out[555] & layer2_out[556]);
     layer3_out[661] <= layer2_out[185] | layer2_out[186];
     layer3_out[662] <= layer2_out[178] & ~layer2_out[179];
     layer3_out[663] <= layer2_out[559];
     layer3_out[664] <= ~layer2_out[598];
     layer3_out[665] <= ~(layer2_out[57] ^ layer2_out[58]);
     layer3_out[666] <= layer2_out[277];
     layer3_out[667] <= ~layer2_out[731];
     layer3_out[668] <= layer2_out[751] & ~layer2_out[750];
     layer3_out[669] <= ~(layer2_out[496] | layer2_out[497]);
     layer3_out[670] <= layer2_out[557] & ~layer2_out[556];
     layer3_out[671] <= 1'b0;
     layer3_out[672] <= layer2_out[754] & ~layer2_out[753];
     layer3_out[673] <= ~layer2_out[241];
     layer3_out[674] <= layer2_out[338];
     layer3_out[675] <= ~layer2_out[63] | layer2_out[62];
     layer3_out[676] <= layer2_out[309] & ~layer2_out[310];
     layer3_out[677] <= layer2_out[619] & ~layer2_out[618];
     layer3_out[678] <= ~layer2_out[183];
     layer3_out[679] <= layer2_out[298];
     layer3_out[680] <= layer2_out[178];
     layer3_out[681] <= ~layer2_out[429];
     layer3_out[682] <= layer2_out[401];
     layer3_out[683] <= ~(layer2_out[731] | layer2_out[732]);
     layer3_out[684] <= layer2_out[289];
     layer3_out[685] <= ~layer2_out[373];
     layer3_out[686] <= ~layer2_out[427];
     layer3_out[687] <= ~layer2_out[486];
     layer3_out[688] <= ~(layer2_out[536] | layer2_out[537]);
     layer3_out[689] <= layer2_out[500];
     layer3_out[690] <= layer2_out[437] & ~layer2_out[438];
     layer3_out[691] <= ~layer2_out[621] | layer2_out[620];
     layer3_out[692] <= layer2_out[693] & ~layer2_out[692];
     layer3_out[693] <= ~(layer2_out[352] | layer2_out[353]);
     layer3_out[694] <= 1'b1;
     layer3_out[695] <= ~layer2_out[184] | layer2_out[183];
     layer3_out[696] <= layer2_out[533] & layer2_out[534];
     layer3_out[697] <= ~layer2_out[562];
     layer3_out[698] <= ~layer2_out[346];
     layer3_out[699] <= layer2_out[312];
     layer3_out[700] <= ~layer2_out[27] | layer2_out[28];
     layer3_out[701] <= layer2_out[419] & ~layer2_out[420];
     layer3_out[702] <= layer2_out[697] | layer2_out[698];
     layer3_out[703] <= ~(layer2_out[232] & layer2_out[233]);
     layer3_out[704] <= layer2_out[105] & ~layer2_out[106];
     layer3_out[705] <= ~(layer2_out[321] | layer2_out[322]);
     layer3_out[706] <= layer2_out[107] & ~layer2_out[106];
     layer3_out[707] <= ~layer2_out[412] | layer2_out[413];
     layer3_out[708] <= layer2_out[7] & ~layer2_out[8];
     layer3_out[709] <= ~(layer2_out[709] | layer2_out[710]);
     layer3_out[710] <= layer2_out[642] & ~layer2_out[643];
     layer3_out[711] <= ~layer2_out[29];
     layer3_out[712] <= ~layer2_out[164];
     layer3_out[713] <= ~layer2_out[626] | layer2_out[625];
     layer3_out[714] <= ~(layer2_out[488] | layer2_out[489]);
     layer3_out[715] <= layer2_out[435];
     layer3_out[716] <= layer2_out[718];
     layer3_out[717] <= ~layer2_out[705] | layer2_out[706];
     layer3_out[718] <= layer2_out[743] & ~layer2_out[742];
     layer3_out[719] <= ~layer2_out[660];
     layer3_out[720] <= ~layer2_out[672];
     layer3_out[721] <= layer2_out[363] | layer2_out[364];
     layer3_out[722] <= layer2_out[479] & ~layer2_out[478];
     layer3_out[723] <= ~layer2_out[724];
     layer3_out[724] <= ~layer2_out[306];
     layer3_out[725] <= ~(layer2_out[466] | layer2_out[467]);
     layer3_out[726] <= layer2_out[144] & ~layer2_out[145];
     layer3_out[727] <= layer2_out[656];
     layer3_out[728] <= ~layer2_out[345];
     layer3_out[729] <= ~(layer2_out[385] ^ layer2_out[386]);
     layer3_out[730] <= ~layer2_out[405];
     layer3_out[731] <= layer2_out[798];
     layer3_out[732] <= layer2_out[450] | layer2_out[451];
     layer3_out[733] <= layer2_out[143];
     layer3_out[734] <= ~layer2_out[393];
     layer3_out[735] <= layer2_out[476] & ~layer2_out[477];
     layer3_out[736] <= ~(layer2_out[765] & layer2_out[766]);
     layer3_out[737] <= ~layer2_out[637];
     layer3_out[738] <= 1'b0;
     layer3_out[739] <= ~layer2_out[65];
     layer3_out[740] <= layer2_out[67] & ~layer2_out[68];
     layer3_out[741] <= layer2_out[486] & ~layer2_out[485];
     layer3_out[742] <= ~layer2_out[361];
     layer3_out[743] <= layer2_out[723] & ~layer2_out[722];
     layer3_out[744] <= layer2_out[128];
     layer3_out[745] <= ~layer2_out[678];
     layer3_out[746] <= ~(layer2_out[104] ^ layer2_out[105]);
     layer3_out[747] <= layer2_out[108] & ~layer2_out[109];
     layer3_out[748] <= ~layer2_out[426];
     layer3_out[749] <= ~layer2_out[137] | layer2_out[138];
     layer3_out[750] <= layer2_out[5] & ~layer2_out[6];
     layer3_out[751] <= layer2_out[117] | layer2_out[118];
     layer3_out[752] <= layer2_out[741] & layer2_out[742];
     layer3_out[753] <= ~layer2_out[775];
     layer3_out[754] <= layer2_out[580];
     layer3_out[755] <= layer2_out[289] & layer2_out[290];
     layer3_out[756] <= layer2_out[300];
     layer3_out[757] <= ~(layer2_out[770] ^ layer2_out[771]);
     layer3_out[758] <= layer2_out[671] | layer2_out[672];
     layer3_out[759] <= ~layer2_out[176];
     layer3_out[760] <= layer2_out[199] & ~layer2_out[200];
     layer3_out[761] <= layer2_out[554] & ~layer2_out[553];
     layer3_out[762] <= ~(layer2_out[675] ^ layer2_out[676]);
     layer3_out[763] <= layer2_out[20];
     layer3_out[764] <= ~layer2_out[18];
     layer3_out[765] <= ~layer2_out[454] | layer2_out[455];
     layer3_out[766] <= ~layer2_out[703];
     layer3_out[767] <= ~(layer2_out[351] | layer2_out[352]);
     layer3_out[768] <= layer2_out[16] ^ layer2_out[17];
     layer3_out[769] <= layer2_out[552];
     layer3_out[770] <= ~layer2_out[716];
     layer3_out[771] <= layer2_out[354] & ~layer2_out[355];
     layer3_out[772] <= layer2_out[747] & layer2_out[748];
     layer3_out[773] <= ~layer2_out[37];
     layer3_out[774] <= layer2_out[424];
     layer3_out[775] <= layer2_out[1] & ~layer2_out[0];
     layer3_out[776] <= layer2_out[542];
     layer3_out[777] <= ~layer2_out[440];
     layer3_out[778] <= layer2_out[551] & ~layer2_out[550];
     layer3_out[779] <= layer2_out[205] | layer2_out[206];
     layer3_out[780] <= ~(layer2_out[77] | layer2_out[78]);
     layer3_out[781] <= layer2_out[76] & layer2_out[77];
     layer3_out[782] <= layer2_out[577] ^ layer2_out[578];
     layer3_out[783] <= layer2_out[727];
     layer3_out[784] <= layer2_out[357] | layer2_out[358];
     layer3_out[785] <= layer2_out[265];
     layer3_out[786] <= ~(layer2_out[175] ^ layer2_out[176]);
     layer3_out[787] <= layer2_out[674];
     layer3_out[788] <= ~(layer2_out[471] & layer2_out[472]);
     layer3_out[789] <= ~layer2_out[261];
     layer3_out[790] <= ~(layer2_out[34] ^ layer2_out[35]);
     layer3_out[791] <= layer2_out[430];
     layer3_out[792] <= ~layer2_out[44];
     layer3_out[793] <= layer2_out[691] | layer2_out[692];
     layer3_out[794] <= layer2_out[649];
     layer3_out[795] <= ~layer2_out[664];
     layer3_out[796] <= layer2_out[750] & ~layer2_out[749];
     layer3_out[797] <= ~layer2_out[763] | layer2_out[762];
     layer3_out[798] <= 1'b1;
     layer3_out[799] <= layer2_out[475];
     layer4_out[0] <= ~(layer3_out[172] & layer3_out[173]);
     layer4_out[1] <= layer3_out[48] & ~layer3_out[47];
     layer4_out[2] <= ~layer3_out[169] | layer3_out[170];
     layer4_out[3] <= ~layer3_out[125];
     layer4_out[4] <= ~layer3_out[76];
     layer4_out[5] <= layer3_out[705];
     layer4_out[6] <= ~layer3_out[117] | layer3_out[116];
     layer4_out[7] <= layer3_out[720] & ~layer3_out[719];
     layer4_out[8] <= ~layer3_out[457] | layer3_out[456];
     layer4_out[9] <= layer3_out[410] & ~layer3_out[411];
     layer4_out[10] <= layer3_out[544] | layer3_out[545];
     layer4_out[11] <= layer3_out[599] & layer3_out[600];
     layer4_out[12] <= layer3_out[529];
     layer4_out[13] <= layer3_out[597] & ~layer3_out[598];
     layer4_out[14] <= 1'b1;
     layer4_out[15] <= ~layer3_out[715];
     layer4_out[16] <= layer3_out[525];
     layer4_out[17] <= layer3_out[91];
     layer4_out[18] <= layer3_out[650] & ~layer3_out[651];
     layer4_out[19] <= ~(layer3_out[373] ^ layer3_out[374]);
     layer4_out[20] <= ~(layer3_out[356] ^ layer3_out[357]);
     layer4_out[21] <= layer3_out[339] & ~layer3_out[338];
     layer4_out[22] <= layer3_out[235];
     layer4_out[23] <= layer3_out[12] ^ layer3_out[13];
     layer4_out[24] <= layer3_out[607] | layer3_out[608];
     layer4_out[25] <= ~layer3_out[250] | layer3_out[249];
     layer4_out[26] <= layer3_out[185];
     layer4_out[27] <= layer3_out[757] ^ layer3_out[758];
     layer4_out[28] <= ~layer3_out[172] | layer3_out[171];
     layer4_out[29] <= ~layer3_out[466] | layer3_out[465];
     layer4_out[30] <= ~layer3_out[390];
     layer4_out[31] <= ~layer3_out[409];
     layer4_out[32] <= ~layer3_out[409];
     layer4_out[33] <= ~layer3_out[540];
     layer4_out[34] <= layer3_out[338];
     layer4_out[35] <= layer3_out[684];
     layer4_out[36] <= layer3_out[368] ^ layer3_out[369];
     layer4_out[37] <= ~layer3_out[330] | layer3_out[331];
     layer4_out[38] <= layer3_out[770];
     layer4_out[39] <= ~layer3_out[300];
     layer4_out[40] <= ~layer3_out[246] | layer3_out[245];
     layer4_out[41] <= layer3_out[711];
     layer4_out[42] <= layer3_out[278] & layer3_out[279];
     layer4_out[43] <= ~layer3_out[290];
     layer4_out[44] <= layer3_out[403];
     layer4_out[45] <= layer3_out[693] & ~layer3_out[692];
     layer4_out[46] <= layer3_out[507] | layer3_out[508];
     layer4_out[47] <= layer3_out[659];
     layer4_out[48] <= ~layer3_out[542] | layer3_out[541];
     layer4_out[49] <= ~layer3_out[433] | layer3_out[432];
     layer4_out[50] <= ~layer3_out[570];
     layer4_out[51] <= layer3_out[70];
     layer4_out[52] <= ~layer3_out[648] | layer3_out[647];
     layer4_out[53] <= ~layer3_out[136] | layer3_out[137];
     layer4_out[54] <= ~layer3_out[199];
     layer4_out[55] <= layer3_out[138] & ~layer3_out[139];
     layer4_out[56] <= layer3_out[351];
     layer4_out[57] <= layer3_out[458];
     layer4_out[58] <= layer3_out[61] | layer3_out[62];
     layer4_out[59] <= ~(layer3_out[9] ^ layer3_out[10]);
     layer4_out[60] <= layer3_out[507];
     layer4_out[61] <= ~layer3_out[559];
     layer4_out[62] <= layer3_out[402] & ~layer3_out[401];
     layer4_out[63] <= ~layer3_out[268];
     layer4_out[64] <= layer3_out[761] & ~layer3_out[760];
     layer4_out[65] <= ~(layer3_out[272] | layer3_out[273]);
     layer4_out[66] <= layer3_out[315] & layer3_out[316];
     layer4_out[67] <= 1'b1;
     layer4_out[68] <= layer3_out[567];
     layer4_out[69] <= layer3_out[424];
     layer4_out[70] <= layer3_out[202];
     layer4_out[71] <= ~layer3_out[105];
     layer4_out[72] <= layer3_out[550];
     layer4_out[73] <= ~layer3_out[605];
     layer4_out[74] <= layer3_out[288];
     layer4_out[75] <= layer3_out[779];
     layer4_out[76] <= layer3_out[752];
     layer4_out[77] <= ~layer3_out[333];
     layer4_out[78] <= layer3_out[366] & ~layer3_out[365];
     layer4_out[79] <= ~layer3_out[451];
     layer4_out[80] <= layer3_out[439];
     layer4_out[81] <= ~layer3_out[238] | layer3_out[237];
     layer4_out[82] <= ~(layer3_out[154] | layer3_out[155]);
     layer4_out[83] <= layer3_out[579] & ~layer3_out[578];
     layer4_out[84] <= ~(layer3_out[319] ^ layer3_out[320]);
     layer4_out[85] <= layer3_out[52] & ~layer3_out[51];
     layer4_out[86] <= ~layer3_out[193] | layer3_out[194];
     layer4_out[87] <= ~layer3_out[96];
     layer4_out[88] <= layer3_out[677] | layer3_out[678];
     layer4_out[89] <= layer3_out[588] & ~layer3_out[587];
     layer4_out[90] <= layer3_out[472] | layer3_out[473];
     layer4_out[91] <= ~layer3_out[648];
     layer4_out[92] <= layer3_out[380];
     layer4_out[93] <= ~layer3_out[424];
     layer4_out[94] <= ~layer3_out[762];
     layer4_out[95] <= ~layer3_out[695] | layer3_out[696];
     layer4_out[96] <= ~layer3_out[669];
     layer4_out[97] <= layer3_out[155] ^ layer3_out[156];
     layer4_out[98] <= ~layer3_out[224];
     layer4_out[99] <= ~(layer3_out[685] & layer3_out[686]);
     layer4_out[100] <= ~(layer3_out[735] & layer3_out[736]);
     layer4_out[101] <= ~layer3_out[394] | layer3_out[393];
     layer4_out[102] <= ~layer3_out[455];
     layer4_out[103] <= layer3_out[577];
     layer4_out[104] <= layer3_out[641];
     layer4_out[105] <= ~layer3_out[128] | layer3_out[127];
     layer4_out[106] <= ~layer3_out[737];
     layer4_out[107] <= layer3_out[264] | layer3_out[265];
     layer4_out[108] <= ~layer3_out[66];
     layer4_out[109] <= layer3_out[382] & layer3_out[383];
     layer4_out[110] <= ~(layer3_out[391] ^ layer3_out[392]);
     layer4_out[111] <= ~layer3_out[655];
     layer4_out[112] <= layer3_out[41];
     layer4_out[113] <= ~(layer3_out[97] | layer3_out[98]);
     layer4_out[114] <= ~layer3_out[788];
     layer4_out[115] <= ~layer3_out[88];
     layer4_out[116] <= ~layer3_out[18];
     layer4_out[117] <= layer3_out[11] & ~layer3_out[10];
     layer4_out[118] <= ~layer3_out[166];
     layer4_out[119] <= ~layer3_out[640] | layer3_out[641];
     layer4_out[120] <= ~layer3_out[335];
     layer4_out[121] <= ~layer3_out[297];
     layer4_out[122] <= layer3_out[676] & layer3_out[677];
     layer4_out[123] <= layer3_out[100];
     layer4_out[124] <= layer3_out[442];
     layer4_out[125] <= layer3_out[561] ^ layer3_out[562];
     layer4_out[126] <= layer3_out[76];
     layer4_out[127] <= ~layer3_out[151] | layer3_out[152];
     layer4_out[128] <= ~layer3_out[252];
     layer4_out[129] <= layer3_out[108] & layer3_out[109];
     layer4_out[130] <= layer3_out[49] & ~layer3_out[48];
     layer4_out[131] <= ~layer3_out[433];
     layer4_out[132] <= layer3_out[443];
     layer4_out[133] <= ~(layer3_out[379] & layer3_out[380]);
     layer4_out[134] <= layer3_out[296] & ~layer3_out[295];
     layer4_out[135] <= layer3_out[769];
     layer4_out[136] <= layer3_out[541] & ~layer3_out[540];
     layer4_out[137] <= layer3_out[43] | layer3_out[44];
     layer4_out[138] <= layer3_out[258] & ~layer3_out[257];
     layer4_out[139] <= layer3_out[791] | layer3_out[792];
     layer4_out[140] <= layer3_out[18] & layer3_out[19];
     layer4_out[141] <= layer3_out[516] & ~layer3_out[515];
     layer4_out[142] <= layer3_out[50];
     layer4_out[143] <= layer3_out[646];
     layer4_out[144] <= ~layer3_out[698];
     layer4_out[145] <= ~layer3_out[558];
     layer4_out[146] <= ~layer3_out[69];
     layer4_out[147] <= ~(layer3_out[81] | layer3_out[82]);
     layer4_out[148] <= layer3_out[483];
     layer4_out[149] <= layer3_out[13] & ~layer3_out[14];
     layer4_out[150] <= ~layer3_out[498];
     layer4_out[151] <= ~(layer3_out[8] ^ layer3_out[9]);
     layer4_out[152] <= ~(layer3_out[709] & layer3_out[710]);
     layer4_out[153] <= ~layer3_out[565] | layer3_out[566];
     layer4_out[154] <= ~layer3_out[396];
     layer4_out[155] <= ~layer3_out[680] | layer3_out[679];
     layer4_out[156] <= layer3_out[107] & layer3_out[108];
     layer4_out[157] <= layer3_out[492];
     layer4_out[158] <= ~layer3_out[785];
     layer4_out[159] <= layer3_out[463] & ~layer3_out[462];
     layer4_out[160] <= layer3_out[232];
     layer4_out[161] <= layer3_out[487] & ~layer3_out[488];
     layer4_out[162] <= ~(layer3_out[202] | layer3_out[203]);
     layer4_out[163] <= layer3_out[482];
     layer4_out[164] <= ~(layer3_out[415] ^ layer3_out[416]);
     layer4_out[165] <= layer3_out[235] | layer3_out[236];
     layer4_out[166] <= ~(layer3_out[233] ^ layer3_out[234]);
     layer4_out[167] <= layer3_out[626];
     layer4_out[168] <= layer3_out[702] & layer3_out[703];
     layer4_out[169] <= ~layer3_out[449];
     layer4_out[170] <= layer3_out[66];
     layer4_out[171] <= layer3_out[635];
     layer4_out[172] <= layer3_out[478] & ~layer3_out[477];
     layer4_out[173] <= ~(layer3_out[693] | layer3_out[694]);
     layer4_out[174] <= ~layer3_out[506] | layer3_out[505];
     layer4_out[175] <= ~layer3_out[388] | layer3_out[389];
     layer4_out[176] <= ~layer3_out[220];
     layer4_out[177] <= layer3_out[666] & layer3_out[667];
     layer4_out[178] <= layer3_out[216];
     layer4_out[179] <= ~(layer3_out[187] & layer3_out[188]);
     layer4_out[180] <= ~layer3_out[763];
     layer4_out[181] <= ~layer3_out[721] | layer3_out[720];
     layer4_out[182] <= ~layer3_out[179] | layer3_out[180];
     layer4_out[183] <= ~layer3_out[495];
     layer4_out[184] <= ~layer3_out[732] | layer3_out[733];
     layer4_out[185] <= layer3_out[95] | layer3_out[96];
     layer4_out[186] <= ~layer3_out[162] | layer3_out[161];
     layer4_out[187] <= layer3_out[652];
     layer4_out[188] <= ~layer3_out[557] | layer3_out[558];
     layer4_out[189] <= ~layer3_out[728] | layer3_out[727];
     layer4_out[190] <= layer3_out[364];
     layer4_out[191] <= ~(layer3_out[521] & layer3_out[522]);
     layer4_out[192] <= layer3_out[267];
     layer4_out[193] <= ~layer3_out[660] | layer3_out[661];
     layer4_out[194] <= layer3_out[89] & layer3_out[90];
     layer4_out[195] <= ~layer3_out[675] | layer3_out[676];
     layer4_out[196] <= ~layer3_out[28];
     layer4_out[197] <= layer3_out[535];
     layer4_out[198] <= layer3_out[397] | layer3_out[398];
     layer4_out[199] <= ~layer3_out[204] | layer3_out[205];
     layer4_out[200] <= ~(layer3_out[113] | layer3_out[114]);
     layer4_out[201] <= layer3_out[372] ^ layer3_out[373];
     layer4_out[202] <= layer3_out[186];
     layer4_out[203] <= ~(layer3_out[215] & layer3_out[216]);
     layer4_out[204] <= layer3_out[691];
     layer4_out[205] <= ~(layer3_out[74] | layer3_out[75]);
     layer4_out[206] <= layer3_out[8] & ~layer3_out[7];
     layer4_out[207] <= ~layer3_out[565];
     layer4_out[208] <= ~layer3_out[59];
     layer4_out[209] <= layer3_out[196] & layer3_out[197];
     layer4_out[210] <= 1'b1;
     layer4_out[211] <= layer3_out[758];
     layer4_out[212] <= ~layer3_out[798] | layer3_out[797];
     layer4_out[213] <= layer3_out[242];
     layer4_out[214] <= layer3_out[137] ^ layer3_out[138];
     layer4_out[215] <= ~layer3_out[644];
     layer4_out[216] <= ~(layer3_out[150] | layer3_out[151]);
     layer4_out[217] <= layer3_out[671] & ~layer3_out[672];
     layer4_out[218] <= ~layer3_out[23] | layer3_out[24];
     layer4_out[219] <= ~(layer3_out[134] ^ layer3_out[135]);
     layer4_out[220] <= layer3_out[406] | layer3_out[407];
     layer4_out[221] <= ~layer3_out[86] | layer3_out[85];
     layer4_out[222] <= ~layer3_out[482];
     layer4_out[223] <= ~layer3_out[303];
     layer4_out[224] <= layer3_out[126];
     layer4_out[225] <= layer3_out[119];
     layer4_out[226] <= ~layer3_out[745];
     layer4_out[227] <= ~layer3_out[230] | layer3_out[231];
     layer4_out[228] <= ~layer3_out[639] | layer3_out[638];
     layer4_out[229] <= ~layer3_out[160];
     layer4_out[230] <= ~(layer3_out[706] | layer3_out[707]);
     layer4_out[231] <= ~(layer3_out[681] ^ layer3_out[682]);
     layer4_out[232] <= layer3_out[596];
     layer4_out[233] <= ~layer3_out[469] | layer3_out[470];
     layer4_out[234] <= ~layer3_out[749];
     layer4_out[235] <= ~layer3_out[377];
     layer4_out[236] <= layer3_out[54];
     layer4_out[237] <= ~layer3_out[326];
     layer4_out[238] <= ~layer3_out[174] | layer3_out[175];
     layer4_out[239] <= layer3_out[582] ^ layer3_out[583];
     layer4_out[240] <= layer3_out[430] & ~layer3_out[429];
     layer4_out[241] <= 1'b1;
     layer4_out[242] <= layer3_out[333] & ~layer3_out[332];
     layer4_out[243] <= ~layer3_out[575];
     layer4_out[244] <= layer3_out[385] | layer3_out[386];
     layer4_out[245] <= ~layer3_out[157];
     layer4_out[246] <= layer3_out[688] & ~layer3_out[687];
     layer4_out[247] <= ~layer3_out[213];
     layer4_out[248] <= layer3_out[519] & layer3_out[520];
     layer4_out[249] <= layer3_out[751] & ~layer3_out[752];
     layer4_out[250] <= layer3_out[227];
     layer4_out[251] <= ~layer3_out[405];
     layer4_out[252] <= layer3_out[207] | layer3_out[208];
     layer4_out[253] <= ~(layer3_out[46] | layer3_out[47]);
     layer4_out[254] <= ~layer3_out[498];
     layer4_out[255] <= layer3_out[84] | layer3_out[85];
     layer4_out[256] <= ~layer3_out[349] | layer3_out[350];
     layer4_out[257] <= layer3_out[357];
     layer4_out[258] <= ~(layer3_out[523] & layer3_out[524]);
     layer4_out[259] <= ~(layer3_out[471] & layer3_out[472]);
     layer4_out[260] <= ~(layer3_out[77] & layer3_out[78]);
     layer4_out[261] <= layer3_out[443] | layer3_out[444];
     layer4_out[262] <= layer3_out[738];
     layer4_out[263] <= ~layer3_out[301] | layer3_out[300];
     layer4_out[264] <= layer3_out[239] & ~layer3_out[240];
     layer4_out[265] <= ~layer3_out[765];
     layer4_out[266] <= layer3_out[612] & ~layer3_out[613];
     layer4_out[267] <= layer3_out[328] & layer3_out[329];
     layer4_out[268] <= layer3_out[730];
     layer4_out[269] <= layer3_out[727] & ~layer3_out[726];
     layer4_out[270] <= layer3_out[718];
     layer4_out[271] <= ~layer3_out[749];
     layer4_out[272] <= layer3_out[690] & ~layer3_out[691];
     layer4_out[273] <= layer3_out[586];
     layer4_out[274] <= ~layer3_out[448] | layer3_out[447];
     layer4_out[275] <= layer3_out[148];
     layer4_out[276] <= layer3_out[273] | layer3_out[274];
     layer4_out[277] <= layer3_out[501] & ~layer3_out[502];
     layer4_out[278] <= ~layer3_out[619];
     layer4_out[279] <= ~layer3_out[683];
     layer4_out[280] <= layer3_out[624] | layer3_out[625];
     layer4_out[281] <= layer3_out[348];
     layer4_out[282] <= ~layer3_out[742];
     layer4_out[283] <= ~layer3_out[15] | layer3_out[16];
     layer4_out[284] <= layer3_out[622];
     layer4_out[285] <= layer3_out[365];
     layer4_out[286] <= layer3_out[67];
     layer4_out[287] <= ~layer3_out[84];
     layer4_out[288] <= layer3_out[34] & ~layer3_out[35];
     layer4_out[289] <= layer3_out[470] & ~layer3_out[471];
     layer4_out[290] <= layer3_out[299] & ~layer3_out[298];
     layer4_out[291] <= ~layer3_out[401];
     layer4_out[292] <= layer3_out[628] | layer3_out[629];
     layer4_out[293] <= layer3_out[304] | layer3_out[305];
     layer4_out[294] <= ~layer3_out[176];
     layer4_out[295] <= layer3_out[139];
     layer4_out[296] <= ~layer3_out[466];
     layer4_out[297] <= ~layer3_out[746];
     layer4_out[298] <= ~layer3_out[675];
     layer4_out[299] <= ~(layer3_out[0] & layer3_out[1]);
     layer4_out[300] <= ~(layer3_out[344] ^ layer3_out[345]);
     layer4_out[301] <= layer3_out[514];
     layer4_out[302] <= ~layer3_out[491];
     layer4_out[303] <= layer3_out[53];
     layer4_out[304] <= layer3_out[493] & layer3_out[494];
     layer4_out[305] <= layer3_out[614] ^ layer3_out[615];
     layer4_out[306] <= ~layer3_out[593];
     layer4_out[307] <= layer3_out[790];
     layer4_out[308] <= layer3_out[522];
     layer4_out[309] <= ~layer3_out[311];
     layer4_out[310] <= ~layer3_out[423];
     layer4_out[311] <= layer3_out[110];
     layer4_out[312] <= ~(layer3_out[238] | layer3_out[239]);
     layer4_out[313] <= ~layer3_out[687];
     layer4_out[314] <= layer3_out[42];
     layer4_out[315] <= layer3_out[634];
     layer4_out[316] <= ~(layer3_out[623] | layer3_out[624]);
     layer4_out[317] <= layer3_out[64];
     layer4_out[318] <= layer3_out[40] & layer3_out[41];
     layer4_out[319] <= layer3_out[225] & layer3_out[226];
     layer4_out[320] <= ~(layer3_out[667] ^ layer3_out[668]);
     layer4_out[321] <= layer3_out[170] & layer3_out[171];
     layer4_out[322] <= ~(layer3_out[189] & layer3_out[190]);
     layer4_out[323] <= layer3_out[457] & ~layer3_out[458];
     layer4_out[324] <= layer3_out[710];
     layer4_out[325] <= layer3_out[735];
     layer4_out[326] <= 1'b0;
     layer4_out[327] <= ~layer3_out[288];
     layer4_out[328] <= 1'b0;
     layer4_out[329] <= layer3_out[217];
     layer4_out[330] <= ~(layer3_out[445] & layer3_out[446]);
     layer4_out[331] <= layer3_out[761] & ~layer3_out[762];
     layer4_out[332] <= ~layer3_out[142];
     layer4_out[333] <= ~(layer3_out[637] | layer3_out[638]);
     layer4_out[334] <= ~layer3_out[123];
     layer4_out[335] <= layer3_out[78] & ~layer3_out[79];
     layer4_out[336] <= ~layer3_out[293];
     layer4_out[337] <= layer3_out[511] & ~layer3_out[512];
     layer4_out[338] <= ~layer3_out[447] | layer3_out[446];
     layer4_out[339] <= layer3_out[243] | layer3_out[244];
     layer4_out[340] <= layer3_out[32];
     layer4_out[341] <= layer3_out[37] | layer3_out[38];
     layer4_out[342] <= layer3_out[645];
     layer4_out[343] <= layer3_out[132] | layer3_out[133];
     layer4_out[344] <= layer3_out[550] & ~layer3_out[549];
     layer4_out[345] <= ~layer3_out[484];
     layer4_out[346] <= ~layer3_out[526];
     layer4_out[347] <= ~(layer3_out[383] & layer3_out[384]);
     layer4_out[348] <= ~(layer3_out[503] & layer3_out[504]);
     layer4_out[349] <= ~(layer3_out[377] & layer3_out[378]);
     layer4_out[350] <= ~layer3_out[141] | layer3_out[140];
     layer4_out[351] <= layer3_out[398] | layer3_out[399];
     layer4_out[352] <= ~layer3_out[223];
     layer4_out[353] <= ~layer3_out[147];
     layer4_out[354] <= ~layer3_out[313] | layer3_out[314];
     layer4_out[355] <= layer3_out[210];
     layer4_out[356] <= layer3_out[33];
     layer4_out[357] <= ~(layer3_out[212] ^ layer3_out[213]);
     layer4_out[358] <= 1'b0;
     layer4_out[359] <= ~layer3_out[253] | layer3_out[254];
     layer4_out[360] <= ~layer3_out[1];
     layer4_out[361] <= layer3_out[616];
     layer4_out[362] <= ~layer3_out[248];
     layer4_out[363] <= layer3_out[31] & ~layer3_out[30];
     layer4_out[364] <= ~layer3_out[121] | layer3_out[120];
     layer4_out[365] <= layer3_out[390] & ~layer3_out[391];
     layer4_out[366] <= ~(layer3_out[743] ^ layer3_out[744]);
     layer4_out[367] <= layer3_out[387];
     layer4_out[368] <= ~layer3_out[0] | layer3_out[2];
     layer4_out[369] <= layer3_out[6] & layer3_out[7];
     layer4_out[370] <= ~layer3_out[26];
     layer4_out[371] <= ~(layer3_out[369] & layer3_out[370]);
     layer4_out[372] <= layer3_out[293] & ~layer3_out[292];
     layer4_out[373] <= layer3_out[787] & ~layer3_out[788];
     layer4_out[374] <= layer3_out[367];
     layer4_out[375] <= layer3_out[347];
     layer4_out[376] <= layer3_out[591] & ~layer3_out[590];
     layer4_out[377] <= layer3_out[755] & layer3_out[756];
     layer4_out[378] <= layer3_out[57];
     layer4_out[379] <= layer3_out[512];
     layer4_out[380] <= layer3_out[26] | layer3_out[27];
     layer4_out[381] <= ~layer3_out[564] | layer3_out[563];
     layer4_out[382] <= ~layer3_out[396] | layer3_out[397];
     layer4_out[383] <= ~(layer3_out[717] | layer3_out[718]);
     layer4_out[384] <= ~(layer3_out[489] ^ layer3_out[490]);
     layer4_out[385] <= layer3_out[104];
     layer4_out[386] <= ~(layer3_out[262] ^ layer3_out[263]);
     layer4_out[387] <= ~layer3_out[613];
     layer4_out[388] <= layer3_out[464];
     layer4_out[389] <= layer3_out[269] | layer3_out[270];
     layer4_out[390] <= layer3_out[554] & ~layer3_out[553];
     layer4_out[391] <= ~layer3_out[5];
     layer4_out[392] <= layer3_out[476] & ~layer3_out[477];
     layer4_out[393] <= ~layer3_out[610];
     layer4_out[394] <= layer3_out[602];
     layer4_out[395] <= layer3_out[376];
     layer4_out[396] <= layer3_out[370] & layer3_out[371];
     layer4_out[397] <= ~(layer3_out[316] ^ layer3_out[317]);
     layer4_out[398] <= ~(layer3_out[780] | layer3_out[781]);
     layer4_out[399] <= ~layer3_out[255];
     layer4_out[400] <= layer3_out[662];
     layer4_out[401] <= layer3_out[414] & ~layer3_out[415];
     layer4_out[402] <= layer3_out[799];
     layer4_out[403] <= layer3_out[781];
     layer4_out[404] <= ~(layer3_out[620] ^ layer3_out[621]);
     layer4_out[405] <= layer3_out[236] & ~layer3_out[237];
     layer4_out[406] <= layer3_out[437] | layer3_out[438];
     layer4_out[407] <= layer3_out[55];
     layer4_out[408] <= layer3_out[580] & layer3_out[581];
     layer4_out[409] <= layer3_out[784];
     layer4_out[410] <= ~layer3_out[707] | layer3_out[708];
     layer4_out[411] <= layer3_out[5] & ~layer3_out[4];
     layer4_out[412] <= layer3_out[562] & layer3_out[563];
     layer4_out[413] <= ~(layer3_out[615] ^ layer3_out[616]);
     layer4_out[414] <= ~layer3_out[537];
     layer4_out[415] <= layer3_out[420] & ~layer3_out[421];
     layer4_out[416] <= ~layer3_out[596];
     layer4_out[417] <= layer3_out[360] & layer3_out[361];
     layer4_out[418] <= ~layer3_out[36];
     layer4_out[419] <= layer3_out[295] & ~layer3_out[294];
     layer4_out[420] <= layer3_out[678] | layer3_out[679];
     layer4_out[421] <= ~layer3_out[438];
     layer4_out[422] <= layer3_out[308];
     layer4_out[423] <= ~layer3_out[627];
     layer4_out[424] <= layer3_out[259] & ~layer3_out[260];
     layer4_out[425] <= ~layer3_out[307] | layer3_out[306];
     layer4_out[426] <= ~(layer3_out[123] & layer3_out[124]);
     layer4_out[427] <= layer3_out[310];
     layer4_out[428] <= layer3_out[747] | layer3_out[748];
     layer4_out[429] <= layer3_out[533] & layer3_out[534];
     layer4_out[430] <= layer3_out[422] & ~layer3_out[421];
     layer4_out[431] <= layer3_out[361] & ~layer3_out[362];
     layer4_out[432] <= layer3_out[567];
     layer4_out[433] <= layer3_out[59] & layer3_out[60];
     layer4_out[434] <= ~layer3_out[342];
     layer4_out[435] <= ~(layer3_out[750] | layer3_out[751]);
     layer4_out[436] <= layer3_out[716];
     layer4_out[437] <= ~layer3_out[796];
     layer4_out[438] <= layer3_out[164];
     layer4_out[439] <= layer3_out[82];
     layer4_out[440] <= layer3_out[111];
     layer4_out[441] <= ~layer3_out[785] | layer3_out[786];
     layer4_out[442] <= ~layer3_out[599];
     layer4_out[443] <= layer3_out[335] & layer3_out[336];
     layer4_out[444] <= layer3_out[731] & layer3_out[732];
     layer4_out[445] <= ~layer3_out[372] | layer3_out[371];
     layer4_out[446] <= ~layer3_out[793];
     layer4_out[447] <= ~(layer3_out[571] ^ layer3_out[572]);
     layer4_out[448] <= layer3_out[36] & ~layer3_out[37];
     layer4_out[449] <= ~layer3_out[496];
     layer4_out[450] <= layer3_out[608];
     layer4_out[451] <= ~(layer3_out[341] ^ layer3_out[342]);
     layer4_out[452] <= ~(layer3_out[551] ^ layer3_out[552]);
     layer4_out[453] <= layer3_out[353] | layer3_out[354];
     layer4_out[454] <= layer3_out[50] | layer3_out[51];
     layer4_out[455] <= layer3_out[362];
     layer4_out[456] <= ~layer3_out[128];
     layer4_out[457] <= ~layer3_out[129];
     layer4_out[458] <= layer3_out[430] & ~layer3_out[431];
     layer4_out[459] <= ~layer3_out[244] | layer3_out[245];
     layer4_out[460] <= ~layer3_out[168];
     layer4_out[461] <= layer3_out[452];
     layer4_out[462] <= layer3_out[429];
     layer4_out[463] <= ~layer3_out[291];
     layer4_out[464] <= layer3_out[115];
     layer4_out[465] <= layer3_out[159];
     layer4_out[466] <= layer3_out[73] & layer3_out[74];
     layer4_out[467] <= 1'b0;
     layer4_out[468] <= ~(layer3_out[80] & layer3_out[81]);
     layer4_out[469] <= layer3_out[585] & ~layer3_out[584];
     layer4_out[470] <= ~layer3_out[662] | layer3_out[661];
     layer4_out[471] <= layer3_out[280];
     layer4_out[472] <= ~layer3_out[713];
     layer4_out[473] <= layer3_out[464];
     layer4_out[474] <= ~layer3_out[532] | layer3_out[533];
     layer4_out[475] <= ~layer3_out[279] | layer3_out[280];
     layer4_out[476] <= layer3_out[453] | layer3_out[454];
     layer4_out[477] <= ~layer3_out[55];
     layer4_out[478] <= layer3_out[122];
     layer4_out[479] <= ~layer3_out[515];
     layer4_out[480] <= layer3_out[723] | layer3_out[724];
     layer4_out[481] <= layer3_out[406];
     layer4_out[482] <= layer3_out[530] & ~layer3_out[529];
     layer4_out[483] <= 1'b0;
     layer4_out[484] <= layer3_out[143] & ~layer3_out[144];
     layer4_out[485] <= layer3_out[434];
     layer4_out[486] <= ~layer3_out[271];
     layer4_out[487] <= layer3_out[14] & ~layer3_out[15];
     layer4_out[488] <= layer3_out[324];
     layer4_out[489] <= layer3_out[152] & layer3_out[153];
     layer4_out[490] <= ~(layer3_out[270] ^ layer3_out[271]);
     layer4_out[491] <= layer3_out[210];
     layer4_out[492] <= ~(layer3_out[777] | layer3_out[778]);
     layer4_out[493] <= ~(layer3_out[91] ^ layer3_out[92]);
     layer4_out[494] <= layer3_out[322] | layer3_out[323];
     layer4_out[495] <= layer3_out[699] & ~layer3_out[700];
     layer4_out[496] <= layer3_out[787];
     layer4_out[497] <= ~layer3_out[142];
     layer4_out[498] <= layer3_out[601];
     layer4_out[499] <= layer3_out[181];
     layer4_out[500] <= ~layer3_out[264] | layer3_out[263];
     layer4_out[501] <= layer3_out[45] ^ layer3_out[46];
     layer4_out[502] <= layer3_out[612] & ~layer3_out[611];
     layer4_out[503] <= layer3_out[632];
     layer4_out[504] <= ~layer3_out[62] | layer3_out[63];
     layer4_out[505] <= ~layer3_out[754];
     layer4_out[506] <= ~layer3_out[149] | layer3_out[150];
     layer4_out[507] <= layer3_out[183] ^ layer3_out[184];
     layer4_out[508] <= layer3_out[22];
     layer4_out[509] <= layer3_out[250];
     layer4_out[510] <= 1'b1;
     layer4_out[511] <= ~layer3_out[568] | layer3_out[569];
     layer4_out[512] <= ~(layer3_out[560] ^ layer3_out[561]);
     layer4_out[513] <= ~(layer3_out[486] ^ layer3_out[487]);
     layer4_out[514] <= ~layer3_out[407];
     layer4_out[515] <= 1'b1;
     layer4_out[516] <= ~(layer3_out[175] ^ layer3_out[176]);
     layer4_out[517] <= layer3_out[556] & ~layer3_out[557];
     layer4_out[518] <= ~layer3_out[469] | layer3_out[468];
     layer4_out[519] <= layer3_out[723];
     layer4_out[520] <= ~(layer3_out[29] | layer3_out[30]);
     layer4_out[521] <= ~layer3_out[531];
     layer4_out[522] <= ~layer3_out[311] | layer3_out[312];
     layer4_out[523] <= layer3_out[223] & ~layer3_out[224];
     layer4_out[524] <= layer3_out[663] & layer3_out[664];
     layer4_out[525] <= ~layer3_out[546] | layer3_out[545];
     layer4_out[526] <= ~layer3_out[113];
     layer4_out[527] <= layer3_out[403];
     layer4_out[528] <= layer3_out[282] ^ layer3_out[283];
     layer4_out[529] <= ~layer3_out[572];
     layer4_out[530] <= layer3_out[291];
     layer4_out[531] <= ~layer3_out[534];
     layer4_out[532] <= layer3_out[592];
     layer4_out[533] <= layer3_out[427] & layer3_out[428];
     layer4_out[534] <= layer3_out[520];
     layer4_out[535] <= layer3_out[502];
     layer4_out[536] <= layer3_out[605];
     layer4_out[537] <= ~layer3_out[330];
     layer4_out[538] <= ~layer3_out[592];
     layer4_out[539] <= ~layer3_out[449] | layer3_out[450];
     layer4_out[540] <= layer3_out[585] & ~layer3_out[586];
     layer4_out[541] <= ~layer3_out[629];
     layer4_out[542] <= layer3_out[548];
     layer4_out[543] <= layer3_out[636] & ~layer3_out[637];
     layer4_out[544] <= ~layer3_out[722];
     layer4_out[545] <= 1'b0;
     layer4_out[546] <= layer3_out[287];
     layer4_out[547] <= layer3_out[724] & layer3_out[725];
     layer4_out[548] <= layer3_out[136] & ~layer3_out[135];
     layer4_out[549] <= ~layer3_out[119];
     layer4_out[550] <= layer3_out[701];
     layer4_out[551] <= layer3_out[57];
     layer4_out[552] <= layer3_out[343] & layer3_out[344];
     layer4_out[553] <= ~layer3_out[669];
     layer4_out[554] <= ~layer3_out[411];
     layer4_out[555] <= ~layer3_out[495];
     layer4_out[556] <= layer3_out[72] & ~layer3_out[73];
     layer4_out[557] <= ~layer3_out[386] | layer3_out[387];
     layer4_out[558] <= ~layer3_out[451];
     layer4_out[559] <= layer3_out[793];
     layer4_out[560] <= ~layer3_out[777];
     layer4_out[561] <= layer3_out[286] & ~layer3_out[285];
     layer4_out[562] <= ~layer3_out[374];
     layer4_out[563] <= layer3_out[791];
     layer4_out[564] <= ~layer3_out[606] | layer3_out[607];
     layer4_out[565] <= layer3_out[783];
     layer4_out[566] <= ~(layer3_out[60] ^ layer3_out[61]);
     layer4_out[567] <= layer3_out[341];
     layer4_out[568] <= layer3_out[670] & ~layer3_out[671];
     layer4_out[569] <= ~layer3_out[588] | layer3_out[589];
     layer4_out[570] <= ~(layer3_out[323] ^ layer3_out[324]);
     layer4_out[571] <= layer3_out[247];
     layer4_out[572] <= layer3_out[28];
     layer4_out[573] <= layer3_out[536] | layer3_out[537];
     layer4_out[574] <= ~(layer3_out[416] & layer3_out[417]);
     layer4_out[575] <= layer3_out[459];
     layer4_out[576] <= layer3_out[603] | layer3_out[604];
     layer4_out[577] <= layer3_out[167] ^ layer3_out[168];
     layer4_out[578] <= layer3_out[547];
     layer4_out[579] <= layer3_out[656] | layer3_out[657];
     layer4_out[580] <= layer3_out[418] | layer3_out[419];
     layer4_out[581] <= ~layer3_out[88];
     layer4_out[582] <= ~(layer3_out[131] & layer3_out[132]);
     layer4_out[583] <= ~layer3_out[740] | layer3_out[739];
     layer4_out[584] <= layer3_out[105];
     layer4_out[585] <= ~layer3_out[544];
     layer4_out[586] <= ~(layer3_out[575] | layer3_out[576]);
     layer4_out[587] <= ~(layer3_out[665] | layer3_out[666]);
     layer4_out[588] <= layer3_out[552];
     layer4_out[589] <= layer3_out[188];
     layer4_out[590] <= layer3_out[16];
     layer4_out[591] <= layer3_out[117] & layer3_out[118];
     layer4_out[592] <= layer3_out[218] ^ layer3_out[219];
     layer4_out[593] <= layer3_out[229] & layer3_out[230];
     layer4_out[594] <= layer3_out[728];
     layer4_out[595] <= layer3_out[425] & ~layer3_out[426];
     layer4_out[596] <= ~layer3_out[277];
     layer4_out[597] <= layer3_out[4];
     layer4_out[598] <= layer3_out[145];
     layer4_out[599] <= ~layer3_out[742];
     layer4_out[600] <= ~layer3_out[261] | layer3_out[260];
     layer4_out[601] <= ~layer3_out[526] | layer3_out[525];
     layer4_out[602] <= ~layer3_out[80];
     layer4_out[603] <= ~layer3_out[426];
     layer4_out[604] <= ~layer3_out[685] | layer3_out[684];
     layer4_out[605] <= layer3_out[716];
     layer4_out[606] <= ~layer3_out[259];
     layer4_out[607] <= layer3_out[160];
     layer4_out[608] <= ~layer3_out[418];
     layer4_out[609] <= ~layer3_out[165] | layer3_out[166];
     layer4_out[610] <= layer3_out[71] & ~layer3_out[72];
     layer4_out[611] <= ~(layer3_out[631] & layer3_out[632]);
     layer4_out[612] <= layer3_out[358] & ~layer3_out[359];
     layer4_out[613] <= layer3_out[577];
     layer4_out[614] <= layer3_out[197] ^ layer3_out[198];
     layer4_out[615] <= ~(layer3_out[22] ^ layer3_out[23]);
     layer4_out[616] <= layer3_out[69] | layer3_out[70];
     layer4_out[617] <= layer3_out[474];
     layer4_out[618] <= ~(layer3_out[740] | layer3_out[741]);
     layer4_out[619] <= ~(layer3_out[654] ^ layer3_out[655]);
     layer4_out[620] <= ~layer3_out[772];
     layer4_out[621] <= ~(layer3_out[359] & layer3_out[360]);
     layer4_out[622] <= ~layer3_out[281];
     layer4_out[623] <= layer3_out[706];
     layer4_out[624] <= ~layer3_out[395];
     layer4_out[625] <= layer3_out[276] & ~layer3_out[275];
     layer4_out[626] <= ~layer3_out[517];
     layer4_out[627] <= layer3_out[475];
     layer4_out[628] <= ~layer3_out[435] | layer3_out[436];
     layer4_out[629] <= layer3_out[24] & ~layer3_out[25];
     layer4_out[630] <= ~layer3_out[519];
     layer4_out[631] <= layer3_out[20];
     layer4_out[632] <= ~layer3_out[569];
     layer4_out[633] <= layer3_out[440] & layer3_out[441];
     layer4_out[634] <= layer3_out[101] & ~layer3_out[100];
     layer4_out[635] <= layer3_out[346] & ~layer3_out[345];
     layer4_out[636] <= layer3_out[659];
     layer4_out[637] <= ~layer3_out[251];
     layer4_out[638] <= layer3_out[555] | layer3_out[556];
     layer4_out[639] <= layer3_out[649] & ~layer3_out[650];
     layer4_out[640] <= ~layer3_out[738];
     layer4_out[641] <= layer3_out[654];
     layer4_out[642] <= ~(layer3_out[538] | layer3_out[539]);
     layer4_out[643] <= ~(layer3_out[308] & layer3_out[309]);
     layer4_out[644] <= layer3_out[315];
     layer4_out[645] <= layer3_out[214];
     layer4_out[646] <= ~(layer3_out[725] & layer3_out[726]);
     layer4_out[647] <= layer3_out[530] & layer3_out[531];
     layer4_out[648] <= layer3_out[313] & ~layer3_out[312];
     layer4_out[649] <= layer3_out[760];
     layer4_out[650] <= layer3_out[437];
     layer4_out[651] <= layer3_out[392];
     layer4_out[652] <= layer3_out[382];
     layer4_out[653] <= ~layer3_out[191];
     layer4_out[654] <= ~layer3_out[232];
     layer4_out[655] <= ~layer3_out[154] | layer3_out[153];
     layer4_out[656] <= layer3_out[630];
     layer4_out[657] <= layer3_out[379] & ~layer3_out[378];
     layer4_out[658] <= ~(layer3_out[38] & layer3_out[39]);
     layer4_out[659] <= layer3_out[674];
     layer4_out[660] <= ~layer3_out[242];
     layer4_out[661] <= ~(layer3_out[200] & layer3_out[201]);
     layer4_out[662] <= ~(layer3_out[32] & layer3_out[33]);
     layer4_out[663] <= layer3_out[331] ^ layer3_out[332];
     layer4_out[664] <= layer3_out[778];
     layer4_out[665] <= layer3_out[657] & layer3_out[658];
     layer4_out[666] <= layer3_out[505] & ~layer3_out[504];
     layer4_out[667] <= ~(layer3_out[771] | layer3_out[772]);
     layer4_out[668] <= ~layer3_out[284];
     layer4_out[669] <= 1'b0;
     layer4_out[670] <= layer3_out[164];
     layer4_out[671] <= layer3_out[255] | layer3_out[256];
     layer4_out[672] <= ~layer3_out[399] | layer3_out[400];
     layer4_out[673] <= ~(layer3_out[180] & layer3_out[181]);
     layer4_out[674] <= layer3_out[645] & ~layer3_out[646];
     layer4_out[675] <= layer3_out[144] & ~layer3_out[145];
     layer4_out[676] <= layer3_out[248];
     layer4_out[677] <= ~(layer3_out[619] & layer3_out[620]);
     layer4_out[678] <= ~layer3_out[321] | layer3_out[320];
     layer4_out[679] <= 1'b1;
     layer4_out[680] <= ~layer3_out[199];
     layer4_out[681] <= ~(layer3_out[366] & layer3_out[367]);
     layer4_out[682] <= ~layer3_out[651];
     layer4_out[683] <= ~layer3_out[510];
     layer4_out[684] <= layer3_out[206] & layer3_out[207];
     layer4_out[685] <= ~layer3_out[509];
     layer4_out[686] <= layer3_out[133] & ~layer3_out[134];
     layer4_out[687] <= ~layer3_out[157];
     layer4_out[688] <= layer3_out[775];
     layer4_out[689] <= layer3_out[211] ^ layer3_out[212];
     layer4_out[690] <= layer3_out[339];
     layer4_out[691] <= ~layer3_out[766] | layer3_out[767];
     layer4_out[692] <= layer3_out[420];
     layer4_out[693] <= ~layer3_out[322];
     layer4_out[694] <= ~layer3_out[87];
     layer4_out[695] <= layer3_out[130] | layer3_out[131];
     layer4_out[696] <= ~layer3_out[774];
     layer4_out[697] <= ~(layer3_out[412] ^ layer3_out[413]);
     layer4_out[698] <= layer3_out[775];
     layer4_out[699] <= ~(layer3_out[492] | layer3_out[493]);
     layer4_out[700] <= ~layer3_out[219];
     layer4_out[701] <= ~(layer3_out[694] ^ layer3_out[695]);
     layer4_out[702] <= ~layer3_out[183];
     layer4_out[703] <= layer3_out[12];
     layer4_out[704] <= ~layer3_out[187];
     layer4_out[705] <= ~layer3_out[509] | layer3_out[508];
     layer4_out[706] <= ~layer3_out[594] | layer3_out[595];
     layer4_out[707] <= ~layer3_out[356] | layer3_out[355];
     layer4_out[708] <= layer3_out[517];
     layer4_out[709] <= layer3_out[618];
     layer4_out[710] <= layer3_out[642] & ~layer3_out[643];
     layer4_out[711] <= layer3_out[228] & ~layer3_out[227];
     layer4_out[712] <= layer3_out[730];
     layer4_out[713] <= ~(layer3_out[413] | layer3_out[414]);
     layer4_out[714] <= layer3_out[45] & ~layer3_out[44];
     layer4_out[715] <= ~layer3_out[468] | layer3_out[467];
     layer4_out[716] <= ~layer3_out[461];
     layer4_out[717] <= ~layer3_out[479] | layer3_out[478];
     layer4_out[718] <= ~(layer3_out[101] | layer3_out[102]);
     layer4_out[719] <= ~layer3_out[240] | layer3_out[241];
     layer4_out[720] <= ~layer3_out[162] | layer3_out[163];
     layer4_out[721] <= ~(layer3_out[703] | layer3_out[704]);
     layer4_out[722] <= ~layer3_out[489] | layer3_out[488];
     layer4_out[723] <= layer3_out[103];
     layer4_out[724] <= ~layer3_out[352];
     layer4_out[725] <= layer3_out[190] & ~layer3_out[191];
     layer4_out[726] <= ~(layer3_out[713] ^ layer3_out[714]);
     layer4_out[727] <= layer3_out[794];
     layer4_out[728] <= ~layer3_out[527] | layer3_out[528];
     layer4_out[729] <= ~layer3_out[208];
     layer4_out[730] <= layer3_out[461] & ~layer3_out[460];
     layer4_out[731] <= layer3_out[474];
     layer4_out[732] <= ~layer3_out[114] | layer3_out[115];
     layer4_out[733] <= layer3_out[796] | layer3_out[797];
     layer4_out[734] <= ~(layer3_out[173] & layer3_out[174]);
     layer4_out[735] <= ~(layer3_out[733] ^ layer3_out[734]);
     layer4_out[736] <= ~(layer3_out[203] ^ layer3_out[204]);
     layer4_out[737] <= ~layer3_out[500];
     layer4_out[738] <= ~layer3_out[746];
     layer4_out[739] <= ~layer3_out[64] | layer3_out[63];
     layer4_out[740] <= ~layer3_out[445] | layer3_out[444];
     layer4_out[741] <= ~layer3_out[767] | layer3_out[768];
     layer4_out[742] <= ~layer3_out[285] | layer3_out[284];
     layer4_out[743] <= 1'b0;
     layer4_out[744] <= ~layer3_out[634] | layer3_out[635];
     layer4_out[745] <= layer3_out[99];
     layer4_out[746] <= layer3_out[177] ^ layer3_out[178];
     layer4_out[747] <= ~(layer3_out[609] | layer3_out[610]);
     layer4_out[748] <= layer3_out[454];
     layer4_out[749] <= ~layer3_out[3] | layer3_out[2];
     layer4_out[750] <= layer3_out[20];
     layer4_out[751] <= ~layer3_out[277] | layer3_out[276];
     layer4_out[752] <= 1'b0;
     layer4_out[753] <= ~(layer3_out[354] | layer3_out[355]);
     layer4_out[754] <= layer3_out[319];
     layer4_out[755] <= layer3_out[305] & layer3_out[306];
     layer4_out[756] <= ~(layer3_out[756] ^ layer3_out[757]);
     layer4_out[757] <= layer3_out[384];
     layer4_out[758] <= layer3_out[701];
     layer4_out[759] <= ~layer3_out[601];
     layer4_out[760] <= layer3_out[125] ^ layer3_out[126];
     layer4_out[761] <= layer3_out[92];
     layer4_out[762] <= ~layer3_out[327];
     layer4_out[763] <= ~layer3_out[639];
     layer4_out[764] <= ~layer3_out[317];
     layer4_out[765] <= layer3_out[697];
     layer4_out[766] <= layer3_out[554] | layer3_out[555];
     layer4_out[767] <= layer3_out[178];
     layer4_out[768] <= layer3_out[274];
     layer4_out[769] <= layer3_out[109] & ~layer3_out[110];
     layer4_out[770] <= ~layer3_out[770];
     layer4_out[771] <= ~(layer3_out[256] & layer3_out[257]);
     layer4_out[772] <= ~layer3_out[486] | layer3_out[485];
     layer4_out[773] <= ~layer3_out[480] | layer3_out[481];
     layer4_out[774] <= layer3_out[149];
     layer4_out[775] <= layer3_out[664] & layer3_out[665];
     layer4_out[776] <= layer3_out[574];
     layer4_out[777] <= layer3_out[347];
     layer4_out[778] <= layer3_out[228];
     layer4_out[779] <= ~layer3_out[622];
     layer4_out[780] <= 1'b0;
     layer4_out[781] <= ~layer3_out[302] | layer3_out[301];
     layer4_out[782] <= ~layer3_out[765];
     layer4_out[783] <= layer3_out[582] & ~layer3_out[581];
     layer4_out[784] <= ~(layer3_out[500] & layer3_out[501]);
     layer4_out[785] <= layer3_out[432] & ~layer3_out[431];
     layer4_out[786] <= ~(layer3_out[689] & layer3_out[690]);
     layer4_out[787] <= ~layer3_out[479];
     layer4_out[788] <= layer3_out[221];
     layer4_out[789] <= layer3_out[304];
     layer4_out[790] <= ~layer3_out[298] | layer3_out[297];
     layer4_out[791] <= ~layer3_out[583];
     layer4_out[792] <= ~layer3_out[351];
     layer4_out[793] <= layer3_out[753] ^ layer3_out[754];
     layer4_out[794] <= ~layer3_out[193];
     layer4_out[795] <= layer3_out[549];
     layer4_out[796] <= layer3_out[327] & ~layer3_out[326];
     layer4_out[797] <= layer3_out[94];
     layer4_out[798] <= layer3_out[268];
     layer4_out[799] <= layer3_out[106];
     layer5_out[0] <= layer4_out[253] & layer4_out[254];
     layer5_out[1] <= ~(layer4_out[117] | layer4_out[118]);
     layer5_out[2] <= layer4_out[645] & ~layer4_out[646];
     layer5_out[3] <= ~(layer4_out[403] ^ layer4_out[404]);
     layer5_out[4] <= layer4_out[345];
     layer5_out[5] <= ~(layer4_out[143] | layer4_out[144]);
     layer5_out[6] <= ~layer4_out[154];
     layer5_out[7] <= layer4_out[196];
     layer5_out[8] <= ~(layer4_out[478] ^ layer4_out[479]);
     layer5_out[9] <= ~layer4_out[687];
     layer5_out[10] <= layer4_out[93];
     layer5_out[11] <= layer4_out[169];
     layer5_out[12] <= ~layer4_out[325];
     layer5_out[13] <= ~layer4_out[372];
     layer5_out[14] <= ~layer4_out[393];
     layer5_out[15] <= ~layer4_out[206];
     layer5_out[16] <= layer4_out[525] & ~layer4_out[526];
     layer5_out[17] <= ~(layer4_out[122] | layer4_out[123]);
     layer5_out[18] <= layer4_out[727] & ~layer4_out[726];
     layer5_out[19] <= ~layer4_out[681] | layer4_out[680];
     layer5_out[20] <= layer4_out[654] & ~layer4_out[655];
     layer5_out[21] <= layer4_out[605];
     layer5_out[22] <= layer4_out[209];
     layer5_out[23] <= layer4_out[784];
     layer5_out[24] <= ~layer4_out[540];
     layer5_out[25] <= layer4_out[610] & ~layer4_out[611];
     layer5_out[26] <= ~layer4_out[510];
     layer5_out[27] <= layer4_out[68];
     layer5_out[28] <= ~layer4_out[449];
     layer5_out[29] <= layer4_out[281] ^ layer4_out[282];
     layer5_out[30] <= layer4_out[403];
     layer5_out[31] <= ~layer4_out[387];
     layer5_out[32] <= ~layer4_out[29];
     layer5_out[33] <= ~(layer4_out[135] | layer4_out[136]);
     layer5_out[34] <= ~layer4_out[455];
     layer5_out[35] <= layer4_out[182] & ~layer4_out[183];
     layer5_out[36] <= ~(layer4_out[452] & layer4_out[453]);
     layer5_out[37] <= ~layer4_out[371];
     layer5_out[38] <= layer4_out[221] ^ layer4_out[222];
     layer5_out[39] <= layer4_out[641];
     layer5_out[40] <= ~layer4_out[340];
     layer5_out[41] <= ~(layer4_out[82] | layer4_out[83]);
     layer5_out[42] <= ~layer4_out[291];
     layer5_out[43] <= ~layer4_out[426];
     layer5_out[44] <= layer4_out[97] & ~layer4_out[98];
     layer5_out[45] <= layer4_out[691] & ~layer4_out[692];
     layer5_out[46] <= layer4_out[799];
     layer5_out[47] <= layer4_out[756] & layer4_out[757];
     layer5_out[48] <= layer4_out[132] & ~layer4_out[133];
     layer5_out[49] <= ~(layer4_out[558] | layer4_out[559]);
     layer5_out[50] <= layer4_out[625];
     layer5_out[51] <= ~layer4_out[265];
     layer5_out[52] <= layer4_out[569];
     layer5_out[53] <= ~layer4_out[477];
     layer5_out[54] <= layer4_out[543] & ~layer4_out[544];
     layer5_out[55] <= ~layer4_out[27];
     layer5_out[56] <= layer4_out[538] ^ layer4_out[539];
     layer5_out[57] <= layer4_out[54] & layer4_out[55];
     layer5_out[58] <= ~layer4_out[378];
     layer5_out[59] <= layer4_out[445] & layer4_out[446];
     layer5_out[60] <= ~layer4_out[440];
     layer5_out[61] <= layer4_out[476];
     layer5_out[62] <= ~(layer4_out[675] & layer4_out[676]);
     layer5_out[63] <= ~layer4_out[140];
     layer5_out[64] <= ~layer4_out[556];
     layer5_out[65] <= ~layer4_out[413];
     layer5_out[66] <= layer4_out[79] & ~layer4_out[78];
     layer5_out[67] <= ~layer4_out[355];
     layer5_out[68] <= layer4_out[668] & layer4_out[669];
     layer5_out[69] <= layer4_out[350] & ~layer4_out[351];
     layer5_out[70] <= layer4_out[0];
     layer5_out[71] <= ~layer4_out[294];
     layer5_out[72] <= layer4_out[728];
     layer5_out[73] <= ~layer4_out[704];
     layer5_out[74] <= ~layer4_out[745];
     layer5_out[75] <= layer4_out[422];
     layer5_out[76] <= layer4_out[534];
     layer5_out[77] <= layer4_out[305] & layer4_out[306];
     layer5_out[78] <= layer4_out[275] & layer4_out[276];
     layer5_out[79] <= layer4_out[494] & layer4_out[495];
     layer5_out[80] <= layer4_out[309] ^ layer4_out[310];
     layer5_out[81] <= ~layer4_out[243];
     layer5_out[82] <= ~layer4_out[145];
     layer5_out[83] <= layer4_out[251] & ~layer4_out[252];
     layer5_out[84] <= layer4_out[597] & layer4_out[598];
     layer5_out[85] <= layer4_out[725] & layer4_out[726];
     layer5_out[86] <= layer4_out[166];
     layer5_out[87] <= ~layer4_out[298];
     layer5_out[88] <= ~layer4_out[332];
     layer5_out[89] <= layer4_out[477] & ~layer4_out[478];
     layer5_out[90] <= layer4_out[487] & layer4_out[488];
     layer5_out[91] <= ~layer4_out[521];
     layer5_out[92] <= layer4_out[613];
     layer5_out[93] <= ~layer4_out[184];
     layer5_out[94] <= layer4_out[479];
     layer5_out[95] <= layer4_out[209] & ~layer4_out[210];
     layer5_out[96] <= layer4_out[160] & ~layer4_out[159];
     layer5_out[97] <= layer4_out[542];
     layer5_out[98] <= ~layer4_out[574];
     layer5_out[99] <= layer4_out[92];
     layer5_out[100] <= ~layer4_out[619];
     layer5_out[101] <= ~layer4_out[789];
     layer5_out[102] <= ~(layer4_out[247] | layer4_out[248]);
     layer5_out[103] <= layer4_out[124] & ~layer4_out[123];
     layer5_out[104] <= layer4_out[288];
     layer5_out[105] <= ~layer4_out[470];
     layer5_out[106] <= layer4_out[167] & ~layer4_out[166];
     layer5_out[107] <= layer4_out[693] & ~layer4_out[694];
     layer5_out[108] <= layer4_out[581];
     layer5_out[109] <= layer4_out[356] & ~layer4_out[357];
     layer5_out[110] <= layer4_out[317] & ~layer4_out[316];
     layer5_out[111] <= layer4_out[49] & ~layer4_out[48];
     layer5_out[112] <= layer4_out[498];
     layer5_out[113] <= layer4_out[357] & layer4_out[358];
     layer5_out[114] <= layer4_out[128] & ~layer4_out[129];
     layer5_out[115] <= layer4_out[115];
     layer5_out[116] <= layer4_out[730] & ~layer4_out[731];
     layer5_out[117] <= layer4_out[445] & ~layer4_out[444];
     layer5_out[118] <= layer4_out[145];
     layer5_out[119] <= layer4_out[233] & ~layer4_out[234];
     layer5_out[120] <= layer4_out[299] & layer4_out[300];
     layer5_out[121] <= ~layer4_out[523];
     layer5_out[122] <= layer4_out[755] & layer4_out[756];
     layer5_out[123] <= layer4_out[519];
     layer5_out[124] <= layer4_out[100];
     layer5_out[125] <= layer4_out[189] & ~layer4_out[188];
     layer5_out[126] <= layer4_out[735] & ~layer4_out[736];
     layer5_out[127] <= layer4_out[426] & ~layer4_out[425];
     layer5_out[128] <= layer4_out[406];
     layer5_out[129] <= layer4_out[774] & ~layer4_out[773];
     layer5_out[130] <= layer4_out[581] & ~layer4_out[582];
     layer5_out[131] <= layer4_out[328];
     layer5_out[132] <= ~layer4_out[647];
     layer5_out[133] <= ~(layer4_out[365] ^ layer4_out[366]);
     layer5_out[134] <= ~layer4_out[527];
     layer5_out[135] <= ~(layer4_out[413] | layer4_out[414]);
     layer5_out[136] <= ~layer4_out[460];
     layer5_out[137] <= ~layer4_out[31];
     layer5_out[138] <= layer4_out[278] & ~layer4_out[277];
     layer5_out[139] <= layer4_out[350] & ~layer4_out[349];
     layer5_out[140] <= layer4_out[493];
     layer5_out[141] <= layer4_out[5] & ~layer4_out[6];
     layer5_out[142] <= layer4_out[321];
     layer5_out[143] <= layer4_out[418] & layer4_out[419];
     layer5_out[144] <= ~(layer4_out[79] | layer4_out[80]);
     layer5_out[145] <= layer4_out[573];
     layer5_out[146] <= layer4_out[528];
     layer5_out[147] <= layer4_out[754] & ~layer4_out[755];
     layer5_out[148] <= layer4_out[753] & ~layer4_out[754];
     layer5_out[149] <= layer4_out[576];
     layer5_out[150] <= layer4_out[294];
     layer5_out[151] <= layer4_out[236];
     layer5_out[152] <= ~(layer4_out[282] | layer4_out[283]);
     layer5_out[153] <= layer4_out[482];
     layer5_out[154] <= ~(layer4_out[186] | layer4_out[187]);
     layer5_out[155] <= layer4_out[23] & layer4_out[24];
     layer5_out[156] <= layer4_out[414];
     layer5_out[157] <= layer4_out[547];
     layer5_out[158] <= ~layer4_out[246];
     layer5_out[159] <= layer4_out[473] & layer4_out[474];
     layer5_out[160] <= layer4_out[714] | layer4_out[715];
     layer5_out[161] <= layer4_out[775] | layer4_out[776];
     layer5_out[162] <= layer4_out[690];
     layer5_out[163] <= layer4_out[352] & ~layer4_out[351];
     layer5_out[164] <= layer4_out[644];
     layer5_out[165] <= layer4_out[59];
     layer5_out[166] <= ~layer4_out[577];
     layer5_out[167] <= ~layer4_out[724];
     layer5_out[168] <= layer4_out[65];
     layer5_out[169] <= layer4_out[782];
     layer5_out[170] <= layer4_out[461];
     layer5_out[171] <= layer4_out[196] & ~layer4_out[195];
     layer5_out[172] <= layer4_out[13] ^ layer4_out[14];
     layer5_out[173] <= layer4_out[168] ^ layer4_out[169];
     layer5_out[174] <= ~layer4_out[473];
     layer5_out[175] <= ~layer4_out[90];
     layer5_out[176] <= ~layer4_out[594];
     layer5_out[177] <= layer4_out[685] & ~layer4_out[686];
     layer5_out[178] <= layer4_out[663];
     layer5_out[179] <= ~layer4_out[330];
     layer5_out[180] <= ~layer4_out[244] | layer4_out[243];
     layer5_out[181] <= ~layer4_out[18];
     layer5_out[182] <= ~layer4_out[566];
     layer5_out[183] <= layer4_out[66];
     layer5_out[184] <= ~(layer4_out[419] ^ layer4_out[420]);
     layer5_out[185] <= ~(layer4_out[508] ^ layer4_out[509]);
     layer5_out[186] <= layer4_out[375];
     layer5_out[187] <= layer4_out[177];
     layer5_out[188] <= ~layer4_out[174];
     layer5_out[189] <= ~layer4_out[617];
     layer5_out[190] <= ~layer4_out[8] | layer4_out[9];
     layer5_out[191] <= layer4_out[401];
     layer5_out[192] <= layer4_out[136] & ~layer4_out[137];
     layer5_out[193] <= layer4_out[367];
     layer5_out[194] <= layer4_out[149];
     layer5_out[195] <= ~layer4_out[207];
     layer5_out[196] <= layer4_out[143] & ~layer4_out[142];
     layer5_out[197] <= layer4_out[549];
     layer5_out[198] <= layer4_out[103] ^ layer4_out[104];
     layer5_out[199] <= layer4_out[734];
     layer5_out[200] <= layer4_out[512];
     layer5_out[201] <= layer4_out[607];
     layer5_out[202] <= ~layer4_out[290];
     layer5_out[203] <= layer4_out[551];
     layer5_out[204] <= layer4_out[651] & ~layer4_out[650];
     layer5_out[205] <= layer4_out[709] & layer4_out[710];
     layer5_out[206] <= layer4_out[323] & ~layer4_out[324];
     layer5_out[207] <= ~layer4_out[749];
     layer5_out[208] <= ~layer4_out[157];
     layer5_out[209] <= layer4_out[723];
     layer5_out[210] <= layer4_out[163] ^ layer4_out[164];
     layer5_out[211] <= layer4_out[435];
     layer5_out[212] <= ~layer4_out[701] | layer4_out[702];
     layer5_out[213] <= ~layer4_out[336];
     layer5_out[214] <= layer4_out[453];
     layer5_out[215] <= ~layer4_out[42];
     layer5_out[216] <= layer4_out[43];
     layer5_out[217] <= layer4_out[524];
     layer5_out[218] <= layer4_out[397];
     layer5_out[219] <= layer4_out[219] & layer4_out[220];
     layer5_out[220] <= ~(layer4_out[324] ^ layer4_out[325]);
     layer5_out[221] <= layer4_out[75];
     layer5_out[222] <= ~layer4_out[616];
     layer5_out[223] <= ~(layer4_out[111] | layer4_out[112]);
     layer5_out[224] <= layer4_out[37];
     layer5_out[225] <= layer4_out[50];
     layer5_out[226] <= layer4_out[732] & layer4_out[733];
     layer5_out[227] <= ~layer4_out[620];
     layer5_out[228] <= ~layer4_out[74];
     layer5_out[229] <= ~layer4_out[4];
     layer5_out[230] <= ~(layer4_out[87] & layer4_out[88]);
     layer5_out[231] <= ~layer4_out[499];
     layer5_out[232] <= layer4_out[722];
     layer5_out[233] <= ~(layer4_out[298] ^ layer4_out[299]);
     layer5_out[234] <= layer4_out[245];
     layer5_out[235] <= layer4_out[567] & ~layer4_out[568];
     layer5_out[236] <= layer4_out[602];
     layer5_out[237] <= ~layer4_out[420];
     layer5_out[238] <= layer4_out[462] & layer4_out[463];
     layer5_out[239] <= ~layer4_out[776];
     layer5_out[240] <= layer4_out[175] & ~layer4_out[174];
     layer5_out[241] <= layer4_out[751] & ~layer4_out[750];
     layer5_out[242] <= layer4_out[163];
     layer5_out[243] <= layer4_out[155];
     layer5_out[244] <= layer4_out[659];
     layer5_out[245] <= layer4_out[649] & layer4_out[650];
     layer5_out[246] <= layer4_out[202] & layer4_out[203];
     layer5_out[247] <= layer4_out[534];
     layer5_out[248] <= ~layer4_out[590];
     layer5_out[249] <= ~(layer4_out[126] | layer4_out[127]);
     layer5_out[250] <= ~layer4_out[91];
     layer5_out[251] <= layer4_out[635] & ~layer4_out[636];
     layer5_out[252] <= ~(layer4_out[689] | layer4_out[690]);
     layer5_out[253] <= layer4_out[492] & ~layer4_out[491];
     layer5_out[254] <= ~layer4_out[360];
     layer5_out[255] <= ~layer4_out[698];
     layer5_out[256] <= ~layer4_out[40];
     layer5_out[257] <= ~(layer4_out[541] ^ layer4_out[542]);
     layer5_out[258] <= layer4_out[424] & ~layer4_out[425];
     layer5_out[259] <= ~layer4_out[593] | layer4_out[592];
     layer5_out[260] <= ~layer4_out[45] | layer4_out[44];
     layer5_out[261] <= ~(layer4_out[599] & layer4_out[600]);
     layer5_out[262] <= ~(layer4_out[201] | layer4_out[202]);
     layer5_out[263] <= ~(layer4_out[745] ^ layer4_out[746]);
     layer5_out[264] <= ~layer4_out[70];
     layer5_out[265] <= ~layer4_out[697];
     layer5_out[266] <= layer4_out[583];
     layer5_out[267] <= ~(layer4_out[245] | layer4_out[246]);
     layer5_out[268] <= ~(layer4_out[623] & layer4_out[624]);
     layer5_out[269] <= layer4_out[172] & ~layer4_out[173];
     layer5_out[270] <= ~(layer4_out[416] ^ layer4_out[417]);
     layer5_out[271] <= layer4_out[536];
     layer5_out[272] <= layer4_out[29] & layer4_out[30];
     layer5_out[273] <= layer4_out[308];
     layer5_out[274] <= layer4_out[747] ^ layer4_out[748];
     layer5_out[275] <= ~layer4_out[67];
     layer5_out[276] <= layer4_out[796];
     layer5_out[277] <= layer4_out[588] & ~layer4_out[589];
     layer5_out[278] <= ~layer4_out[600];
     layer5_out[279] <= ~(layer4_out[797] | layer4_out[798]);
     layer5_out[280] <= layer4_out[597] & ~layer4_out[596];
     layer5_out[281] <= layer4_out[560] & layer4_out[561];
     layer5_out[282] <= ~layer4_out[82];
     layer5_out[283] <= ~layer4_out[505];
     layer5_out[284] <= layer4_out[36] & layer4_out[37];
     layer5_out[285] <= layer4_out[720];
     layer5_out[286] <= ~layer4_out[794];
     layer5_out[287] <= layer4_out[557] & ~layer4_out[558];
     layer5_out[288] <= ~layer4_out[348];
     layer5_out[289] <= ~layer4_out[133];
     layer5_out[290] <= layer4_out[484] & ~layer4_out[485];
     layer5_out[291] <= ~(layer4_out[258] | layer4_out[259]);
     layer5_out[292] <= layer4_out[653] ^ layer4_out[654];
     layer5_out[293] <= ~layer4_out[606];
     layer5_out[294] <= ~(layer4_out[375] ^ layer4_out[376]);
     layer5_out[295] <= ~layer4_out[380];
     layer5_out[296] <= layer4_out[694];
     layer5_out[297] <= layer4_out[340] & layer4_out[341];
     layer5_out[298] <= ~(layer4_out[658] | layer4_out[659]);
     layer5_out[299] <= layer4_out[22];
     layer5_out[300] <= layer4_out[362];
     layer5_out[301] <= ~layer4_out[679];
     layer5_out[302] <= layer4_out[583];
     layer5_out[303] <= ~(layer4_out[254] | layer4_out[255]);
     layer5_out[304] <= layer4_out[344] & ~layer4_out[343];
     layer5_out[305] <= layer4_out[217] & ~layer4_out[218];
     layer5_out[306] <= ~layer4_out[666];
     layer5_out[307] <= ~layer4_out[337];
     layer5_out[308] <= layer4_out[194];
     layer5_out[309] <= ~layer4_out[85];
     layer5_out[310] <= ~layer4_out[657] | layer4_out[658];
     layer5_out[311] <= layer4_out[382] & ~layer4_out[381];
     layer5_out[312] <= layer4_out[267] & ~layer4_out[266];
     layer5_out[313] <= layer4_out[17];
     layer5_out[314] <= layer4_out[287];
     layer5_out[315] <= layer4_out[96] ^ layer4_out[97];
     layer5_out[316] <= layer4_out[372];
     layer5_out[317] <= layer4_out[353];
     layer5_out[318] <= layer4_out[302];
     layer5_out[319] <= layer4_out[223];
     layer5_out[320] <= layer4_out[490] & layer4_out[491];
     layer5_out[321] <= ~layer4_out[624];
     layer5_out[322] <= layer4_out[436] & ~layer4_out[435];
     layer5_out[323] <= layer4_out[218] ^ layer4_out[219];
     layer5_out[324] <= layer4_out[191];
     layer5_out[325] <= ~layer4_out[562];
     layer5_out[326] <= layer4_out[43] & ~layer4_out[42];
     layer5_out[327] <= layer4_out[516] & ~layer4_out[517];
     layer5_out[328] <= layer4_out[285] & ~layer4_out[284];
     layer5_out[329] <= layer4_out[767];
     layer5_out[330] <= layer4_out[407] ^ layer4_out[408];
     layer5_out[331] <= layer4_out[180];
     layer5_out[332] <= layer4_out[609] & ~layer4_out[610];
     layer5_out[333] <= ~layer4_out[93];
     layer5_out[334] <= layer4_out[523];
     layer5_out[335] <= ~(layer4_out[235] | layer4_out[236]);
     layer5_out[336] <= layer4_out[652] & ~layer4_out[651];
     layer5_out[337] <= ~layer4_out[88];
     layer5_out[338] <= ~layer4_out[778];
     layer5_out[339] <= layer4_out[432];
     layer5_out[340] <= layer4_out[544];
     layer5_out[341] <= ~layer4_out[227];
     layer5_out[342] <= layer4_out[766];
     layer5_out[343] <= layer4_out[252] & ~layer4_out[253];
     layer5_out[344] <= layer4_out[187] & layer4_out[188];
     layer5_out[345] <= layer4_out[592];
     layer5_out[346] <= ~layer4_out[238];
     layer5_out[347] <= layer4_out[182] & ~layer4_out[181];
     layer5_out[348] <= layer4_out[305];
     layer5_out[349] <= layer4_out[789] | layer4_out[790];
     layer5_out[350] <= layer4_out[670] & ~layer4_out[671];
     layer5_out[351] <= layer4_out[128];
     layer5_out[352] <= ~layer4_out[157];
     layer5_out[353] <= ~layer4_out[232];
     layer5_out[354] <= layer4_out[763] & layer4_out[764];
     layer5_out[355] <= ~(layer4_out[193] & layer4_out[194]);
     layer5_out[356] <= layer4_out[536] & layer4_out[537];
     layer5_out[357] <= layer4_out[769];
     layer5_out[358] <= ~layer4_out[332];
     layer5_out[359] <= ~layer4_out[378] | layer4_out[377];
     layer5_out[360] <= layer4_out[199] & ~layer4_out[198];
     layer5_out[361] <= ~layer4_out[705];
     layer5_out[362] <= layer4_out[433];
     layer5_out[363] <= layer4_out[199];
     layer5_out[364] <= ~(layer4_out[306] ^ layer4_out[307]);
     layer5_out[365] <= layer4_out[2];
     layer5_out[366] <= ~layer4_out[210];
     layer5_out[367] <= layer4_out[739] & layer4_out[740];
     layer5_out[368] <= ~layer4_out[159];
     layer5_out[369] <= layer4_out[444] & ~layer4_out[443];
     layer5_out[370] <= ~layer4_out[629];
     layer5_out[371] <= ~layer4_out[458];
     layer5_out[372] <= layer4_out[343];
     layer5_out[373] <= ~layer4_out[192];
     layer5_out[374] <= ~(layer4_out[51] | layer4_out[52]);
     layer5_out[375] <= layer4_out[502] & ~layer4_out[503];
     layer5_out[376] <= ~(layer4_out[447] ^ layer4_out[448]);
     layer5_out[377] <= ~(layer4_out[481] | layer4_out[482]);
     layer5_out[378] <= layer4_out[622] & ~layer4_out[623];
     layer5_out[379] <= layer4_out[432];
     layer5_out[380] <= layer4_out[399] & layer4_out[400];
     layer5_out[381] <= ~layer4_out[767];
     layer5_out[382] <= layer4_out[470] & ~layer4_out[469];
     layer5_out[383] <= layer4_out[540];
     layer5_out[384] <= layer4_out[26] & ~layer4_out[25];
     layer5_out[385] <= layer4_out[784];
     layer5_out[386] <= ~layer4_out[287];
     layer5_out[387] <= layer4_out[116] & layer4_out[117];
     layer5_out[388] <= layer4_out[752] & layer4_out[753];
     layer5_out[389] <= ~layer4_out[284];
     layer5_out[390] <= ~layer4_out[679];
     layer5_out[391] <= layer4_out[6] | layer4_out[7];
     layer5_out[392] <= layer4_out[242] & ~layer4_out[241];
     layer5_out[393] <= layer4_out[446] & ~layer4_out[447];
     layer5_out[394] <= ~layer4_out[762] | layer4_out[761];
     layer5_out[395] <= layer4_out[637];
     layer5_out[396] <= ~layer4_out[303];
     layer5_out[397] <= ~(layer4_out[466] ^ layer4_out[467]);
     layer5_out[398] <= layer4_out[203] & layer4_out[204];
     layer5_out[399] <= ~(layer4_out[388] | layer4_out[389]);
     layer5_out[400] <= ~layer4_out[731];
     layer5_out[401] <= layer4_out[409] & ~layer4_out[410];
     layer5_out[402] <= ~layer4_out[630] | layer4_out[629];
     layer5_out[403] <= ~layer4_out[500];
     layer5_out[404] <= layer4_out[369] & ~layer4_out[370];
     layer5_out[405] <= ~(layer4_out[229] ^ layer4_out[230]);
     layer5_out[406] <= ~layer4_out[464];
     layer5_out[407] <= ~(layer4_out[333] | layer4_out[334]);
     layer5_out[408] <= layer4_out[461];
     layer5_out[409] <= layer4_out[442] & ~layer4_out[441];
     layer5_out[410] <= ~layer4_out[172];
     layer5_out[411] <= ~layer4_out[63];
     layer5_out[412] <= layer4_out[25] & ~layer4_out[24];
     layer5_out[413] <= ~layer4_out[423];
     layer5_out[414] <= layer4_out[258] & ~layer4_out[257];
     layer5_out[415] <= ~layer4_out[589];
     layer5_out[416] <= layer4_out[279] & layer4_out[280];
     layer5_out[417] <= ~(layer4_out[708] ^ layer4_out[709]);
     layer5_out[418] <= ~(layer4_out[206] ^ layer4_out[207]);
     layer5_out[419] <= layer4_out[518] | layer4_out[519];
     layer5_out[420] <= layer4_out[23] & ~layer4_out[22];
     layer5_out[421] <= layer4_out[330] & layer4_out[331];
     layer5_out[422] <= layer4_out[40];
     layer5_out[423] <= layer4_out[220] & layer4_out[221];
     layer5_out[424] <= layer4_out[632] & ~layer4_out[631];
     layer5_out[425] <= layer4_out[606] & ~layer4_out[607];
     layer5_out[426] <= ~(layer4_out[272] | layer4_out[273]);
     layer5_out[427] <= ~(layer4_out[471] & layer4_out[472]);
     layer5_out[428] <= layer4_out[177];
     layer5_out[429] <= ~layer4_out[239] | layer4_out[238];
     layer5_out[430] <= layer4_out[102];
     layer5_out[431] <= ~layer4_out[545];
     layer5_out[432] <= layer4_out[699];
     layer5_out[433] <= ~layer4_out[249];
     layer5_out[434] <= layer4_out[125];
     layer5_out[435] <= layer4_out[132];
     layer5_out[436] <= ~layer4_out[495];
     layer5_out[437] <= layer4_out[667];
     layer5_out[438] <= ~(layer4_out[411] | layer4_out[412]);
     layer5_out[439] <= layer4_out[717];
     layer5_out[440] <= ~layer4_out[111];
     layer5_out[441] <= ~layer4_out[503] | layer4_out[504];
     layer5_out[442] <= layer4_out[733] | layer4_out[734];
     layer5_out[443] <= layer4_out[347];
     layer5_out[444] <= ~(layer4_out[640] | layer4_out[641]);
     layer5_out[445] <= ~layer4_out[150];
     layer5_out[446] <= layer4_out[436];
     layer5_out[447] <= ~layer4_out[687];
     layer5_out[448] <= ~(layer4_out[230] | layer4_out[231]);
     layer5_out[449] <= layer4_out[256] & layer4_out[257];
     layer5_out[450] <= layer4_out[662];
     layer5_out[451] <= ~(layer4_out[30] | layer4_out[31]);
     layer5_out[452] <= layer4_out[137];
     layer5_out[453] <= ~layer4_out[684] | layer4_out[685];
     layer5_out[454] <= ~layer4_out[139];
     layer5_out[455] <= ~layer4_out[718];
     layer5_out[456] <= ~layer4_out[643];
     layer5_out[457] <= ~(layer4_out[105] ^ layer4_out[106]);
     layer5_out[458] <= layer4_out[632] & layer4_out[633];
     layer5_out[459] <= layer4_out[53];
     layer5_out[460] <= ~layer4_out[313];
     layer5_out[461] <= layer4_out[379];
     layer5_out[462] <= layer4_out[587] ^ layer4_out[588];
     layer5_out[463] <= layer4_out[678];
     layer5_out[464] <= ~(layer4_out[531] | layer4_out[532]);
     layer5_out[465] <= layer4_out[769] & layer4_out[770];
     layer5_out[466] <= layer4_out[421] & ~layer4_out[422];
     layer5_out[467] <= ~(layer4_out[729] | layer4_out[730]);
     layer5_out[468] <= ~layer4_out[100];
     layer5_out[469] <= ~(layer4_out[506] & layer4_out[507]);
     layer5_out[470] <= ~(layer4_out[771] & layer4_out[772]);
     layer5_out[471] <= ~layer4_out[585];
     layer5_out[472] <= ~(layer4_out[664] ^ layer4_out[665]);
     layer5_out[473] <= ~(layer4_out[215] ^ layer4_out[216]);
     layer5_out[474] <= ~layer4_out[270];
     layer5_out[475] <= ~(layer4_out[161] & layer4_out[162]);
     layer5_out[476] <= ~layer4_out[58];
     layer5_out[477] <= ~layer4_out[649];
     layer5_out[478] <= ~(layer4_out[315] | layer4_out[316]);
     layer5_out[479] <= layer4_out[226] & ~layer4_out[225];
     layer5_out[480] <= ~(layer4_out[311] ^ layer4_out[312]);
     layer5_out[481] <= ~layer4_out[771];
     layer5_out[482] <= ~layer4_out[368];
     layer5_out[483] <= layer4_out[9] & ~layer4_out[10];
     layer5_out[484] <= layer4_out[786];
     layer5_out[485] <= ~(layer4_out[451] & layer4_out[452]);
     layer5_out[486] <= layer4_out[19] | layer4_out[20];
     layer5_out[487] <= ~layer4_out[699] | layer4_out[700];
     layer5_out[488] <= ~(layer4_out[118] & layer4_out[119]);
     layer5_out[489] <= layer4_out[507];
     layer5_out[490] <= ~(layer4_out[240] | layer4_out[241]);
     layer5_out[491] <= ~(layer4_out[58] & layer4_out[59]);
     layer5_out[492] <= layer4_out[168];
     layer5_out[493] <= layer4_out[672] & layer4_out[673];
     layer5_out[494] <= ~layer4_out[669];
     layer5_out[495] <= ~layer4_out[779];
     layer5_out[496] <= layer4_out[160];
     layer5_out[497] <= layer4_out[792];
     layer5_out[498] <= ~layer4_out[201];
     layer5_out[499] <= layer4_out[384];
     layer5_out[500] <= ~layer4_out[278] | layer4_out[279];
     layer5_out[501] <= layer4_out[190];
     layer5_out[502] <= layer4_out[280] & ~layer4_out[281];
     layer5_out[503] <= layer4_out[300] & ~layer4_out[301];
     layer5_out[504] <= layer4_out[384] & layer4_out[385];
     layer5_out[505] <= ~(layer4_out[262] | layer4_out[263]);
     layer5_out[506] <= layer4_out[485] ^ layer4_out[486];
     layer5_out[507] <= ~layer4_out[83];
     layer5_out[508] <= ~layer4_out[63];
     layer5_out[509] <= ~layer4_out[81];
     layer5_out[510] <= layer4_out[418];
     layer5_out[511] <= ~layer4_out[69];
     layer5_out[512] <= ~layer4_out[255] | layer4_out[256];
     layer5_out[513] <= layer4_out[549] & layer4_out[550];
     layer5_out[514] <= ~layer4_out[796];
     layer5_out[515] <= layer4_out[500] & layer4_out[501];
     layer5_out[516] <= ~layer4_out[788];
     layer5_out[517] <= ~layer4_out[392];
     layer5_out[518] <= layer4_out[151] & ~layer4_out[152];
     layer5_out[519] <= layer4_out[393] & layer4_out[394];
     layer5_out[520] <= ~layer4_out[587];
     layer5_out[521] <= layer4_out[439] | layer4_out[440];
     layer5_out[522] <= layer4_out[382] & layer4_out[383];
     layer5_out[523] <= layer4_out[405];
     layer5_out[524] <= layer4_out[765];
     layer5_out[525] <= ~layer4_out[141];
     layer5_out[526] <= ~(layer4_out[496] ^ layer4_out[497]);
     layer5_out[527] <= ~layer4_out[14];
     layer5_out[528] <= layer4_out[688] & ~layer4_out[689];
     layer5_out[529] <= ~layer4_out[781];
     layer5_out[530] <= layer4_out[609];
     layer5_out[531] <= ~layer4_out[335];
     layer5_out[532] <= ~(layer4_out[612] & layer4_out[613]);
     layer5_out[533] <= layer4_out[311] & ~layer4_out[310];
     layer5_out[534] <= layer4_out[716] & ~layer4_out[715];
     layer5_out[535] <= ~layer4_out[511];
     layer5_out[536] <= ~layer4_out[703] | layer4_out[704];
     layer5_out[537] <= layer4_out[113];
     layer5_out[538] <= ~layer4_out[437];
     layer5_out[539] <= layer4_out[743];
     layer5_out[540] <= ~(layer4_out[95] | layer4_out[96]);
     layer5_out[541] <= layer4_out[759] ^ layer4_out[760];
     layer5_out[542] <= layer4_out[751];
     layer5_out[543] <= ~(layer4_out[727] | layer4_out[728]);
     layer5_out[544] <= layer4_out[323];
     layer5_out[545] <= ~(layer4_out[291] | layer4_out[292]);
     layer5_out[546] <= layer4_out[338];
     layer5_out[547] <= ~layer4_out[562];
     layer5_out[548] <= layer4_out[319] & ~layer4_out[318];
     layer5_out[549] <= layer4_out[793] & ~layer4_out[792];
     layer5_out[550] <= ~layer4_out[51];
     layer5_out[551] <= ~layer4_out[480];
     layer5_out[552] <= layer4_out[725];
     layer5_out[553] <= layer4_out[104] & ~layer4_out[105];
     layer5_out[554] <= layer4_out[530] & ~layer4_out[529];
     layer5_out[555] <= ~layer4_out[603];
     layer5_out[556] <= ~layer4_out[555] | layer4_out[554];
     layer5_out[557] <= layer4_out[676] & layer4_out[677];
     layer5_out[558] <= layer4_out[328] & ~layer4_out[327];
     layer5_out[559] <= ~(layer4_out[4] & layer4_out[5]);
     layer5_out[560] <= layer4_out[563];
     layer5_out[561] <= ~layer4_out[750];
     layer5_out[562] <= layer4_out[618];
     layer5_out[563] <= layer4_out[638] & layer4_out[639];
     layer5_out[564] <= ~(layer4_out[449] | layer4_out[450]);
     layer5_out[565] <= layer4_out[130] & ~layer4_out[131];
     layer5_out[566] <= ~layer4_out[389];
     layer5_out[567] <= ~layer4_out[204];
     layer5_out[568] <= layer4_out[454] & layer4_out[455];
     layer5_out[569] <= layer4_out[616];
     layer5_out[570] <= layer4_out[214] & layer4_out[215];
     layer5_out[571] <= layer4_out[565] & layer4_out[566];
     layer5_out[572] <= ~layer4_out[35];
     layer5_out[573] <= layer4_out[573] & layer4_out[574];
     layer5_out[574] <= ~layer4_out[391];
     layer5_out[575] <= layer4_out[653] & ~layer4_out[652];
     layer5_out[576] <= ~layer4_out[268];
     layer5_out[577] <= ~layer4_out[647];
     layer5_out[578] <= layer4_out[682];
     layer5_out[579] <= layer4_out[711] & ~layer4_out[712];
     layer5_out[580] <= ~layer4_out[364];
     layer5_out[581] <= layer4_out[191] | layer4_out[192];
     layer5_out[582] <= layer4_out[577];
     layer5_out[583] <= layer4_out[313];
     layer5_out[584] <= layer4_out[261] & ~layer4_out[260];
     layer5_out[585] <= ~layer4_out[701] | layer4_out[700];
     layer5_out[586] <= layer4_out[484];
     layer5_out[587] <= layer4_out[612] & ~layer4_out[611];
     layer5_out[588] <= layer4_out[95];
     layer5_out[589] <= layer4_out[416];
     layer5_out[590] <= layer4_out[550] & layer4_out[551];
     layer5_out[591] <= layer4_out[274] & layer4_out[275];
     layer5_out[592] <= ~(layer4_out[320] | layer4_out[321]);
     layer5_out[593] <= layer4_out[3];
     layer5_out[594] <= layer4_out[232];
     layer5_out[595] <= layer4_out[531] & ~layer4_out[530];
     layer5_out[596] <= ~layer4_out[77];
     layer5_out[597] <= ~layer4_out[490] | layer4_out[489];
     layer5_out[598] <= layer4_out[376];
     layer5_out[599] <= layer4_out[7] & ~layer4_out[8];
     layer5_out[600] <= ~(layer4_out[780] ^ layer4_out[781]);
     layer5_out[601] <= ~layer4_out[790];
     layer5_out[602] <= ~layer4_out[667];
     layer5_out[603] <= ~layer4_out[411];
     layer5_out[604] <= layer4_out[710];
     layer5_out[605] <= layer4_out[53] & layer4_out[54];
     layer5_out[606] <= layer4_out[120] & layer4_out[121];
     layer5_out[607] <= ~(layer4_out[644] | layer4_out[645]);
     layer5_out[608] <= layer4_out[584] ^ layer4_out[585];
     layer5_out[609] <= ~layer4_out[319];
     layer5_out[610] <= layer4_out[134];
     layer5_out[611] <= ~layer4_out[401];
     layer5_out[612] <= layer4_out[664] & ~layer4_out[663];
     layer5_out[613] <= ~layer4_out[693];
     layer5_out[614] <= layer4_out[292] & layer4_out[293];
     layer5_out[615] <= layer4_out[374] & ~layer4_out[373];
     layer5_out[616] <= ~(layer4_out[430] | layer4_out[431]);
     layer5_out[617] <= layer4_out[352] & layer4_out[353];
     layer5_out[618] <= layer4_out[489];
     layer5_out[619] <= ~layer4_out[65];
     layer5_out[620] <= ~(layer4_out[98] ^ layer4_out[99]);
     layer5_out[621] <= ~(layer4_out[317] | layer4_out[318]);
     layer5_out[622] <= layer4_out[226] & layer4_out[227];
     layer5_out[623] <= layer4_out[492];
     layer5_out[624] <= ~layer4_out[273];
     layer5_out[625] <= layer4_out[626] | layer4_out[627];
     layer5_out[626] <= ~(layer4_out[595] | layer4_out[596]);
     layer5_out[627] <= layer4_out[265] & layer4_out[266];
     layer5_out[628] <= layer4_out[639];
     layer5_out[629] <= ~layer4_out[296] | layer4_out[297];
     layer5_out[630] <= layer4_out[580] & ~layer4_out[579];
     layer5_out[631] <= ~layer4_out[356];
     layer5_out[632] <= ~layer4_out[259];
     layer5_out[633] <= layer4_out[385] ^ layer4_out[386];
     layer5_out[634] <= ~(layer4_out[307] | layer4_out[308]);
     layer5_out[635] <= layer4_out[674] & ~layer4_out[673];
     layer5_out[636] <= layer4_out[261] & layer4_out[262];
     layer5_out[637] <= layer4_out[512] & layer4_out[513];
     layer5_out[638] <= layer4_out[603];
     layer5_out[639] <= ~layer4_out[695];
     layer5_out[640] <= ~layer4_out[251];
     layer5_out[641] <= layer4_out[180] & ~layer4_out[181];
     layer5_out[642] <= layer4_out[706] & layer4_out[707];
     layer5_out[643] <= ~layer4_out[240];
     layer5_out[644] <= layer4_out[228] & ~layer4_out[229];
     layer5_out[645] <= layer4_out[268] | layer4_out[269];
     layer5_out[646] <= layer4_out[718] & ~layer4_out[717];
     layer5_out[647] <= layer4_out[11] & layer4_out[12];
     layer5_out[648] <= ~(layer4_out[302] | layer4_out[303]);
     layer5_out[649] <= ~(layer4_out[428] & layer4_out[429]);
     layer5_out[650] <= layer4_out[615] & ~layer4_out[614];
     layer5_out[651] <= layer4_out[73] & ~layer4_out[72];
     layer5_out[652] <= layer4_out[314] ^ layer4_out[315];
     layer5_out[653] <= layer4_out[599] & ~layer4_out[598];
     layer5_out[654] <= layer4_out[164] & ~layer4_out[165];
     layer5_out[655] <= layer4_out[358] ^ layer4_out[359];
     layer5_out[656] <= ~(layer4_out[211] | layer4_out[212]);
     layer5_out[657] <= layer4_out[513] ^ layer4_out[514];
     layer5_out[658] <= layer4_out[772] & layer4_out[773];
     layer5_out[659] <= ~layer4_out[570];
     layer5_out[660] <= ~(layer4_out[10] | layer4_out[11]);
     layer5_out[661] <= layer4_out[438];
     layer5_out[662] <= layer4_out[366] & ~layer4_out[367];
     layer5_out[663] <= layer4_out[578];
     layer5_out[664] <= layer4_out[777] & layer4_out[778];
     layer5_out[665] <= layer4_out[78];
     layer5_out[666] <= layer4_out[276] & ~layer4_out[277];
     layer5_out[667] <= layer4_out[660];
     layer5_out[668] <= layer4_out[295];
     layer5_out[669] <= layer4_out[474] & layer4_out[475];
     layer5_out[670] <= ~layer4_out[271];
     layer5_out[671] <= ~layer4_out[546];
     layer5_out[672] <= layer4_out[153];
     layer5_out[673] <= layer4_out[342];
     layer5_out[674] <= layer4_out[537];
     layer5_out[675] <= layer4_out[33] ^ layer4_out[34];
     layer5_out[676] <= ~(layer4_out[760] ^ layer4_out[761]);
     layer5_out[677] <= layer4_out[737] & ~layer4_out[736];
     layer5_out[678] <= ~(layer4_out[442] | layer4_out[443]);
     layer5_out[679] <= layer4_out[214] & ~layer4_out[213];
     layer5_out[680] <= ~(layer4_out[553] ^ layer4_out[554]);
     layer5_out[681] <= ~(layer4_out[464] ^ layer4_out[465]);
     layer5_out[682] <= layer4_out[785];
     layer5_out[683] <= layer4_out[520] & ~layer4_out[521];
     layer5_out[684] <= ~layer4_out[683] | layer4_out[682];
     layer5_out[685] <= ~(layer4_out[86] | layer4_out[87]);
     layer5_out[686] <= layer4_out[121];
     layer5_out[687] <= ~layer4_out[468];
     layer5_out[688] <= layer4_out[637] & ~layer4_out[636];
     layer5_out[689] <= layer4_out[185] & ~layer4_out[186];
     layer5_out[690] <= ~layer4_out[564];
     layer5_out[691] <= ~(layer4_out[450] | layer4_out[451]);
     layer5_out[692] <= ~(layer4_out[46] ^ layer4_out[47]);
     layer5_out[693] <= layer4_out[630] & layer4_out[631];
     layer5_out[694] <= layer4_out[427] & ~layer4_out[428];
     layer5_out[695] <= layer4_out[27];
     layer5_out[696] <= ~layer4_out[16];
     layer5_out[697] <= layer4_out[271] & ~layer4_out[272];
     layer5_out[698] <= layer4_out[758] | layer4_out[759];
     layer5_out[699] <= ~layer4_out[502];
     layer5_out[700] <= ~(layer4_out[627] & layer4_out[628]);
     layer5_out[701] <= ~(layer4_out[743] | layer4_out[744]);
     layer5_out[702] <= ~layer4_out[458] | layer4_out[457];
     layer5_out[703] <= ~(layer4_out[138] ^ layer4_out[139]);
     layer5_out[704] <= layer4_out[409];
     layer5_out[705] <= ~layer4_out[486];
     layer5_out[706] <= ~layer4_out[703] | layer4_out[702];
     layer5_out[707] <= layer4_out[148] & ~layer4_out[147];
     layer5_out[708] <= ~layer4_out[285];
     layer5_out[709] <= layer4_out[20] | layer4_out[21];
     layer5_out[710] <= ~layer4_out[107];
     layer5_out[711] <= ~layer4_out[45];
     layer5_out[712] <= layer4_out[528];
     layer5_out[713] <= layer4_out[35] ^ layer4_out[36];
     layer5_out[714] <= ~(layer4_out[762] | layer4_out[763]);
     layer5_out[715] <= layer4_out[793];
     layer5_out[716] <= layer4_out[198] & ~layer4_out[197];
     layer5_out[717] <= layer4_out[683];
     layer5_out[718] <= ~layer4_out[0];
     layer5_out[719] <= ~(layer4_out[119] & layer4_out[120]);
     layer5_out[720] <= layer4_out[223] & layer4_out[224];
     layer5_out[721] <= layer4_out[514];
     layer5_out[722] <= layer4_out[465];
     layer5_out[723] <= layer4_out[719] & ~layer4_out[720];
     layer5_out[724] <= layer4_out[572] & ~layer4_out[571];
     layer5_out[725] <= ~layer4_out[216];
     layer5_out[726] <= ~(layer4_out[396] | layer4_out[397]);
     layer5_out[727] <= layer4_out[741] & layer4_out[742];
     layer5_out[728] <= layer4_out[126] & ~layer4_out[125];
     layer5_out[729] <= layer4_out[60] & ~layer4_out[61];
     layer5_out[730] <= layer4_out[518];
     layer5_out[731] <= layer4_out[16] ^ layer4_out[17];
     layer5_out[732] <= layer4_out[129];
     layer5_out[733] <= layer4_out[184] & ~layer4_out[185];
     layer5_out[734] <= ~(layer4_out[249] | layer4_out[250]);
     layer5_out[735] <= ~(layer4_out[738] ^ layer4_out[739]);
     layer5_out[736] <= layer4_out[657] & ~layer4_out[656];
     layer5_out[737] <= ~(layer4_out[594] | layer4_out[595]);
     layer5_out[738] <= layer4_out[360] & ~layer4_out[359];
     layer5_out[739] <= ~layer4_out[364] | layer4_out[365];
     layer5_out[740] <= ~(layer4_out[38] | layer4_out[39]);
     layer5_out[741] <= layer4_out[671] & layer4_out[672];
     layer5_out[742] <= layer4_out[170] & ~layer4_out[171];
     layer5_out[743] <= layer4_out[456] ^ layer4_out[457];
     layer5_out[744] <= layer4_out[109] & layer4_out[110];
     layer5_out[745] <= ~layer4_out[62] | layer4_out[61];
     layer5_out[746] <= layer4_out[12];
     layer5_out[747] <= layer4_out[395];
     layer5_out[748] <= ~layer4_out[741];
     layer5_out[749] <= layer4_out[516];
     layer5_out[750] <= layer4_out[338];
     layer5_out[751] <= layer4_out[707];
     layer5_out[752] <= ~(layer4_out[153] ^ layer4_out[154]);
     layer5_out[753] <= layer4_out[151];
     layer5_out[754] <= layer4_out[635];
     layer5_out[755] <= layer4_out[504];
     layer5_out[756] <= layer4_out[398] & ~layer4_out[399];
     layer5_out[757] <= layer4_out[552];
     layer5_out[758] <= layer4_out[674] & layer4_out[675];
     layer5_out[759] <= layer4_out[347] & ~layer4_out[346];
     layer5_out[760] <= layer4_out[55] & ~layer4_out[56];
     layer5_out[761] <= ~(layer4_out[556] | layer4_out[557]);
     layer5_out[762] <= ~layer4_out[570];
     layer5_out[763] <= layer4_out[112];
     layer5_out[764] <= layer4_out[212] ^ layer4_out[213];
     layer5_out[765] <= layer4_out[533];
     layer5_out[766] <= ~(layer4_out[344] | layer4_out[345]);
     layer5_out[767] <= ~layer4_out[712];
     layer5_out[768] <= ~layer4_out[386];
     layer5_out[769] <= ~layer4_out[147];
     layer5_out[770] <= layer4_out[362] & ~layer4_out[361];
     layer5_out[771] <= ~layer4_out[179];
     layer5_out[772] <= ~layer4_out[775];
     layer5_out[773] <= ~(layer4_out[71] | layer4_out[72]);
     layer5_out[774] <= layer4_out[101] & layer4_out[102];
     layer5_out[775] <= ~(layer4_out[633] | layer4_out[634]);
     layer5_out[776] <= ~layer4_out[175];
     layer5_out[777] <= layer4_out[225];
     layer5_out[778] <= layer4_out[714] & ~layer4_out[713];
     layer5_out[779] <= layer4_out[56] & layer4_out[57];
     layer5_out[780] <= layer4_out[48];
     layer5_out[781] <= ~layer4_out[326];
     layer5_out[782] <= layer4_out[757];
     layer5_out[783] <= ~layer4_out[747];
     layer5_out[784] <= layer4_out[429] & layer4_out[430];
     layer5_out[785] <= layer4_out[468] & ~layer4_out[469];
     layer5_out[786] <= ~layer4_out[33];
     layer5_out[787] <= ~layer4_out[560];
     layer5_out[788] <= layer4_out[738] & ~layer4_out[737];
     layer5_out[789] <= layer4_out[234] ^ layer4_out[235];
     layer5_out[790] <= layer4_out[86];
     layer5_out[791] <= layer4_out[74] & ~layer4_out[75];
     layer5_out[792] <= layer4_out[621] & ~layer4_out[622];
     layer5_out[793] <= layer4_out[115] & ~layer4_out[114];
     layer5_out[794] <= layer4_out[263] & ~layer4_out[264];
     layer5_out[795] <= ~(layer4_out[655] ^ layer4_out[656]);
     layer5_out[796] <= layer4_out[108];
     layer5_out[797] <= layer4_out[107] & ~layer4_out[108];
     layer5_out[798] <= layer4_out[396];
     layer5_out[799] <= ~layer4_out[405];
      last_layer_output <= layer5_out;

      result[0] <= last_layer_output[0] + last_layer_output[1] + last_layer_output[2] + last_layer_output[3] + last_layer_output[4] + last_layer_output[5] + last_layer_output[6] + last_layer_output[7] + last_layer_output[8] + last_layer_output[9] + last_layer_output[10] + last_layer_output[11] + last_layer_output[12] + last_layer_output[13] + last_layer_output[14] + last_layer_output[15] + last_layer_output[16] + last_layer_output[17] + last_layer_output[18] + last_layer_output[19] + last_layer_output[20] + last_layer_output[21] + last_layer_output[22] + last_layer_output[23] + last_layer_output[24] + last_layer_output[25] + last_layer_output[26] + last_layer_output[27] + last_layer_output[28] + last_layer_output[29] + last_layer_output[30] + last_layer_output[31] + last_layer_output[32] + last_layer_output[33] + last_layer_output[34] + last_layer_output[35] + last_layer_output[36] + last_layer_output[37] + last_layer_output[38] + last_layer_output[39] + last_layer_output[40] + last_layer_output[41] + last_layer_output[42] + last_layer_output[43] + last_layer_output[44] + last_layer_output[45] + last_layer_output[46] + last_layer_output[47] + last_layer_output[48] + last_layer_output[49] + last_layer_output[50] + last_layer_output[51] + last_layer_output[52] + last_layer_output[53] + last_layer_output[54] + last_layer_output[55] + last_layer_output[56] + last_layer_output[57] + last_layer_output[58] + last_layer_output[59] + last_layer_output[60] + last_layer_output[61] + last_layer_output[62] + last_layer_output[63] + last_layer_output[64] + last_layer_output[65] + last_layer_output[66] + last_layer_output[67] + last_layer_output[68] + last_layer_output[69] + last_layer_output[70] + last_layer_output[71] + last_layer_output[72] + last_layer_output[73] + last_layer_output[74] + last_layer_output[75] + last_layer_output[76] + last_layer_output[77] + last_layer_output[78] + last_layer_output[79];
      result[1] <= last_layer_output[80] + last_layer_output[81] + last_layer_output[82] + last_layer_output[83] + last_layer_output[84] + last_layer_output[85] + last_layer_output[86] + last_layer_output[87] + last_layer_output[88] + last_layer_output[89] + last_layer_output[90] + last_layer_output[91] + last_layer_output[92] + last_layer_output[93] + last_layer_output[94] + last_layer_output[95] + last_layer_output[96] + last_layer_output[97] + last_layer_output[98] + last_layer_output[99] + last_layer_output[100] + last_layer_output[101] + last_layer_output[102] + last_layer_output[103] + last_layer_output[104] + last_layer_output[105] + last_layer_output[106] + last_layer_output[107] + last_layer_output[108] + last_layer_output[109] + last_layer_output[110] + last_layer_output[111] + last_layer_output[112] + last_layer_output[113] + last_layer_output[114] + last_layer_output[115] + last_layer_output[116] + last_layer_output[117] + last_layer_output[118] + last_layer_output[119] + last_layer_output[120] + last_layer_output[121] + last_layer_output[122] + last_layer_output[123] + last_layer_output[124] + last_layer_output[125] + last_layer_output[126] + last_layer_output[127] + last_layer_output[128] + last_layer_output[129] + last_layer_output[130] + last_layer_output[131] + last_layer_output[132] + last_layer_output[133] + last_layer_output[134] + last_layer_output[135] + last_layer_output[136] + last_layer_output[137] + last_layer_output[138] + last_layer_output[139] + last_layer_output[140] + last_layer_output[141] + last_layer_output[142] + last_layer_output[143] + last_layer_output[144] + last_layer_output[145] + last_layer_output[146] + last_layer_output[147] + last_layer_output[148] + last_layer_output[149] + last_layer_output[150] + last_layer_output[151] + last_layer_output[152] + last_layer_output[153] + last_layer_output[154] + last_layer_output[155] + last_layer_output[156] + last_layer_output[157] + last_layer_output[158] + last_layer_output[159];
      result[2] <= last_layer_output[160] + last_layer_output[161] + last_layer_output[162] + last_layer_output[163] + last_layer_output[164] + last_layer_output[165] + last_layer_output[166] + last_layer_output[167] + last_layer_output[168] + last_layer_output[169] + last_layer_output[170] + last_layer_output[171] + last_layer_output[172] + last_layer_output[173] + last_layer_output[174] + last_layer_output[175] + last_layer_output[176] + last_layer_output[177] + last_layer_output[178] + last_layer_output[179] + last_layer_output[180] + last_layer_output[181] + last_layer_output[182] + last_layer_output[183] + last_layer_output[184] + last_layer_output[185] + last_layer_output[186] + last_layer_output[187] + last_layer_output[188] + last_layer_output[189] + last_layer_output[190] + last_layer_output[191] + last_layer_output[192] + last_layer_output[193] + last_layer_output[194] + last_layer_output[195] + last_layer_output[196] + last_layer_output[197] + last_layer_output[198] + last_layer_output[199] + last_layer_output[200] + last_layer_output[201] + last_layer_output[202] + last_layer_output[203] + last_layer_output[204] + last_layer_output[205] + last_layer_output[206] + last_layer_output[207] + last_layer_output[208] + last_layer_output[209] + last_layer_output[210] + last_layer_output[211] + last_layer_output[212] + last_layer_output[213] + last_layer_output[214] + last_layer_output[215] + last_layer_output[216] + last_layer_output[217] + last_layer_output[218] + last_layer_output[219] + last_layer_output[220] + last_layer_output[221] + last_layer_output[222] + last_layer_output[223] + last_layer_output[224] + last_layer_output[225] + last_layer_output[226] + last_layer_output[227] + last_layer_output[228] + last_layer_output[229] + last_layer_output[230] + last_layer_output[231] + last_layer_output[232] + last_layer_output[233] + last_layer_output[234] + last_layer_output[235] + last_layer_output[236] + last_layer_output[237] + last_layer_output[238] + last_layer_output[239];
      result[3] <= last_layer_output[240] + last_layer_output[241] + last_layer_output[242] + last_layer_output[243] + last_layer_output[244] + last_layer_output[245] + last_layer_output[246] + last_layer_output[247] + last_layer_output[248] + last_layer_output[249] + last_layer_output[250] + last_layer_output[251] + last_layer_output[252] + last_layer_output[253] + last_layer_output[254] + last_layer_output[255] + last_layer_output[256] + last_layer_output[257] + last_layer_output[258] + last_layer_output[259] + last_layer_output[260] + last_layer_output[261] + last_layer_output[262] + last_layer_output[263] + last_layer_output[264] + last_layer_output[265] + last_layer_output[266] + last_layer_output[267] + last_layer_output[268] + last_layer_output[269] + last_layer_output[270] + last_layer_output[271] + last_layer_output[272] + last_layer_output[273] + last_layer_output[274] + last_layer_output[275] + last_layer_output[276] + last_layer_output[277] + last_layer_output[278] + last_layer_output[279] + last_layer_output[280] + last_layer_output[281] + last_layer_output[282] + last_layer_output[283] + last_layer_output[284] + last_layer_output[285] + last_layer_output[286] + last_layer_output[287] + last_layer_output[288] + last_layer_output[289] + last_layer_output[290] + last_layer_output[291] + last_layer_output[292] + last_layer_output[293] + last_layer_output[294] + last_layer_output[295] + last_layer_output[296] + last_layer_output[297] + last_layer_output[298] + last_layer_output[299] + last_layer_output[300] + last_layer_output[301] + last_layer_output[302] + last_layer_output[303] + last_layer_output[304] + last_layer_output[305] + last_layer_output[306] + last_layer_output[307] + last_layer_output[308] + last_layer_output[309] + last_layer_output[310] + last_layer_output[311] + last_layer_output[312] + last_layer_output[313] + last_layer_output[314] + last_layer_output[315] + last_layer_output[316] + last_layer_output[317] + last_layer_output[318] + last_layer_output[319];
      result[4] <= last_layer_output[320] + last_layer_output[321] + last_layer_output[322] + last_layer_output[323] + last_layer_output[324] + last_layer_output[325] + last_layer_output[326] + last_layer_output[327] + last_layer_output[328] + last_layer_output[329] + last_layer_output[330] + last_layer_output[331] + last_layer_output[332] + last_layer_output[333] + last_layer_output[334] + last_layer_output[335] + last_layer_output[336] + last_layer_output[337] + last_layer_output[338] + last_layer_output[339] + last_layer_output[340] + last_layer_output[341] + last_layer_output[342] + last_layer_output[343] + last_layer_output[344] + last_layer_output[345] + last_layer_output[346] + last_layer_output[347] + last_layer_output[348] + last_layer_output[349] + last_layer_output[350] + last_layer_output[351] + last_layer_output[352] + last_layer_output[353] + last_layer_output[354] + last_layer_output[355] + last_layer_output[356] + last_layer_output[357] + last_layer_output[358] + last_layer_output[359] + last_layer_output[360] + last_layer_output[361] + last_layer_output[362] + last_layer_output[363] + last_layer_output[364] + last_layer_output[365] + last_layer_output[366] + last_layer_output[367] + last_layer_output[368] + last_layer_output[369] + last_layer_output[370] + last_layer_output[371] + last_layer_output[372] + last_layer_output[373] + last_layer_output[374] + last_layer_output[375] + last_layer_output[376] + last_layer_output[377] + last_layer_output[378] + last_layer_output[379] + last_layer_output[380] + last_layer_output[381] + last_layer_output[382] + last_layer_output[383] + last_layer_output[384] + last_layer_output[385] + last_layer_output[386] + last_layer_output[387] + last_layer_output[388] + last_layer_output[389] + last_layer_output[390] + last_layer_output[391] + last_layer_output[392] + last_layer_output[393] + last_layer_output[394] + last_layer_output[395] + last_layer_output[396] + last_layer_output[397] + last_layer_output[398] + last_layer_output[399];
      result[5] <= last_layer_output[400] + last_layer_output[401] + last_layer_output[402] + last_layer_output[403] + last_layer_output[404] + last_layer_output[405] + last_layer_output[406] + last_layer_output[407] + last_layer_output[408] + last_layer_output[409] + last_layer_output[410] + last_layer_output[411] + last_layer_output[412] + last_layer_output[413] + last_layer_output[414] + last_layer_output[415] + last_layer_output[416] + last_layer_output[417] + last_layer_output[418] + last_layer_output[419] + last_layer_output[420] + last_layer_output[421] + last_layer_output[422] + last_layer_output[423] + last_layer_output[424] + last_layer_output[425] + last_layer_output[426] + last_layer_output[427] + last_layer_output[428] + last_layer_output[429] + last_layer_output[430] + last_layer_output[431] + last_layer_output[432] + last_layer_output[433] + last_layer_output[434] + last_layer_output[435] + last_layer_output[436] + last_layer_output[437] + last_layer_output[438] + last_layer_output[439] + last_layer_output[440] + last_layer_output[441] + last_layer_output[442] + last_layer_output[443] + last_layer_output[444] + last_layer_output[445] + last_layer_output[446] + last_layer_output[447] + last_layer_output[448] + last_layer_output[449] + last_layer_output[450] + last_layer_output[451] + last_layer_output[452] + last_layer_output[453] + last_layer_output[454] + last_layer_output[455] + last_layer_output[456] + last_layer_output[457] + last_layer_output[458] + last_layer_output[459] + last_layer_output[460] + last_layer_output[461] + last_layer_output[462] + last_layer_output[463] + last_layer_output[464] + last_layer_output[465] + last_layer_output[466] + last_layer_output[467] + last_layer_output[468] + last_layer_output[469] + last_layer_output[470] + last_layer_output[471] + last_layer_output[472] + last_layer_output[473] + last_layer_output[474] + last_layer_output[475] + last_layer_output[476] + last_layer_output[477] + last_layer_output[478] + last_layer_output[479];
      result[6] <= last_layer_output[480] + last_layer_output[481] + last_layer_output[482] + last_layer_output[483] + last_layer_output[484] + last_layer_output[485] + last_layer_output[486] + last_layer_output[487] + last_layer_output[488] + last_layer_output[489] + last_layer_output[490] + last_layer_output[491] + last_layer_output[492] + last_layer_output[493] + last_layer_output[494] + last_layer_output[495] + last_layer_output[496] + last_layer_output[497] + last_layer_output[498] + last_layer_output[499] + last_layer_output[500] + last_layer_output[501] + last_layer_output[502] + last_layer_output[503] + last_layer_output[504] + last_layer_output[505] + last_layer_output[506] + last_layer_output[507] + last_layer_output[508] + last_layer_output[509] + last_layer_output[510] + last_layer_output[511] + last_layer_output[512] + last_layer_output[513] + last_layer_output[514] + last_layer_output[515] + last_layer_output[516] + last_layer_output[517] + last_layer_output[518] + last_layer_output[519] + last_layer_output[520] + last_layer_output[521] + last_layer_output[522] + last_layer_output[523] + last_layer_output[524] + last_layer_output[525] + last_layer_output[526] + last_layer_output[527] + last_layer_output[528] + last_layer_output[529] + last_layer_output[530] + last_layer_output[531] + last_layer_output[532] + last_layer_output[533] + last_layer_output[534] + last_layer_output[535] + last_layer_output[536] + last_layer_output[537] + last_layer_output[538] + last_layer_output[539] + last_layer_output[540] + last_layer_output[541] + last_layer_output[542] + last_layer_output[543] + last_layer_output[544] + last_layer_output[545] + last_layer_output[546] + last_layer_output[547] + last_layer_output[548] + last_layer_output[549] + last_layer_output[550] + last_layer_output[551] + last_layer_output[552] + last_layer_output[553] + last_layer_output[554] + last_layer_output[555] + last_layer_output[556] + last_layer_output[557] + last_layer_output[558] + last_layer_output[559];
      result[7] <= last_layer_output[560] + last_layer_output[561] + last_layer_output[562] + last_layer_output[563] + last_layer_output[564] + last_layer_output[565] + last_layer_output[566] + last_layer_output[567] + last_layer_output[568] + last_layer_output[569] + last_layer_output[570] + last_layer_output[571] + last_layer_output[572] + last_layer_output[573] + last_layer_output[574] + last_layer_output[575] + last_layer_output[576] + last_layer_output[577] + last_layer_output[578] + last_layer_output[579] + last_layer_output[580] + last_layer_output[581] + last_layer_output[582] + last_layer_output[583] + last_layer_output[584] + last_layer_output[585] + last_layer_output[586] + last_layer_output[587] + last_layer_output[588] + last_layer_output[589] + last_layer_output[590] + last_layer_output[591] + last_layer_output[592] + last_layer_output[593] + last_layer_output[594] + last_layer_output[595] + last_layer_output[596] + last_layer_output[597] + last_layer_output[598] + last_layer_output[599] + last_layer_output[600] + last_layer_output[601] + last_layer_output[602] + last_layer_output[603] + last_layer_output[604] + last_layer_output[605] + last_layer_output[606] + last_layer_output[607] + last_layer_output[608] + last_layer_output[609] + last_layer_output[610] + last_layer_output[611] + last_layer_output[612] + last_layer_output[613] + last_layer_output[614] + last_layer_output[615] + last_layer_output[616] + last_layer_output[617] + last_layer_output[618] + last_layer_output[619] + last_layer_output[620] + last_layer_output[621] + last_layer_output[622] + last_layer_output[623] + last_layer_output[624] + last_layer_output[625] + last_layer_output[626] + last_layer_output[627] + last_layer_output[628] + last_layer_output[629] + last_layer_output[630] + last_layer_output[631] + last_layer_output[632] + last_layer_output[633] + last_layer_output[634] + last_layer_output[635] + last_layer_output[636] + last_layer_output[637] + last_layer_output[638] + last_layer_output[639];
      result[8] <= last_layer_output[640] + last_layer_output[641] + last_layer_output[642] + last_layer_output[643] + last_layer_output[644] + last_layer_output[645] + last_layer_output[646] + last_layer_output[647] + last_layer_output[648] + last_layer_output[649] + last_layer_output[650] + last_layer_output[651] + last_layer_output[652] + last_layer_output[653] + last_layer_output[654] + last_layer_output[655] + last_layer_output[656] + last_layer_output[657] + last_layer_output[658] + last_layer_output[659] + last_layer_output[660] + last_layer_output[661] + last_layer_output[662] + last_layer_output[663] + last_layer_output[664] + last_layer_output[665] + last_layer_output[666] + last_layer_output[667] + last_layer_output[668] + last_layer_output[669] + last_layer_output[670] + last_layer_output[671] + last_layer_output[672] + last_layer_output[673] + last_layer_output[674] + last_layer_output[675] + last_layer_output[676] + last_layer_output[677] + last_layer_output[678] + last_layer_output[679] + last_layer_output[680] + last_layer_output[681] + last_layer_output[682] + last_layer_output[683] + last_layer_output[684] + last_layer_output[685] + last_layer_output[686] + last_layer_output[687] + last_layer_output[688] + last_layer_output[689] + last_layer_output[690] + last_layer_output[691] + last_layer_output[692] + last_layer_output[693] + last_layer_output[694] + last_layer_output[695] + last_layer_output[696] + last_layer_output[697] + last_layer_output[698] + last_layer_output[699] + last_layer_output[700] + last_layer_output[701] + last_layer_output[702] + last_layer_output[703] + last_layer_output[704] + last_layer_output[705] + last_layer_output[706] + last_layer_output[707] + last_layer_output[708] + last_layer_output[709] + last_layer_output[710] + last_layer_output[711] + last_layer_output[712] + last_layer_output[713] + last_layer_output[714] + last_layer_output[715] + last_layer_output[716] + last_layer_output[717] + last_layer_output[718] + last_layer_output[719];
      result[9] <= last_layer_output[720] + last_layer_output[721] + last_layer_output[722] + last_layer_output[723] + last_layer_output[724] + last_layer_output[725] + last_layer_output[726] + last_layer_output[727] + last_layer_output[728] + last_layer_output[729] + last_layer_output[730] + last_layer_output[731] + last_layer_output[732] + last_layer_output[733] + last_layer_output[734] + last_layer_output[735] + last_layer_output[736] + last_layer_output[737] + last_layer_output[738] + last_layer_output[739] + last_layer_output[740] + last_layer_output[741] + last_layer_output[742] + last_layer_output[743] + last_layer_output[744] + last_layer_output[745] + last_layer_output[746] + last_layer_output[747] + last_layer_output[748] + last_layer_output[749] + last_layer_output[750] + last_layer_output[751] + last_layer_output[752] + last_layer_output[753] + last_layer_output[754] + last_layer_output[755] + last_layer_output[756] + last_layer_output[757] + last_layer_output[758] + last_layer_output[759] + last_layer_output[760] + last_layer_output[761] + last_layer_output[762] + last_layer_output[763] + last_layer_output[764] + last_layer_output[765] + last_layer_output[766] + last_layer_output[767] + last_layer_output[768] + last_layer_output[769] + last_layer_output[770] + last_layer_output[771] + last_layer_output[772] + last_layer_output[773] + last_layer_output[774] + last_layer_output[775] + last_layer_output[776] + last_layer_output[777] + last_layer_output[778] + last_layer_output[779] + last_layer_output[780] + last_layer_output[781] + last_layer_output[782] + last_layer_output[783] + last_layer_output[784] + last_layer_output[785] + last_layer_output[786] + last_layer_output[787] + last_layer_output[788] + last_layer_output[789] + last_layer_output[790] + last_layer_output[791] + last_layer_output[792] + last_layer_output[793] + last_layer_output[794] + last_layer_output[795] + last_layer_output[796] + last_layer_output[797] + last_layer_output[798] + last_layer_output[799];
end
      assign y[69:63]=result[0];
      assign y[62:56]=result[1];
      assign y[55:49]=result[2];
      assign y[48:42]=result[3];
      assign y[41:35]=result[4];
      assign y[34:28]=result[5];
      assign y[27:21]=result[6];
      assign y[20:14]=result[7];
      assign y[13:7]=result[8];
      assign y[6:0]=result[9];
endmodule