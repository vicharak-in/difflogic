module logic_network (    input clk,
    input wire [399:0] x,
    output wire [49:0] y
);
      reg [299:0] layer0_out = 0;
      reg [299:0] layer1_out = 0;
      reg [299:0] layer2_out = 0;
      reg [299:0] layer3_out = 0;
      reg [299:0] last_layer_output = 0;
      reg [4:0] result [9:0];
      always @(posedge clk) begin
     layer0_out[0] <= ~(x[106] | x[107]);
     layer0_out[1] <= x[194];
     layer0_out[2] <= ~x[91];
     layer0_out[3] <= x[198];
     layer0_out[4] <= ~x[235];
     layer0_out[5] <= ~(x[181] | x[182]);
     layer0_out[6] <= ~x[189];
     layer0_out[7] <= 1'b0;
     layer0_out[8] <= x[153] | x[154];
     layer0_out[9] <= x[308];
     layer0_out[10] <= ~(x[174] | x[175]);
     layer0_out[11] <= x[193] | x[194];
     layer0_out[12] <= ~(x[76] | x[77]);
     layer0_out[13] <= 1'b1;
     layer0_out[14] <= ~(x[268] | x[269]);
     layer0_out[15] <= ~(x[65] & x[66]);
     layer0_out[16] <= ~(x[107] | x[108]);
     layer0_out[17] <= x[127];
     layer0_out[18] <= ~(x[384] | x[385]);
     layer0_out[19] <= ~x[210] | x[211];
     layer0_out[20] <= x[129] | x[130];
     layer0_out[21] <= ~x[139];
     layer0_out[22] <= ~x[74];
     layer0_out[23] <= x[250] | x[251];
     layer0_out[24] <= 1'b1;
     layer0_out[25] <= 1'b0;
     layer0_out[26] <= x[332] | x[333];
     layer0_out[27] <= ~x[78];
     layer0_out[28] <= ~x[102] | x[101];
     layer0_out[29] <= 1'b0;
     layer0_out[30] <= 1'b0;
     layer0_out[31] <= ~x[177];
     layer0_out[32] <= x[156] | x[157];
     layer0_out[33] <= x[192];
     layer0_out[34] <= x[164] | x[165];
     layer0_out[35] <= x[105] | x[106];
     layer0_out[36] <= x[121] | x[122];
     layer0_out[37] <= ~(x[147] | x[148]);
     layer0_out[38] <= x[5] & ~x[6];
     layer0_out[39] <= ~(x[158] | x[159]);
     layer0_out[40] <= x[216] | x[217];
     layer0_out[41] <= ~(x[82] | x[83]);
     layer0_out[42] <= x[87] | x[88];
     layer0_out[43] <= x[8] | x[9];
     layer0_out[44] <= ~x[12] | x[13];
     layer0_out[45] <= x[241];
     layer0_out[46] <= x[157] | x[158];
     layer0_out[47] <= 1'b0;
     layer0_out[48] <= x[373] & ~x[372];
     layer0_out[49] <= x[316] | x[317];
     layer0_out[50] <= ~(x[378] | x[379]);
     layer0_out[51] <= ~x[27];
     layer0_out[52] <= ~(x[34] | x[35]);
     layer0_out[53] <= ~(x[318] | x[319]);
     layer0_out[54] <= ~(x[354] | x[355]);
     layer0_out[55] <= x[381] & ~x[380];
     layer0_out[56] <= ~x[365];
     layer0_out[57] <= x[288] | x[289];
     layer0_out[58] <= x[30] | x[31];
     layer0_out[59] <= ~(x[151] | x[152]);
     layer0_out[60] <= x[141] | x[142];
     layer0_out[61] <= x[128];
     layer0_out[62] <= x[146] | x[147];
     layer0_out[63] <= x[134];
     layer0_out[64] <= 1'b1;
     layer0_out[65] <= x[144] | x[145];
     layer0_out[66] <= x[382] & ~x[383];
     layer0_out[67] <= x[151];
     layer0_out[68] <= ~x[346];
     layer0_out[69] <= x[275];
     layer0_out[70] <= x[68] | x[69];
     layer0_out[71] <= x[226];
     layer0_out[72] <= 1'b0;
     layer0_out[73] <= x[114];
     layer0_out[74] <= ~x[1];
     layer0_out[75] <= ~x[218];
     layer0_out[76] <= ~x[370];
     layer0_out[77] <= x[83] | x[84];
     layer0_out[78] <= x[160];
     layer0_out[79] <= 1'b1;
     layer0_out[80] <= x[324] | x[325];
     layer0_out[81] <= ~(x[262] | x[263]);
     layer0_out[82] <= x[222] & ~x[223];
     layer0_out[83] <= 1'b0;
     layer0_out[84] <= ~(x[246] | x[247]);
     layer0_out[85] <= ~(x[276] | x[277]);
     layer0_out[86] <= x[230] | x[231];
     layer0_out[87] <= x[273];
     layer0_out[88] <= x[252];
     layer0_out[89] <= ~x[97] | x[98];
     layer0_out[90] <= x[190];
     layer0_out[91] <= 1'b1;
     layer0_out[92] <= x[51];
     layer0_out[93] <= 1'b1;
     layer0_out[94] <= ~x[108];
     layer0_out[95] <= x[61] | x[62];
     layer0_out[96] <= 1'b1;
     layer0_out[97] <= x[160] & x[161];
     layer0_out[98] <= ~(x[166] | x[167]);
     layer0_out[99] <= x[135] | x[136];
     layer0_out[100] <= ~(x[96] | x[97]);
     layer0_out[101] <= ~(x[356] | x[357]);
     layer0_out[102] <= x[291] & ~x[290];
     layer0_out[103] <= 1'b1;
     layer0_out[104] <= ~(x[238] | x[239]);
     layer0_out[105] <= ~(x[183] | x[184]);
     layer0_out[106] <= ~(x[212] | x[213]);
     layer0_out[107] <= ~(x[70] & x[71]);
     layer0_out[108] <= x[336] | x[337];
     layer0_out[109] <= x[293];
     layer0_out[110] <= ~x[86];
     layer0_out[111] <= x[45] | x[46];
     layer0_out[112] <= 1'b0;
     layer0_out[113] <= x[79] & ~x[78];
     layer0_out[114] <= ~x[6] | x[7];
     layer0_out[115] <= ~(x[44] ^ x[45]);
     layer0_out[116] <= x[282] | x[283];
     layer0_out[117] <= ~x[399] | x[398];
     layer0_out[118] <= 1'b0;
     layer0_out[119] <= x[193] & ~x[192];
     layer0_out[120] <= ~(x[236] | x[237]);
     layer0_out[121] <= ~x[11];
     layer0_out[122] <= ~(x[228] | x[229]);
     layer0_out[123] <= ~x[270];
     layer0_out[124] <= ~x[120];
     layer0_out[125] <= ~x[111] | x[112];
     layer0_out[126] <= ~(x[131] | x[132]);
     layer0_out[127] <= x[334] | x[335];
     layer0_out[128] <= x[58] | x[59];
     layer0_out[129] <= x[16];
     layer0_out[130] <= x[13] & ~x[14];
     layer0_out[131] <= ~(x[322] | x[323]);
     layer0_out[132] <= ~(x[340] | x[341]);
     layer0_out[133] <= ~(x[182] | x[183]);
     layer0_out[134] <= x[99] & ~x[98];
     layer0_out[135] <= ~x[117];
     layer0_out[136] <= ~(x[50] & x[51]);
     layer0_out[137] <= ~(x[202] | x[203]);
     layer0_out[138] <= ~(x[56] | x[57]);
     layer0_out[139] <= x[360] | x[361];
     layer0_out[140] <= x[259];
     layer0_out[141] <= ~x[33];
     layer0_out[142] <= ~x[123] | x[122];
     layer0_out[143] <= x[138] | x[139];
     layer0_out[144] <= x[142] | x[143];
     layer0_out[145] <= 1'b0;
     layer0_out[146] <= ~(x[88] | x[89]);
     layer0_out[147] <= ~(x[21] | x[22]);
     layer0_out[148] <= 1'b1;
     layer0_out[149] <= ~x[167];
     layer0_out[150] <= x[279];
     layer0_out[151] <= ~x[2];
     layer0_out[152] <= ~x[133];
     layer0_out[153] <= x[95] ^ x[96];
     layer0_out[154] <= x[314] | x[315];
     layer0_out[155] <= x[342] | x[343];
     layer0_out[156] <= ~x[29];
     layer0_out[157] <= 1'b0;
     layer0_out[158] <= ~(x[362] | x[363]);
     layer0_out[159] <= x[124] | x[125];
     layer0_out[160] <= x[295];
     layer0_out[161] <= x[19] | x[20];
     layer0_out[162] <= x[155] ^ x[156];
     layer0_out[163] <= x[162] | x[163];
     layer0_out[164] <= ~(x[114] & x[115]);
     layer0_out[165] <= ~(x[74] | x[75]);
     layer0_out[166] <= ~x[196];
     layer0_out[167] <= x[67] & x[68];
     layer0_out[168] <= x[84] | x[85];
     layer0_out[169] <= x[70];
     layer0_out[170] <= 1'b0;
     layer0_out[171] <= x[125] | x[126];
     layer0_out[172] <= ~(x[32] & x[33]);
     layer0_out[173] <= ~x[168];
     layer0_out[174] <= ~x[175];
     layer0_out[175] <= x[39] ^ x[40];
     layer0_out[176] <= x[313];
     layer0_out[177] <= ~(x[256] | x[257]);
     layer0_out[178] <= x[187] | x[188];
     layer0_out[179] <= ~x[15];
     layer0_out[180] <= ~x[25];
     layer0_out[181] <= ~(x[171] | x[172]);
     layer0_out[182] <= x[109] | x[110];
     layer0_out[183] <= 1'b1;
     layer0_out[184] <= ~(x[224] | x[225]);
     layer0_out[185] <= ~(x[366] & x[367]);
     layer0_out[186] <= 1'b1;
     layer0_out[187] <= 1'b0;
     layer0_out[188] <= x[352] | x[353];
     layer0_out[189] <= x[163] | x[164];
     layer0_out[190] <= 1'b0;
     layer0_out[191] <= ~(x[184] | x[185]);
     layer0_out[192] <= 1'b0;
     layer0_out[193] <= x[59] | x[60];
     layer0_out[194] <= ~(x[161] | x[162]);
     layer0_out[195] <= x[26] | x[27];
     layer0_out[196] <= 1'b0;
     layer0_out[197] <= 1'b0;
     layer0_out[198] <= x[186] | x[187];
     layer0_out[199] <= x[197] & ~x[196];
     layer0_out[200] <= x[23] | x[24];
     layer0_out[201] <= x[4] & ~x[3];
     layer0_out[202] <= ~x[103];
     layer0_out[203] <= ~x[43];
     layer0_out[204] <= ~(x[81] ^ x[82]);
     layer0_out[205] <= ~(x[358] | x[359]);
     layer0_out[206] <= ~(x[93] | x[94]);
     layer0_out[207] <= ~(x[254] | x[255]);
     layer0_out[208] <= x[130] | x[131];
     layer0_out[209] <= x[181] & ~x[180];
     layer0_out[210] <= x[284] | x[285];
     layer0_out[211] <= 1'b1;
     layer0_out[212] <= x[63];
     layer0_out[213] <= x[176] & ~x[177];
     layer0_out[214] <= ~(x[214] | x[215]);
     layer0_out[215] <= ~(x[396] | x[397]);
     layer0_out[216] <= ~x[26];
     layer0_out[217] <= ~x[54];
     layer0_out[218] <= ~(x[388] | x[389]);
     layer0_out[219] <= x[79] & ~x[80];
     layer0_out[220] <= x[90] | x[91];
     layer0_out[221] <= ~(x[104] | x[105]);
     layer0_out[222] <= ~(x[99] | x[100]);
     layer0_out[223] <= x[172] | x[173];
     layer0_out[224] <= ~x[170];
     layer0_out[225] <= ~(x[152] | x[153]);
     layer0_out[226] <= ~x[339] | x[338];
     layer0_out[227] <= x[326] | x[327];
     layer0_out[228] <= x[248] | x[249];
     layer0_out[229] <= x[126] | x[127];
     layer0_out[230] <= 1'b0;
     layer0_out[231] <= 1'b0;
     layer0_out[232] <= ~x[208];
     layer0_out[233] <= x[296] | x[297];
     layer0_out[234] <= ~(x[115] | x[116]);
     layer0_out[235] <= ~(x[94] | x[95]);
     layer0_out[236] <= ~x[207];
     layer0_out[237] <= x[112] | x[113];
     layer0_out[238] <= ~(x[9] & x[10]);
     layer0_out[239] <= x[72] & ~x[71];
     layer0_out[240] <= x[242] | x[243];
     layer0_out[241] <= x[18] & ~x[17];
     layer0_out[242] <= ~x[116];
     layer0_out[243] <= ~x[110];
     layer0_out[244] <= ~x[31];
     layer0_out[245] <= ~(x[260] & x[261]);
     layer0_out[246] <= 1'b0;
     layer0_out[247] <= ~(x[48] | x[49]);
     layer0_out[248] <= x[66] | x[67];
     layer0_out[249] <= ~(x[386] | x[387]);
     layer0_out[250] <= 1'b0;
     layer0_out[251] <= ~(x[123] | x[124]);
     layer0_out[252] <= ~(x[49] & x[50]);
     layer0_out[253] <= 1'b0;
     layer0_out[254] <= x[280] | x[281];
     layer0_out[255] <= x[320] | x[321];
     layer0_out[256] <= 1'b0;
     layer0_out[257] <= x[204] | x[205];
     layer0_out[258] <= ~(x[350] & x[351]);
     layer0_out[259] <= x[55] & ~x[54];
     layer0_out[260] <= x[145] | x[146];
     layer0_out[261] <= ~x[56];
     layer0_out[262] <= x[149] & ~x[148];
     layer0_out[263] <= x[221];
     layer0_out[264] <= ~x[306];
     layer0_out[265] <= ~x[80] | x[81];
     layer0_out[266] <= x[244] | x[245];
     layer0_out[267] <= x[377];
     layer0_out[268] <= ~(x[188] | x[189]);
     layer0_out[269] <= 1'b1;
     layer0_out[270] <= 1'b0;
     layer0_out[271] <= 1'b0;
     layer0_out[272] <= x[72] & ~x[73];
     layer0_out[273] <= 1'b0;
     layer0_out[274] <= ~x[40] | x[41];
     layer0_out[275] <= x[302] | x[303];
     layer0_out[276] <= ~x[149];
     layer0_out[277] <= x[344] | x[345];
     layer0_out[278] <= ~(x[46] | x[47]);
     layer0_out[279] <= ~(x[137] ^ x[138]);
     layer0_out[280] <= 1'b0;
     layer0_out[281] <= 1'b0;
     layer0_out[282] <= 1'b1;
     layer0_out[283] <= x[197] | x[198];
     layer0_out[284] <= ~(x[185] | x[186]);
     layer0_out[285] <= x[92] | x[93];
     layer0_out[286] <= ~(x[368] & x[369]);
     layer0_out[287] <= x[137];
     layer0_out[288] <= ~(x[36] | x[37]);
     layer0_out[289] <= 1'b0;
     layer0_out[290] <= x[199] | x[200];
     layer0_out[291] <= 1'b1;
     layer0_out[292] <= ~(x[165] | x[166]);
     layer0_out[293] <= 1'b1;
     layer0_out[294] <= x[264] | x[265];
     layer0_out[295] <= x[22];
     layer0_out[296] <= 1'b1;
     layer0_out[297] <= x[38];
     layer0_out[298] <= ~(x[154] | x[155]);
     layer0_out[299] <= x[169] | x[170];
     layer1_out[0] <= ~layer0_out[90];
     layer1_out[1] <= layer0_out[202];
     layer1_out[2] <= layer0_out[47] & ~layer0_out[48];
     layer1_out[3] <= layer0_out[5];
     layer1_out[4] <= ~layer0_out[6];
     layer1_out[5] <= layer0_out[266] | layer0_out[267];
     layer1_out[6] <= ~layer0_out[84];
     layer1_out[7] <= layer0_out[105];
     layer1_out[8] <= ~layer0_out[168];
     layer1_out[9] <= layer0_out[198];
     layer1_out[10] <= layer0_out[133];
     layer1_out[11] <= layer0_out[232] & ~layer0_out[233];
     layer1_out[12] <= ~(layer0_out[189] ^ layer0_out[190]);
     layer1_out[13] <= ~(layer0_out[193] | layer0_out[194]);
     layer1_out[14] <= ~(layer0_out[44] & layer0_out[45]);
     layer1_out[15] <= layer0_out[184];
     layer1_out[16] <= ~(layer0_out[234] | layer0_out[235]);
     layer1_out[17] <= ~layer0_out[258];
     layer1_out[18] <= ~layer0_out[101] | layer0_out[100];
     layer1_out[19] <= layer0_out[30] | layer0_out[31];
     layer1_out[20] <= ~(layer0_out[278] & layer0_out[279]);
     layer1_out[21] <= layer0_out[28] & ~layer0_out[29];
     layer1_out[22] <= layer0_out[288];
     layer1_out[23] <= ~layer0_out[214] | layer0_out[215];
     layer1_out[24] <= ~(layer0_out[36] | layer0_out[37]);
     layer1_out[25] <= layer0_out[107] & ~layer0_out[108];
     layer1_out[26] <= 1'b1;
     layer1_out[27] <= ~layer0_out[59];
     layer1_out[28] <= layer0_out[39];
     layer1_out[29] <= ~(layer0_out[114] | layer0_out[115]);
     layer1_out[30] <= ~layer0_out[127];
     layer1_out[31] <= ~layer0_out[298] | layer0_out[297];
     layer1_out[32] <= ~layer0_out[98];
     layer1_out[33] <= layer0_out[141];
     layer1_out[34] <= ~layer0_out[26];
     layer1_out[35] <= 1'b1;
     layer1_out[36] <= layer0_out[98] & ~layer0_out[99];
     layer1_out[37] <= ~layer0_out[270] | layer0_out[269];
     layer1_out[38] <= layer0_out[295] | layer0_out[296];
     layer1_out[39] <= 1'b0;
     layer1_out[40] <= layer0_out[161] & ~layer0_out[162];
     layer1_out[41] <= ~layer0_out[17];
     layer1_out[42] <= layer0_out[249];
     layer1_out[43] <= layer0_out[256] & ~layer0_out[255];
     layer1_out[44] <= layer0_out[277] | layer0_out[278];
     layer1_out[45] <= 1'b0;
     layer1_out[46] <= ~layer0_out[159];
     layer1_out[47] <= ~(layer0_out[104] & layer0_out[105]);
     layer1_out[48] <= 1'b1;
     layer1_out[49] <= layer0_out[120];
     layer1_out[50] <= layer0_out[53] & layer0_out[54];
     layer1_out[51] <= ~(layer0_out[175] | layer0_out[176]);
     layer1_out[52] <= ~layer0_out[198];
     layer1_out[53] <= ~(layer0_out[13] ^ layer0_out[14]);
     layer1_out[54] <= layer0_out[54];
     layer1_out[55] <= ~layer0_out[119] | layer0_out[118];
     layer1_out[56] <= ~layer0_out[126];
     layer1_out[57] <= layer0_out[123] & ~layer0_out[124];
     layer1_out[58] <= layer0_out[254] | layer0_out[255];
     layer1_out[59] <= layer0_out[135] | layer0_out[136];
     layer1_out[60] <= 1'b1;
     layer1_out[61] <= ~layer0_out[280];
     layer1_out[62] <= layer0_out[58];
     layer1_out[63] <= 1'b1;
     layer1_out[64] <= layer0_out[260];
     layer1_out[65] <= layer0_out[257];
     layer1_out[66] <= ~layer0_out[62] | layer0_out[63];
     layer1_out[67] <= layer0_out[126];
     layer1_out[68] <= layer0_out[240];
     layer1_out[69] <= ~(layer0_out[210] ^ layer0_out[211]);
     layer1_out[70] <= ~layer0_out[41] | layer0_out[40];
     layer1_out[71] <= ~layer0_out[122];
     layer1_out[72] <= ~layer0_out[208];
     layer1_out[73] <= layer0_out[24] ^ layer0_out[25];
     layer1_out[74] <= layer0_out[116];
     layer1_out[75] <= ~layer0_out[120] | layer0_out[121];
     layer1_out[76] <= layer0_out[56] & ~layer0_out[55];
     layer1_out[77] <= layer0_out[101] | layer0_out[102];
     layer1_out[78] <= layer0_out[75] & ~layer0_out[76];
     layer1_out[79] <= layer0_out[48] & layer0_out[49];
     layer1_out[80] <= ~layer0_out[143];
     layer1_out[81] <= ~layer0_out[111];
     layer1_out[82] <= ~layer0_out[232];
     layer1_out[83] <= ~layer0_out[185];
     layer1_out[84] <= ~layer0_out[110] | layer0_out[111];
     layer1_out[85] <= layer0_out[92];
     layer1_out[86] <= 1'b1;
     layer1_out[87] <= ~(layer0_out[294] | layer0_out[295]);
     layer1_out[88] <= 1'b1;
     layer1_out[89] <= ~layer0_out[266];
     layer1_out[90] <= ~(layer0_out[227] & layer0_out[228]);
     layer1_out[91] <= layer0_out[206] & ~layer0_out[205];
     layer1_out[92] <= layer0_out[144] & layer0_out[145];
     layer1_out[93] <= layer0_out[92];
     layer1_out[94] <= layer0_out[283];
     layer1_out[95] <= ~layer0_out[133];
     layer1_out[96] <= layer0_out[130] | layer0_out[131];
     layer1_out[97] <= layer0_out[287] | layer0_out[288];
     layer1_out[98] <= ~layer0_out[261] | layer0_out[262];
     layer1_out[99] <= ~layer0_out[222] | layer0_out[223];
     layer1_out[100] <= ~layer0_out[10] | layer0_out[11];
     layer1_out[101] <= layer0_out[56] | layer0_out[57];
     layer1_out[102] <= layer0_out[290];
     layer1_out[103] <= ~layer0_out[207];
     layer1_out[104] <= layer0_out[177] & ~layer0_out[178];
     layer1_out[105] <= layer0_out[67] | layer0_out[68];
     layer1_out[106] <= layer0_out[281] & ~layer0_out[282];
     layer1_out[107] <= layer0_out[200];
     layer1_out[108] <= ~layer0_out[27] | layer0_out[26];
     layer1_out[109] <= ~layer0_out[248] | layer0_out[247];
     layer1_out[110] <= layer0_out[109];
     layer1_out[111] <= layer0_out[0];
     layer1_out[112] <= ~(layer0_out[147] ^ layer0_out[148]);
     layer1_out[113] <= layer0_out[238];
     layer1_out[114] <= layer0_out[220] & ~layer0_out[219];
     layer1_out[115] <= ~layer0_out[236];
     layer1_out[116] <= ~layer0_out[81] | layer0_out[82];
     layer1_out[117] <= layer0_out[221];
     layer1_out[118] <= layer0_out[93] | layer0_out[94];
     layer1_out[119] <= layer0_out[292];
     layer1_out[120] <= layer0_out[280] & ~layer0_out[279];
     layer1_out[121] <= layer0_out[220] & layer0_out[221];
     layer1_out[122] <= layer0_out[63] | layer0_out[64];
     layer1_out[123] <= layer0_out[286];
     layer1_out[124] <= layer0_out[140] & layer0_out[141];
     layer1_out[125] <= layer0_out[267] | layer0_out[268];
     layer1_out[126] <= layer0_out[88] & layer0_out[89];
     layer1_out[127] <= ~layer0_out[176];
     layer1_out[128] <= layer0_out[299];
     layer1_out[129] <= ~layer0_out[202];
     layer1_out[130] <= layer0_out[271] & layer0_out[272];
     layer1_out[131] <= ~layer0_out[110] | layer0_out[109];
     layer1_out[132] <= ~layer0_out[242] | layer0_out[243];
     layer1_out[133] <= ~(layer0_out[35] | layer0_out[36]);
     layer1_out[134] <= ~(layer0_out[128] | layer0_out[129]);
     layer1_out[135] <= layer0_out[1];
     layer1_out[136] <= ~layer0_out[181];
     layer1_out[137] <= layer0_out[62];
     layer1_out[138] <= ~layer0_out[65];
     layer1_out[139] <= layer0_out[72] & layer0_out[73];
     layer1_out[140] <= ~(layer0_out[148] & layer0_out[149]);
     layer1_out[141] <= layer0_out[163] & ~layer0_out[162];
     layer1_out[142] <= 1'b1;
     layer1_out[143] <= ~layer0_out[12];
     layer1_out[144] <= ~layer0_out[100] | layer0_out[99];
     layer1_out[145] <= layer0_out[166];
     layer1_out[146] <= layer0_out[290];
     layer1_out[147] <= layer0_out[65];
     layer1_out[148] <= ~(layer0_out[192] & layer0_out[193]);
     layer1_out[149] <= ~layer0_out[247];
     layer1_out[150] <= layer0_out[46];
     layer1_out[151] <= ~layer0_out[37];
     layer1_out[152] <= layer0_out[81];
     layer1_out[153] <= 1'b1;
     layer1_out[154] <= layer0_out[129] & layer0_out[130];
     layer1_out[155] <= layer0_out[8] | layer0_out[9];
     layer1_out[156] <= ~layer0_out[166] | layer0_out[165];
     layer1_out[157] <= ~(layer0_out[174] | layer0_out[175]);
     layer1_out[158] <= layer0_out[249];
     layer1_out[159] <= 1'b1;
     layer1_out[160] <= layer0_out[139];
     layer1_out[161] <= ~layer0_out[151] | layer0_out[150];
     layer1_out[162] <= ~layer0_out[114];
     layer1_out[163] <= ~(layer0_out[212] ^ layer0_out[213]);
     layer1_out[164] <= layer0_out[189] & ~layer0_out[188];
     layer1_out[165] <= layer0_out[31] | layer0_out[32];
     layer1_out[166] <= 1'b1;
     layer1_out[167] <= layer0_out[13];
     layer1_out[168] <= layer0_out[227];
     layer1_out[169] <= layer0_out[137];
     layer1_out[170] <= layer0_out[51] | layer0_out[52];
     layer1_out[171] <= ~layer0_out[163] | layer0_out[164];
     layer1_out[172] <= layer0_out[42] ^ layer0_out[43];
     layer1_out[173] <= layer0_out[179] ^ layer0_out[180];
     layer1_out[174] <= layer0_out[276];
     layer1_out[175] <= layer0_out[224];
     layer1_out[176] <= ~(layer0_out[15] & layer0_out[16]);
     layer1_out[177] <= layer0_out[86] & ~layer0_out[87];
     layer1_out[178] <= layer0_out[154] | layer0_out[155];
     layer1_out[179] <= ~(layer0_out[187] | layer0_out[188]);
     layer1_out[180] <= layer0_out[144];
     layer1_out[181] <= layer0_out[113];
     layer1_out[182] <= ~layer0_out[214] | layer0_out[213];
     layer1_out[183] <= 1'b1;
     layer1_out[184] <= 1'b0;
     layer1_out[185] <= layer0_out[194] & layer0_out[195];
     layer1_out[186] <= ~layer0_out[211];
     layer1_out[187] <= layer0_out[217] & ~layer0_out[218];
     layer1_out[188] <= ~layer0_out[234] | layer0_out[233];
     layer1_out[189] <= layer0_out[236];
     layer1_out[190] <= ~layer0_out[264];
     layer1_out[191] <= ~layer0_out[158];
     layer1_out[192] <= ~layer0_out[137];
     layer1_out[193] <= ~(layer0_out[122] & layer0_out[123]);
     layer1_out[194] <= ~layer0_out[103];
     layer1_out[195] <= ~layer0_out[251];
     layer1_out[196] <= layer0_out[3] & ~layer0_out[4];
     layer1_out[197] <= ~(layer0_out[20] & layer0_out[21]);
     layer1_out[198] <= ~layer0_out[238] | layer0_out[237];
     layer1_out[199] <= 1'b1;
     layer1_out[200] <= ~layer0_out[218];
     layer1_out[201] <= layer0_out[196] & layer0_out[197];
     layer1_out[202] <= 1'b1;
     layer1_out[203] <= layer0_out[85];
     layer1_out[204] <= 1'b1;
     layer1_out[205] <= layer0_out[181] & layer0_out[182];
     layer1_out[206] <= layer0_out[200] | layer0_out[201];
     layer1_out[207] <= layer0_out[156] & ~layer0_out[155];
     layer1_out[208] <= ~layer0_out[15] | layer0_out[14];
     layer1_out[209] <= layer0_out[286];
     layer1_out[210] <= layer0_out[69];
     layer1_out[211] <= ~(layer0_out[216] & layer0_out[217]);
     layer1_out[212] <= ~layer0_out[0] | layer0_out[1];
     layer1_out[213] <= 1'b1;
     layer1_out[214] <= ~layer0_out[116];
     layer1_out[215] <= layer0_out[2] & ~layer0_out[3];
     layer1_out[216] <= ~(layer0_out[224] | layer0_out[225]);
     layer1_out[217] <= layer0_out[49] & layer0_out[50];
     layer1_out[218] <= 1'b0;
     layer1_out[219] <= layer0_out[283] | layer0_out[284];
     layer1_out[220] <= layer0_out[228] | layer0_out[229];
     layer1_out[221] <= layer0_out[50] & ~layer0_out[51];
     layer1_out[222] <= 1'b1;
     layer1_out[223] <= ~layer0_out[245] | layer0_out[244];
     layer1_out[224] <= ~layer0_out[284];
     layer1_out[225] <= layer0_out[124] | layer0_out[125];
     layer1_out[226] <= layer0_out[80];
     layer1_out[227] <= ~layer0_out[52] | layer0_out[53];
     layer1_out[228] <= layer0_out[23];
     layer1_out[229] <= ~(layer0_out[59] & layer0_out[60]);
     layer1_out[230] <= layer0_out[210];
     layer1_out[231] <= ~layer0_out[76];
     layer1_out[232] <= ~layer0_out[154];
     layer1_out[233] <= ~layer0_out[74] | layer0_out[73];
     layer1_out[234] <= ~layer0_out[18];
     layer1_out[235] <= ~layer0_out[184];
     layer1_out[236] <= layer0_out[103] & ~layer0_out[104];
     layer1_out[237] <= layer0_out[147] & ~layer0_out[146];
     layer1_out[238] <= ~layer0_out[88];
     layer1_out[239] <= ~(layer0_out[215] & layer0_out[216]);
     layer1_out[240] <= layer0_out[106];
     layer1_out[241] <= layer0_out[187];
     layer1_out[242] <= ~layer0_out[275];
     layer1_out[243] <= layer0_out[171];
     layer1_out[244] <= layer0_out[196] & ~layer0_out[195];
     layer1_out[245] <= ~layer0_out[8];
     layer1_out[246] <= 1'b1;
     layer1_out[247] <= layer0_out[169] | layer0_out[170];
     layer1_out[248] <= ~(layer0_out[241] ^ layer0_out[242]);
     layer1_out[249] <= ~layer0_out[229];
     layer1_out[250] <= ~(layer0_out[90] & layer0_out[91]);
     layer1_out[251] <= layer0_out[84] & layer0_out[85];
     layer1_out[252] <= ~layer0_out[168];
     layer1_out[253] <= ~(layer0_out[160] ^ layer0_out[161]);
     layer1_out[254] <= layer0_out[243] & ~layer0_out[244];
     layer1_out[255] <= ~(layer0_out[29] & layer0_out[30]);
     layer1_out[256] <= layer0_out[131] & layer0_out[132];
     layer1_out[257] <= 1'b1;
     layer1_out[258] <= layer0_out[263];
     layer1_out[259] <= layer0_out[149];
     layer1_out[260] <= ~(layer0_out[74] | layer0_out[75]);
     layer1_out[261] <= ~layer0_out[79];
     layer1_out[262] <= layer0_out[240] & ~layer0_out[241];
     layer1_out[263] <= layer0_out[292];
     layer1_out[264] <= ~layer0_out[32] | layer0_out[33];
     layer1_out[265] <= ~layer0_out[34];
     layer1_out[266] <= layer0_out[23];
     layer1_out[267] <= layer0_out[257] & layer0_out[258];
     layer1_out[268] <= layer0_out[297] & ~layer0_out[296];
     layer1_out[269] <= ~layer0_out[146];
     layer1_out[270] <= 1'b1;
     layer1_out[271] <= ~layer0_out[264] | layer0_out[263];
     layer1_out[272] <= ~layer0_out[260];
     layer1_out[273] <= layer0_out[95];
     layer1_out[274] <= ~layer0_out[191];
     layer1_out[275] <= ~layer0_out[60];
     layer1_out[276] <= ~layer0_out[159];
     layer1_out[277] <= layer0_out[19];
     layer1_out[278] <= ~layer0_out[277];
     layer1_out[279] <= 1'b0;
     layer1_out[280] <= layer0_out[173];
     layer1_out[281] <= ~(layer0_out[21] & layer0_out[22]);
     layer1_out[282] <= ~layer0_out[138] | layer0_out[139];
     layer1_out[283] <= layer0_out[251];
     layer1_out[284] <= layer0_out[152];
     layer1_out[285] <= layer0_out[294];
     layer1_out[286] <= layer0_out[71];
     layer1_out[287] <= ~layer0_out[34];
     layer1_out[288] <= ~layer0_out[208] | layer0_out[209];
     layer1_out[289] <= ~layer0_out[77];
     layer1_out[290] <= ~layer0_out[172];
     layer1_out[291] <= ~(layer0_out[43] | layer0_out[44]);
     layer1_out[292] <= ~(layer0_out[9] & layer0_out[10]);
     layer1_out[293] <= layer0_out[66] | layer0_out[67];
     layer1_out[294] <= ~layer0_out[273] | layer0_out[272];
     layer1_out[295] <= ~(layer0_out[190] | layer0_out[191]);
     layer1_out[296] <= layer0_out[152] & ~layer0_out[153];
     layer1_out[297] <= 1'b1;
     layer1_out[298] <= ~layer0_out[268];
     layer1_out[299] <= layer0_out[205] & ~layer0_out[204];
     layer2_out[0] <= layer1_out[255] & ~layer1_out[254];
     layer2_out[1] <= layer1_out[155];
     layer2_out[2] <= ~layer1_out[38];
     layer2_out[3] <= ~layer1_out[128] | layer1_out[129];
     layer2_out[4] <= ~layer1_out[283] | layer1_out[282];
     layer2_out[5] <= ~layer1_out[174];
     layer2_out[6] <= layer1_out[86];
     layer2_out[7] <= ~layer1_out[44];
     layer2_out[8] <= layer1_out[0];
     layer2_out[9] <= ~layer1_out[151];
     layer2_out[10] <= layer1_out[218];
     layer2_out[11] <= layer1_out[276];
     layer2_out[12] <= ~layer1_out[195];
     layer2_out[13] <= layer1_out[131] | layer1_out[132];
     layer2_out[14] <= layer1_out[28] & ~layer1_out[27];
     layer2_out[15] <= layer1_out[118] & layer1_out[119];
     layer2_out[16] <= ~layer1_out[171];
     layer2_out[17] <= layer1_out[150];
     layer2_out[18] <= layer1_out[182];
     layer2_out[19] <= layer1_out[123];
     layer2_out[20] <= 1'b0;
     layer2_out[21] <= layer1_out[25];
     layer2_out[22] <= ~layer1_out[65] | layer1_out[66];
     layer2_out[23] <= ~layer1_out[183];
     layer2_out[24] <= ~layer1_out[133];
     layer2_out[25] <= ~layer1_out[190];
     layer2_out[26] <= layer1_out[136] & ~layer1_out[135];
     layer2_out[27] <= ~layer1_out[203];
     layer2_out[28] <= layer1_out[156];
     layer2_out[29] <= ~layer1_out[169];
     layer2_out[30] <= layer1_out[147] ^ layer1_out[148];
     layer2_out[31] <= ~layer1_out[17];
     layer2_out[32] <= ~layer1_out[41];
     layer2_out[33] <= ~layer1_out[113] | layer1_out[114];
     layer2_out[34] <= layer1_out[140];
     layer2_out[35] <= ~layer1_out[196] | layer1_out[197];
     layer2_out[36] <= ~layer1_out[175];
     layer2_out[37] <= ~layer1_out[256];
     layer2_out[38] <= layer1_out[292];
     layer2_out[39] <= ~layer1_out[67] | layer1_out[68];
     layer2_out[40] <= layer1_out[249] | layer1_out[250];
     layer2_out[41] <= ~layer1_out[104];
     layer2_out[42] <= ~layer1_out[237];
     layer2_out[43] <= ~layer1_out[56];
     layer2_out[44] <= layer1_out[250];
     layer2_out[45] <= layer1_out[278] | layer1_out[279];
     layer2_out[46] <= ~layer1_out[189] | layer1_out[190];
     layer2_out[47] <= layer1_out[39] & layer1_out[40];
     layer2_out[48] <= layer1_out[105] ^ layer1_out[106];
     layer2_out[49] <= ~layer1_out[251];
     layer2_out[50] <= layer1_out[227];
     layer2_out[51] <= layer1_out[71];
     layer2_out[52] <= layer1_out[200] & layer1_out[201];
     layer2_out[53] <= ~layer1_out[66];
     layer2_out[54] <= ~layer1_out[59];
     layer2_out[55] <= ~layer1_out[131];
     layer2_out[56] <= layer1_out[143] | layer1_out[144];
     layer2_out[57] <= ~layer1_out[127] | layer1_out[126];
     layer2_out[58] <= layer1_out[160] | layer1_out[161];
     layer2_out[59] <= ~(layer1_out[172] | layer1_out[173]);
     layer2_out[60] <= ~layer1_out[243];
     layer2_out[61] <= ~layer1_out[74];
     layer2_out[62] <= ~layer1_out[3];
     layer2_out[63] <= ~layer1_out[137] | layer1_out[136];
     layer2_out[64] <= layer1_out[146];
     layer2_out[65] <= ~layer1_out[266];
     layer2_out[66] <= ~layer1_out[231] | layer1_out[232];
     layer2_out[67] <= layer1_out[249] & ~layer1_out[248];
     layer2_out[68] <= layer1_out[121];
     layer2_out[69] <= layer1_out[37] & ~layer1_out[36];
     layer2_out[70] <= ~layer1_out[260];
     layer2_out[71] <= ~layer1_out[149];
     layer2_out[72] <= ~layer1_out[205];
     layer2_out[73] <= layer1_out[215];
     layer2_out[74] <= layer1_out[127] & layer1_out[128];
     layer2_out[75] <= ~layer1_out[207];
     layer2_out[76] <= ~layer1_out[23];
     layer2_out[77] <= layer1_out[197];
     layer2_out[78] <= ~(layer1_out[193] & layer1_out[194]);
     layer2_out[79] <= layer1_out[225] & ~layer1_out[226];
     layer2_out[80] <= ~layer1_out[290];
     layer2_out[81] <= layer1_out[179] | layer1_out[180];
     layer2_out[82] <= ~layer1_out[48];
     layer2_out[83] <= layer1_out[63] ^ layer1_out[64];
     layer2_out[84] <= layer1_out[223];
     layer2_out[85] <= ~layer1_out[138] | layer1_out[137];
     layer2_out[86] <= ~(layer1_out[98] | layer1_out[99]);
     layer2_out[87] <= layer1_out[60] | layer1_out[61];
     layer2_out[88] <= ~layer1_out[198];
     layer2_out[89] <= layer1_out[24];
     layer2_out[90] <= ~layer1_out[195];
     layer2_out[91] <= layer1_out[183] | layer1_out[184];
     layer2_out[92] <= layer1_out[295];
     layer2_out[93] <= 1'b0;
     layer2_out[94] <= layer1_out[88] & ~layer1_out[89];
     layer2_out[95] <= layer1_out[272];
     layer2_out[96] <= ~layer1_out[111];
     layer2_out[97] <= ~layer1_out[252];
     layer2_out[98] <= layer1_out[84];
     layer2_out[99] <= layer1_out[176] | layer1_out[177];
     layer2_out[100] <= layer1_out[154] & ~layer1_out[153];
     layer2_out[101] <= layer1_out[176] & ~layer1_out[175];
     layer2_out[102] <= layer1_out[259];
     layer2_out[103] <= layer1_out[31];
     layer2_out[104] <= layer1_out[163];
     layer2_out[105] <= layer1_out[152] & layer1_out[153];
     layer2_out[106] <= ~layer1_out[65];
     layer2_out[107] <= 1'b0;
     layer2_out[108] <= ~(layer1_out[45] ^ layer1_out[46]);
     layer2_out[109] <= ~layer1_out[8] | layer1_out[9];
     layer2_out[110] <= ~layer1_out[232];
     layer2_out[111] <= ~layer1_out[178];
     layer2_out[112] <= layer1_out[289] & ~layer1_out[288];
     layer2_out[113] <= 1'b1;
     layer2_out[114] <= ~(layer1_out[241] ^ layer1_out[242]);
     layer2_out[115] <= ~layer1_out[203];
     layer2_out[116] <= layer1_out[91] & layer1_out[92];
     layer2_out[117] <= ~(layer1_out[226] ^ layer1_out[227]);
     layer2_out[118] <= layer1_out[97];
     layer2_out[119] <= ~(layer1_out[236] & layer1_out[237]);
     layer2_out[120] <= ~layer1_out[62];
     layer2_out[121] <= ~layer1_out[219] | layer1_out[218];
     layer2_out[122] <= ~(layer1_out[245] ^ layer1_out[246]);
     layer2_out[123] <= layer1_out[68] | layer1_out[69];
     layer2_out[124] <= ~layer1_out[185];
     layer2_out[125] <= layer1_out[158];
     layer2_out[126] <= ~layer1_out[298];
     layer2_out[127] <= ~layer1_out[234];
     layer2_out[128] <= layer1_out[19] & ~layer1_out[20];
     layer2_out[129] <= layer1_out[42] & ~layer1_out[43];
     layer2_out[130] <= layer1_out[164];
     layer2_out[131] <= ~layer1_out[15];
     layer2_out[132] <= layer1_out[44];
     layer2_out[133] <= ~layer1_out[171];
     layer2_out[134] <= layer1_out[116] | layer1_out[117];
     layer2_out[135] <= layer1_out[52] & ~layer1_out[53];
     layer2_out[136] <= layer1_out[242];
     layer2_out[137] <= layer1_out[118];
     layer2_out[138] <= layer1_out[266] & ~layer1_out[267];
     layer2_out[139] <= layer1_out[170];
     layer2_out[140] <= layer1_out[209];
     layer2_out[141] <= layer1_out[144];
     layer2_out[142] <= ~layer1_out[110];
     layer2_out[143] <= layer1_out[158] & layer1_out[159];
     layer2_out[144] <= ~layer1_out[220] | layer1_out[221];
     layer2_out[145] <= ~layer1_out[224];
     layer2_out[146] <= layer1_out[210] & layer1_out[211];
     layer2_out[147] <= layer1_out[200];
     layer2_out[148] <= layer1_out[57];
     layer2_out[149] <= ~(layer1_out[54] & layer1_out[55]);
     layer2_out[150] <= ~layer1_out[264];
     layer2_out[151] <= layer1_out[115];
     layer2_out[152] <= layer1_out[273] ^ layer1_out[274];
     layer2_out[153] <= layer1_out[33];
     layer2_out[154] <= ~layer1_out[138];
     layer2_out[155] <= layer1_out[280];
     layer2_out[156] <= ~layer1_out[28];
     layer2_out[157] <= layer1_out[188];
     layer2_out[158] <= layer1_out[155] & ~layer1_out[154];
     layer2_out[159] <= ~layer1_out[36];
     layer2_out[160] <= layer1_out[287] | layer1_out[288];
     layer2_out[161] <= ~layer1_out[267];
     layer2_out[162] <= 1'b0;
     layer2_out[163] <= layer1_out[10] & ~layer1_out[11];
     layer2_out[164] <= ~layer1_out[221];
     layer2_out[165] <= ~(layer1_out[163] | layer1_out[164]);
     layer2_out[166] <= layer1_out[97];
     layer2_out[167] <= layer1_out[191] | layer1_out[192];
     layer2_out[168] <= layer1_out[113];
     layer2_out[169] <= ~layer1_out[87];
     layer2_out[170] <= layer1_out[207];
     layer2_out[171] <= ~layer1_out[278];
     layer2_out[172] <= layer1_out[160];
     layer2_out[173] <= layer1_out[100];
     layer2_out[174] <= ~layer1_out[240];
     layer2_out[175] <= layer1_out[290];
     layer2_out[176] <= ~(layer1_out[292] & layer1_out[293]);
     layer2_out[177] <= ~layer1_out[216];
     layer2_out[178] <= ~layer1_out[296] | layer1_out[295];
     layer2_out[179] <= layer1_out[93];
     layer2_out[180] <= layer1_out[233] & ~layer1_out[234];
     layer2_out[181] <= layer1_out[50] & layer1_out[51];
     layer2_out[182] <= layer1_out[16] & ~layer1_out[15];
     layer2_out[183] <= ~layer1_out[230];
     layer2_out[184] <= layer1_out[13];
     layer2_out[185] <= ~(layer1_out[89] & layer1_out[90]);
     layer2_out[186] <= layer1_out[52] & ~layer1_out[51];
     layer2_out[187] <= ~layer1_out[209];
     layer2_out[188] <= ~layer1_out[32];
     layer2_out[189] <= layer1_out[293] & ~layer1_out[294];
     layer2_out[190] <= layer1_out[287] & ~layer1_out[286];
     layer2_out[191] <= layer1_out[109] & ~layer1_out[108];
     layer2_out[192] <= ~layer1_out[123] | layer1_out[124];
     layer2_out[193] <= layer1_out[47];
     layer2_out[194] <= layer1_out[133];
     layer2_out[195] <= 1'b0;
     layer2_out[196] <= layer1_out[6];
     layer2_out[197] <= ~(layer1_out[134] & layer1_out[135]);
     layer2_out[198] <= ~layer1_out[72] | layer1_out[71];
     layer2_out[199] <= layer1_out[3] & ~layer1_out[4];
     layer2_out[200] <= layer1_out[165] | layer1_out[166];
     layer2_out[201] <= layer1_out[62] ^ layer1_out[63];
     layer2_out[202] <= ~layer1_out[70];
     layer2_out[203] <= layer1_out[235];
     layer2_out[204] <= ~layer1_out[74];
     layer2_out[205] <= ~layer1_out[193];
     layer2_out[206] <= layer1_out[85];
     layer2_out[207] <= layer1_out[214] & ~layer1_out[213];
     layer2_out[208] <= ~layer1_out[298];
     layer2_out[209] <= ~(layer1_out[148] & layer1_out[149]);
     layer2_out[210] <= layer1_out[260] & layer1_out[261];
     layer2_out[211] <= layer1_out[253] & layer1_out[254];
     layer2_out[212] <= ~(layer1_out[262] | layer1_out[263]);
     layer2_out[213] <= layer1_out[78];
     layer2_out[214] <= layer1_out[142] & ~layer1_out[143];
     layer2_out[215] <= layer1_out[94];
     layer2_out[216] <= layer1_out[268] & ~layer1_out[269];
     layer2_out[217] <= layer1_out[187];
     layer2_out[218] <= layer1_out[34];
     layer2_out[219] <= 1'b1;
     layer2_out[220] <= layer1_out[125];
     layer2_out[221] <= ~layer1_out[101] | layer1_out[102];
     layer2_out[222] <= ~layer1_out[141];
     layer2_out[223] <= ~(layer1_out[124] | layer1_out[125]);
     layer2_out[224] <= 1'b0;
     layer2_out[225] <= ~layer1_out[280];
     layer2_out[226] <= ~(layer1_out[146] | layer1_out[147]);
     layer2_out[227] <= 1'b0;
     layer2_out[228] <= layer1_out[56];
     layer2_out[229] <= layer1_out[40] ^ layer1_out[41];
     layer2_out[230] <= layer1_out[104];
     layer2_out[231] <= ~layer1_out[229];
     layer2_out[232] <= ~(layer1_out[0] | layer1_out[2]);
     layer2_out[233] <= ~layer1_out[1];
     layer2_out[234] <= layer1_out[257] & layer1_out[258];
     layer2_out[235] <= layer1_out[81];
     layer2_out[236] <= layer1_out[167];
     layer2_out[237] <= layer1_out[121] & ~layer1_out[120];
     layer2_out[238] <= ~layer1_out[7] | layer1_out[6];
     layer2_out[239] <= ~layer1_out[27];
     layer2_out[240] <= layer1_out[214] & layer1_out[215];
     layer2_out[241] <= ~layer1_out[5];
     layer2_out[242] <= layer1_out[19];
     layer2_out[243] <= layer1_out[9] & layer1_out[10];
     layer2_out[244] <= layer1_out[275] & ~layer1_out[274];
     layer2_out[245] <= ~layer1_out[245];
     layer2_out[246] <= layer1_out[206];
     layer2_out[247] <= ~(layer1_out[46] | layer1_out[47]);
     layer2_out[248] <= layer1_out[283];
     layer2_out[249] <= layer1_out[50];
     layer2_out[250] <= layer1_out[262];
     layer2_out[251] <= layer1_out[100];
     layer2_out[252] <= layer1_out[23] ^ layer1_out[24];
     layer2_out[253] <= layer1_out[239];
     layer2_out[254] <= layer1_out[7];
     layer2_out[255] <= 1'b0;
     layer2_out[256] <= ~layer1_out[230];
     layer2_out[257] <= ~(layer1_out[94] | layer1_out[95]);
     layer2_out[258] <= ~layer1_out[178] | layer1_out[179];
     layer2_out[259] <= layer1_out[272];
     layer2_out[260] <= 1'b0;
     layer2_out[261] <= ~(layer1_out[119] ^ layer1_out[120]);
     layer2_out[262] <= ~layer1_out[219];
     layer2_out[263] <= 1'b1;
     layer2_out[264] <= layer1_out[212];
     layer2_out[265] <= ~layer1_out[296];
     layer2_out[266] <= layer1_out[58];
     layer2_out[267] <= layer1_out[82] | layer1_out[83];
     layer2_out[268] <= layer1_out[12] & ~layer1_out[11];
     layer2_out[269] <= ~layer1_out[81];
     layer2_out[270] <= ~layer1_out[285];
     layer2_out[271] <= ~layer1_out[116];
     layer2_out[272] <= ~layer1_out[78];
     layer2_out[273] <= layer1_out[246] ^ layer1_out[247];
     layer2_out[274] <= ~layer1_out[75];
     layer2_out[275] <= ~(layer1_out[102] | layer1_out[103]);
     layer2_out[276] <= layer1_out[22];
     layer2_out[277] <= ~(layer1_out[76] & layer1_out[77]);
     layer2_out[278] <= layer1_out[275] & layer1_out[276];
     layer2_out[279] <= layer1_out[255] & ~layer1_out[256];
     layer2_out[280] <= layer1_out[223];
     layer2_out[281] <= layer1_out[168];
     layer2_out[282] <= ~layer1_out[112];
     layer2_out[283] <= layer1_out[281] | layer1_out[282];
     layer2_out[284] <= layer1_out[95] & layer1_out[96];
     layer2_out[285] <= layer1_out[247] & ~layer1_out[248];
     layer2_out[286] <= 1'b0;
     layer2_out[287] <= ~(layer1_out[107] | layer1_out[108]);
     layer2_out[288] <= 1'b0;
     layer2_out[289] <= layer1_out[212];
     layer2_out[290] <= ~(layer1_out[201] & layer1_out[202]);
     layer2_out[291] <= layer1_out[17] ^ layer1_out[18];
     layer2_out[292] <= ~(layer1_out[185] & layer1_out[186]);
     layer2_out[293] <= layer1_out[140] | layer1_out[141];
     layer2_out[294] <= ~layer1_out[87] | layer1_out[88];
     layer2_out[295] <= ~layer1_out[239];
     layer2_out[296] <= ~layer1_out[80];
     layer2_out[297] <= layer1_out[34];
     layer2_out[298] <= ~(layer1_out[161] & layer1_out[162]);
     layer2_out[299] <= layer1_out[189];
     layer3_out[0] <= layer2_out[117];
     layer3_out[1] <= ~layer2_out[183] | layer2_out[184];
     layer3_out[2] <= layer2_out[41] & ~layer2_out[42];
     layer3_out[3] <= layer2_out[221];
     layer3_out[4] <= ~layer2_out[73];
     layer3_out[5] <= layer2_out[250];
     layer3_out[6] <= layer2_out[8] & ~layer2_out[7];
     layer3_out[7] <= layer2_out[205] & ~layer2_out[204];
     layer3_out[8] <= ~layer2_out[143];
     layer3_out[9] <= ~(layer2_out[274] | layer2_out[275]);
     layer3_out[10] <= layer2_out[220];
     layer3_out[11] <= layer2_out[208];
     layer3_out[12] <= ~layer2_out[105];
     layer3_out[13] <= ~layer2_out[136];
     layer3_out[14] <= ~layer2_out[31];
     layer3_out[15] <= layer2_out[94];
     layer3_out[16] <= layer2_out[65];
     layer3_out[17] <= ~(layer2_out[51] | layer2_out[52]);
     layer3_out[18] <= layer2_out[215] & ~layer2_out[216];
     layer3_out[19] <= layer2_out[69];
     layer3_out[20] <= layer2_out[29];
     layer3_out[21] <= layer2_out[150];
     layer3_out[22] <= layer2_out[52] | layer2_out[53];
     layer3_out[23] <= ~(layer2_out[223] ^ layer2_out[224]);
     layer3_out[24] <= layer2_out[157];
     layer3_out[25] <= ~(layer2_out[120] & layer2_out[121]);
     layer3_out[26] <= layer2_out[65];
     layer3_out[27] <= layer2_out[17];
     layer3_out[28] <= ~(layer2_out[47] ^ layer2_out[48]);
     layer3_out[29] <= layer2_out[141];
     layer3_out[30] <= layer2_out[194] & ~layer2_out[193];
     layer3_out[31] <= ~(layer2_out[172] | layer2_out[173]);
     layer3_out[32] <= ~layer2_out[284];
     layer3_out[33] <= layer2_out[15];
     layer3_out[34] <= layer2_out[218];
     layer3_out[35] <= layer2_out[113] & ~layer2_out[114];
     layer3_out[36] <= layer2_out[111] & layer2_out[112];
     layer3_out[37] <= ~layer2_out[264];
     layer3_out[38] <= ~layer2_out[178];
     layer3_out[39] <= ~layer2_out[173];
     layer3_out[40] <= layer2_out[287];
     layer3_out[41] <= layer2_out[71];
     layer3_out[42] <= layer2_out[74];
     layer3_out[43] <= ~(layer2_out[109] | layer2_out[110]);
     layer3_out[44] <= ~layer2_out[77];
     layer3_out[45] <= layer2_out[278];
     layer3_out[46] <= layer2_out[190] & layer2_out[191];
     layer3_out[47] <= layer2_out[55] & ~layer2_out[54];
     layer3_out[48] <= layer2_out[0];
     layer3_out[49] <= layer2_out[12] & ~layer2_out[13];
     layer3_out[50] <= ~layer2_out[157];
     layer3_out[51] <= layer2_out[181] & ~layer2_out[180];
     layer3_out[52] <= layer2_out[51];
     layer3_out[53] <= ~layer2_out[69];
     layer3_out[54] <= layer2_out[202] & ~layer2_out[203];
     layer3_out[55] <= layer2_out[138];
     layer3_out[56] <= layer2_out[67] & layer2_out[68];
     layer3_out[57] <= ~(layer2_out[3] | layer2_out[4]);
     layer3_out[58] <= ~layer2_out[167];
     layer3_out[59] <= layer2_out[256] & layer2_out[257];
     layer3_out[60] <= ~layer2_out[295];
     layer3_out[61] <= layer2_out[266];
     layer3_out[62] <= layer2_out[58];
     layer3_out[63] <= layer2_out[226] ^ layer2_out[227];
     layer3_out[64] <= layer2_out[248] & ~layer2_out[247];
     layer3_out[65] <= ~layer2_out[85];
     layer3_out[66] <= layer2_out[285];
     layer3_out[67] <= layer2_out[76] | layer2_out[77];
     layer3_out[68] <= layer2_out[229] & layer2_out[230];
     layer3_out[69] <= layer2_out[186];
     layer3_out[70] <= layer2_out[229] & ~layer2_out[228];
     layer3_out[71] <= layer2_out[135];
     layer3_out[72] <= ~layer2_out[241];
     layer3_out[73] <= ~(layer2_out[182] | layer2_out[183]);
     layer3_out[74] <= ~(layer2_out[26] ^ layer2_out[27]);
     layer3_out[75] <= layer2_out[139] & layer2_out[140];
     layer3_out[76] <= ~layer2_out[159];
     layer3_out[77] <= layer2_out[155] & ~layer2_out[154];
     layer3_out[78] <= ~layer2_out[5];
     layer3_out[79] <= layer2_out[9];
     layer3_out[80] <= layer2_out[254];
     layer3_out[81] <= layer2_out[90] & ~layer2_out[89];
     layer3_out[82] <= layer2_out[57];
     layer3_out[83] <= layer2_out[9];
     layer3_out[84] <= layer2_out[214] ^ layer2_out[215];
     layer3_out[85] <= layer2_out[222] & ~layer2_out[223];
     layer3_out[86] <= ~layer2_out[79];
     layer3_out[87] <= layer2_out[149] & ~layer2_out[148];
     layer3_out[88] <= layer2_out[129] & ~layer2_out[128];
     layer3_out[89] <= layer2_out[289] ^ layer2_out[290];
     layer3_out[90] <= ~layer2_out[3];
     layer3_out[91] <= layer2_out[60] & ~layer2_out[59];
     layer3_out[92] <= ~layer2_out[280];
     layer3_out[93] <= layer2_out[232];
     layer3_out[94] <= ~layer2_out[177];
     layer3_out[95] <= layer2_out[115];
     layer3_out[96] <= layer2_out[147];
     layer3_out[97] <= ~(layer2_out[96] | layer2_out[97]);
     layer3_out[98] <= ~(layer2_out[99] ^ layer2_out[100]);
     layer3_out[99] <= ~layer2_out[287];
     layer3_out[100] <= ~layer2_out[153];
     layer3_out[101] <= layer2_out[90];
     layer3_out[102] <= layer2_out[115] | layer2_out[116];
     layer3_out[103] <= ~layer2_out[185];
     layer3_out[104] <= layer2_out[146];
     layer3_out[105] <= ~layer2_out[81];
     layer3_out[106] <= layer2_out[36];
     layer3_out[107] <= ~layer2_out[201];
     layer3_out[108] <= layer2_out[268];
     layer3_out[109] <= ~layer2_out[164] | layer2_out[165];
     layer3_out[110] <= ~(layer2_out[294] & layer2_out[295]);
     layer3_out[111] <= layer2_out[11];
     layer3_out[112] <= ~layer2_out[238];
     layer3_out[113] <= ~(layer2_out[93] ^ layer2_out[94]);
     layer3_out[114] <= layer2_out[244];
     layer3_out[115] <= ~layer2_out[44];
     layer3_out[116] <= layer2_out[253];
     layer3_out[117] <= ~layer2_out[108];
     layer3_out[118] <= layer2_out[27];
     layer3_out[119] <= ~layer2_out[218];
     layer3_out[120] <= layer2_out[71];
     layer3_out[121] <= layer2_out[130];
     layer3_out[122] <= layer2_out[19] | layer2_out[20];
     layer3_out[123] <= ~layer2_out[192] | layer2_out[191];
     layer3_out[124] <= ~(layer2_out[146] | layer2_out[147]);
     layer3_out[125] <= layer2_out[297];
     layer3_out[126] <= ~layer2_out[206];
     layer3_out[127] <= layer2_out[97];
     layer3_out[128] <= layer2_out[240];
     layer3_out[129] <= layer2_out[73];
     layer3_out[130] <= layer2_out[170];
     layer3_out[131] <= layer2_out[24];
     layer3_out[132] <= layer2_out[284];
     layer3_out[133] <= ~layer2_out[161];
     layer3_out[134] <= layer2_out[174] & ~layer2_out[175];
     layer3_out[135] <= ~layer2_out[75];
     layer3_out[136] <= layer2_out[261];
     layer3_out[137] <= layer2_out[92];
     layer3_out[138] <= layer2_out[238];
     layer3_out[139] <= ~layer2_out[226];
     layer3_out[140] <= ~layer2_out[83];
     layer3_out[141] <= layer2_out[119] & layer2_out[120];
     layer3_out[142] <= ~layer2_out[206];
     layer3_out[143] <= layer2_out[201];
     layer3_out[144] <= layer2_out[233] | layer2_out[234];
     layer3_out[145] <= layer2_out[178] & ~layer2_out[179];
     layer3_out[146] <= ~layer2_out[281];
     layer3_out[147] <= layer2_out[66];
     layer3_out[148] <= ~layer2_out[244];
     layer3_out[149] <= layer2_out[195] ^ layer2_out[196];
     layer3_out[150] <= ~layer2_out[291];
     layer3_out[151] <= ~layer2_out[254];
     layer3_out[152] <= layer2_out[88];
     layer3_out[153] <= layer2_out[293];
     layer3_out[154] <= layer2_out[37];
     layer3_out[155] <= ~layer2_out[39];
     layer3_out[156] <= ~(layer2_out[227] ^ layer2_out[228]);
     layer3_out[157] <= ~layer2_out[95];
     layer3_out[158] <= ~layer2_out[166];
     layer3_out[159] <= ~layer2_out[1];
     layer3_out[160] <= layer2_out[14];
     layer3_out[161] <= ~layer2_out[123];
     layer3_out[162] <= layer2_out[85];
     layer3_out[163] <= ~(layer2_out[155] | layer2_out[156]);
     layer3_out[164] <= layer2_out[168] & ~layer2_out[169];
     layer3_out[165] <= layer2_out[24];
     layer3_out[166] <= layer2_out[32];
     layer3_out[167] <= layer2_out[224] ^ layer2_out[225];
     layer3_out[168] <= ~layer2_out[259];
     layer3_out[169] <= ~layer2_out[135];
     layer3_out[170] <= ~layer2_out[158];
     layer3_out[171] <= layer2_out[122] & ~layer2_out[123];
     layer3_out[172] <= layer2_out[212];
     layer3_out[173] <= ~layer2_out[63] | layer2_out[62];
     layer3_out[174] <= ~layer2_out[60];
     layer3_out[175] <= layer2_out[61] & layer2_out[62];
     layer3_out[176] <= layer2_out[53];
     layer3_out[177] <= ~layer2_out[39];
     layer3_out[178] <= ~(layer2_out[194] ^ layer2_out[195]);
     layer3_out[179] <= ~layer2_out[102];
     layer3_out[180] <= layer2_out[149] & ~layer2_out[150];
     layer3_out[181] <= layer2_out[262];
     layer3_out[182] <= layer2_out[44] & ~layer2_out[45];
     layer3_out[183] <= ~(layer2_out[33] ^ layer2_out[34]);
     layer3_out[184] <= layer2_out[217];
     layer3_out[185] <= ~layer2_out[103];
     layer3_out[186] <= ~layer2_out[283];
     layer3_out[187] <= ~layer2_out[269];
     layer3_out[188] <= ~(layer2_out[140] | layer2_out[141]);
     layer3_out[189] <= layer2_out[185];
     layer3_out[190] <= layer2_out[234] | layer2_out[235];
     layer3_out[191] <= ~layer2_out[275];
     layer3_out[192] <= ~layer2_out[106];
     layer3_out[193] <= ~(layer2_out[246] | layer2_out[247]);
     layer3_out[194] <= ~layer2_out[258];
     layer3_out[195] <= layer2_out[57] & ~layer2_out[56];
     layer3_out[196] <= layer2_out[187];
     layer3_out[197] <= layer2_out[280];
     layer3_out[198] <= ~layer2_out[98];
     layer3_out[199] <= ~layer2_out[63];
     layer3_out[200] <= layer2_out[122];
     layer3_out[201] <= layer2_out[86];
     layer3_out[202] <= ~(layer2_out[25] | layer2_out[26]);
     layer3_out[203] <= layer2_out[171] & ~layer2_out[172];
     layer3_out[204] <= ~layer2_out[38];
     layer3_out[205] <= layer2_out[131] & ~layer2_out[130];
     layer3_out[206] <= layer2_out[92] ^ layer2_out[93];
     layer3_out[207] <= layer2_out[293];
     layer3_out[208] <= ~layer2_out[22];
     layer3_out[209] <= ~layer2_out[45] | layer2_out[46];
     layer3_out[210] <= ~(layer2_out[46] ^ layer2_out[47]);
     layer3_out[211] <= layer2_out[111];
     layer3_out[212] <= layer2_out[179];
     layer3_out[213] <= ~(layer2_out[209] ^ layer2_out[210]);
     layer3_out[214] <= layer2_out[42] & layer2_out[43];
     layer3_out[215] <= ~layer2_out[235];
     layer3_out[216] <= ~layer2_out[267];
     layer3_out[217] <= layer2_out[249];
     layer3_out[218] <= ~layer2_out[124];
     layer3_out[219] <= ~layer2_out[193];
     layer3_out[220] <= layer2_out[175];
     layer3_out[221] <= ~layer2_out[214];
     layer3_out[222] <= layer2_out[15];
     layer3_out[223] <= layer2_out[19];
     layer3_out[224] <= ~layer2_out[167];
     layer3_out[225] <= layer2_out[103];
     layer3_out[226] <= layer2_out[81];
     layer3_out[227] <= ~layer2_out[171];
     layer3_out[228] <= layer2_out[246];
     layer3_out[229] <= layer2_out[112] ^ layer2_out[113];
     layer3_out[230] <= layer2_out[144] & layer2_out[145];
     layer3_out[231] <= ~layer2_out[108] | layer2_out[107];
     layer3_out[232] <= layer2_out[220];
     layer3_out[233] <= layer2_out[199];
     layer3_out[234] <= layer2_out[230];
     layer3_out[235] <= ~layer2_out[49];
     layer3_out[236] <= ~layer2_out[139];
     layer3_out[237] <= layer2_out[199] & ~layer2_out[198];
     layer3_out[238] <= layer2_out[190];
     layer3_out[239] <= layer2_out[278] & ~layer2_out[279];
     layer3_out[240] <= layer2_out[5];
     layer3_out[241] <= ~layer2_out[239];
     layer3_out[242] <= layer2_out[117];
     layer3_out[243] <= layer2_out[265];
     layer3_out[244] <= ~layer2_out[270];
     layer3_out[245] <= ~layer2_out[272];
     layer3_out[246] <= ~layer2_out[11];
     layer3_out[247] <= ~layer2_out[88];
     layer3_out[248] <= ~(layer2_out[17] ^ layer2_out[18]);
     layer3_out[249] <= layer2_out[151];
     layer3_out[250] <= ~layer2_out[126];
     layer3_out[251] <= layer2_out[101];
     layer3_out[252] <= ~layer2_out[40];
     layer3_out[253] <= ~layer2_out[299];
     layer3_out[254] <= layer2_out[236] & ~layer2_out[237];
     layer3_out[255] <= ~layer2_out[0];
     layer3_out[256] <= layer2_out[56];
     layer3_out[257] <= ~layer2_out[256];
     layer3_out[258] <= ~layer2_out[259];
     layer3_out[259] <= ~layer2_out[143];
     layer3_out[260] <= ~layer2_out[291];
     layer3_out[261] <= layer2_out[163];
     layer3_out[262] <= layer2_out[21];
     layer3_out[263] <= layer2_out[232];
     layer3_out[264] <= layer2_out[181];
     layer3_out[265] <= ~layer2_out[105];
     layer3_out[266] <= ~layer2_out[208];
     layer3_out[267] <= layer2_out[243];
     layer3_out[268] <= layer2_out[211];
     layer3_out[269] <= ~layer2_out[84];
     layer3_out[270] <= ~(layer2_out[28] | layer2_out[29]);
     layer3_out[271] <= layer2_out[274];
     layer3_out[272] <= layer2_out[251] & ~layer2_out[250];
     layer3_out[273] <= layer2_out[204];
     layer3_out[274] <= layer2_out[34];
     layer3_out[275] <= ~layer2_out[134];
     layer3_out[276] <= layer2_out[262];
     layer3_out[277] <= ~layer2_out[197];
     layer3_out[278] <= ~layer2_out[188];
     layer3_out[279] <= layer2_out[160] ^ layer2_out[161];
     layer3_out[280] <= layer2_out[7];
     layer3_out[281] <= ~(layer2_out[118] ^ layer2_out[119]);
     layer3_out[282] <= layer2_out[127];
     layer3_out[283] <= layer2_out[297] & layer2_out[298];
     layer3_out[284] <= layer2_out[271] & layer2_out[272];
     layer3_out[285] <= ~layer2_out[196];
     layer3_out[286] <= ~layer2_out[30];
     layer3_out[287] <= layer2_out[211];
     layer3_out[288] <= layer2_out[289];
     layer3_out[289] <= layer2_out[50] & ~layer2_out[49];
     layer3_out[290] <= layer2_out[251];
     layer3_out[291] <= layer2_out[276] & ~layer2_out[277];
     layer3_out[292] <= layer2_out[21] & layer2_out[22];
     layer3_out[293] <= layer2_out[270];
     layer3_out[294] <= ~layer2_out[132];
     layer3_out[295] <= ~(layer2_out[162] ^ layer2_out[163]);
     layer3_out[296] <= layer2_out[154] & ~layer2_out[153];
     layer3_out[297] <= ~layer2_out[132];
     layer3_out[298] <= layer2_out[79];
     layer3_out[299] <= layer2_out[127] & ~layer2_out[128];
      last_layer_output <= layer3_out;

      result[0] <= last_layer_output[0] + last_layer_output[1] + last_layer_output[2] + last_layer_output[3] + last_layer_output[4] + last_layer_output[5] + last_layer_output[6] + last_layer_output[7] + last_layer_output[8] + last_layer_output[9] + last_layer_output[10] + last_layer_output[11] + last_layer_output[12] + last_layer_output[13] + last_layer_output[14] + last_layer_output[15] + last_layer_output[16] + last_layer_output[17] + last_layer_output[18] + last_layer_output[19] + last_layer_output[20] + last_layer_output[21] + last_layer_output[22] + last_layer_output[23] + last_layer_output[24] + last_layer_output[25] + last_layer_output[26] + last_layer_output[27] + last_layer_output[28] + last_layer_output[29];
      result[1] <= last_layer_output[30] + last_layer_output[31] + last_layer_output[32] + last_layer_output[33] + last_layer_output[34] + last_layer_output[35] + last_layer_output[36] + last_layer_output[37] + last_layer_output[38] + last_layer_output[39] + last_layer_output[40] + last_layer_output[41] + last_layer_output[42] + last_layer_output[43] + last_layer_output[44] + last_layer_output[45] + last_layer_output[46] + last_layer_output[47] + last_layer_output[48] + last_layer_output[49] + last_layer_output[50] + last_layer_output[51] + last_layer_output[52] + last_layer_output[53] + last_layer_output[54] + last_layer_output[55] + last_layer_output[56] + last_layer_output[57] + last_layer_output[58] + last_layer_output[59];
      result[2] <= last_layer_output[60] + last_layer_output[61] + last_layer_output[62] + last_layer_output[63] + last_layer_output[64] + last_layer_output[65] + last_layer_output[66] + last_layer_output[67] + last_layer_output[68] + last_layer_output[69] + last_layer_output[70] + last_layer_output[71] + last_layer_output[72] + last_layer_output[73] + last_layer_output[74] + last_layer_output[75] + last_layer_output[76] + last_layer_output[77] + last_layer_output[78] + last_layer_output[79] + last_layer_output[80] + last_layer_output[81] + last_layer_output[82] + last_layer_output[83] + last_layer_output[84] + last_layer_output[85] + last_layer_output[86] + last_layer_output[87] + last_layer_output[88] + last_layer_output[89];
      result[3] <= last_layer_output[90] + last_layer_output[91] + last_layer_output[92] + last_layer_output[93] + last_layer_output[94] + last_layer_output[95] + last_layer_output[96] + last_layer_output[97] + last_layer_output[98] + last_layer_output[99] + last_layer_output[100] + last_layer_output[101] + last_layer_output[102] + last_layer_output[103] + last_layer_output[104] + last_layer_output[105] + last_layer_output[106] + last_layer_output[107] + last_layer_output[108] + last_layer_output[109] + last_layer_output[110] + last_layer_output[111] + last_layer_output[112] + last_layer_output[113] + last_layer_output[114] + last_layer_output[115] + last_layer_output[116] + last_layer_output[117] + last_layer_output[118] + last_layer_output[119];
      result[4] <= last_layer_output[120] + last_layer_output[121] + last_layer_output[122] + last_layer_output[123] + last_layer_output[124] + last_layer_output[125] + last_layer_output[126] + last_layer_output[127] + last_layer_output[128] + last_layer_output[129] + last_layer_output[130] + last_layer_output[131] + last_layer_output[132] + last_layer_output[133] + last_layer_output[134] + last_layer_output[135] + last_layer_output[136] + last_layer_output[137] + last_layer_output[138] + last_layer_output[139] + last_layer_output[140] + last_layer_output[141] + last_layer_output[142] + last_layer_output[143] + last_layer_output[144] + last_layer_output[145] + last_layer_output[146] + last_layer_output[147] + last_layer_output[148] + last_layer_output[149];
      result[5] <= last_layer_output[150] + last_layer_output[151] + last_layer_output[152] + last_layer_output[153] + last_layer_output[154] + last_layer_output[155] + last_layer_output[156] + last_layer_output[157] + last_layer_output[158] + last_layer_output[159] + last_layer_output[160] + last_layer_output[161] + last_layer_output[162] + last_layer_output[163] + last_layer_output[164] + last_layer_output[165] + last_layer_output[166] + last_layer_output[167] + last_layer_output[168] + last_layer_output[169] + last_layer_output[170] + last_layer_output[171] + last_layer_output[172] + last_layer_output[173] + last_layer_output[174] + last_layer_output[175] + last_layer_output[176] + last_layer_output[177] + last_layer_output[178] + last_layer_output[179];
      result[6] <= last_layer_output[180] + last_layer_output[181] + last_layer_output[182] + last_layer_output[183] + last_layer_output[184] + last_layer_output[185] + last_layer_output[186] + last_layer_output[187] + last_layer_output[188] + last_layer_output[189] + last_layer_output[190] + last_layer_output[191] + last_layer_output[192] + last_layer_output[193] + last_layer_output[194] + last_layer_output[195] + last_layer_output[196] + last_layer_output[197] + last_layer_output[198] + last_layer_output[199] + last_layer_output[200] + last_layer_output[201] + last_layer_output[202] + last_layer_output[203] + last_layer_output[204] + last_layer_output[205] + last_layer_output[206] + last_layer_output[207] + last_layer_output[208] + last_layer_output[209];
      result[7] <= last_layer_output[210] + last_layer_output[211] + last_layer_output[212] + last_layer_output[213] + last_layer_output[214] + last_layer_output[215] + last_layer_output[216] + last_layer_output[217] + last_layer_output[218] + last_layer_output[219] + last_layer_output[220] + last_layer_output[221] + last_layer_output[222] + last_layer_output[223] + last_layer_output[224] + last_layer_output[225] + last_layer_output[226] + last_layer_output[227] + last_layer_output[228] + last_layer_output[229] + last_layer_output[230] + last_layer_output[231] + last_layer_output[232] + last_layer_output[233] + last_layer_output[234] + last_layer_output[235] + last_layer_output[236] + last_layer_output[237] + last_layer_output[238] + last_layer_output[239];
      result[8] <= last_layer_output[240] + last_layer_output[241] + last_layer_output[242] + last_layer_output[243] + last_layer_output[244] + last_layer_output[245] + last_layer_output[246] + last_layer_output[247] + last_layer_output[248] + last_layer_output[249] + last_layer_output[250] + last_layer_output[251] + last_layer_output[252] + last_layer_output[253] + last_layer_output[254] + last_layer_output[255] + last_layer_output[256] + last_layer_output[257] + last_layer_output[258] + last_layer_output[259] + last_layer_output[260] + last_layer_output[261] + last_layer_output[262] + last_layer_output[263] + last_layer_output[264] + last_layer_output[265] + last_layer_output[266] + last_layer_output[267] + last_layer_output[268] + last_layer_output[269];
      result[9] <= last_layer_output[270] + last_layer_output[271] + last_layer_output[272] + last_layer_output[273] + last_layer_output[274] + last_layer_output[275] + last_layer_output[276] + last_layer_output[277] + last_layer_output[278] + last_layer_output[279] + last_layer_output[280] + last_layer_output[281] + last_layer_output[282] + last_layer_output[283] + last_layer_output[284] + last_layer_output[285] + last_layer_output[286] + last_layer_output[287] + last_layer_output[288] + last_layer_output[289] + last_layer_output[290] + last_layer_output[291] + last_layer_output[292] + last_layer_output[293] + last_layer_output[294] + last_layer_output[295] + last_layer_output[296] + last_layer_output[297] + last_layer_output[298] + last_layer_output[299];
end
      assign y[49:45]=result[0];
      assign y[44:40]=result[1];
      assign y[39:35]=result[2];
      assign y[34:30]=result[3];
      assign y[29:25]=result[4];
      assign y[24:20]=result[5];
      assign y[19:15]=result[6];
      assign y[14:10]=result[7];
      assign y[9:5]=result[8];
      assign y[4:0]=result[9];
endmodule
