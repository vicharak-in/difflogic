module logic_network (    input clk,
    input wire [9215:0] x,
    output wire [109:0] y
);
      reg [11999:0] layer0_out = 0;
      reg [11999:0] layer1_out = 0;
      reg [11999:0] layer2_out = 0;
      reg [11999:0] layer3_out = 0;
      reg [11999:0] last_layer_output = 0;
      reg [10:0] result [9:0];
      always @(posedge clk) begin
     layer0_out[0] <= ~(x[160] ^ x[161]);
     layer0_out[1] <= ~(x[5594] & x[5595]);
     layer0_out[2] <= ~x[4073];
     layer0_out[3] <= ~(x[2259] & x[2261]);
     layer0_out[4] <= ~(x[859] & x[860]);
     layer0_out[5] <= x[149] & x[150];
     layer0_out[6] <= ~x[4197];
     layer0_out[7] <= x[6760] & ~x[6759];
     layer0_out[8] <= x[5433] & x[5434];
     layer0_out[9] <= ~(x[2045] & x[2047]);
     layer0_out[10] <= x[1382] & x[1384];
     layer0_out[11] <= ~(x[2555] ^ x[2557]);
     layer0_out[12] <= x[3728];
     layer0_out[13] <= ~x[464];
     layer0_out[14] <= x[5744] & x[5745];
     layer0_out[15] <= ~x[70];
     layer0_out[16] <= x[281];
     layer0_out[17] <= x[8407];
     layer0_out[18] <= ~x[2353];
     layer0_out[19] <= x[3548] | x[3549];
     layer0_out[20] <= x[5251] & x[5252];
     layer0_out[21] <= ~x[3376];
     layer0_out[22] <= ~(x[8958] & x[8959]);
     layer0_out[23] <= x[5457] | x[5458];
     layer0_out[24] <= ~x[9087];
     layer0_out[25] <= ~x[2602];
     layer0_out[26] <= x[3666] | x[3667];
     layer0_out[27] <= ~x[7736];
     layer0_out[28] <= ~(x[4492] & x[4493]);
     layer0_out[29] <= x[6999] ^ x[7000];
     layer0_out[30] <= x[7254] ^ x[7255];
     layer0_out[31] <= ~(x[2235] ^ x[2236]);
     layer0_out[32] <= x[2156] & x[2158];
     layer0_out[33] <= 1'b0;
     layer0_out[34] <= x[753] & x[754];
     layer0_out[35] <= x[6321] | x[6322];
     layer0_out[36] <= ~x[247];
     layer0_out[37] <= ~(x[1905] & x[1907]);
     layer0_out[38] <= x[968] ^ x[970];
     layer0_out[39] <= x[5456] & x[5457];
     layer0_out[40] <= x[8758] & x[8759];
     layer0_out[41] <= x[3042] & ~x[3041];
     layer0_out[42] <= x[2343] & x[2344];
     layer0_out[43] <= x[4213] ^ x[4214];
     layer0_out[44] <= x[6057] & x[6058];
     layer0_out[45] <= x[3034] & x[3035];
     layer0_out[46] <= x[1377] & x[1378];
     layer0_out[47] <= ~(x[191] & x[192]);
     layer0_out[48] <= x[8693];
     layer0_out[49] <= x[5717];
     layer0_out[50] <= ~x[4912];
     layer0_out[51] <= ~x[6473];
     layer0_out[52] <= x[2277];
     layer0_out[53] <= ~(x[8521] | x[8522]);
     layer0_out[54] <= ~(x[148] & x[150]);
     layer0_out[55] <= ~(x[2607] & x[2608]);
     layer0_out[56] <= ~(x[4785] | x[4786]);
     layer0_out[57] <= ~x[2337];
     layer0_out[58] <= ~(x[3390] & x[3391]);
     layer0_out[59] <= ~x[4090];
     layer0_out[60] <= x[5762] | x[5763];
     layer0_out[61] <= x[7421];
     layer0_out[62] <= 1'b0;
     layer0_out[63] <= x[8526] & x[8527];
     layer0_out[64] <= ~x[8511];
     layer0_out[65] <= x[1942] | x[1943];
     layer0_out[66] <= x[2452] & x[2453];
     layer0_out[67] <= x[4364] ^ x[4365];
     layer0_out[68] <= ~(x[7165] & x[7166]);
     layer0_out[69] <= x[2213] | x[2215];
     layer0_out[70] <= x[1815];
     layer0_out[71] <= ~(x[1345] & x[1347]);
     layer0_out[72] <= x[6351] | x[6352];
     layer0_out[73] <= ~(x[4063] & x[4064]);
     layer0_out[74] <= x[3574] & x[3575];
     layer0_out[75] <= ~x[7137];
     layer0_out[76] <= ~(x[4284] & x[4285]);
     layer0_out[77] <= x[8117] & x[8118];
     layer0_out[78] <= x[6588] & x[6589];
     layer0_out[79] <= ~x[5742];
     layer0_out[80] <= x[1106] & x[1108];
     layer0_out[81] <= ~x[3795];
     layer0_out[82] <= 1'b0;
     layer0_out[83] <= ~(x[6567] & x[6568]);
     layer0_out[84] <= x[5718] & x[5719];
     layer0_out[85] <= ~(x[1056] & x[1057]);
     layer0_out[86] <= x[3485] | x[3486];
     layer0_out[87] <= ~(x[5116] ^ x[5117]);
     layer0_out[88] <= x[2034] ^ x[2035];
     layer0_out[89] <= ~(x[1742] ^ x[1744]);
     layer0_out[90] <= 1'b1;
     layer0_out[91] <= ~(x[8249] | x[8250]);
     layer0_out[92] <= x[7965] & x[7966];
     layer0_out[93] <= ~(x[1481] & x[1482]);
     layer0_out[94] <= x[6944] & ~x[6943];
     layer0_out[95] <= x[1164] & x[1166];
     layer0_out[96] <= x[71] & x[72];
     layer0_out[97] <= x[4004] | x[4005];
     layer0_out[98] <= ~(x[1131] ^ x[1133]);
     layer0_out[99] <= x[6724] & x[6725];
     layer0_out[100] <= x[3462] & ~x[3463];
     layer0_out[101] <= ~x[5204];
     layer0_out[102] <= x[2398] | x[2400];
     layer0_out[103] <= ~(x[5311] & x[5312]);
     layer0_out[104] <= ~(x[5111] ^ x[5112]);
     layer0_out[105] <= ~(x[135] ^ x[137]);
     layer0_out[106] <= ~x[7044];
     layer0_out[107] <= ~(x[2126] & x[2127]);
     layer0_out[108] <= ~x[73];
     layer0_out[109] <= x[5231] | x[5232];
     layer0_out[110] <= ~x[6229] | x[6230];
     layer0_out[111] <= x[1575];
     layer0_out[112] <= ~(x[2414] & x[2415]);
     layer0_out[113] <= ~(x[2981] & x[2982]);
     layer0_out[114] <= x[7384] | x[7385];
     layer0_out[115] <= x[2697] & x[2698];
     layer0_out[116] <= x[5112] | x[5113];
     layer0_out[117] <= ~x[1716];
     layer0_out[118] <= x[7279] ^ x[7280];
     layer0_out[119] <= x[7098] & x[7099];
     layer0_out[120] <= ~(x[5078] ^ x[5079]);
     layer0_out[121] <= ~(x[4934] | x[4935]);
     layer0_out[122] <= x[3869] & x[3870];
     layer0_out[123] <= x[6398];
     layer0_out[124] <= x[3375] | x[3376];
     layer0_out[125] <= x[5532] ^ x[5533];
     layer0_out[126] <= 1'b0;
     layer0_out[127] <= x[1591] & x[1593];
     layer0_out[128] <= ~(x[2142] & x[2143]);
     layer0_out[129] <= x[390] | x[392];
     layer0_out[130] <= x[605] & x[607];
     layer0_out[131] <= x[6133] & x[6134];
     layer0_out[132] <= x[977] & x[979];
     layer0_out[133] <= ~(x[282] & x[283]);
     layer0_out[134] <= x[5365] & x[5366];
     layer0_out[135] <= x[434] | x[435];
     layer0_out[136] <= ~(x[4983] | x[4984]);
     layer0_out[137] <= ~(x[6864] & x[6865]);
     layer0_out[138] <= ~(x[2048] & x[2050]);
     layer0_out[139] <= 1'b0;
     layer0_out[140] <= ~(x[1624] & x[1626]);
     layer0_out[141] <= x[7423] | x[7424];
     layer0_out[142] <= x[425] | x[426];
     layer0_out[143] <= x[2330] ^ x[2332];
     layer0_out[144] <= x[9107] | x[9108];
     layer0_out[145] <= x[8306] | x[8307];
     layer0_out[146] <= ~x[6724] | x[6723];
     layer0_out[147] <= x[137] | x[138];
     layer0_out[148] <= x[2772] ^ x[2774];
     layer0_out[149] <= ~x[707] | x[709];
     layer0_out[150] <= ~(x[8251] & x[8252]);
     layer0_out[151] <= x[176] ^ x[178];
     layer0_out[152] <= ~(x[6319] & x[6320]);
     layer0_out[153] <= ~x[2135] | x[2133];
     layer0_out[154] <= x[4948] | x[4949];
     layer0_out[155] <= ~(x[4024] | x[4025]);
     layer0_out[156] <= ~(x[3175] ^ x[3176]);
     layer0_out[157] <= 1'b1;
     layer0_out[158] <= ~(x[8834] ^ x[8835]);
     layer0_out[159] <= x[9188] & x[9189];
     layer0_out[160] <= ~(x[8307] & x[8308]);
     layer0_out[161] <= ~x[4307];
     layer0_out[162] <= x[5389] | x[5390];
     layer0_out[163] <= 1'b1;
     layer0_out[164] <= ~(x[1813] & x[1814]);
     layer0_out[165] <= ~(x[5551] | x[5552]);
     layer0_out[166] <= ~(x[2461] ^ x[2462]);
     layer0_out[167] <= x[3013];
     layer0_out[168] <= 1'b0;
     layer0_out[169] <= ~x[8634] | x[8635];
     layer0_out[170] <= ~(x[2826] ^ x[2827]);
     layer0_out[171] <= ~(x[2254] | x[2255]);
     layer0_out[172] <= ~(x[4359] & x[4360]);
     layer0_out[173] <= ~x[3199];
     layer0_out[174] <= ~(x[3368] ^ x[3369]);
     layer0_out[175] <= ~(x[2528] | x[2529]);
     layer0_out[176] <= x[8938] | x[8939];
     layer0_out[177] <= ~(x[8962] | x[8963]);
     layer0_out[178] <= ~(x[8895] & x[8896]);
     layer0_out[179] <= ~x[6293] | x[6292];
     layer0_out[180] <= ~x[3685];
     layer0_out[181] <= 1'b1;
     layer0_out[182] <= ~(x[805] & x[806]);
     layer0_out[183] <= ~(x[3542] ^ x[3543]);
     layer0_out[184] <= ~(x[2384] & x[2385]);
     layer0_out[185] <= x[5984];
     layer0_out[186] <= ~(x[140] | x[141]);
     layer0_out[187] <= x[5216] | x[5217];
     layer0_out[188] <= x[6465] ^ x[6466];
     layer0_out[189] <= x[5636] ^ x[5637];
     layer0_out[190] <= ~x[3535];
     layer0_out[191] <= ~(x[5090] & x[5091]);
     layer0_out[192] <= x[4995] | x[4996];
     layer0_out[193] <= x[7431] & x[7432];
     layer0_out[194] <= ~x[512];
     layer0_out[195] <= ~x[268];
     layer0_out[196] <= ~(x[6539] & x[6540]);
     layer0_out[197] <= ~(x[1301] & x[1303]);
     layer0_out[198] <= x[3320];
     layer0_out[199] <= 1'b1;
     layer0_out[200] <= x[8681] | x[8682];
     layer0_out[201] <= 1'b0;
     layer0_out[202] <= x[1888] & x[1890];
     layer0_out[203] <= x[7431];
     layer0_out[204] <= x[807] | x[808];
     layer0_out[205] <= ~(x[990] | x[991]);
     layer0_out[206] <= 1'b1;
     layer0_out[207] <= ~(x[2133] & x[2134]);
     layer0_out[208] <= ~x[4734];
     layer0_out[209] <= x[8763] & ~x[8762];
     layer0_out[210] <= ~x[9136];
     layer0_out[211] <= x[5317] & x[5318];
     layer0_out[212] <= ~(x[62] ^ x[64]);
     layer0_out[213] <= ~(x[1347] & x[1348]);
     layer0_out[214] <= ~x[1374];
     layer0_out[215] <= ~(x[7146] & x[7147]);
     layer0_out[216] <= ~(x[9097] | x[9098]);
     layer0_out[217] <= x[1319] & ~x[1321];
     layer0_out[218] <= ~x[5523];
     layer0_out[219] <= 1'b0;
     layer0_out[220] <= ~x[8931];
     layer0_out[221] <= x[8936] & ~x[8935];
     layer0_out[222] <= x[604] | x[606];
     layer0_out[223] <= x[8054];
     layer0_out[224] <= ~(x[691] | x[692]);
     layer0_out[225] <= x[453] & ~x[455];
     layer0_out[226] <= ~(x[8613] ^ x[8614]);
     layer0_out[227] <= ~(x[182] & x[183]);
     layer0_out[228] <= x[1510] | x[1511];
     layer0_out[229] <= x[2626] ^ x[2628];
     layer0_out[230] <= x[2503] & ~x[2505];
     layer0_out[231] <= ~(x[2381] & x[2382]);
     layer0_out[232] <= ~(x[2928] | x[2929]);
     layer0_out[233] <= x[969] | x[971];
     layer0_out[234] <= x[8976] | x[8977];
     layer0_out[235] <= ~(x[3277] & x[3278]);
     layer0_out[236] <= x[8146] ^ x[8147];
     layer0_out[237] <= x[4490] & ~x[4491];
     layer0_out[238] <= ~(x[2562] & x[2564]);
     layer0_out[239] <= ~(x[5721] | x[5722]);
     layer0_out[240] <= ~(x[2732] ^ x[2734]);
     layer0_out[241] <= x[692];
     layer0_out[242] <= x[6299] & x[6300];
     layer0_out[243] <= ~(x[4329] | x[4330]);
     layer0_out[244] <= x[377] ^ x[378];
     layer0_out[245] <= x[2780];
     layer0_out[246] <= x[4061] | x[4062];
     layer0_out[247] <= ~(x[891] ^ x[892]);
     layer0_out[248] <= x[377] & x[379];
     layer0_out[249] <= ~(x[3630] & x[3631]);
     layer0_out[250] <= 1'b1;
     layer0_out[251] <= ~(x[2518] & x[2519]);
     layer0_out[252] <= ~(x[8098] | x[8099]);
     layer0_out[253] <= ~(x[7960] | x[7961]);
     layer0_out[254] <= x[7215];
     layer0_out[255] <= x[432] & x[434];
     layer0_out[256] <= ~(x[995] & x[996]);
     layer0_out[257] <= ~x[1127];
     layer0_out[258] <= x[1561] ^ x[1563];
     layer0_out[259] <= ~(x[1488] & x[1489]);
     layer0_out[260] <= 1'b1;
     layer0_out[261] <= ~(x[5559] & x[5560]);
     layer0_out[262] <= ~(x[2985] & x[2986]);
     layer0_out[263] <= x[6157] | x[6158];
     layer0_out[264] <= ~(x[3252] ^ x[3253]);
     layer0_out[265] <= x[607] ^ x[609];
     layer0_out[266] <= x[8356];
     layer0_out[267] <= x[2714] ^ x[2716];
     layer0_out[268] <= ~(x[6303] ^ x[6304]);
     layer0_out[269] <= x[3687] & ~x[3688];
     layer0_out[270] <= x[1210] & ~x[1209];
     layer0_out[271] <= x[6090] ^ x[6091];
     layer0_out[272] <= ~(x[2725] & x[2726]);
     layer0_out[273] <= x[2679];
     layer0_out[274] <= x[1829] & x[1830];
     layer0_out[275] <= x[8774] & x[8775];
     layer0_out[276] <= ~(x[6130] & x[6131]);
     layer0_out[277] <= x[4877] ^ x[4878];
     layer0_out[278] <= ~(x[5295] & x[5296]);
     layer0_out[279] <= x[7840] ^ x[7841];
     layer0_out[280] <= x[8678];
     layer0_out[281] <= x[565] & ~x[567];
     layer0_out[282] <= x[1322] & x[1323];
     layer0_out[283] <= ~(x[6045] & x[6046]);
     layer0_out[284] <= ~(x[5257] | x[5258]);
     layer0_out[285] <= x[7897] | x[7898];
     layer0_out[286] <= ~(x[866] | x[868]);
     layer0_out[287] <= x[3542] & ~x[3541];
     layer0_out[288] <= ~(x[8082] ^ x[8083]);
     layer0_out[289] <= x[1091] & x[1093];
     layer0_out[290] <= ~x[1848];
     layer0_out[291] <= 1'b1;
     layer0_out[292] <= x[1011] | x[1012];
     layer0_out[293] <= x[8658] & x[8659];
     layer0_out[294] <= ~(x[3581] & x[3582]);
     layer0_out[295] <= ~(x[1554] ^ x[1556]);
     layer0_out[296] <= ~(x[1640] ^ x[1642]);
     layer0_out[297] <= x[924];
     layer0_out[298] <= x[4720] ^ x[4721];
     layer0_out[299] <= x[4744] & x[4745];
     layer0_out[300] <= x[9041] | x[9042];
     layer0_out[301] <= ~(x[6364] | x[6365]);
     layer0_out[302] <= x[2404] & ~x[2403];
     layer0_out[303] <= x[2573] & x[2575];
     layer0_out[304] <= ~(x[3284] | x[3285]);
     layer0_out[305] <= x[6005] & x[6006];
     layer0_out[306] <= ~x[1990];
     layer0_out[307] <= x[8868] ^ x[8869];
     layer0_out[308] <= x[8366] ^ x[8367];
     layer0_out[309] <= x[5181] & x[5182];
     layer0_out[310] <= x[2470] & ~x[2471];
     layer0_out[311] <= x[6542] | x[6543];
     layer0_out[312] <= ~(x[806] | x[808]);
     layer0_out[313] <= x[7176] & ~x[7177];
     layer0_out[314] <= ~(x[1684] & x[1686]);
     layer0_out[315] <= ~x[2705];
     layer0_out[316] <= x[1337] & x[1338];
     layer0_out[317] <= x[8109];
     layer0_out[318] <= ~x[2247];
     layer0_out[319] <= ~(x[7166] | x[7167]);
     layer0_out[320] <= ~(x[717] & x[719]);
     layer0_out[321] <= ~x[6648];
     layer0_out[322] <= 1'b0;
     layer0_out[323] <= x[3233] | x[3234];
     layer0_out[324] <= x[2803] | x[2804];
     layer0_out[325] <= x[5525] | x[5526];
     layer0_out[326] <= x[6893];
     layer0_out[327] <= ~(x[6971] & x[6972]);
     layer0_out[328] <= ~(x[3648] & x[3649]);
     layer0_out[329] <= x[2679] & ~x[2677];
     layer0_out[330] <= x[2298];
     layer0_out[331] <= ~(x[5536] & x[5537]);
     layer0_out[332] <= x[4669] & x[4670];
     layer0_out[333] <= x[4849] ^ x[4850];
     layer0_out[334] <= ~(x[5995] ^ x[5996]);
     layer0_out[335] <= x[5410];
     layer0_out[336] <= ~(x[1382] & x[1383]);
     layer0_out[337] <= x[7808] ^ x[7809];
     layer0_out[338] <= x[5580] & x[5581];
     layer0_out[339] <= x[1489] & x[1490];
     layer0_out[340] <= x[3200];
     layer0_out[341] <= ~x[5894];
     layer0_out[342] <= x[4756] ^ x[4757];
     layer0_out[343] <= x[7935] ^ x[7936];
     layer0_out[344] <= x[77] & x[79];
     layer0_out[345] <= ~x[74];
     layer0_out[346] <= x[2660] & x[2661];
     layer0_out[347] <= ~(x[6533] | x[6534]);
     layer0_out[348] <= x[7736] ^ x[7737];
     layer0_out[349] <= x[6658];
     layer0_out[350] <= x[8883] & ~x[8882];
     layer0_out[351] <= ~(x[5885] & x[5886]);
     layer0_out[352] <= x[8371] | x[8372];
     layer0_out[353] <= x[5962] | x[5963];
     layer0_out[354] <= ~(x[4906] | x[4907]);
     layer0_out[355] <= x[1764] & x[1766];
     layer0_out[356] <= ~(x[1658] & x[1660]);
     layer0_out[357] <= x[4969] & ~x[4968];
     layer0_out[358] <= x[112] ^ x[114];
     layer0_out[359] <= ~(x[8939] | x[8940]);
     layer0_out[360] <= ~(x[1953] & x[1954]);
     layer0_out[361] <= ~(x[2068] & x[2070]);
     layer0_out[362] <= x[808] | x[810];
     layer0_out[363] <= x[457] | x[459];
     layer0_out[364] <= 1'b1;
     layer0_out[365] <= x[4683];
     layer0_out[366] <= ~(x[4418] & x[4419]);
     layer0_out[367] <= x[152] | x[153];
     layer0_out[368] <= ~x[99];
     layer0_out[369] <= ~(x[1657] & x[1658]);
     layer0_out[370] <= x[3678];
     layer0_out[371] <= ~x[6455];
     layer0_out[372] <= x[876] & x[877];
     layer0_out[373] <= ~x[3996] | x[3995];
     layer0_out[374] <= x[7604] | x[7605];
     layer0_out[375] <= ~x[4080] | x[4081];
     layer0_out[376] <= x[6565];
     layer0_out[377] <= ~x[1792] | x[1790];
     layer0_out[378] <= ~x[7689];
     layer0_out[379] <= ~(x[2272] | x[2274]);
     layer0_out[380] <= ~x[4267];
     layer0_out[381] <= x[5961] ^ x[5962];
     layer0_out[382] <= ~x[1983] | x[1982];
     layer0_out[383] <= x[7328] & x[7329];
     layer0_out[384] <= ~(x[2031] | x[2032]);
     layer0_out[385] <= x[902];
     layer0_out[386] <= ~(x[1645] & x[1647]);
     layer0_out[387] <= ~(x[7310] | x[7311]);
     layer0_out[388] <= ~(x[5388] & x[5389]);
     layer0_out[389] <= x[3667];
     layer0_out[390] <= x[4635] & x[4636];
     layer0_out[391] <= x[1322];
     layer0_out[392] <= x[1826] & ~x[1827];
     layer0_out[393] <= x[1921];
     layer0_out[394] <= x[2716] ^ x[2717];
     layer0_out[395] <= ~x[703] | x[701];
     layer0_out[396] <= x[5396] & x[5397];
     layer0_out[397] <= ~(x[1049] & x[1050]);
     layer0_out[398] <= 1'b0;
     layer0_out[399] <= x[821] | x[823];
     layer0_out[400] <= x[3460] & ~x[3459];
     layer0_out[401] <= x[132];
     layer0_out[402] <= ~(x[341] & x[343]);
     layer0_out[403] <= ~x[5622];
     layer0_out[404] <= ~(x[2704] & x[2705]);
     layer0_out[405] <= x[5382] & ~x[5383];
     layer0_out[406] <= ~(x[299] & x[301]);
     layer0_out[407] <= x[5948] & x[5949];
     layer0_out[408] <= x[4019] & x[4020];
     layer0_out[409] <= ~(x[3142] ^ x[3143]);
     layer0_out[410] <= ~(x[9096] & x[9097]);
     layer0_out[411] <= ~(x[5818] & x[5819]);
     layer0_out[412] <= ~(x[6081] | x[6082]);
     layer0_out[413] <= x[2091] & ~x[2092];
     layer0_out[414] <= ~(x[8234] | x[8235]);
     layer0_out[415] <= ~x[8380];
     layer0_out[416] <= x[8281];
     layer0_out[417] <= ~(x[3998] | x[3999]);
     layer0_out[418] <= ~(x[8219] | x[8220]);
     layer0_out[419] <= x[1557] & ~x[1559];
     layer0_out[420] <= ~(x[1814] | x[1816]);
     layer0_out[421] <= x[7616] ^ x[7617];
     layer0_out[422] <= ~x[1127];
     layer0_out[423] <= ~x[6094] | x[6095];
     layer0_out[424] <= ~(x[4578] ^ x[4579]);
     layer0_out[425] <= ~x[6386] | x[6387];
     layer0_out[426] <= ~(x[2659] ^ x[2660]);
     layer0_out[427] <= ~(x[5262] & x[5263]);
     layer0_out[428] <= 1'b1;
     layer0_out[429] <= ~(x[8235] & x[8236]);
     layer0_out[430] <= x[2158] & x[2159];
     layer0_out[431] <= ~(x[835] | x[836]);
     layer0_out[432] <= ~(x[8058] | x[8059]);
     layer0_out[433] <= ~(x[8141] ^ x[8142]);
     layer0_out[434] <= x[2413];
     layer0_out[435] <= ~x[8805];
     layer0_out[436] <= x[7714];
     layer0_out[437] <= ~(x[779] & x[781]);
     layer0_out[438] <= ~(x[4917] | x[4918]);
     layer0_out[439] <= x[2218] & x[2220];
     layer0_out[440] <= x[4596] & ~x[4597];
     layer0_out[441] <= 1'b0;
     layer0_out[442] <= x[653] & x[655];
     layer0_out[443] <= 1'b0;
     layer0_out[444] <= ~x[6280];
     layer0_out[445] <= 1'b1;
     layer0_out[446] <= x[560] & x[561];
     layer0_out[447] <= x[2880] | x[2881];
     layer0_out[448] <= ~(x[4901] & x[4902]);
     layer0_out[449] <= x[5239] & x[5240];
     layer0_out[450] <= x[8164];
     layer0_out[451] <= x[5379] | x[5380];
     layer0_out[452] <= ~(x[9143] | x[9144]);
     layer0_out[453] <= x[4366];
     layer0_out[454] <= x[2];
     layer0_out[455] <= ~(x[1794] & x[1795]);
     layer0_out[456] <= x[1896] & x[1898];
     layer0_out[457] <= ~(x[6016] & x[6017]);
     layer0_out[458] <= ~x[1920];
     layer0_out[459] <= ~(x[728] & x[730]);
     layer0_out[460] <= x[4696];
     layer0_out[461] <= ~x[4278];
     layer0_out[462] <= ~(x[1102] | x[1104]);
     layer0_out[463] <= x[5770];
     layer0_out[464] <= x[845];
     layer0_out[465] <= x[4303] & x[4304];
     layer0_out[466] <= x[6298] | x[6299];
     layer0_out[467] <= x[3345] | x[3346];
     layer0_out[468] <= 1'b0;
     layer0_out[469] <= x[2028] ^ x[2030];
     layer0_out[470] <= ~x[5362] | x[5363];
     layer0_out[471] <= ~(x[272] & x[273]);
     layer0_out[472] <= ~(x[2006] ^ x[2008]);
     layer0_out[473] <= ~(x[1594] & x[1596]);
     layer0_out[474] <= 1'b1;
     layer0_out[475] <= x[697] | x[698];
     layer0_out[476] <= x[6921] | x[6922];
     layer0_out[477] <= x[7525] ^ x[7526];
     layer0_out[478] <= ~(x[9036] | x[9037]);
     layer0_out[479] <= x[1703] & x[1704];
     layer0_out[480] <= ~(x[9082] & x[9083]);
     layer0_out[481] <= x[655] ^ x[657];
     layer0_out[482] <= 1'b1;
     layer0_out[483] <= ~(x[8496] | x[8497]);
     layer0_out[484] <= x[914];
     layer0_out[485] <= ~x[98];
     layer0_out[486] <= x[8869] & x[8870];
     layer0_out[487] <= x[3799] & ~x[3800];
     layer0_out[488] <= ~(x[591] & x[593]);
     layer0_out[489] <= ~(x[1809] | x[1810]);
     layer0_out[490] <= x[7231] & x[7232];
     layer0_out[491] <= ~(x[9201] & x[9202]);
     layer0_out[492] <= ~(x[6549] | x[6550]);
     layer0_out[493] <= x[944];
     layer0_out[494] <= x[894] & x[896];
     layer0_out[495] <= ~x[6189] | x[6188];
     layer0_out[496] <= ~(x[511] & x[513]);
     layer0_out[497] <= ~x[6214] | x[6215];
     layer0_out[498] <= x[909] & x[911];
     layer0_out[499] <= x[5405] | x[5406];
     layer0_out[500] <= ~(x[161] ^ x[163]);
     layer0_out[501] <= x[7974] ^ x[7975];
     layer0_out[502] <= ~x[2354] | x[2356];
     layer0_out[503] <= ~(x[1325] & x[1326]);
     layer0_out[504] <= ~x[6608];
     layer0_out[505] <= x[5611] & x[5612];
     layer0_out[506] <= ~(x[2053] | x[2054]);
     layer0_out[507] <= ~(x[1432] & x[1433]);
     layer0_out[508] <= 1'b1;
     layer0_out[509] <= ~(x[8772] | x[8773]);
     layer0_out[510] <= x[6305];
     layer0_out[511] <= x[1743] & x[1744];
     layer0_out[512] <= x[6326] & ~x[6327];
     layer0_out[513] <= x[2256] & x[2258];
     layer0_out[514] <= x[8860] | x[8861];
     layer0_out[515] <= ~(x[5008] | x[5009]);
     layer0_out[516] <= x[8776] | x[8777];
     layer0_out[517] <= ~x[5283] | x[5284];
     layer0_out[518] <= x[4299] & x[4300];
     layer0_out[519] <= ~x[1704];
     layer0_out[520] <= x[8690] & x[8691];
     layer0_out[521] <= ~x[6002];
     layer0_out[522] <= ~x[537];
     layer0_out[523] <= ~(x[1611] & x[1613]);
     layer0_out[524] <= x[1866] & x[1868];
     layer0_out[525] <= x[938];
     layer0_out[526] <= x[1001] & x[1002];
     layer0_out[527] <= ~x[7893] | x[7894];
     layer0_out[528] <= ~(x[2471] ^ x[2473]);
     layer0_out[529] <= ~(x[3594] ^ x[3595]);
     layer0_out[530] <= ~(x[3871] ^ x[3872]);
     layer0_out[531] <= ~(x[1884] & x[1885]);
     layer0_out[532] <= x[5546] & x[5547];
     layer0_out[533] <= x[4241] & ~x[4240];
     layer0_out[534] <= x[2552] & x[2554];
     layer0_out[535] <= x[50] & x[51];
     layer0_out[536] <= x[9005] | x[9006];
     layer0_out[537] <= ~(x[1255] & x[1256]);
     layer0_out[538] <= x[385];
     layer0_out[539] <= ~(x[3593] & x[3594]);
     layer0_out[540] <= x[168] & x[170];
     layer0_out[541] <= x[5056] & x[5057];
     layer0_out[542] <= x[8890];
     layer0_out[543] <= ~(x[2195] & x[2197]);
     layer0_out[544] <= x[2207] ^ x[2208];
     layer0_out[545] <= x[261] & ~x[259];
     layer0_out[546] <= ~(x[462] & x[463]);
     layer0_out[547] <= x[716] ^ x[718];
     layer0_out[548] <= x[1738] ^ x[1739];
     layer0_out[549] <= ~(x[3694] | x[3695]);
     layer0_out[550] <= ~x[8946];
     layer0_out[551] <= ~(x[8527] | x[8528]);
     layer0_out[552] <= ~x[7650] | x[7649];
     layer0_out[553] <= x[399] | x[400];
     layer0_out[554] <= x[7968] | x[7969];
     layer0_out[555] <= ~(x[3754] | x[3755]);
     layer0_out[556] <= ~(x[870] & x[872]);
     layer0_out[557] <= 1'b1;
     layer0_out[558] <= ~x[7474];
     layer0_out[559] <= ~(x[8422] ^ x[8423]);
     layer0_out[560] <= x[2729] & x[2731];
     layer0_out[561] <= x[1264] | x[1266];
     layer0_out[562] <= x[9025];
     layer0_out[563] <= 1'b1;
     layer0_out[564] <= x[3411] | x[3412];
     layer0_out[565] <= x[6168];
     layer0_out[566] <= ~x[265] | x[263];
     layer0_out[567] <= ~(x[5459] | x[5460]);
     layer0_out[568] <= x[646] & ~x[648];
     layer0_out[569] <= 1'b0;
     layer0_out[570] <= 1'b1;
     layer0_out[571] <= x[4477] | x[4478];
     layer0_out[572] <= x[1945] & x[1947];
     layer0_out[573] <= x[5818];
     layer0_out[574] <= x[1];
     layer0_out[575] <= x[506] & x[507];
     layer0_out[576] <= x[337] & x[338];
     layer0_out[577] <= ~(x[4594] & x[4595]);
     layer0_out[578] <= x[4165] ^ x[4166];
     layer0_out[579] <= ~(x[3037] | x[3038]);
     layer0_out[580] <= x[1245] & x[1247];
     layer0_out[581] <= ~(x[673] ^ x[675]);
     layer0_out[582] <= x[2515] & x[2516];
     layer0_out[583] <= ~(x[9074] & x[9075]);
     layer0_out[584] <= x[2508] & x[2509];
     layer0_out[585] <= ~x[2042] | x[2040];
     layer0_out[586] <= ~(x[812] ^ x[814]);
     layer0_out[587] <= x[2132] & x[2133];
     layer0_out[588] <= x[3625] & x[3626];
     layer0_out[589] <= ~(x[6730] & x[6731]);
     layer0_out[590] <= ~x[4095];
     layer0_out[591] <= ~(x[2729] & x[2730]);
     layer0_out[592] <= ~(x[1159] & x[1161]);
     layer0_out[593] <= x[423] & x[424];
     layer0_out[594] <= ~(x[1404] & x[1406]);
     layer0_out[595] <= 1'b1;
     layer0_out[596] <= x[7946] | x[7947];
     layer0_out[597] <= x[3264];
     layer0_out[598] <= ~x[2620];
     layer0_out[599] <= ~(x[6159] ^ x[6160]);
     layer0_out[600] <= ~(x[4499] & x[4500]);
     layer0_out[601] <= x[2109] | x[2110];
     layer0_out[602] <= x[1409] ^ x[1411];
     layer0_out[603] <= ~(x[1922] & x[1924]);
     layer0_out[604] <= x[2189] ^ x[2191];
     layer0_out[605] <= x[1237];
     layer0_out[606] <= ~(x[1741] & x[1742]);
     layer0_out[607] <= x[4055];
     layer0_out[608] <= 1'b0;
     layer0_out[609] <= x[6667] & x[6668];
     layer0_out[610] <= x[1022];
     layer0_out[611] <= ~(x[1180] & x[1182]);
     layer0_out[612] <= ~(x[7276] ^ x[7277]);
     layer0_out[613] <= ~x[3831];
     layer0_out[614] <= x[939] | x[941];
     layer0_out[615] <= ~x[2960];
     layer0_out[616] <= x[8426];
     layer0_out[617] <= ~(x[6129] & x[6130]);
     layer0_out[618] <= ~x[2313];
     layer0_out[619] <= x[6249] | x[6250];
     layer0_out[620] <= x[5675] & x[5676];
     layer0_out[621] <= 1'b0;
     layer0_out[622] <= x[2346] & x[2348];
     layer0_out[623] <= x[7963] | x[7964];
     layer0_out[624] <= x[2096] & x[2098];
     layer0_out[625] <= ~x[3490];
     layer0_out[626] <= 1'b0;
     layer0_out[627] <= 1'b1;
     layer0_out[628] <= ~(x[648] & x[649]);
     layer0_out[629] <= ~(x[2416] & x[2417]);
     layer0_out[630] <= x[632] & ~x[634];
     layer0_out[631] <= ~(x[7462] ^ x[7463]);
     layer0_out[632] <= x[8957] & x[8958];
     layer0_out[633] <= ~(x[1671] ^ x[1672]);
     layer0_out[634] <= 1'b1;
     layer0_out[635] <= ~(x[7229] | x[7230]);
     layer0_out[636] <= ~(x[8642] | x[8643]);
     layer0_out[637] <= ~(x[1472] & x[1474]);
     layer0_out[638] <= x[1373] ^ x[1375];
     layer0_out[639] <= 1'b1;
     layer0_out[640] <= ~x[9118];
     layer0_out[641] <= ~x[4748];
     layer0_out[642] <= x[8682] | x[8683];
     layer0_out[643] <= x[4590] & ~x[4589];
     layer0_out[644] <= ~(x[4287] ^ x[4288]);
     layer0_out[645] <= x[409];
     layer0_out[646] <= x[1131] & x[1132];
     layer0_out[647] <= x[8338];
     layer0_out[648] <= ~(x[8042] | x[8043]);
     layer0_out[649] <= ~(x[6237] & x[6238]);
     layer0_out[650] <= ~x[7584];
     layer0_out[651] <= x[2015] & x[2017];
     layer0_out[652] <= 1'b1;
     layer0_out[653] <= ~(x[2913] & x[2914]);
     layer0_out[654] <= x[113] & ~x[115];
     layer0_out[655] <= ~(x[1482] & x[1484]);
     layer0_out[656] <= ~(x[660] & x[661]);
     layer0_out[657] <= ~(x[1672] & x[1674]);
     layer0_out[658] <= ~(x[4] & x[6]);
     layer0_out[659] <= ~x[2492] | x[2493];
     layer0_out[660] <= x[8327];
     layer0_out[661] <= ~(x[5036] ^ x[5037]);
     layer0_out[662] <= ~x[3225];
     layer0_out[663] <= ~x[754] | x[752];
     layer0_out[664] <= ~(x[1822] | x[1823]);
     layer0_out[665] <= ~x[8032];
     layer0_out[666] <= ~(x[2456] & x[2457]);
     layer0_out[667] <= x[274] & x[276];
     layer0_out[668] <= ~(x[949] & x[950]);
     layer0_out[669] <= x[1273];
     layer0_out[670] <= ~(x[1031] & x[1032]);
     layer0_out[671] <= x[8156] | x[8157];
     layer0_out[672] <= 1'b1;
     layer0_out[673] <= x[2510];
     layer0_out[674] <= x[4078] | x[4079];
     layer0_out[675] <= ~(x[2642] & x[2644]);
     layer0_out[676] <= 1'b0;
     layer0_out[677] <= 1'b0;
     layer0_out[678] <= ~(x[1873] & x[1875]);
     layer0_out[679] <= x[4778] & ~x[4777];
     layer0_out[680] <= 1'b0;
     layer0_out[681] <= ~x[1886];
     layer0_out[682] <= ~(x[862] & x[864]);
     layer0_out[683] <= x[8709] & ~x[8710];
     layer0_out[684] <= ~x[879];
     layer0_out[685] <= x[5945] & x[5946];
     layer0_out[686] <= ~x[8385];
     layer0_out[687] <= x[276];
     layer0_out[688] <= x[750] & x[752];
     layer0_out[689] <= x[583] & x[584];
     layer0_out[690] <= x[4969] | x[4970];
     layer0_out[691] <= ~(x[1822] & x[1824]);
     layer0_out[692] <= 1'b0;
     layer0_out[693] <= x[1869] & x[1871];
     layer0_out[694] <= 1'b1;
     layer0_out[695] <= ~(x[2323] & x[2325]);
     layer0_out[696] <= ~(x[1720] & x[1721]);
     layer0_out[697] <= ~x[4177];
     layer0_out[698] <= ~(x[679] & x[681]);
     layer0_out[699] <= x[3843] & x[3844];
     layer0_out[700] <= 1'b0;
     layer0_out[701] <= ~(x[1280] | x[1281]);
     layer0_out[702] <= ~(x[6985] ^ x[6986]);
     layer0_out[703] <= x[4257];
     layer0_out[704] <= x[7852];
     layer0_out[705] <= ~(x[6662] | x[6663]);
     layer0_out[706] <= x[8622] | x[8623];
     layer0_out[707] <= ~(x[5065] ^ x[5066]);
     layer0_out[708] <= ~(x[6107] | x[6108]);
     layer0_out[709] <= x[2025] & x[2027];
     layer0_out[710] <= x[3373];
     layer0_out[711] <= 1'b1;
     layer0_out[712] <= x[3584] & x[3585];
     layer0_out[713] <= x[7796];
     layer0_out[714] <= x[4690] | x[4691];
     layer0_out[715] <= ~x[1788];
     layer0_out[716] <= ~(x[6959] | x[6960]);
     layer0_out[717] <= x[1954];
     layer0_out[718] <= x[7082] & x[7083];
     layer0_out[719] <= x[5634] | x[5635];
     layer0_out[720] <= ~(x[3955] | x[3956]);
     layer0_out[721] <= x[925];
     layer0_out[722] <= ~x[4268];
     layer0_out[723] <= ~(x[1630] & x[1632]);
     layer0_out[724] <= x[1828] & x[1829];
     layer0_out[725] <= ~x[5755] | x[5756];
     layer0_out[726] <= x[8540];
     layer0_out[727] <= ~x[1222];
     layer0_out[728] <= ~(x[9028] & x[9029]);
     layer0_out[729] <= ~(x[1396] | x[1398]);
     layer0_out[730] <= x[1591];
     layer0_out[731] <= x[819];
     layer0_out[732] <= ~(x[237] & x[239]);
     layer0_out[733] <= ~(x[617] & x[618]);
     layer0_out[734] <= ~x[7813] | x[7812];
     layer0_out[735] <= x[1094];
     layer0_out[736] <= x[228] | x[229];
     layer0_out[737] <= x[2230] & x[2232];
     layer0_out[738] <= ~(x[6818] & x[6819]);
     layer0_out[739] <= 1'b0;
     layer0_out[740] <= x[5851] & x[5852];
     layer0_out[741] <= ~x[833];
     layer0_out[742] <= x[7851] | x[7852];
     layer0_out[743] <= x[8469] & x[8470];
     layer0_out[744] <= ~(x[4579] & x[4580]);
     layer0_out[745] <= ~(x[6989] ^ x[6990]);
     layer0_out[746] <= x[6245] & x[6246];
     layer0_out[747] <= ~x[204] | x[206];
     layer0_out[748] <= 1'b0;
     layer0_out[749] <= x[5144] & x[5145];
     layer0_out[750] <= ~(x[1225] & x[1226]);
     layer0_out[751] <= ~(x[4468] & x[4469]);
     layer0_out[752] <= ~x[8533];
     layer0_out[753] <= x[2278] | x[2279];
     layer0_out[754] <= ~x[3422];
     layer0_out[755] <= ~(x[1863] & x[1865]);
     layer0_out[756] <= ~x[6362];
     layer0_out[757] <= ~(x[485] ^ x[486]);
     layer0_out[758] <= ~(x[1872] & x[1873]);
     layer0_out[759] <= x[3988] ^ x[3989];
     layer0_out[760] <= ~(x[7831] ^ x[7832]);
     layer0_out[761] <= x[8431] | x[8432];
     layer0_out[762] <= x[7627] | x[7628];
     layer0_out[763] <= x[1454] & x[1455];
     layer0_out[764] <= 1'b1;
     layer0_out[765] <= x[1583] & x[1585];
     layer0_out[766] <= x[770] | x[772];
     layer0_out[767] <= x[2369] & x[2370];
     layer0_out[768] <= x[645] & x[647];
     layer0_out[769] <= x[8081];
     layer0_out[770] <= ~(x[8805] & x[8806]);
     layer0_out[771] <= ~(x[1295] & x[1297]);
     layer0_out[772] <= ~(x[4332] & x[4333]);
     layer0_out[773] <= ~(x[8829] ^ x[8830]);
     layer0_out[774] <= ~(x[1308] | x[1309]);
     layer0_out[775] <= ~x[455];
     layer0_out[776] <= 1'b1;
     layer0_out[777] <= 1'b1;
     layer0_out[778] <= ~(x[2097] & x[2098]);
     layer0_out[779] <= ~x[6803] | x[6802];
     layer0_out[780] <= ~(x[3131] & x[3132]);
     layer0_out[781] <= x[2693] ^ x[2694];
     layer0_out[782] <= x[643] & x[644];
     layer0_out[783] <= ~x[3620];
     layer0_out[784] <= ~x[339];
     layer0_out[785] <= x[1202] & x[1204];
     layer0_out[786] <= x[2737] ^ x[2738];
     layer0_out[787] <= x[2727] ^ x[2728];
     layer0_out[788] <= x[6240] | x[6241];
     layer0_out[789] <= x[4787];
     layer0_out[790] <= ~(x[1418] & x[1419]);
     layer0_out[791] <= x[1831] & x[1832];
     layer0_out[792] <= 1'b0;
     layer0_out[793] <= x[2555] ^ x[2556];
     layer0_out[794] <= ~(x[5992] & x[5993]);
     layer0_out[795] <= ~x[9054];
     layer0_out[796] <= ~(x[4970] | x[4971]);
     layer0_out[797] <= x[6571] ^ x[6572];
     layer0_out[798] <= ~(x[6300] | x[6301]);
     layer0_out[799] <= ~x[6331];
     layer0_out[800] <= ~(x[1085] | x[1086]);
     layer0_out[801] <= ~x[2142];
     layer0_out[802] <= x[8212] | x[8213];
     layer0_out[803] <= 1'b1;
     layer0_out[804] <= x[6231];
     layer0_out[805] <= ~x[830] | x[829];
     layer0_out[806] <= x[2588] & x[2590];
     layer0_out[807] <= x[3236] | x[3237];
     layer0_out[808] <= x[321];
     layer0_out[809] <= x[7999] ^ x[8000];
     layer0_out[810] <= ~x[8375];
     layer0_out[811] <= x[1361] | x[1363];
     layer0_out[812] <= x[8731] | x[8732];
     layer0_out[813] <= x[4789] | x[4790];
     layer0_out[814] <= x[1602] & x[1603];
     layer0_out[815] <= x[8562] & x[8563];
     layer0_out[816] <= x[5402] & x[5403];
     layer0_out[817] <= ~(x[1370] & x[1371]);
     layer0_out[818] <= ~(x[1063] ^ x[1065]);
     layer0_out[819] <= 1'b0;
     layer0_out[820] <= ~(x[4731] & x[4732]);
     layer0_out[821] <= ~(x[5754] & x[5755]);
     layer0_out[822] <= x[4029];
     layer0_out[823] <= x[2462] ^ x[2464];
     layer0_out[824] <= x[2330] & x[2331];
     layer0_out[825] <= x[3669] & x[3670];
     layer0_out[826] <= x[1712];
     layer0_out[827] <= 1'b1;
     layer0_out[828] <= x[211] & x[213];
     layer0_out[829] <= ~(x[4569] ^ x[4570]);
     layer0_out[830] <= x[8326] & ~x[8325];
     layer0_out[831] <= 1'b1;
     layer0_out[832] <= x[260] ^ x[261];
     layer0_out[833] <= x[6935] ^ x[6936];
     layer0_out[834] <= x[9014] & x[9015];
     layer0_out[835] <= x[494];
     layer0_out[836] <= x[4448] | x[4449];
     layer0_out[837] <= ~x[8026] | x[8027];
     layer0_out[838] <= 1'b1;
     layer0_out[839] <= x[2571] & x[2572];
     layer0_out[840] <= x[1924] & ~x[1925];
     layer0_out[841] <= ~(x[349] & x[351]);
     layer0_out[842] <= ~(x[4728] | x[4729]);
     layer0_out[843] <= 1'b1;
     layer0_out[844] <= x[535] & x[537];
     layer0_out[845] <= x[777] & x[778];
     layer0_out[846] <= ~(x[538] & x[539]);
     layer0_out[847] <= x[1419] & x[1420];
     layer0_out[848] <= ~(x[8196] & x[8197]);
     layer0_out[849] <= ~(x[8456] ^ x[8457]);
     layer0_out[850] <= x[6709] & x[6710];
     layer0_out[851] <= x[7261] | x[7262];
     layer0_out[852] <= x[6151] | x[6152];
     layer0_out[853] <= ~x[1071];
     layer0_out[854] <= ~x[1638];
     layer0_out[855] <= ~(x[9099] & x[9100]);
     layer0_out[856] <= ~x[454];
     layer0_out[857] <= x[2184] & x[2186];
     layer0_out[858] <= x[2658];
     layer0_out[859] <= x[7175];
     layer0_out[860] <= ~(x[2275] | x[2277]);
     layer0_out[861] <= ~(x[1718] & x[1719]);
     layer0_out[862] <= ~(x[3993] | x[3994]);
     layer0_out[863] <= ~(x[8559] | x[8560]);
     layer0_out[864] <= x[1435] | x[1437];
     layer0_out[865] <= ~x[1379];
     layer0_out[866] <= ~(x[8879] | x[8880]);
     layer0_out[867] <= x[2029] & x[2030];
     layer0_out[868] <= x[8338];
     layer0_out[869] <= x[78] & ~x[77];
     layer0_out[870] <= x[4443] & x[4444];
     layer0_out[871] <= x[1802] & x[1803];
     layer0_out[872] <= ~(x[8330] | x[8331]);
     layer0_out[873] <= x[1569] & x[1571];
     layer0_out[874] <= ~(x[2931] & x[2932]);
     layer0_out[875] <= 1'b0;
     layer0_out[876] <= ~(x[6836] & x[6837]);
     layer0_out[877] <= x[2376] & x[2378];
     layer0_out[878] <= 1'b0;
     layer0_out[879] <= x[1642] | x[1644];
     layer0_out[880] <= x[9114];
     layer0_out[881] <= 1'b0;
     layer0_out[882] <= x[264] & ~x[266];
     layer0_out[883] <= ~x[7209];
     layer0_out[884] <= x[2674] & ~x[2672];
     layer0_out[885] <= x[1603] ^ x[1605];
     layer0_out[886] <= ~(x[109] & x[110]);
     layer0_out[887] <= x[215] & x[217];
     layer0_out[888] <= 1'b1;
     layer0_out[889] <= ~(x[3209] | x[3210]);
     layer0_out[890] <= x[216] ^ x[217];
     layer0_out[891] <= ~x[6575];
     layer0_out[892] <= ~(x[279] & x[280]);
     layer0_out[893] <= x[7837] | x[7838];
     layer0_out[894] <= x[2092] & x[2094];
     layer0_out[895] <= ~(x[4184] | x[4185]);
     layer0_out[896] <= ~(x[3022] & x[3023]);
     layer0_out[897] <= ~(x[96] & x[98]);
     layer0_out[898] <= x[4914] & x[4915];
     layer0_out[899] <= x[1656] | x[1657];
     layer0_out[900] <= x[6378];
     layer0_out[901] <= ~(x[2390] & x[2391]);
     layer0_out[902] <= ~x[2173];
     layer0_out[903] <= x[4945] ^ x[4946];
     layer0_out[904] <= x[2546] & x[2547];
     layer0_out[905] <= ~x[1761] | x[1760];
     layer0_out[906] <= x[839];
     layer0_out[907] <= ~(x[1730] & x[1731]);
     layer0_out[908] <= ~(x[7017] & x[7018]);
     layer0_out[909] <= ~(x[7345] | x[7346]);
     layer0_out[910] <= x[7705] | x[7706];
     layer0_out[911] <= ~(x[6329] ^ x[6330]);
     layer0_out[912] <= x[2139] & x[2141];
     layer0_out[913] <= ~(x[6572] | x[6573]);
     layer0_out[914] <= x[3725];
     layer0_out[915] <= ~(x[3905] | x[3906]);
     layer0_out[916] <= x[1653] ^ x[1655];
     layer0_out[917] <= x[638];
     layer0_out[918] <= ~(x[586] & x[588]);
     layer0_out[919] <= x[7174];
     layer0_out[920] <= 1'b0;
     layer0_out[921] <= x[3697] | x[3698];
     layer0_out[922] <= ~(x[2943] | x[2944]);
     layer0_out[923] <= x[4702] & x[4703];
     layer0_out[924] <= x[8114] & ~x[8113];
     layer0_out[925] <= x[702] & x[704];
     layer0_out[926] <= ~(x[2436] | x[2438]);
     layer0_out[927] <= x[3577] & ~x[3576];
     layer0_out[928] <= x[2689] ^ x[2691];
     layer0_out[929] <= x[8404] & x[8405];
     layer0_out[930] <= ~(x[943] | x[945]);
     layer0_out[931] <= ~x[296];
     layer0_out[932] <= x[2782] ^ x[2783];
     layer0_out[933] <= ~(x[1090] ^ x[1091]);
     layer0_out[934] <= x[1956] | x[1958];
     layer0_out[935] <= 1'b1;
     layer0_out[936] <= x[2348] & x[2349];
     layer0_out[937] <= ~(x[3759] & x[3760]);
     layer0_out[938] <= x[4745] | x[4746];
     layer0_out[939] <= x[1046] & ~x[1048];
     layer0_out[940] <= ~(x[2258] | x[2259]);
     layer0_out[941] <= ~(x[3336] ^ x[3337]);
     layer0_out[942] <= ~(x[2492] & x[2494]);
     layer0_out[943] <= x[1303] & x[1305];
     layer0_out[944] <= ~(x[1474] & x[1475]);
     layer0_out[945] <= ~x[862];
     layer0_out[946] <= x[2199] ^ x[2200];
     layer0_out[947] <= x[1005] & x[1006];
     layer0_out[948] <= ~(x[7088] ^ x[7089]);
     layer0_out[949] <= x[2017] ^ x[2018];
     layer0_out[950] <= ~x[4967];
     layer0_out[951] <= x[9177] ^ x[9178];
     layer0_out[952] <= x[535] ^ x[536];
     layer0_out[953] <= x[8362];
     layer0_out[954] <= ~(x[706] ^ x[708]);
     layer0_out[955] <= x[5225] & x[5226];
     layer0_out[956] <= ~(x[5586] & x[5587]);
     layer0_out[957] <= x[1356] & x[1358];
     layer0_out[958] <= x[6366] | x[6367];
     layer0_out[959] <= ~(x[5740] & x[5741]);
     layer0_out[960] <= ~x[94];
     layer0_out[961] <= ~(x[1756] & x[1757]);
     layer0_out[962] <= x[8336] | x[8337];
     layer0_out[963] <= x[2137] & x[2138];
     layer0_out[964] <= ~x[2417];
     layer0_out[965] <= 1'b0;
     layer0_out[966] <= x[86] & x[88];
     layer0_out[967] <= x[6275];
     layer0_out[968] <= ~(x[2125] & x[2126]);
     layer0_out[969] <= ~x[1993];
     layer0_out[970] <= x[6918] ^ x[6919];
     layer0_out[971] <= x[544] ^ x[546];
     layer0_out[972] <= ~(x[5131] | x[5132]);
     layer0_out[973] <= ~(x[8262] & x[8263]);
     layer0_out[974] <= x[268] & x[269];
     layer0_out[975] <= ~x[1876];
     layer0_out[976] <= x[809];
     layer0_out[977] <= ~(x[1350] & x[1352]);
     layer0_out[978] <= ~(x[457] & x[458]);
     layer0_out[979] <= ~x[527];
     layer0_out[980] <= ~(x[84] | x[86]);
     layer0_out[981] <= x[3306];
     layer0_out[982] <= ~x[654];
     layer0_out[983] <= ~(x[2520] ^ x[2522]);
     layer0_out[984] <= x[5850] & x[5851];
     layer0_out[985] <= ~(x[5714] | x[5715]);
     layer0_out[986] <= 1'b1;
     layer0_out[987] <= ~(x[5174] & x[5175]);
     layer0_out[988] <= ~(x[2127] & x[2128]);
     layer0_out[989] <= ~(x[8771] | x[8772]);
     layer0_out[990] <= x[2096];
     layer0_out[991] <= x[4911] | x[4912];
     layer0_out[992] <= ~(x[2649] & x[2651]);
     layer0_out[993] <= ~(x[1705] & x[1706]);
     layer0_out[994] <= ~x[3971] | x[3970];
     layer0_out[995] <= x[8564] & x[8565];
     layer0_out[996] <= ~x[2145];
     layer0_out[997] <= x[946] & x[948];
     layer0_out[998] <= x[621] & x[622];
     layer0_out[999] <= x[3858] ^ x[3859];
     layer0_out[1000] <= ~(x[997] & x[998]);
     layer0_out[1001] <= x[5149] & x[5150];
     layer0_out[1002] <= x[7] ^ x[8];
     layer0_out[1003] <= ~(x[4572] & x[4573]);
     layer0_out[1004] <= ~(x[7116] & x[7117]);
     layer0_out[1005] <= x[2923] & ~x[2924];
     layer0_out[1006] <= x[5193];
     layer0_out[1007] <= x[125] | x[126];
     layer0_out[1008] <= ~(x[5363] & x[5364]);
     layer0_out[1009] <= ~(x[5807] & x[5808]);
     layer0_out[1010] <= x[768];
     layer0_out[1011] <= x[2424];
     layer0_out[1012] <= ~x[1670];
     layer0_out[1013] <= ~(x[2138] & x[2139]);
     layer0_out[1014] <= ~(x[7517] ^ x[7518]);
     layer0_out[1015] <= x[2432] & x[2434];
     layer0_out[1016] <= x[7502] ^ x[7503];
     layer0_out[1017] <= x[6125] & x[6126];
     layer0_out[1018] <= ~(x[3907] ^ x[3908]);
     layer0_out[1019] <= x[4413];
     layer0_out[1020] <= ~(x[4705] | x[4706]);
     layer0_out[1021] <= ~(x[300] ^ x[301]);
     layer0_out[1022] <= x[1059] | x[1061];
     layer0_out[1023] <= ~x[4734];
     layer0_out[1024] <= x[3247];
     layer0_out[1025] <= ~x[3746];
     layer0_out[1026] <= 1'b0;
     layer0_out[1027] <= x[7658];
     layer0_out[1028] <= 1'b1;
     layer0_out[1029] <= 1'b0;
     layer0_out[1030] <= x[7570];
     layer0_out[1031] <= x[4289] & x[4290];
     layer0_out[1032] <= x[6886];
     layer0_out[1033] <= ~(x[4442] | x[4443]);
     layer0_out[1034] <= 1'b1;
     layer0_out[1035] <= x[611] ^ x[612];
     layer0_out[1036] <= x[4754] | x[4755];
     layer0_out[1037] <= ~(x[6597] & x[6598]);
     layer0_out[1038] <= x[8894] & x[8895];
     layer0_out[1039] <= ~x[1660];
     layer0_out[1040] <= ~x[5604];
     layer0_out[1041] <= ~x[1456] | x[1458];
     layer0_out[1042] <= ~(x[6801] | x[6802]);
     layer0_out[1043] <= ~x[2607] | x[2606];
     layer0_out[1044] <= x[9159] ^ x[9160];
     layer0_out[1045] <= x[296] & ~x[298];
     layer0_out[1046] <= 1'b0;
     layer0_out[1047] <= x[6486] | x[6487];
     layer0_out[1048] <= ~x[7581];
     layer0_out[1049] <= ~x[7854];
     layer0_out[1050] <= 1'b0;
     layer0_out[1051] <= ~(x[1436] & x[1438]);
     layer0_out[1052] <= x[5004] ^ x[5005];
     layer0_out[1053] <= ~x[8796] | x[8795];
     layer0_out[1054] <= ~(x[2383] & x[2385]);
     layer0_out[1055] <= x[8742] ^ x[8743];
     layer0_out[1056] <= x[4883] | x[4884];
     layer0_out[1057] <= x[6095] & x[6096];
     layer0_out[1058] <= 1'b0;
     layer0_out[1059] <= ~(x[2407] & x[2408]);
     layer0_out[1060] <= x[379] | x[381];
     layer0_out[1061] <= x[1961] | x[1962];
     layer0_out[1062] <= ~(x[2314] & x[2316]);
     layer0_out[1063] <= x[1939];
     layer0_out[1064] <= ~x[2046];
     layer0_out[1065] <= ~x[7482];
     layer0_out[1066] <= x[520] & x[521];
     layer0_out[1067] <= ~(x[75] & x[76]);
     layer0_out[1068] <= ~(x[314] | x[315]);
     layer0_out[1069] <= 1'b0;
     layer0_out[1070] <= x[7031] & ~x[7030];
     layer0_out[1071] <= x[7609] & x[7610];
     layer0_out[1072] <= ~(x[1302] & x[1303]);
     layer0_out[1073] <= x[921] | x[922];
     layer0_out[1074] <= x[6489] & x[6490];
     layer0_out[1075] <= ~x[1923] | x[1924];
     layer0_out[1076] <= x[8290] | x[8291];
     layer0_out[1077] <= x[2389] ^ x[2391];
     layer0_out[1078] <= x[672] ^ x[673];
     layer0_out[1079] <= x[3947] | x[3948];
     layer0_out[1080] <= x[1702] | x[1703];
     layer0_out[1081] <= x[6526] & ~x[6525];
     layer0_out[1082] <= x[7101];
     layer0_out[1083] <= ~(x[633] ^ x[635]);
     layer0_out[1084] <= ~(x[7820] | x[7821]);
     layer0_out[1085] <= ~(x[1950] & x[1951]);
     layer0_out[1086] <= ~(x[2076] | x[2077]);
     layer0_out[1087] <= ~(x[3730] ^ x[3731]);
     layer0_out[1088] <= x[7627];
     layer0_out[1089] <= x[4262] ^ x[4263];
     layer0_out[1090] <= x[2032] & ~x[2034];
     layer0_out[1091] <= x[7700] & x[7701];
     layer0_out[1092] <= ~(x[2218] & x[2219]);
     layer0_out[1093] <= ~(x[9011] ^ x[9012]);
     layer0_out[1094] <= ~(x[318] & x[319]);
     layer0_out[1095] <= x[9063] & ~x[9062];
     layer0_out[1096] <= ~(x[722] & x[723]);
     layer0_out[1097] <= ~(x[6983] ^ x[6984]);
     layer0_out[1098] <= ~(x[8181] | x[8182]);
     layer0_out[1099] <= ~x[2577] | x[2576];
     layer0_out[1100] <= ~x[530];
     layer0_out[1101] <= x[670] | x[672];
     layer0_out[1102] <= ~(x[1848] & x[1849]);
     layer0_out[1103] <= x[1081] & x[1083];
     layer0_out[1104] <= x[8072] ^ x[8073];
     layer0_out[1105] <= ~(x[2085] & x[2087]);
     layer0_out[1106] <= ~x[565] | x[564];
     layer0_out[1107] <= ~x[1523];
     layer0_out[1108] <= x[1650] & x[1651];
     layer0_out[1109] <= ~(x[4394] & x[4395]);
     layer0_out[1110] <= ~(x[17] & x[19]);
     layer0_out[1111] <= ~(x[889] ^ x[890]);
     layer0_out[1112] <= x[5535] & x[5536];
     layer0_out[1113] <= x[4340] | x[4341];
     layer0_out[1114] <= ~(x[6416] | x[6417]);
     layer0_out[1115] <= 1'b0;
     layer0_out[1116] <= 1'b1;
     layer0_out[1117] <= ~(x[5452] & x[5453]);
     layer0_out[1118] <= ~x[8510] | x[8509];
     layer0_out[1119] <= x[1139];
     layer0_out[1120] <= ~(x[2299] ^ x[2301]);
     layer0_out[1121] <= ~(x[4420] & x[4421]);
     layer0_out[1122] <= x[1576];
     layer0_out[1123] <= x[7102] | x[7103];
     layer0_out[1124] <= ~x[8474];
     layer0_out[1125] <= ~(x[7050] ^ x[7051]);
     layer0_out[1126] <= x[6354] | x[6355];
     layer0_out[1127] <= ~(x[5761] & x[5762]);
     layer0_out[1128] <= ~(x[8352] & x[8353]);
     layer0_out[1129] <= x[3703] & ~x[3702];
     layer0_out[1130] <= x[5443] & x[5444];
     layer0_out[1131] <= ~(x[1124] & x[1126]);
     layer0_out[1132] <= x[7438] | x[7439];
     layer0_out[1133] <= x[7491] | x[7492];
     layer0_out[1134] <= ~x[3009];
     layer0_out[1135] <= x[2391] & x[2393];
     layer0_out[1136] <= x[982] | x[984];
     layer0_out[1137] <= x[8850] & x[8851];
     layer0_out[1138] <= ~(x[392] | x[393]);
     layer0_out[1139] <= x[4333] & x[4334];
     layer0_out[1140] <= ~(x[1406] ^ x[1407]);
     layer0_out[1141] <= x[738] | x[739];
     layer0_out[1142] <= ~(x[2260] & x[2261]);
     layer0_out[1143] <= ~(x[861] & x[863]);
     layer0_out[1144] <= ~(x[814] & x[815]);
     layer0_out[1145] <= ~(x[5477] & x[5478]);
     layer0_out[1146] <= x[3638] ^ x[3639];
     layer0_out[1147] <= ~(x[2030] & x[2032]);
     layer0_out[1148] <= x[2375] & ~x[2376];
     layer0_out[1149] <= 1'b0;
     layer0_out[1150] <= ~(x[9137] | x[9138]);
     layer0_out[1151] <= ~(x[5210] & x[5211]);
     layer0_out[1152] <= ~(x[246] & x[247]);
     layer0_out[1153] <= ~x[306];
     layer0_out[1154] <= ~(x[8345] & x[8346]);
     layer0_out[1155] <= x[2314] & x[2315];
     layer0_out[1156] <= ~x[6325] | x[6326];
     layer0_out[1157] <= x[8011] & ~x[8012];
     layer0_out[1158] <= ~(x[3729] & x[3730]);
     layer0_out[1159] <= x[690];
     layer0_out[1160] <= x[589] & x[591];
     layer0_out[1161] <= x[1969] & x[1971];
     layer0_out[1162] <= ~(x[568] | x[569]);
     layer0_out[1163] <= ~(x[2044] & x[2045]);
     layer0_out[1164] <= ~(x[822] ^ x[823]);
     layer0_out[1165] <= x[5534];
     layer0_out[1166] <= ~(x[1625] & x[1627]);
     layer0_out[1167] <= ~(x[2706] & x[2707]);
     layer0_out[1168] <= x[1295] & x[1296];
     layer0_out[1169] <= x[2715] ^ x[2716];
     layer0_out[1170] <= ~(x[1086] & x[1087]);
     layer0_out[1171] <= ~(x[2821] & x[2822]);
     layer0_out[1172] <= ~x[3890];
     layer0_out[1173] <= ~(x[7650] | x[7651]);
     layer0_out[1174] <= x[2014] & x[2015];
     layer0_out[1175] <= ~(x[3329] ^ x[3330]);
     layer0_out[1176] <= x[1771] ^ x[1773];
     layer0_out[1177] <= x[852] | x[854];
     layer0_out[1178] <= 1'b0;
     layer0_out[1179] <= ~(x[4782] | x[4783]);
     layer0_out[1180] <= x[2462] | x[2463];
     layer0_out[1181] <= x[1646];
     layer0_out[1182] <= x[813] & x[814];
     layer0_out[1183] <= ~x[2630] | x[2632];
     layer0_out[1184] <= ~x[5766];
     layer0_out[1185] <= x[3636];
     layer0_out[1186] <= ~x[7755];
     layer0_out[1187] <= ~(x[4406] & x[4407]);
     layer0_out[1188] <= x[8309];
     layer0_out[1189] <= ~(x[3238] | x[3239]);
     layer0_out[1190] <= x[8414] & x[8415];
     layer0_out[1191] <= x[6701];
     layer0_out[1192] <= ~x[6076] | x[6077];
     layer0_out[1193] <= ~x[1977] | x[1978];
     layer0_out[1194] <= x[490] | x[492];
     layer0_out[1195] <= x[6524] | x[6525];
     layer0_out[1196] <= x[3614] ^ x[3615];
     layer0_out[1197] <= ~(x[1351] ^ x[1352]);
     layer0_out[1198] <= ~(x[4120] | x[4121]);
     layer0_out[1199] <= 1'b0;
     layer0_out[1200] <= x[353] | x[354];
     layer0_out[1201] <= x[3758] | x[3759];
     layer0_out[1202] <= 1'b1;
     layer0_out[1203] <= x[3902] & ~x[3903];
     layer0_out[1204] <= x[5526];
     layer0_out[1205] <= ~(x[1124] ^ x[1125]);
     layer0_out[1206] <= x[5245] & x[5246];
     layer0_out[1207] <= x[6803] | x[6804];
     layer0_out[1208] <= x[952] | x[953];
     layer0_out[1209] <= x[6807] ^ x[6808];
     layer0_out[1210] <= ~(x[8432] | x[8433]);
     layer0_out[1211] <= x[7541] | x[7542];
     layer0_out[1212] <= x[2684] & x[2685];
     layer0_out[1213] <= 1'b1;
     layer0_out[1214] <= ~(x[2840] & x[2841]);
     layer0_out[1215] <= ~x[7130] | x[7131];
     layer0_out[1216] <= ~(x[2968] | x[2969]);
     layer0_out[1217] <= ~(x[8888] ^ x[8889]);
     layer0_out[1218] <= ~x[448];
     layer0_out[1219] <= x[2022] & x[2024];
     layer0_out[1220] <= x[1549];
     layer0_out[1221] <= x[1677] ^ x[1679];
     layer0_out[1222] <= ~(x[3032] & x[3033]);
     layer0_out[1223] <= ~(x[5583] & x[5584]);
     layer0_out[1224] <= x[432] & ~x[431];
     layer0_out[1225] <= ~(x[7026] & x[7027]);
     layer0_out[1226] <= ~x[6674] | x[6675];
     layer0_out[1227] <= ~x[8852];
     layer0_out[1228] <= x[4314] | x[4315];
     layer0_out[1229] <= ~(x[4461] | x[4462]);
     layer0_out[1230] <= x[7763] | x[7764];
     layer0_out[1231] <= x[2251] ^ x[2253];
     layer0_out[1232] <= ~(x[6449] | x[6450]);
     layer0_out[1233] <= x[6889] | x[6890];
     layer0_out[1234] <= x[5584] & x[5585];
     layer0_out[1235] <= ~(x[8512] ^ x[8513]);
     layer0_out[1236] <= x[5887] | x[5888];
     layer0_out[1237] <= ~(x[4974] ^ x[4975]);
     layer0_out[1238] <= ~(x[4186] | x[4187]);
     layer0_out[1239] <= x[7578];
     layer0_out[1240] <= ~x[2069];
     layer0_out[1241] <= x[3248] | x[3249];
     layer0_out[1242] <= ~(x[6585] | x[6586]);
     layer0_out[1243] <= ~x[3166];
     layer0_out[1244] <= x[1931] | x[1932];
     layer0_out[1245] <= ~(x[9146] | x[9147]);
     layer0_out[1246] <= ~(x[2025] & x[2026]);
     layer0_out[1247] <= x[7600] | x[7601];
     layer0_out[1248] <= ~(x[7951] ^ x[7952]);
     layer0_out[1249] <= ~(x[2507] & x[2509]);
     layer0_out[1250] <= ~(x[7474] | x[7475]);
     layer0_out[1251] <= x[4603] & ~x[4602];
     layer0_out[1252] <= x[2304] & x[2305];
     layer0_out[1253] <= ~x[93];
     layer0_out[1254] <= x[6255];
     layer0_out[1255] <= ~x[2186];
     layer0_out[1256] <= ~(x[1998] & x[2000]);
     layer0_out[1257] <= x[5505] & x[5506];
     layer0_out[1258] <= x[8287] & x[8288];
     layer0_out[1259] <= ~(x[1757] | x[1758]);
     layer0_out[1260] <= ~x[8024] | x[8023];
     layer0_out[1261] <= x[5218] & x[5219];
     layer0_out[1262] <= ~(x[7311] | x[7312]);
     layer0_out[1263] <= ~(x[127] & x[128]);
     layer0_out[1264] <= x[5103] | x[5104];
     layer0_out[1265] <= x[1355] & x[1357];
     layer0_out[1266] <= 1'b1;
     layer0_out[1267] <= ~(x[1617] & x[1618]);
     layer0_out[1268] <= x[5682] & x[5683];
     layer0_out[1269] <= x[6072] & x[6073];
     layer0_out[1270] <= ~x[1074];
     layer0_out[1271] <= x[5871] & x[5872];
     layer0_out[1272] <= ~x[6916];
     layer0_out[1273] <= x[2549] & x[2550];
     layer0_out[1274] <= x[4051] | x[4052];
     layer0_out[1275] <= 1'b0;
     layer0_out[1276] <= x[6378] | x[6379];
     layer0_out[1277] <= x[4001] | x[4002];
     layer0_out[1278] <= ~(x[2306] & x[2308]);
     layer0_out[1279] <= x[8657] & x[8658];
     layer0_out[1280] <= x[5825] & x[5826];
     layer0_out[1281] <= ~(x[6655] & x[6656]);
     layer0_out[1282] <= x[8377] & x[8378];
     layer0_out[1283] <= ~(x[1214] | x[1216]);
     layer0_out[1284] <= ~x[621] | x[623];
     layer0_out[1285] <= ~(x[1563] & x[1564]);
     layer0_out[1286] <= ~(x[89] & x[91]);
     layer0_out[1287] <= ~(x[8402] | x[8403]);
     layer0_out[1288] <= x[7283] & ~x[7282];
     layer0_out[1289] <= x[7129];
     layer0_out[1290] <= ~(x[1254] & x[1256]);
     layer0_out[1291] <= x[1968] & x[1970];
     layer0_out[1292] <= 1'b0;
     layer0_out[1293] <= x[5266];
     layer0_out[1294] <= x[8197] | x[8198];
     layer0_out[1295] <= ~(x[8918] & x[8919]);
     layer0_out[1296] <= 1'b1;
     layer0_out[1297] <= 1'b1;
     layer0_out[1298] <= ~(x[4581] & x[4582]);
     layer0_out[1299] <= x[2554] & x[2556];
     layer0_out[1300] <= ~(x[718] | x[720]);
     layer0_out[1301] <= 1'b0;
     layer0_out[1302] <= ~(x[624] & x[625]);
     layer0_out[1303] <= ~(x[255] | x[257]);
     layer0_out[1304] <= x[4978] | x[4979];
     layer0_out[1305] <= ~x[4896];
     layer0_out[1306] <= 1'b0;
     layer0_out[1307] <= x[5484] & x[5485];
     layer0_out[1308] <= 1'b0;
     layer0_out[1309] <= ~(x[1656] & x[1658]);
     layer0_out[1310] <= x[269] & x[270];
     layer0_out[1311] <= ~(x[8725] | x[8726]);
     layer0_out[1312] <= 1'b1;
     layer0_out[1313] <= 1'b0;
     layer0_out[1314] <= ~(x[1595] & x[1597]);
     layer0_out[1315] <= ~x[4597] | x[4598];
     layer0_out[1316] <= ~x[240];
     layer0_out[1317] <= x[4244] ^ x[4245];
     layer0_out[1318] <= x[8574] & x[8575];
     layer0_out[1319] <= ~x[2106];
     layer0_out[1320] <= ~(x[681] ^ x[683]);
     layer0_out[1321] <= ~(x[1006] | x[1008]);
     layer0_out[1322] <= x[1257];
     layer0_out[1323] <= x[7950];
     layer0_out[1324] <= x[7494] & x[7495];
     layer0_out[1325] <= x[2480] & x[2481];
     layer0_out[1326] <= x[699] | x[701];
     layer0_out[1327] <= ~(x[5939] & x[5940]);
     layer0_out[1328] <= x[825];
     layer0_out[1329] <= ~x[4417];
     layer0_out[1330] <= ~(x[4530] | x[4531]);
     layer0_out[1331] <= ~x[2043];
     layer0_out[1332] <= ~(x[1313] & x[1315]);
     layer0_out[1333] <= ~x[6439];
     layer0_out[1334] <= ~x[1446];
     layer0_out[1335] <= ~x[3005];
     layer0_out[1336] <= ~x[6236];
     layer0_out[1337] <= x[2733];
     layer0_out[1338] <= ~(x[1700] & x[1701]);
     layer0_out[1339] <= ~(x[1891] & x[1892]);
     layer0_out[1340] <= 1'b0;
     layer0_out[1341] <= ~(x[150] ^ x[152]);
     layer0_out[1342] <= ~(x[7156] | x[7157]);
     layer0_out[1343] <= x[1975] ^ x[1977];
     layer0_out[1344] <= x[136] ^ x[137];
     layer0_out[1345] <= x[610] ^ x[612];
     layer0_out[1346] <= x[513] ^ x[514];
     layer0_out[1347] <= ~x[1867];
     layer0_out[1348] <= ~(x[722] | x[724]);
     layer0_out[1349] <= x[5067] ^ x[5068];
     layer0_out[1350] <= ~(x[1805] ^ x[1806]);
     layer0_out[1351] <= x[1307] | x[1309];
     layer0_out[1352] <= ~x[5495];
     layer0_out[1353] <= 1'b0;
     layer0_out[1354] <= x[5516] | x[5517];
     layer0_out[1355] <= ~(x[4803] & x[4804]);
     layer0_out[1356] <= x[135] | x[136];
     layer0_out[1357] <= x[282] ^ x[284];
     layer0_out[1358] <= x[1097] | x[1099];
     layer0_out[1359] <= ~(x[6339] | x[6340]);
     layer0_out[1360] <= ~(x[1161] & x[1162]);
     layer0_out[1361] <= x[4798] | x[4799];
     layer0_out[1362] <= ~(x[4280] & x[4281]);
     layer0_out[1363] <= x[5455];
     layer0_out[1364] <= ~(x[447] & x[449]);
     layer0_out[1365] <= x[2122] ^ x[2123];
     layer0_out[1366] <= ~(x[5624] & x[5625]);
     layer0_out[1367] <= x[6945];
     layer0_out[1368] <= x[1457] ^ x[1459];
     layer0_out[1369] <= ~(x[23] & x[25]);
     layer0_out[1370] <= ~x[3354];
     layer0_out[1371] <= 1'b0;
     layer0_out[1372] <= ~(x[1385] & x[1386]);
     layer0_out[1373] <= ~(x[1697] ^ x[1699]);
     layer0_out[1374] <= ~(x[3080] ^ x[3081]);
     layer0_out[1375] <= x[3852] ^ x[3853];
     layer0_out[1376] <= 1'b1;
     layer0_out[1377] <= ~(x[4562] ^ x[4563]);
     layer0_out[1378] <= ~(x[3128] | x[3129]);
     layer0_out[1379] <= ~(x[1181] ^ x[1182]);
     layer0_out[1380] <= ~x[7192];
     layer0_out[1381] <= ~(x[2091] & x[2093]);
     layer0_out[1382] <= ~(x[4773] | x[4774]);
     layer0_out[1383] <= x[7769];
     layer0_out[1384] <= ~(x[275] ^ x[276]);
     layer0_out[1385] <= ~x[8179];
     layer0_out[1386] <= ~x[6242];
     layer0_out[1387] <= ~x[6577];
     layer0_out[1388] <= ~x[2523];
     layer0_out[1389] <= x[2644] & x[2645];
     layer0_out[1390] <= ~x[6039];
     layer0_out[1391] <= x[2037] | x[2038];
     layer0_out[1392] <= x[201] | x[202];
     layer0_out[1393] <= ~(x[7890] & x[7891]);
     layer0_out[1394] <= ~(x[6846] | x[6847]);
     layer0_out[1395] <= ~(x[551] ^ x[552]);
     layer0_out[1396] <= ~(x[5474] ^ x[5475]);
     layer0_out[1397] <= x[249] | x[250];
     layer0_out[1398] <= ~(x[239] & x[241]);
     layer0_out[1399] <= 1'b1;
     layer0_out[1400] <= x[2449] & x[2451];
     layer0_out[1401] <= ~x[5501];
     layer0_out[1402] <= ~(x[2242] & x[2243]);
     layer0_out[1403] <= ~(x[2572] & x[2574]);
     layer0_out[1404] <= 1'b0;
     layer0_out[1405] <= x[7195];
     layer0_out[1406] <= ~x[552] | x[554];
     layer0_out[1407] <= ~(x[1936] & x[1938]);
     layer0_out[1408] <= x[1410] & x[1411];
     layer0_out[1409] <= ~(x[3575] ^ x[3576]);
     layer0_out[1410] <= x[8192];
     layer0_out[1411] <= ~(x[4074] ^ x[4075]);
     layer0_out[1412] <= ~x[779] | x[778];
     layer0_out[1413] <= ~x[5110];
     layer0_out[1414] <= ~(x[445] & x[447]);
     layer0_out[1415] <= x[6740] & x[6741];
     layer0_out[1416] <= x[1080];
     layer0_out[1417] <= x[3337] ^ x[3338];
     layer0_out[1418] <= x[9087] & x[9088];
     layer0_out[1419] <= ~x[3821];
     layer0_out[1420] <= x[8401] & x[8402];
     layer0_out[1421] <= ~(x[2623] & x[2625]);
     layer0_out[1422] <= x[2829] & x[2830];
     layer0_out[1423] <= ~(x[6725] & x[6726]);
     layer0_out[1424] <= x[2197] ^ x[2199];
     layer0_out[1425] <= x[4011] ^ x[4012];
     layer0_out[1426] <= x[7245] & x[7246];
     layer0_out[1427] <= ~(x[7982] | x[7983]);
     layer0_out[1428] <= x[1108] ^ x[1109];
     layer0_out[1429] <= x[2780] ^ x[2782];
     layer0_out[1430] <= ~x[8295];
     layer0_out[1431] <= x[666] ^ x[668];
     layer0_out[1432] <= ~(x[3191] ^ x[3192]);
     layer0_out[1433] <= ~x[4066];
     layer0_out[1434] <= x[4131] & x[4132];
     layer0_out[1435] <= x[19] & x[21];
     layer0_out[1436] <= ~(x[2519] & x[2520]);
     layer0_out[1437] <= x[8904];
     layer0_out[1438] <= x[576];
     layer0_out[1439] <= ~(x[5401] ^ x[5402]);
     layer0_out[1440] <= x[299] & ~x[298];
     layer0_out[1441] <= ~(x[2553] & x[2555]);
     layer0_out[1442] <= ~(x[4605] | x[4606]);
     layer0_out[1443] <= x[643] ^ x[645];
     layer0_out[1444] <= x[1745];
     layer0_out[1445] <= ~(x[8614] & x[8615]);
     layer0_out[1446] <= ~(x[6305] | x[6306]);
     layer0_out[1447] <= ~(x[2320] & x[2322]);
     layer0_out[1448] <= x[5779] | x[5780];
     layer0_out[1449] <= x[5243];
     layer0_out[1450] <= x[5499];
     layer0_out[1451] <= x[6758];
     layer0_out[1452] <= 1'b1;
     layer0_out[1453] <= ~(x[3926] ^ x[3927]);
     layer0_out[1454] <= ~(x[6677] & x[6678]);
     layer0_out[1455] <= ~(x[4674] ^ x[4675]);
     layer0_out[1456] <= ~(x[582] & x[584]);
     layer0_out[1457] <= x[1400] ^ x[1402];
     layer0_out[1458] <= x[14];
     layer0_out[1459] <= ~x[4018];
     layer0_out[1460] <= ~(x[3940] ^ x[3941]);
     layer0_out[1461] <= x[2681];
     layer0_out[1462] <= x[8013];
     layer0_out[1463] <= ~(x[1927] & x[1929]);
     layer0_out[1464] <= x[2192];
     layer0_out[1465] <= ~(x[741] & x[742]);
     layer0_out[1466] <= 1'b1;
     layer0_out[1467] <= ~(x[4710] & x[4711]);
     layer0_out[1468] <= ~x[3101];
     layer0_out[1469] <= x[22] & x[24];
     layer0_out[1470] <= x[5972] & ~x[5971];
     layer0_out[1471] <= ~(x[4824] | x[4825]);
     layer0_out[1472] <= x[8924] | x[8925];
     layer0_out[1473] <= x[2362] & ~x[2364];
     layer0_out[1474] <= ~(x[5358] ^ x[5359]);
     layer0_out[1475] <= x[5870];
     layer0_out[1476] <= x[1236] ^ x[1237];
     layer0_out[1477] <= x[7123] | x[7124];
     layer0_out[1478] <= x[1284] & x[1286];
     layer0_out[1479] <= ~(x[2366] | x[2368]);
     layer0_out[1480] <= ~x[1294];
     layer0_out[1481] <= ~x[2029] | x[2031];
     layer0_out[1482] <= x[1721] & x[1723];
     layer0_out[1483] <= ~(x[835] & x[837]);
     layer0_out[1484] <= ~(x[6685] | x[6686]);
     layer0_out[1485] <= ~x[2269];
     layer0_out[1486] <= x[8120];
     layer0_out[1487] <= ~(x[3408] | x[3409]);
     layer0_out[1488] <= ~x[7010];
     layer0_out[1489] <= x[3712] ^ x[3713];
     layer0_out[1490] <= x[5059] | x[5060];
     layer0_out[1491] <= ~(x[885] | x[886]);
     layer0_out[1492] <= ~(x[372] | x[374]);
     layer0_out[1493] <= ~(x[8789] | x[8790]);
     layer0_out[1494] <= x[6262] & ~x[6263];
     layer0_out[1495] <= ~(x[1708] & x[1709]);
     layer0_out[1496] <= x[2165] & ~x[2163];
     layer0_out[1497] <= 1'b0;
     layer0_out[1498] <= ~(x[2431] ^ x[2432]);
     layer0_out[1499] <= ~(x[300] | x[302]);
     layer0_out[1500] <= ~x[804] | x[806];
     layer0_out[1501] <= x[2342];
     layer0_out[1502] <= x[191] & ~x[189];
     layer0_out[1503] <= x[8059] & x[8060];
     layer0_out[1504] <= x[3241] | x[3242];
     layer0_out[1505] <= ~(x[361] & x[363]);
     layer0_out[1506] <= x[2490];
     layer0_out[1507] <= ~x[325];
     layer0_out[1508] <= x[5228] & x[5229];
     layer0_out[1509] <= x[1780] & x[1781];
     layer0_out[1510] <= x[3278] ^ x[3279];
     layer0_out[1511] <= ~(x[5331] & x[5332]);
     layer0_out[1512] <= ~(x[944] | x[946]);
     layer0_out[1513] <= ~(x[8268] & x[8269]);
     layer0_out[1514] <= x[4603] & x[4604];
     layer0_out[1515] <= ~(x[991] & x[993]);
     layer0_out[1516] <= x[1868] ^ x[1870];
     layer0_out[1517] <= ~(x[7058] | x[7059]);
     layer0_out[1518] <= ~x[6264];
     layer0_out[1519] <= x[1181] & x[1183];
     layer0_out[1520] <= ~(x[4046] | x[4047]);
     layer0_out[1521] <= x[4054] ^ x[4055];
     layer0_out[1522] <= 1'b1;
     layer0_out[1523] <= ~(x[8080] ^ x[8081]);
     layer0_out[1524] <= ~x[1677] | x[1678];
     layer0_out[1525] <= x[8823];
     layer0_out[1526] <= x[8803] | x[8804];
     layer0_out[1527] <= x[6306] & x[6307];
     layer0_out[1528] <= ~x[7844];
     layer0_out[1529] <= ~x[8689] | x[8690];
     layer0_out[1530] <= ~x[3916];
     layer0_out[1531] <= ~(x[6811] | x[6812]);
     layer0_out[1532] <= ~x[2013];
     layer0_out[1533] <= x[2531] & x[2533];
     layer0_out[1534] <= ~(x[5869] ^ x[5870]);
     layer0_out[1535] <= ~(x[2379] | x[2381]);
     layer0_out[1536] <= ~x[6089];
     layer0_out[1537] <= x[517];
     layer0_out[1538] <= x[3801] & x[3802];
     layer0_out[1539] <= ~(x[7067] | x[7068]);
     layer0_out[1540] <= x[3388] & ~x[3389];
     layer0_out[1541] <= ~x[7446];
     layer0_out[1542] <= x[850] & x[851];
     layer0_out[1543] <= x[2755] ^ x[2757];
     layer0_out[1544] <= x[3845];
     layer0_out[1545] <= ~(x[2008] ^ x[2010]);
     layer0_out[1546] <= ~x[5516];
     layer0_out[1547] <= x[3296] | x[3297];
     layer0_out[1548] <= ~x[1831] | x[1829];
     layer0_out[1549] <= ~(x[1203] | x[1204]);
     layer0_out[1550] <= ~(x[2087] & x[2089]);
     layer0_out[1551] <= ~(x[3079] ^ x[3080]);
     layer0_out[1552] <= x[8313] | x[8314];
     layer0_out[1553] <= ~(x[4929] ^ x[4930]);
     layer0_out[1554] <= x[2577] & ~x[2579];
     layer0_out[1555] <= x[1833] & x[1835];
     layer0_out[1556] <= x[8210] ^ x[8211];
     layer0_out[1557] <= x[2989] ^ x[2990];
     layer0_out[1558] <= x[5378] & x[5379];
     layer0_out[1559] <= ~(x[5162] & x[5163]);
     layer0_out[1560] <= 1'b1;
     layer0_out[1561] <= x[4844];
     layer0_out[1562] <= x[4350];
     layer0_out[1563] <= ~(x[331] & x[333]);
     layer0_out[1564] <= x[2881] & x[2882];
     layer0_out[1565] <= x[715] & x[716];
     layer0_out[1566] <= x[5808] & x[5809];
     layer0_out[1567] <= ~(x[6281] ^ x[6282]);
     layer0_out[1568] <= x[5890] | x[5891];
     layer0_out[1569] <= ~(x[3027] & x[3028]);
     layer0_out[1570] <= x[41] | x[42];
     layer0_out[1571] <= ~(x[2371] & x[2372]);
     layer0_out[1572] <= x[7368];
     layer0_out[1573] <= x[902];
     layer0_out[1574] <= 1'b0;
     layer0_out[1575] <= ~(x[3468] ^ x[3469]);
     layer0_out[1576] <= ~x[2845];
     layer0_out[1577] <= x[7783] & x[7784];
     layer0_out[1578] <= ~x[1023];
     layer0_out[1579] <= ~(x[2183] | x[2184]);
     layer0_out[1580] <= x[2465] ^ x[2467];
     layer0_out[1581] <= ~(x[1878] ^ x[1879]);
     layer0_out[1582] <= x[1991];
     layer0_out[1583] <= ~(x[6136] | x[6137]);
     layer0_out[1584] <= ~(x[3156] & x[3157]);
     layer0_out[1585] <= ~x[7460] | x[7461];
     layer0_out[1586] <= x[774] | x[775];
     layer0_out[1587] <= 1'b1;
     layer0_out[1588] <= x[1760] | x[1762];
     layer0_out[1589] <= x[383];
     layer0_out[1590] <= ~(x[5462] & x[5463]);
     layer0_out[1591] <= ~(x[1712] | x[1713]);
     layer0_out[1592] <= 1'b1;
     layer0_out[1593] <= x[2497];
     layer0_out[1594] <= x[2343] | x[2345];
     layer0_out[1595] <= ~x[8038];
     layer0_out[1596] <= ~(x[8413] | x[8414]);
     layer0_out[1597] <= ~(x[5983] | x[5984]);
     layer0_out[1598] <= x[2129] | x[2130];
     layer0_out[1599] <= x[2224] & ~x[2225];
     layer0_out[1600] <= ~(x[5711] | x[5712]);
     layer0_out[1601] <= x[1434] ^ x[1436];
     layer0_out[1602] <= ~(x[1066] ^ x[1067]);
     layer0_out[1603] <= ~(x[3488] & x[3489]);
     layer0_out[1604] <= ~x[7757] | x[7758];
     layer0_out[1605] <= x[1964] & x[1965];
     layer0_out[1606] <= x[2541] ^ x[2542];
     layer0_out[1607] <= ~(x[4315] | x[4316]);
     layer0_out[1608] <= x[6739] ^ x[6740];
     layer0_out[1609] <= ~(x[687] & x[689]);
     layer0_out[1610] <= x[2967];
     layer0_out[1611] <= x[8506] | x[8507];
     layer0_out[1612] <= ~x[686] | x[687];
     layer0_out[1613] <= 1'b0;
     layer0_out[1614] <= x[4339] | x[4340];
     layer0_out[1615] <= x[9039];
     layer0_out[1616] <= ~(x[9100] | x[9101]);
     layer0_out[1617] <= x[1106];
     layer0_out[1618] <= ~x[2610];
     layer0_out[1619] <= ~x[5821] | x[5822];
     layer0_out[1620] <= 1'b1;
     layer0_out[1621] <= 1'b1;
     layer0_out[1622] <= ~(x[8068] | x[8069]);
     layer0_out[1623] <= x[336] & x[338];
     layer0_out[1624] <= ~(x[5258] & x[5259]);
     layer0_out[1625] <= ~(x[3164] ^ x[3165]);
     layer0_out[1626] <= ~x[371] | x[372];
     layer0_out[1627] <= x[4732] & x[4733];
     layer0_out[1628] <= ~(x[427] & x[429]);
     layer0_out[1629] <= ~(x[5529] & x[5530]);
     layer0_out[1630] <= ~(x[1555] | x[1556]);
     layer0_out[1631] <= x[2203] & x[2205];
     layer0_out[1632] <= 1'b1;
     layer0_out[1633] <= 1'b1;
     layer0_out[1634] <= ~(x[8348] & x[8349]);
     layer0_out[1635] <= ~(x[5060] ^ x[5061]);
     layer0_out[1636] <= x[3031] ^ x[3032];
     layer0_out[1637] <= ~(x[7872] ^ x[7873]);
     layer0_out[1638] <= 1'b0;
     layer0_out[1639] <= ~(x[4909] | x[4910]);
     layer0_out[1640] <= x[2361] ^ x[2362];
     layer0_out[1641] <= ~(x[961] & x[963]);
     layer0_out[1642] <= x[3657] ^ x[3658];
     layer0_out[1643] <= x[1941];
     layer0_out[1644] <= x[2209] & x[2211];
     layer0_out[1645] <= x[289] & ~x[288];
     layer0_out[1646] <= x[2193] & x[2195];
     layer0_out[1647] <= ~(x[8861] & x[8862]);
     layer0_out[1648] <= ~x[1281];
     layer0_out[1649] <= ~(x[7749] ^ x[7750]);
     layer0_out[1650] <= ~x[381] | x[382];
     layer0_out[1651] <= ~(x[1033] & x[1034]);
     layer0_out[1652] <= ~(x[4198] & x[4199]);
     layer0_out[1653] <= ~(x[2565] & x[2567]);
     layer0_out[1654] <= ~(x[289] ^ x[291]);
     layer0_out[1655] <= x[1841] ^ x[1843];
     layer0_out[1656] <= x[3930];
     layer0_out[1657] <= x[1752] & x[1754];
     layer0_out[1658] <= 1'b1;
     layer0_out[1659] <= x[4356] & x[4357];
     layer0_out[1660] <= ~(x[652] & x[654]);
     layer0_out[1661] <= x[1501] ^ x[1503];
     layer0_out[1662] <= ~(x[1910] | x[1912]);
     layer0_out[1663] <= ~x[956] | x[954];
     layer0_out[1664] <= x[1497];
     layer0_out[1665] <= x[2835];
     layer0_out[1666] <= x[2234] & x[2236];
     layer0_out[1667] <= ~x[6505] | x[6504];
     layer0_out[1668] <= ~(x[458] & x[460]);
     layer0_out[1669] <= x[5435] | x[5436];
     layer0_out[1670] <= ~(x[6340] | x[6341]);
     layer0_out[1671] <= ~(x[1046] | x[1047]);
     layer0_out[1672] <= ~x[3514] | x[3515];
     layer0_out[1673] <= 1'b1;
     layer0_out[1674] <= x[538] & x[540];
     layer0_out[1675] <= ~(x[3432] | x[3433]);
     layer0_out[1676] <= x[6984] & ~x[6985];
     layer0_out[1677] <= 1'b0;
     layer0_out[1678] <= x[3168] & x[3169];
     layer0_out[1679] <= x[2499];
     layer0_out[1680] <= ~(x[2700] ^ x[2701]);
     layer0_out[1681] <= ~x[6986];
     layer0_out[1682] <= ~(x[6557] | x[6558]);
     layer0_out[1683] <= x[1253] & ~x[1255];
     layer0_out[1684] <= ~x[244];
     layer0_out[1685] <= 1'b1;
     layer0_out[1686] <= ~(x[575] & x[576]);
     layer0_out[1687] <= x[2261] & x[2262];
     layer0_out[1688] <= ~(x[6563] ^ x[6564]);
     layer0_out[1689] <= ~(x[1734] | x[1736]);
     layer0_out[1690] <= ~(x[5344] & x[5345]);
     layer0_out[1691] <= x[2355] & x[2356];
     layer0_out[1692] <= x[6602];
     layer0_out[1693] <= x[5565] | x[5566];
     layer0_out[1694] <= x[1825] ^ x[1826];
     layer0_out[1695] <= ~(x[14] & x[16]);
     layer0_out[1696] <= x[5381] & x[5382];
     layer0_out[1697] <= x[3870] ^ x[3871];
     layer0_out[1698] <= x[1676] & x[1677];
     layer0_out[1699] <= ~x[1242];
     layer0_out[1700] <= x[8292] ^ x[8293];
     layer0_out[1701] <= ~(x[5902] & x[5903]);
     layer0_out[1702] <= ~(x[7014] ^ x[7015]);
     layer0_out[1703] <= ~x[8802];
     layer0_out[1704] <= x[8473];
     layer0_out[1705] <= x[4658];
     layer0_out[1706] <= ~x[2085];
     layer0_out[1707] <= ~(x[8769] | x[8770]);
     layer0_out[1708] <= 1'b0;
     layer0_out[1709] <= ~(x[1835] & x[1837]);
     layer0_out[1710] <= x[2222];
     layer0_out[1711] <= x[8735] & x[8736];
     layer0_out[1712] <= ~(x[3887] ^ x[3888]);
     layer0_out[1713] <= x[4021] | x[4022];
     layer0_out[1714] <= 1'b1;
     layer0_out[1715] <= x[5835] & x[5836];
     layer0_out[1716] <= x[8785] | x[8786];
     layer0_out[1717] <= ~(x[1048] & x[1050]);
     layer0_out[1718] <= ~(x[1373] & x[1374]);
     layer0_out[1719] <= ~(x[2768] & x[2769]);
     layer0_out[1720] <= x[6716];
     layer0_out[1721] <= ~(x[6172] | x[6173]);
     layer0_out[1722] <= x[987];
     layer0_out[1723] <= x[389] & x[391];
     layer0_out[1724] <= ~x[495];
     layer0_out[1725] <= x[6392] | x[6393];
     layer0_out[1726] <= x[9126] ^ x[9127];
     layer0_out[1727] <= ~(x[1906] & x[1907]);
     layer0_out[1728] <= x[7193];
     layer0_out[1729] <= ~x[2596];
     layer0_out[1730] <= ~(x[265] & x[267]);
     layer0_out[1731] <= x[3324] ^ x[3325];
     layer0_out[1732] <= x[8] & ~x[6];
     layer0_out[1733] <= x[514] ^ x[515];
     layer0_out[1734] <= x[685] & x[686];
     layer0_out[1735] <= x[5176] & ~x[5175];
     layer0_out[1736] <= x[4135] ^ x[4136];
     layer0_out[1737] <= x[5427] & x[5428];
     layer0_out[1738] <= ~(x[3309] & x[3310]);
     layer0_out[1739] <= x[2984] | x[2985];
     layer0_out[1740] <= ~(x[1531] ^ x[1532]);
     layer0_out[1741] <= ~(x[4319] & x[4320]);
     layer0_out[1742] <= x[3388] & ~x[3387];
     layer0_out[1743] <= x[1086] ^ x[1088];
     layer0_out[1744] <= ~x[3751] | x[3752];
     layer0_out[1745] <= x[5648];
     layer0_out[1746] <= ~x[1732] | x[1730];
     layer0_out[1747] <= ~(x[174] ^ x[175]);
     layer0_out[1748] <= x[3585] ^ x[3586];
     layer0_out[1749] <= x[546] & ~x[548];
     layer0_out[1750] <= x[313] & x[314];
     layer0_out[1751] <= ~(x[1567] ^ x[1568]);
     layer0_out[1752] <= x[710] | x[711];
     layer0_out[1753] <= x[3096] | x[3097];
     layer0_out[1754] <= 1'b0;
     layer0_out[1755] <= ~(x[1585] & x[1586]);
     layer0_out[1756] <= x[1403] | x[1405];
     layer0_out[1757] <= ~(x[334] & x[335]);
     layer0_out[1758] <= 1'b0;
     layer0_out[1759] <= x[1486] & x[1488];
     layer0_out[1760] <= 1'b1;
     layer0_out[1761] <= x[1971] & x[1973];
     layer0_out[1762] <= x[844] & x[846];
     layer0_out[1763] <= x[4611] & x[4612];
     layer0_out[1764] <= ~(x[907] | x[909]);
     layer0_out[1765] <= x[1756] & ~x[1758];
     layer0_out[1766] <= x[3108] | x[3109];
     layer0_out[1767] <= x[8265] & ~x[8264];
     layer0_out[1768] <= ~(x[816] ^ x[817]);
     layer0_out[1769] <= ~x[2139] | x[2137];
     layer0_out[1770] <= ~(x[7911] & x[7912]);
     layer0_out[1771] <= x[1764] | x[1765];
     layer0_out[1772] <= ~x[7304];
     layer0_out[1773] <= x[4400] ^ x[4401];
     layer0_out[1774] <= ~(x[4955] | x[4956]);
     layer0_out[1775] <= ~(x[2702] ^ x[2704]);
     layer0_out[1776] <= 1'b0;
     layer0_out[1777] <= ~(x[1383] | x[1385]);
     layer0_out[1778] <= ~(x[1424] & x[1425]);
     layer0_out[1779] <= x[562] & ~x[564];
     layer0_out[1780] <= x[3019] & x[3020];
     layer0_out[1781] <= x[5361] & x[5362];
     layer0_out[1782] <= x[1596] ^ x[1597];
     layer0_out[1783] <= x[7358];
     layer0_out[1784] <= x[401] & x[402];
     layer0_out[1785] <= ~x[8786];
     layer0_out[1786] <= x[6341] & x[6342];
     layer0_out[1787] <= ~x[6150];
     layer0_out[1788] <= x[1387] & x[1388];
     layer0_out[1789] <= ~x[7427];
     layer0_out[1790] <= ~x[461] | x[460];
     layer0_out[1791] <= x[5729] & x[5730];
     layer0_out[1792] <= ~(x[2542] & x[2544]);
     layer0_out[1793] <= x[1005];
     layer0_out[1794] <= ~(x[2538] | x[2539]);
     layer0_out[1795] <= ~(x[6628] & x[6629]);
     layer0_out[1796] <= x[3218];
     layer0_out[1797] <= 1'b0;
     layer0_out[1798] <= x[7887];
     layer0_out[1799] <= ~(x[728] & x[729]);
     layer0_out[1800] <= ~(x[1344] & x[1345]);
     layer0_out[1801] <= ~(x[2081] | x[2083]);
     layer0_out[1802] <= ~(x[799] & x[801]);
     layer0_out[1803] <= 1'b1;
     layer0_out[1804] <= ~(x[1765] & x[1767]);
     layer0_out[1805] <= ~(x[1880] ^ x[1881]);
     layer0_out[1806] <= x[5521] | x[5522];
     layer0_out[1807] <= ~x[1229];
     layer0_out[1808] <= x[7061] | x[7062];
     layer0_out[1809] <= ~x[1137];
     layer0_out[1810] <= x[155] | x[156];
     layer0_out[1811] <= ~(x[8644] | x[8645]);
     layer0_out[1812] <= ~(x[771] & x[772]);
     layer0_out[1813] <= ~(x[2280] & x[2282]);
     layer0_out[1814] <= ~x[106];
     layer0_out[1815] <= x[6503] | x[6504];
     layer0_out[1816] <= x[831];
     layer0_out[1817] <= ~x[3569];
     layer0_out[1818] <= ~x[2721];
     layer0_out[1819] <= x[3005] & x[3006];
     layer0_out[1820] <= 1'b1;
     layer0_out[1821] <= ~x[4423] | x[4422];
     layer0_out[1822] <= x[4726] & x[4727];
     layer0_out[1823] <= x[462] & x[464];
     layer0_out[1824] <= x[3496];
     layer0_out[1825] <= x[86] & ~x[85];
     layer0_out[1826] <= x[5118] ^ x[5119];
     layer0_out[1827] <= x[2479];
     layer0_out[1828] <= ~(x[477] | x[478]);
     layer0_out[1829] <= x[6058] & x[6059];
     layer0_out[1830] <= 1'b0;
     layer0_out[1831] <= x[3500];
     layer0_out[1832] <= ~x[2508];
     layer0_out[1833] <= 1'b0;
     layer0_out[1834] <= 1'b1;
     layer0_out[1835] <= ~(x[6387] | x[6388]);
     layer0_out[1836] <= x[9197] & ~x[9196];
     layer0_out[1837] <= ~(x[8579] | x[8580]);
     layer0_out[1838] <= x[3735] | x[3736];
     layer0_out[1839] <= x[3137];
     layer0_out[1840] <= x[3138] | x[3139];
     layer0_out[1841] <= x[7070] & x[7071];
     layer0_out[1842] <= ~x[2378] | x[2379];
     layer0_out[1843] <= x[2292] & ~x[2291];
     layer0_out[1844] <= ~(x[3952] | x[3953]);
     layer0_out[1845] <= x[4302] | x[4303];
     layer0_out[1846] <= x[339] & x[341];
     layer0_out[1847] <= 1'b1;
     layer0_out[1848] <= x[7801];
     layer0_out[1849] <= ~(x[7526] | x[7527]);
     layer0_out[1850] <= x[5804] ^ x[5805];
     layer0_out[1851] <= ~(x[8427] | x[8428]);
     layer0_out[1852] <= ~x[2203] | x[2204];
     layer0_out[1853] <= ~(x[2479] & x[2480]);
     layer0_out[1854] <= x[2866];
     layer0_out[1855] <= x[8173] ^ x[8174];
     layer0_out[1856] <= x[3663] & x[3664];
     layer0_out[1857] <= ~(x[2558] ^ x[2559]);
     layer0_out[1858] <= ~x[6964];
     layer0_out[1859] <= x[5538] & x[5539];
     layer0_out[1860] <= ~(x[7475] ^ x[7476]);
     layer0_out[1861] <= x[6855] ^ x[6856];
     layer0_out[1862] <= x[8820] | x[8821];
     layer0_out[1863] <= x[5774] & x[5775];
     layer0_out[1864] <= ~x[209];
     layer0_out[1865] <= ~x[428];
     layer0_out[1866] <= ~(x[791] | x[793]);
     layer0_out[1867] <= ~x[7396] | x[7397];
     layer0_out[1868] <= ~(x[5640] & x[5641]);
     layer0_out[1869] <= x[1995];
     layer0_out[1870] <= ~x[4457] | x[4456];
     layer0_out[1871] <= ~(x[1796] ^ x[1798]);
     layer0_out[1872] <= ~x[664] | x[665];
     layer0_out[1873] <= ~x[1051] | x[1049];
     layer0_out[1874] <= x[8676];
     layer0_out[1875] <= ~x[1789];
     layer0_out[1876] <= ~(x[7915] & x[7916]);
     layer0_out[1877] <= x[7893];
     layer0_out[1878] <= ~(x[5673] | x[5674]);
     layer0_out[1879] <= x[2063] ^ x[2064];
     layer0_out[1880] <= x[382] ^ x[384];
     layer0_out[1881] <= ~x[8994];
     layer0_out[1882] <= ~(x[5571] & x[5572]);
     layer0_out[1883] <= ~(x[6718] ^ x[6719]);
     layer0_out[1884] <= ~(x[1629] & x[1631]);
     layer0_out[1885] <= ~(x[1626] & x[1628]);
     layer0_out[1886] <= ~(x[2184] ^ x[2185]);
     layer0_out[1887] <= ~(x[2701] ^ x[2702]);
     layer0_out[1888] <= x[5229] & x[5230];
     layer0_out[1889] <= 1'b1;
     layer0_out[1890] <= ~(x[7039] ^ x[7040]);
     layer0_out[1891] <= x[3742];
     layer0_out[1892] <= x[2073] & x[2075];
     layer0_out[1893] <= x[1876];
     layer0_out[1894] <= ~(x[2657] ^ x[2659]);
     layer0_out[1895] <= x[2830] ^ x[2831];
     layer0_out[1896] <= ~(x[1103] & x[1105]);
     layer0_out[1897] <= x[4248];
     layer0_out[1898] <= ~(x[7621] | x[7622]);
     layer0_out[1899] <= x[6520];
     layer0_out[1900] <= ~(x[1767] | x[1768]);
     layer0_out[1901] <= x[5084] | x[5085];
     layer0_out[1902] <= x[2207] & x[2209];
     layer0_out[1903] <= ~(x[1924] & x[1926]);
     layer0_out[1904] <= ~(x[8109] & x[8110]);
     layer0_out[1905] <= x[4156] & x[4157];
     layer0_out[1906] <= x[1460] & x[1461];
     layer0_out[1907] <= 1'b0;
     layer0_out[1908] <= ~(x[2342] & x[2344]);
     layer0_out[1909] <= x[2249] & x[2250];
     layer0_out[1910] <= x[5107] ^ x[5108];
     layer0_out[1911] <= x[1684] & x[1685];
     layer0_out[1912] <= x[660] & x[662];
     layer0_out[1913] <= ~(x[3951] | x[3952]);
     layer0_out[1914] <= x[1459];
     layer0_out[1915] <= x[698] | x[700];
     layer0_out[1916] <= x[4567] & x[4568];
     layer0_out[1917] <= ~(x[116] ^ x[118]);
     layer0_out[1918] <= 1'b1;
     layer0_out[1919] <= x[5959] | x[5960];
     layer0_out[1920] <= ~(x[743] & x[745]);
     layer0_out[1921] <= 1'b0;
     layer0_out[1922] <= ~x[3567];
     layer0_out[1923] <= x[2090] & x[2091];
     layer0_out[1924] <= ~(x[6390] | x[6391]);
     layer0_out[1925] <= 1'b1;
     layer0_out[1926] <= ~(x[2681] & x[2682]);
     layer0_out[1927] <= x[4377] & x[4378];
     layer0_out[1928] <= 1'b1;
     layer0_out[1929] <= ~x[8489];
     layer0_out[1930] <= 1'b1;
     layer0_out[1931] <= x[757] ^ x[758];
     layer0_out[1932] <= x[3343];
     layer0_out[1933] <= x[1166] & ~x[1167];
     layer0_out[1934] <= ~(x[8395] & x[8396]);
     layer0_out[1935] <= ~(x[5809] & x[5810]);
     layer0_out[1936] <= ~(x[116] ^ x[117]);
     layer0_out[1937] <= ~(x[6178] | x[6179]);
     layer0_out[1938] <= x[6176] | x[6177];
     layer0_out[1939] <= x[1030] & ~x[1028];
     layer0_out[1940] <= ~(x[5075] ^ x[5076]);
     layer0_out[1941] <= ~(x[6158] | x[6159]);
     layer0_out[1942] <= x[5823] & x[5824];
     layer0_out[1943] <= ~(x[6997] | x[6998]);
     layer0_out[1944] <= ~(x[1158] & x[1159]);
     layer0_out[1945] <= ~x[6461];
     layer0_out[1946] <= ~(x[5985] | x[5986]);
     layer0_out[1947] <= x[8237];
     layer0_out[1948] <= x[4962] ^ x[4963];
     layer0_out[1949] <= x[7860] ^ x[7861];
     layer0_out[1950] <= x[1874] | x[1875];
     layer0_out[1951] <= ~(x[8561] | x[8562]);
     layer0_out[1952] <= x[316] | x[318];
     layer0_out[1953] <= x[7274] & x[7275];
     layer0_out[1954] <= ~(x[1556] ^ x[1558]);
     layer0_out[1955] <= x[1882] | x[1884];
     layer0_out[1956] <= ~(x[4430] & x[4431]);
     layer0_out[1957] <= x[5776];
     layer0_out[1958] <= x[3348];
     layer0_out[1959] <= ~(x[6166] | x[6167]);
     layer0_out[1960] <= x[1848] | x[1850];
     layer0_out[1961] <= x[7] & x[9];
     layer0_out[1962] <= ~(x[1214] & x[1215]);
     layer0_out[1963] <= x[1631];
     layer0_out[1964] <= x[5127] & x[5128];
     layer0_out[1965] <= x[2380] | x[2382];
     layer0_out[1966] <= ~(x[5074] ^ x[5075]);
     layer0_out[1967] <= ~(x[8913] | x[8914]);
     layer0_out[1968] <= ~x[1211];
     layer0_out[1969] <= ~x[7065] | x[7064];
     layer0_out[1970] <= ~(x[8984] & x[8985]);
     layer0_out[1971] <= ~x[2247];
     layer0_out[1972] <= x[138];
     layer0_out[1973] <= ~(x[7752] ^ x[7753]);
     layer0_out[1974] <= x[2710] & x[2711];
     layer0_out[1975] <= x[8495] | x[8496];
     layer0_out[1976] <= ~(x[1032] | x[1034]);
     layer0_out[1977] <= ~(x[2065] | x[2066]);
     layer0_out[1978] <= ~(x[187] | x[188]);
     layer0_out[1979] <= ~x[69];
     layer0_out[1980] <= ~x[2804];
     layer0_out[1981] <= ~x[2294] | x[2295];
     layer0_out[1982] <= x[4838] | x[4839];
     layer0_out[1983] <= ~(x[7025] ^ x[7026]);
     layer0_out[1984] <= x[1695] & x[1697];
     layer0_out[1985] <= x[4548] & x[4549];
     layer0_out[1986] <= x[3400] ^ x[3401];
     layer0_out[1987] <= ~(x[6327] ^ x[6328]);
     layer0_out[1988] <= x[2541] & x[2543];
     layer0_out[1989] <= x[2988] & x[2989];
     layer0_out[1990] <= ~(x[3938] | x[3939]);
     layer0_out[1991] <= x[1045] & ~x[1046];
     layer0_out[1992] <= x[730] & x[732];
     layer0_out[1993] <= x[7835] ^ x[7836];
     layer0_out[1994] <= x[2562] & x[2563];
     layer0_out[1995] <= x[348];
     layer0_out[1996] <= ~(x[2978] | x[2979]);
     layer0_out[1997] <= ~(x[2165] & x[2166]);
     layer0_out[1998] <= x[37];
     layer0_out[1999] <= 1'b1;
     layer0_out[2000] <= x[8073] & x[8074];
     layer0_out[2001] <= ~x[2279] | x[2281];
     layer0_out[2002] <= ~(x[5724] ^ x[5725]);
     layer0_out[2003] <= x[1809];
     layer0_out[2004] <= ~(x[2249] & x[2251]);
     layer0_out[2005] <= ~(x[981] | x[982]);
     layer0_out[2006] <= x[4012] & x[4013];
     layer0_out[2007] <= ~(x[2550] & x[2552]);
     layer0_out[2008] <= x[1054];
     layer0_out[2009] <= ~x[1696] | x[1694];
     layer0_out[2010] <= x[7532] | x[7533];
     layer0_out[2011] <= ~(x[1069] & x[1071]);
     layer0_out[2012] <= x[1948];
     layer0_out[2013] <= x[7240];
     layer0_out[2014] <= x[7485];
     layer0_out[2015] <= x[2638] & ~x[2640];
     layer0_out[2016] <= ~(x[9021] & x[9022]);
     layer0_out[2017] <= ~(x[3385] & x[3386]);
     layer0_out[2018] <= ~(x[2412] & x[2413]);
     layer0_out[2019] <= ~(x[6748] | x[6749]);
     layer0_out[2020] <= ~(x[7454] | x[7455]);
     layer0_out[2021] <= ~(x[871] & x[872]);
     layer0_out[2022] <= x[9015] & x[9016];
     layer0_out[2023] <= x[6202] | x[6203];
     layer0_out[2024] <= x[2615] & x[2617];
     layer0_out[2025] <= x[2217];
     layer0_out[2026] <= 1'b0;
     layer0_out[2027] <= ~(x[667] & x[668]);
     layer0_out[2028] <= x[1168] & x[1170];
     layer0_out[2029] <= x[6546] & x[6547];
     layer0_out[2030] <= x[8215] ^ x[8216];
     layer0_out[2031] <= x[5554] | x[5555];
     layer0_out[2032] <= ~(x[813] ^ x[815]);
     layer0_out[2033] <= x[7224];
     layer0_out[2034] <= ~x[8450];
     layer0_out[2035] <= x[230] & x[232];
     layer0_out[2036] <= ~(x[2393] & x[2394]);
     layer0_out[2037] <= ~x[6065] | x[6064];
     layer0_out[2038] <= x[2506] & x[2507];
     layer0_out[2039] <= ~x[8335];
     layer0_out[2040] <= ~(x[8736] & x[8737]);
     layer0_out[2041] <= ~(x[5645] & x[5646]);
     layer0_out[2042] <= x[2005] ^ x[2007];
     layer0_out[2043] <= x[1135];
     layer0_out[2044] <= ~(x[3613] & x[3614]);
     layer0_out[2045] <= ~x[7788] | x[7787];
     layer0_out[2046] <= ~(x[888] | x[889]);
     layer0_out[2047] <= x[7189] | x[7190];
     layer0_out[2048] <= x[1838] ^ x[1840];
     layer0_out[2049] <= x[6276] | x[6277];
     layer0_out[2050] <= x[5012];
     layer0_out[2051] <= x[7941] ^ x[7942];
     layer0_out[2052] <= x[1864] | x[1866];
     layer0_out[2053] <= x[5227] & x[5228];
     layer0_out[2054] <= x[7712] & ~x[7711];
     layer0_out[2055] <= ~(x[4020] | x[4021]);
     layer0_out[2056] <= ~(x[454] ^ x[455]);
     layer0_out[2057] <= x[508] | x[509];
     layer0_out[2058] <= x[745] | x[746];
     layer0_out[2059] <= 1'b0;
     layer0_out[2060] <= ~(x[1996] | x[1998]);
     layer0_out[2061] <= ~(x[7152] & x[7153]);
     layer0_out[2062] <= x[7414] ^ x[7415];
     layer0_out[2063] <= ~(x[461] & x[463]);
     layer0_out[2064] <= ~(x[7809] | x[7810]);
     layer0_out[2065] <= ~(x[4030] & x[4031]);
     layer0_out[2066] <= ~(x[4599] ^ x[4600]);
     layer0_out[2067] <= x[1450] | x[1452];
     layer0_out[2068] <= ~x[1526];
     layer0_out[2069] <= ~x[288];
     layer0_out[2070] <= 1'b1;
     layer0_out[2071] <= ~(x[1393] ^ x[1394]);
     layer0_out[2072] <= x[3284];
     layer0_out[2073] <= x[776] & x[777];
     layer0_out[2074] <= x[1414];
     layer0_out[2075] <= ~(x[8311] & x[8312]);
     layer0_out[2076] <= x[2202];
     layer0_out[2077] <= x[7009];
     layer0_out[2078] <= ~(x[2912] & x[2913]);
     layer0_out[2079] <= ~(x[5511] & x[5512]);
     layer0_out[2080] <= x[1444] | x[1445];
     layer0_out[2081] <= ~x[3];
     layer0_out[2082] <= ~(x[1542] & x[1544]);
     layer0_out[2083] <= ~(x[7162] ^ x[7163]);
     layer0_out[2084] <= ~(x[2220] & x[2221]);
     layer0_out[2085] <= 1'b0;
     layer0_out[2086] <= x[510] & ~x[511];
     layer0_out[2087] <= x[1615] & x[1617];
     layer0_out[2088] <= ~(x[8315] & x[8316]);
     layer0_out[2089] <= ~(x[2730] ^ x[2731]);
     layer0_out[2090] <= x[1932] ^ x[1934];
     layer0_out[2091] <= ~(x[4172] ^ x[4173]);
     layer0_out[2092] <= x[3910] ^ x[3911];
     layer0_out[2093] <= ~x[5853];
     layer0_out[2094] <= ~(x[4489] | x[4490]);
     layer0_out[2095] <= ~(x[2685] & x[2687]);
     layer0_out[2096] <= x[6060] & x[6061];
     layer0_out[2097] <= ~x[7588] | x[7589];
     layer0_out[2098] <= x[5998] & x[5999];
     layer0_out[2099] <= ~(x[3111] & x[3112]);
     layer0_out[2100] <= ~(x[4828] & x[4829]);
     layer0_out[2101] <= x[559] & x[560];
     layer0_out[2102] <= x[7] & ~x[5];
     layer0_out[2103] <= ~(x[3996] | x[3997]);
     layer0_out[2104] <= x[4738] & x[4739];
     layer0_out[2105] <= ~(x[2132] & x[2134]);
     layer0_out[2106] <= x[6822] & x[6823];
     layer0_out[2107] <= x[4916] & x[4917];
     layer0_out[2108] <= x[1223] ^ x[1225];
     layer0_out[2109] <= ~(x[1713] ^ x[1715]);
     layer0_out[2110] <= x[2694];
     layer0_out[2111] <= x[577] & ~x[575];
     layer0_out[2112] <= 1'b0;
     layer0_out[2113] <= ~x[5987];
     layer0_out[2114] <= 1'b0;
     layer0_out[2115] <= ~(x[325] ^ x[327]);
     layer0_out[2116] <= x[572] & ~x[571];
     layer0_out[2117] <= ~(x[2365] & x[2366]);
     layer0_out[2118] <= ~(x[2406] & x[2407]);
     layer0_out[2119] <= ~(x[2841] ^ x[2842]);
     layer0_out[2120] <= x[5853] | x[5854];
     layer0_out[2121] <= ~(x[2457] & x[2459]);
     layer0_out[2122] <= x[2387] & x[2389];
     layer0_out[2123] <= ~(x[304] & x[305]);
     layer0_out[2124] <= x[2265] & x[2267];
     layer0_out[2125] <= x[1473] & ~x[1471];
     layer0_out[2126] <= ~x[2336] | x[2334];
     layer0_out[2127] <= x[2147] & x[2148];
     layer0_out[2128] <= ~(x[6313] | x[6314]);
     layer0_out[2129] <= ~(x[9012] | x[9013]);
     layer0_out[2130] <= ~(x[2743] & x[2744]);
     layer0_out[2131] <= x[4353] & x[4354];
     layer0_out[2132] <= x[7289];
     layer0_out[2133] <= x[2779] ^ x[2781];
     layer0_out[2134] <= ~(x[2447] & x[2449]);
     layer0_out[2135] <= x[1598] & x[1599];
     layer0_out[2136] <= ~(x[1271] & x[1272]);
     layer0_out[2137] <= ~(x[196] & x[197]);
     layer0_out[2138] <= ~x[4666] | x[4665];
     layer0_out[2139] <= ~x[7302];
     layer0_out[2140] <= ~x[956];
     layer0_out[2141] <= x[1343] | x[1345];
     layer0_out[2142] <= ~(x[3800] & x[3801]);
     layer0_out[2143] <= ~(x[803] ^ x[804]);
     layer0_out[2144] <= x[2594] & x[2596];
     layer0_out[2145] <= ~(x[3246] & x[3247]);
     layer0_out[2146] <= ~(x[2536] & x[2538]);
     layer0_out[2147] <= x[27] & ~x[26];
     layer0_out[2148] <= ~(x[917] & x[919]);
     layer0_out[2149] <= x[4226] & x[4227];
     layer0_out[2150] <= x[5776] | x[5777];
     layer0_out[2151] <= ~x[2416];
     layer0_out[2152] <= ~(x[2325] & x[2326]);
     layer0_out[2153] <= x[3617] ^ x[3618];
     layer0_out[2154] <= ~(x[1744] & x[1745]);
     layer0_out[2155] <= 1'b0;
     layer0_out[2156] <= ~(x[5420] & x[5421]);
     layer0_out[2157] <= ~(x[7762] & x[7763]);
     layer0_out[2158] <= ~x[5137];
     layer0_out[2159] <= ~x[5769];
     layer0_out[2160] <= ~(x[5791] | x[5792]);
     layer0_out[2161] <= x[6370] | x[6371];
     layer0_out[2162] <= ~(x[4618] & x[4619]);
     layer0_out[2163] <= x[1463] & x[1465];
     layer0_out[2164] <= ~(x[9047] ^ x[9048]);
     layer0_out[2165] <= 1'b0;
     layer0_out[2166] <= ~x[6995];
     layer0_out[2167] <= x[2339] & ~x[2341];
     layer0_out[2168] <= ~(x[6596] | x[6597]);
     layer0_out[2169] <= ~(x[4391] & x[4392]);
     layer0_out[2170] <= 1'b1;
     layer0_out[2171] <= x[3811] | x[3812];
     layer0_out[2172] <= x[379] & ~x[378];
     layer0_out[2173] <= ~x[5476];
     layer0_out[2174] <= x[5139] & x[5140];
     layer0_out[2175] <= ~(x[8979] | x[8980]);
     layer0_out[2176] <= ~(x[6774] & x[6775]);
     layer0_out[2177] <= ~(x[4739] & x[4740]);
     layer0_out[2178] <= 1'b0;
     layer0_out[2179] <= ~(x[8457] & x[8458]);
     layer0_out[2180] <= x[4809] | x[4810];
     layer0_out[2181] <= x[841];
     layer0_out[2182] <= x[7259] & ~x[7260];
     layer0_out[2183] <= ~(x[8155] | x[8156]);
     layer0_out[2184] <= ~(x[2566] & x[2567]);
     layer0_out[2185] <= ~(x[6980] | x[6981]);
     layer0_out[2186] <= 1'b1;
     layer0_out[2187] <= ~x[2311];
     layer0_out[2188] <= x[8584] & ~x[8583];
     layer0_out[2189] <= x[26] ^ x[28];
     layer0_out[2190] <= x[4281] & ~x[4282];
     layer0_out[2191] <= ~(x[8969] | x[8970]);
     layer0_out[2192] <= ~(x[4090] ^ x[4091]);
     layer0_out[2193] <= ~(x[7327] | x[7328]);
     layer0_out[2194] <= x[1336] ^ x[1338];
     layer0_out[2195] <= ~(x[1783] & x[1785]);
     layer0_out[2196] <= ~x[870];
     layer0_out[2197] <= x[1765] & x[1766];
     layer0_out[2198] <= x[988];
     layer0_out[2199] <= x[1549] & x[1550];
     layer0_out[2200] <= x[4959];
     layer0_out[2201] <= ~(x[5630] | x[5631]);
     layer0_out[2202] <= x[7505] | x[7506];
     layer0_out[2203] <= x[577] | x[578];
     layer0_out[2204] <= x[3812] & x[3813];
     layer0_out[2205] <= ~(x[794] & x[795]);
     layer0_out[2206] <= x[504] | x[506];
     layer0_out[2207] <= ~(x[3516] | x[3517]);
     layer0_out[2208] <= x[5574];
     layer0_out[2209] <= ~(x[576] ^ x[578]);
     layer0_out[2210] <= 1'b1;
     layer0_out[2211] <= ~(x[1769] & x[1770]);
     layer0_out[2212] <= ~(x[2901] & x[2902]);
     layer0_out[2213] <= ~(x[6126] & x[6127]);
     layer0_out[2214] <= ~x[1952];
     layer0_out[2215] <= x[1872] & x[1874];
     layer0_out[2216] <= ~x[2347] | x[2345];
     layer0_out[2217] <= ~(x[874] & x[876]);
     layer0_out[2218] <= ~x[4551] | x[4552];
     layer0_out[2219] <= x[2752] | x[2753];
     layer0_out[2220] <= x[6618] | x[6619];
     layer0_out[2221] <= x[8435] | x[8436];
     layer0_out[2222] <= x[599];
     layer0_out[2223] <= ~x[6466];
     layer0_out[2224] <= x[2144] & x[2145];
     layer0_out[2225] <= ~(x[1056] | x[1058]);
     layer0_out[2226] <= ~(x[607] ^ x[608]);
     layer0_out[2227] <= ~(x[8625] | x[8626]);
     layer0_out[2228] <= x[6863] | x[6864];
     layer0_out[2229] <= x[761] ^ x[762];
     layer0_out[2230] <= ~(x[6044] ^ x[6045]);
     layer0_out[2231] <= ~x[7594] | x[7595];
     layer0_out[2232] <= ~(x[4763] & x[4764]);
     layer0_out[2233] <= x[818] & x[820];
     layer0_out[2234] <= x[7759] | x[7760];
     layer0_out[2235] <= ~x[4925] | x[4924];
     layer0_out[2236] <= x[6584] | x[6585];
     layer0_out[2237] <= ~x[7212];
     layer0_out[2238] <= x[236] & x[238];
     layer0_out[2239] <= ~(x[6371] & x[6372]);
     layer0_out[2240] <= ~(x[6346] & x[6347]);
     layer0_out[2241] <= ~(x[4370] & x[4371]);
     layer0_out[2242] <= ~x[4317];
     layer0_out[2243] <= ~(x[441] & x[442]);
     layer0_out[2244] <= x[2477] & x[2479];
     layer0_out[2245] <= ~(x[6182] | x[6183]);
     layer0_out[2246] <= ~x[106];
     layer0_out[2247] <= x[7322] & x[7323];
     layer0_out[2248] <= x[386] & ~x[385];
     layer0_out[2249] <= x[2692] ^ x[2693];
     layer0_out[2250] <= x[665];
     layer0_out[2251] <= ~(x[2039] ^ x[2041]);
     layer0_out[2252] <= ~(x[8781] | x[8782]);
     layer0_out[2253] <= x[2688] & x[2689];
     layer0_out[2254] <= ~(x[7048] & x[7049]);
     layer0_out[2255] <= ~(x[1354] ^ x[1355]);
     layer0_out[2256] <= ~(x[1176] | x[1177]);
     layer0_out[2257] <= ~x[6636];
     layer0_out[2258] <= ~(x[3721] | x[3722]);
     layer0_out[2259] <= ~(x[3643] ^ x[3644]);
     layer0_out[2260] <= 1'b0;
     layer0_out[2261] <= x[8925] & x[8926];
     layer0_out[2262] <= ~x[4922];
     layer0_out[2263] <= ~(x[2102] & x[2103]);
     layer0_out[2264] <= ~(x[4408] ^ x[4409]);
     layer0_out[2265] <= ~(x[6429] | x[6430]);
     layer0_out[2266] <= ~(x[2194] & x[2195]);
     layer0_out[2267] <= x[2425] & x[2426];
     layer0_out[2268] <= ~(x[7991] ^ x[7992]);
     layer0_out[2269] <= ~x[8453];
     layer0_out[2270] <= ~(x[2488] & x[2490]);
     layer0_out[2271] <= ~x[640];
     layer0_out[2272] <= x[6038] & x[6039];
     layer0_out[2273] <= ~x[106];
     layer0_out[2274] <= ~x[1269];
     layer0_out[2275] <= ~(x[4149] & x[4150]);
     layer0_out[2276] <= x[5027] & x[5028];
     layer0_out[2277] <= x[5607];
     layer0_out[2278] <= ~(x[2995] & x[2996]);
     layer0_out[2279] <= 1'b0;
     layer0_out[2280] <= x[6804] | x[6805];
     layer0_out[2281] <= ~(x[3402] | x[3403]);
     layer0_out[2282] <= x[1252] | x[1253];
     layer0_out[2283] <= x[5072] | x[5073];
     layer0_out[2284] <= x[7828] ^ x[7829];
     layer0_out[2285] <= ~(x[1590] & x[1591]);
     layer0_out[2286] <= ~(x[4676] & x[4677]);
     layer0_out[2287] <= ~(x[380] ^ x[381]);
     layer0_out[2288] <= ~(x[11] & x[13]);
     layer0_out[2289] <= ~(x[6153] | x[6154]);
     layer0_out[2290] <= x[3360] & ~x[3359];
     layer0_out[2291] <= ~(x[3294] | x[3295]);
     layer0_out[2292] <= ~(x[2671] & x[2672]);
     layer0_out[2293] <= ~(x[5024] | x[5025]);
     layer0_out[2294] <= x[9046];
     layer0_out[2295] <= x[1812] | x[1814];
     layer0_out[2296] <= 1'b0;
     layer0_out[2297] <= x[1477] & ~x[1479];
     layer0_out[2298] <= x[7501] ^ x[7502];
     layer0_out[2299] <= ~(x[5446] & x[5447]);
     layer0_out[2300] <= x[6451];
     layer0_out[2301] <= x[5515];
     layer0_out[2302] <= ~x[375] | x[373];
     layer0_out[2303] <= ~x[7860];
     layer0_out[2304] <= x[2426] | x[2427];
     layer0_out[2305] <= x[7149] ^ x[7150];
     layer0_out[2306] <= x[1621];
     layer0_out[2307] <= x[5105];
     layer0_out[2308] <= ~(x[2147] & x[2149]);
     layer0_out[2309] <= x[5757] & x[5758];
     layer0_out[2310] <= x[3589] & ~x[3588];
     layer0_out[2311] <= ~(x[4662] ^ x[4663]);
     layer0_out[2312] <= x[4928] | x[4929];
     layer0_out[2313] <= ~(x[2677] & x[2678]);
     layer0_out[2314] <= x[6902] | x[6903];
     layer0_out[2315] <= ~x[1229];
     layer0_out[2316] <= ~(x[7722] & x[7723]);
     layer0_out[2317] <= ~x[294];
     layer0_out[2318] <= x[2143] | x[2144];
     layer0_out[2319] <= x[2646] & x[2648];
     layer0_out[2320] <= x[1246] & ~x[1244];
     layer0_out[2321] <= ~(x[2953] & x[2954]);
     layer0_out[2322] <= x[2182];
     layer0_out[2323] <= x[8415] | x[8416];
     layer0_out[2324] <= ~(x[2664] | x[2665]);
     layer0_out[2325] <= ~(x[5451] & x[5452]);
     layer0_out[2326] <= x[302];
     layer0_out[2327] <= ~x[7170];
     layer0_out[2328] <= ~(x[213] | x[215]);
     layer0_out[2329] <= x[8666] | x[8667];
     layer0_out[2330] <= ~(x[3419] | x[3420]);
     layer0_out[2331] <= ~x[436] | x[438];
     layer0_out[2332] <= ~x[2724];
     layer0_out[2333] <= ~(x[8782] | x[8783]);
     layer0_out[2334] <= ~x[4435];
     layer0_out[2335] <= ~(x[8531] | x[8532]);
     layer0_out[2336] <= ~(x[808] ^ x[809]);
     layer0_out[2337] <= ~x[6693];
     layer0_out[2338] <= ~(x[5273] & x[5274]);
     layer0_out[2339] <= ~(x[5354] & x[5355]);
     layer0_out[2340] <= x[1724] & x[1725];
     layer0_out[2341] <= ~(x[1051] & x[1053]);
     layer0_out[2342] <= ~(x[6772] | x[6773]);
     layer0_out[2343] <= ~x[7653] | x[7654];
     layer0_out[2344] <= ~x[1144] | x[1143];
     layer0_out[2345] <= ~(x[3530] & x[3531]);
     layer0_out[2346] <= ~x[3604];
     layer0_out[2347] <= ~x[1916] | x[1915];
     layer0_out[2348] <= ~(x[1068] & x[1069]);
     layer0_out[2349] <= ~(x[7411] | x[7412]);
     layer0_out[2350] <= ~x[1440];
     layer0_out[2351] <= x[542] | x[543];
     layer0_out[2352] <= ~(x[3386] | x[3387]);
     layer0_out[2353] <= x[4373] ^ x[4374];
     layer0_out[2354] <= ~(x[2407] & x[2409]);
     layer0_out[2355] <= ~(x[6402] | x[6403]);
     layer0_out[2356] <= x[8388];
     layer0_out[2357] <= x[8517] & ~x[8516];
     layer0_out[2358] <= ~x[4791];
     layer0_out[2359] <= ~(x[2915] ^ x[2916]);
     layer0_out[2360] <= x[2090] & x[2092];
     layer0_out[2361] <= ~(x[1167] & x[1168]);
     layer0_out[2362] <= x[4815] & x[4816];
     layer0_out[2363] <= x[2049] & x[2051];
     layer0_out[2364] <= ~(x[1221] ^ x[1223]);
     layer0_out[2365] <= ~(x[4434] & x[4435]);
     layer0_out[2366] <= x[2113];
     layer0_out[2367] <= x[1535] & x[1536];
     layer0_out[2368] <= 1'b1;
     layer0_out[2369] <= ~(x[2177] & x[2179]);
     layer0_out[2370] <= x[6969];
     layer0_out[2371] <= ~(x[1881] ^ x[1882]);
     layer0_out[2372] <= x[950] | x[952];
     layer0_out[2373] <= ~(x[1122] & x[1123]);
     layer0_out[2374] <= x[2523] ^ x[2525];
     layer0_out[2375] <= x[4421];
     layer0_out[2376] <= x[2404] & x[2405];
     layer0_out[2377] <= x[1678] & x[1680];
     layer0_out[2378] <= x[102] | x[104];
     layer0_out[2379] <= ~x[2731];
     layer0_out[2380] <= ~(x[5222] & x[5223]);
     layer0_out[2381] <= ~(x[5508] & x[5509]);
     layer0_out[2382] <= x[1887];
     layer0_out[2383] <= ~x[3933] | x[3932];
     layer0_out[2384] <= ~(x[2861] ^ x[2862]);
     layer0_out[2385] <= x[959] & x[960];
     layer0_out[2386] <= ~(x[4318] | x[4319]);
     layer0_out[2387] <= 1'b1;
     layer0_out[2388] <= ~x[467];
     layer0_out[2389] <= x[2087] & x[2088];
     layer0_out[2390] <= 1'b1;
     layer0_out[2391] <= ~x[5653];
     layer0_out[2392] <= x[1320] & x[1322];
     layer0_out[2393] <= x[7530] | x[7531];
     layer0_out[2394] <= x[1073];
     layer0_out[2395] <= ~(x[3883] ^ x[3884]);
     layer0_out[2396] <= ~(x[4069] | x[4070]);
     layer0_out[2397] <= x[2663] ^ x[2664];
     layer0_out[2398] <= x[5213] & x[5214];
     layer0_out[2399] <= ~(x[2364] & x[2366]);
     layer0_out[2400] <= x[6161] & ~x[6160];
     layer0_out[2401] <= x[8107];
     layer0_out[2402] <= ~(x[6991] | x[6992]);
     layer0_out[2403] <= ~(x[4325] & x[4326]);
     layer0_out[2404] <= x[6396] | x[6397];
     layer0_out[2405] <= ~(x[1125] & x[1126]);
     layer0_out[2406] <= ~(x[1440] & x[1441]);
     layer0_out[2407] <= x[1867] | x[1868];
     layer0_out[2408] <= ~x[1237] | x[1235];
     layer0_out[2409] <= x[5574] | x[5575];
     layer0_out[2410] <= x[5195] & x[5196];
     layer0_out[2411] <= ~(x[721] ^ x[722]);
     layer0_out[2412] <= ~x[5685];
     layer0_out[2413] <= x[6189] | x[6190];
     layer0_out[2414] <= x[1875];
     layer0_out[2415] <= ~(x[2966] & x[2967]);
     layer0_out[2416] <= ~x[5672];
     layer0_out[2417] <= x[6853] & ~x[6854];
     layer0_out[2418] <= ~x[1043];
     layer0_out[2419] <= x[7113] ^ x[7114];
     layer0_out[2420] <= x[1840] ^ x[1842];
     layer0_out[2421] <= x[1415];
     layer0_out[2422] <= x[6634];
     layer0_out[2423] <= x[6776] & x[6777];
     layer0_out[2424] <= ~(x[1685] | x[1686]);
     layer0_out[2425] <= x[2281] ^ x[2283];
     layer0_out[2426] <= x[1146] & ~x[1145];
     layer0_out[2427] <= ~x[9007];
     layer0_out[2428] <= x[8149] & x[8150];
     layer0_out[2429] <= ~(x[1323] & x[1324]);
     layer0_out[2430] <= ~(x[5690] & x[5691]);
     layer0_out[2431] <= x[4363];
     layer0_out[2432] <= x[1710];
     layer0_out[2433] <= 1'b1;
     layer0_out[2434] <= ~x[1403];
     layer0_out[2435] <= x[290] ^ x[292];
     layer0_out[2436] <= ~x[7539];
     layer0_out[2437] <= ~(x[7408] | x[7409]);
     layer0_out[2438] <= x[1824] | x[1826];
     layer0_out[2439] <= ~(x[3154] & x[3155]);
     layer0_out[2440] <= ~(x[7052] & x[7053]);
     layer0_out[2441] <= ~(x[4716] ^ x[4717]);
     layer0_out[2442] <= x[1432] ^ x[1434];
     layer0_out[2443] <= x[6427] | x[6428];
     layer0_out[2444] <= ~(x[5518] | x[5519]);
     layer0_out[2445] <= ~(x[899] & x[901]);
     layer0_out[2446] <= ~x[1931];
     layer0_out[2447] <= ~(x[1425] & x[1426]);
     layer0_out[2448] <= x[375] & ~x[374];
     layer0_out[2449] <= ~(x[7225] | x[7226]);
     layer0_out[2450] <= ~(x[287] ^ x[289]);
     layer0_out[2451] <= ~x[828] | x[829];
     layer0_out[2452] <= 1'b0;
     layer0_out[2453] <= ~x[7441];
     layer0_out[2454] <= x[5908] & x[5909];
     layer0_out[2455] <= x[478] & ~x[479];
     layer0_out[2456] <= x[3814] & x[3815];
     layer0_out[2457] <= x[2680] & x[2682];
     layer0_out[2458] <= ~x[7008];
     layer0_out[2459] <= x[7196] & ~x[7195];
     layer0_out[2460] <= ~(x[761] & x[763]);
     layer0_out[2461] <= ~(x[2599] ^ x[2600]);
     layer0_out[2462] <= x[691] ^ x[693];
     layer0_out[2463] <= x[1958] ^ x[1959];
     layer0_out[2464] <= ~(x[4774] | x[4775]);
     layer0_out[2465] <= 1'b1;
     layer0_out[2466] <= ~(x[7085] ^ x[7086]);
     layer0_out[2467] <= x[5224] & x[5225];
     layer0_out[2468] <= ~x[7443];
     layer0_out[2469] <= x[882] | x[883];
     layer0_out[2470] <= x[4075];
     layer0_out[2471] <= x[803] & x[805];
     layer0_out[2472] <= x[7679];
     layer0_out[2473] <= ~(x[66] | x[67]);
     layer0_out[2474] <= ~x[3452] | x[3451];
     layer0_out[2475] <= ~(x[6625] | x[6626]);
     layer0_out[2476] <= x[2200] & x[2202];
     layer0_out[2477] <= x[7433] ^ x[7434];
     layer0_out[2478] <= ~x[3752];
     layer0_out[2479] <= ~x[1573] | x[1574];
     layer0_out[2480] <= x[8328] | x[8329];
     layer0_out[2481] <= ~(x[9079] & x[9080]);
     layer0_out[2482] <= ~(x[413] & x[414]);
     layer0_out[2483] <= x[4921];
     layer0_out[2484] <= x[1100] & x[1102];
     layer0_out[2485] <= x[2041] & x[2042];
     layer0_out[2486] <= x[7081] & ~x[7082];
     layer0_out[2487] <= x[10] ^ x[11];
     layer0_out[2488] <= x[6295];
     layer0_out[2489] <= ~(x[9002] & x[9003]);
     layer0_out[2490] <= ~(x[4167] | x[4168]);
     layer0_out[2491] <= ~(x[6566] & x[6567]);
     layer0_out[2492] <= ~(x[620] | x[621]);
     layer0_out[2493] <= ~x[6697] | x[6698];
     layer0_out[2494] <= x[342] & x[344];
     layer0_out[2495] <= ~(x[9023] & x[9024]);
     layer0_out[2496] <= 1'b0;
     layer0_out[2497] <= x[1536] & x[1538];
     layer0_out[2498] <= x[4244];
     layer0_out[2499] <= ~x[8050];
     layer0_out[2500] <= ~(x[6444] | x[6445]);
     layer0_out[2501] <= 1'b0;
     layer0_out[2502] <= ~(x[4977] | x[4978]);
     layer0_out[2503] <= ~(x[4158] & x[4159]);
     layer0_out[2504] <= x[254] & x[255];
     layer0_out[2505] <= ~x[162];
     layer0_out[2506] <= ~(x[2378] & x[2380]);
     layer0_out[2507] <= x[5301] | x[5302];
     layer0_out[2508] <= ~(x[7556] | x[7557]);
     layer0_out[2509] <= ~(x[733] ^ x[735]);
     layer0_out[2510] <= x[128] & x[129];
     layer0_out[2511] <= ~x[7023] | x[7024];
     layer0_out[2512] <= x[695] & x[696];
     layer0_out[2513] <= ~(x[4624] | x[4625]);
     layer0_out[2514] <= 1'b0;
     layer0_out[2515] <= 1'b1;
     layer0_out[2516] <= x[1632] & x[1633];
     layer0_out[2517] <= ~(x[5981] | x[5982]);
     layer0_out[2518] <= 1'b1;
     layer0_out[2519] <= ~(x[1539] ^ x[1540]);
     layer0_out[2520] <= x[2616] & x[2618];
     layer0_out[2521] <= ~x[1338];
     layer0_out[2522] <= x[2867] & x[2868];
     layer0_out[2523] <= ~(x[3590] ^ x[3591]);
     layer0_out[2524] <= ~(x[9064] | x[9065]);
     layer0_out[2525] <= ~(x[523] & x[525]);
     layer0_out[2526] <= ~(x[3650] & x[3651]);
     layer0_out[2527] <= 1'b0;
     layer0_out[2528] <= 1'b0;
     layer0_out[2529] <= x[5087] | x[5088];
     layer0_out[2530] <= x[9018];
     layer0_out[2531] <= x[2794] | x[2795];
     layer0_out[2532] <= x[151] & x[153];
     layer0_out[2533] <= x[4915] | x[4916];
     layer0_out[2534] <= ~(x[7032] | x[7033]);
     layer0_out[2535] <= x[7875] ^ x[7876];
     layer0_out[2536] <= x[5226] & x[5227];
     layer0_out[2537] <= ~(x[1886] | x[1887]);
     layer0_out[2538] <= x[650] ^ x[652];
     layer0_out[2539] <= x[141];
     layer0_out[2540] <= ~(x[3749] | x[3750]);
     layer0_out[2541] <= x[1186] & x[1188];
     layer0_out[2542] <= x[7258];
     layer0_out[2543] <= ~(x[7129] | x[7130]);
     layer0_out[2544] <= ~(x[1890] ^ x[1891]);
     layer0_out[2545] <= x[145] & x[147];
     layer0_out[2546] <= ~(x[1976] | x[1978]);
     layer0_out[2547] <= x[2921];
     layer0_out[2548] <= x[6685] & ~x[6684];
     layer0_out[2549] <= x[3635] | x[3636];
     layer0_out[2550] <= x[3232] & ~x[3233];
     layer0_out[2551] <= 1'b1;
     layer0_out[2552] <= x[8797];
     layer0_out[2553] <= x[28] & x[29];
     layer0_out[2554] <= x[2586] & ~x[2588];
     layer0_out[2555] <= ~x[277];
     layer0_out[2556] <= x[5206];
     layer0_out[2557] <= x[8520];
     layer0_out[2558] <= ~x[4780] | x[4781];
     layer0_out[2559] <= x[986] & ~x[988];
     layer0_out[2560] <= ~(x[4017] | x[4018]);
     layer0_out[2561] <= ~(x[1182] & x[1184]);
     layer0_out[2562] <= x[2273] ^ x[2275];
     layer0_out[2563] <= x[3583] & x[3584];
     layer0_out[2564] <= x[4656] | x[4657];
     layer0_out[2565] <= x[2615] & x[2616];
     layer0_out[2566] <= ~(x[3331] & x[3332]);
     layer0_out[2567] <= ~x[8877];
     layer0_out[2568] <= x[2960] & x[2961];
     layer0_out[2569] <= ~(x[3502] & x[3503]);
     layer0_out[2570] <= x[414];
     layer0_out[2571] <= x[6865] ^ x[6866];
     layer0_out[2572] <= x[2261] & x[2263];
     layer0_out[2573] <= x[3859] ^ x[3860];
     layer0_out[2574] <= x[5752] ^ x[5753];
     layer0_out[2575] <= x[6647] | x[6648];
     layer0_out[2576] <= ~(x[6285] & x[6286]);
     layer0_out[2577] <= x[982] & x[983];
     layer0_out[2578] <= ~(x[4813] | x[4814]);
     layer0_out[2579] <= ~x[7349];
     layer0_out[2580] <= x[7489] & ~x[7488];
     layer0_out[2581] <= ~x[2661] | x[2663];
     layer0_out[2582] <= ~x[8632] | x[8631];
     layer0_out[2583] <= x[1265] & x[1267];
     layer0_out[2584] <= ~(x[7074] | x[7075]);
     layer0_out[2585] <= x[6243];
     layer0_out[2586] <= x[7405] | x[7406];
     layer0_out[2587] <= ~(x[2160] & x[2161]);
     layer0_out[2588] <= ~(x[4473] & x[4474]);
     layer0_out[2589] <= x[1313] ^ x[1314];
     layer0_out[2590] <= ~x[59] | x[61];
     layer0_out[2591] <= x[8137];
     layer0_out[2592] <= x[4549];
     layer0_out[2593] <= ~(x[8260] & x[8261]);
     layer0_out[2594] <= x[5066] | x[5067];
     layer0_out[2595] <= x[3743] & ~x[3744];
     layer0_out[2596] <= ~(x[5376] & x[5377]);
     layer0_out[2597] <= ~x[536];
     layer0_out[2598] <= x[4412] & x[4413];
     layer0_out[2599] <= ~(x[2050] | x[2051]);
     layer0_out[2600] <= x[7711];
     layer0_out[2601] <= ~x[1071];
     layer0_out[2602] <= ~(x[3850] | x[3851]);
     layer0_out[2603] <= ~(x[6573] | x[6574]);
     layer0_out[2604] <= x[2757] ^ x[2759];
     layer0_out[2605] <= x[1276];
     layer0_out[2606] <= ~(x[2589] | x[2590]);
     layer0_out[2607] <= ~(x[528] & x[529]);
     layer0_out[2608] <= x[5723] & x[5724];
     layer0_out[2609] <= x[6085];
     layer0_out[2610] <= x[2165] & x[2167];
     layer0_out[2611] <= x[6541] & ~x[6540];
     layer0_out[2612] <= x[2167] & x[2169];
     layer0_out[2613] <= ~(x[2719] & x[2721]);
     layer0_out[2614] <= x[2571] & x[2573];
     layer0_out[2615] <= 1'b1;
     layer0_out[2616] <= 1'b1;
     layer0_out[2617] <= x[3351] | x[3352];
     layer0_out[2618] <= x[99] | x[101];
     layer0_out[2619] <= ~x[8542];
     layer0_out[2620] <= ~x[1721];
     layer0_out[2621] <= ~(x[5898] & x[5899]);
     layer0_out[2622] <= ~x[2037];
     layer0_out[2623] <= ~(x[5502] & x[5503]);
     layer0_out[2624] <= ~(x[8719] | x[8720]);
     layer0_out[2625] <= 1'b1;
     layer0_out[2626] <= x[6289] | x[6290];
     layer0_out[2627] <= x[6811];
     layer0_out[2628] <= x[3350];
     layer0_out[2629] <= ~(x[3849] | x[3850]);
     layer0_out[2630] <= x[4477] & ~x[4476];
     layer0_out[2631] <= x[6364] & ~x[6363];
     layer0_out[2632] <= 1'b1;
     layer0_out[2633] <= x[6357];
     layer0_out[2634] <= x[1500] & x[1502];
     layer0_out[2635] <= x[3450] | x[3451];
     layer0_out[2636] <= x[4546] & ~x[4547];
     layer0_out[2637] <= x[3518] ^ x[3519];
     layer0_out[2638] <= x[5013] | x[5014];
     layer0_out[2639] <= ~(x[657] ^ x[658]);
     layer0_out[2640] <= ~(x[2308] & x[2310]);
     layer0_out[2641] <= ~(x[8160] ^ x[8161]);
     layer0_out[2642] <= ~(x[9067] | x[9068]);
     layer0_out[2643] <= ~x[1887];
     layer0_out[2644] <= ~x[8968];
     layer0_out[2645] <= x[4681] | x[4682];
     layer0_out[2646] <= x[8147];
     layer0_out[2647] <= x[3691] & x[3692];
     layer0_out[2648] <= ~x[3305];
     layer0_out[2649] <= ~x[2877];
     layer0_out[2650] <= ~(x[2367] & x[2368]);
     layer0_out[2651] <= x[6036];
     layer0_out[2652] <= ~(x[3807] ^ x[3808]);
     layer0_out[2653] <= x[8133] & ~x[8132];
     layer0_out[2654] <= ~(x[2827] | x[2828]);
     layer0_out[2655] <= ~(x[1758] | x[1760]);
     layer0_out[2656] <= ~(x[8950] & x[8951]);
     layer0_out[2657] <= x[24] & x[25];
     layer0_out[2658] <= x[4645] & ~x[4644];
     layer0_out[2659] <= ~(x[5550] | x[5551]);
     layer0_out[2660] <= ~(x[2518] ^ x[2520]);
     layer0_out[2661] <= x[4717] & x[4718];
     layer0_out[2662] <= ~(x[2459] ^ x[2461]);
     layer0_out[2663] <= ~x[7447];
     layer0_out[2664] <= ~(x[3363] & x[3364]);
     layer0_out[2665] <= x[1609] & x[1611];
     layer0_out[2666] <= ~(x[5544] | x[5545]);
     layer0_out[2667] <= x[6806] & x[6807];
     layer0_out[2668] <= x[1460] & ~x[1462];
     layer0_out[2669] <= ~(x[8998] & x[8999]);
     layer0_out[2670] <= ~x[1008];
     layer0_out[2671] <= x[2188] & x[2189];
     layer0_out[2672] <= ~(x[4146] | x[4147]);
     layer0_out[2673] <= ~x[987];
     layer0_out[2674] <= 1'b0;
     layer0_out[2675] <= x[1663] & x[1664];
     layer0_out[2676] <= x[259] & ~x[257];
     layer0_out[2677] <= x[5598] & ~x[5597];
     layer0_out[2678] <= ~(x[6234] | x[6235]);
     layer0_out[2679] <= x[2413] & x[2414];
     layer0_out[2680] <= x[1720] & x[1722];
     layer0_out[2681] <= x[5043] ^ x[5044];
     layer0_out[2682] <= x[960];
     layer0_out[2683] <= x[1387] & ~x[1385];
     layer0_out[2684] <= ~x[1367];
     layer0_out[2685] <= ~x[2463];
     layer0_out[2686] <= ~(x[2519] & x[2521]);
     layer0_out[2687] <= ~(x[2634] & x[2635]);
     layer0_out[2688] <= ~x[356];
     layer0_out[2689] <= ~(x[3261] | x[3262]);
     layer0_out[2690] <= x[551] & x[553];
     layer0_out[2691] <= ~(x[7063] | x[7064]);
     layer0_out[2692] <= ~(x[1314] & x[1315]);
     layer0_out[2693] <= ~(x[4963] & x[4964]);
     layer0_out[2694] <= x[251] & ~x[249];
     layer0_out[2695] <= x[6649] | x[6650];
     layer0_out[2696] <= ~(x[175] & x[176]);
     layer0_out[2697] <= x[4004] & ~x[4003];
     layer0_out[2698] <= ~(x[8507] & x[8508]);
     layer0_out[2699] <= x[4976] ^ x[4977];
     layer0_out[2700] <= ~x[7824];
     layer0_out[2701] <= ~x[2230];
     layer0_out[2702] <= ~(x[4767] & x[4768]);
     layer0_out[2703] <= 1'b1;
     layer0_out[2704] <= x[8574];
     layer0_out[2705] <= ~(x[526] & x[527]);
     layer0_out[2706] <= ~(x[1192] | x[1194]);
     layer0_out[2707] <= ~(x[683] & x[685]);
     layer0_out[2708] <= x[910] & x[912];
     layer0_out[2709] <= ~(x[6068] & x[6069]);
     layer0_out[2710] <= ~(x[1542] & x[1543]);
     layer0_out[2711] <= ~(x[1352] & x[1353]);
     layer0_out[2712] <= ~(x[6348] | x[6349]);
     layer0_out[2713] <= ~x[419] | x[421];
     layer0_out[2714] <= x[9209] | x[9210];
     layer0_out[2715] <= ~(x[3026] & x[3027]);
     layer0_out[2716] <= x[6913];
     layer0_out[2717] <= x[4620] | x[4621];
     layer0_out[2718] <= ~x[4162];
     layer0_out[2719] <= ~x[4657];
     layer0_out[2720] <= ~(x[7487] ^ x[7488]);
     layer0_out[2721] <= ~x[1907];
     layer0_out[2722] <= ~x[957] | x[959];
     layer0_out[2723] <= 1'b0;
     layer0_out[2724] <= x[3173];
     layer0_out[2725] <= x[2686] & x[2688];
     layer0_out[2726] <= ~(x[6896] | x[6897]);
     layer0_out[2727] <= ~(x[8051] & x[8052]);
     layer0_out[2728] <= ~x[1248];
     layer0_out[2729] <= ~x[2371];
     layer0_out[2730] <= x[6727];
     layer0_out[2731] <= x[5260] | x[5261];
     layer0_out[2732] <= 1'b1;
     layer0_out[2733] <= ~(x[4999] | x[5000]);
     layer0_out[2734] <= x[873];
     layer0_out[2735] <= ~x[1923];
     layer0_out[2736] <= x[4362] ^ x[4363];
     layer0_out[2737] <= ~(x[1970] | x[1971]);
     layer0_out[2738] <= x[6221] ^ x[6222];
     layer0_out[2739] <= x[5997];
     layer0_out[2740] <= x[6476];
     layer0_out[2741] <= x[758];
     layer0_out[2742] <= x[2329] & ~x[2327];
     layer0_out[2743] <= x[3703] & x[3704];
     layer0_out[2744] <= x[5976] | x[5977];
     layer0_out[2745] <= 1'b0;
     layer0_out[2746] <= 1'b1;
     layer0_out[2747] <= ~(x[7022] | x[7023]);
     layer0_out[2748] <= x[7106] | x[7107];
     layer0_out[2749] <= ~(x[6177] | x[6178]);
     layer0_out[2750] <= x[9004];
     layer0_out[2751] <= x[4775] ^ x[4776];
     layer0_out[2752] <= x[6905];
     layer0_out[2753] <= x[1757] | x[1759];
     layer0_out[2754] <= x[8974] & x[8975];
     layer0_out[2755] <= x[5025] | x[5026];
     layer0_out[2756] <= ~(x[7340] & x[7341]);
     layer0_out[2757] <= x[7992] ^ x[7993];
     layer0_out[2758] <= x[2800] & ~x[2801];
     layer0_out[2759] <= ~x[2211];
     layer0_out[2760] <= ~x[7429] | x[7430];
     layer0_out[2761] <= x[5569] & x[5570];
     layer0_out[2762] <= x[3059] & x[3060];
     layer0_out[2763] <= ~(x[4419] ^ x[4420]);
     layer0_out[2764] <= ~x[7573];
     layer0_out[2765] <= x[122] ^ x[123];
     layer0_out[2766] <= ~(x[5836] & x[5837]);
     layer0_out[2767] <= ~x[7781];
     layer0_out[2768] <= x[427] & ~x[426];
     layer0_out[2769] <= x[5194] & x[5195];
     layer0_out[2770] <= ~(x[8445] ^ x[8446]);
     layer0_out[2771] <= x[2432];
     layer0_out[2772] <= x[3777] ^ x[3778];
     layer0_out[2773] <= x[54] & x[55];
     layer0_out[2774] <= x[5590];
     layer0_out[2775] <= 1'b0;
     layer0_out[2776] <= x[7942] | x[7943];
     layer0_out[2777] <= x[3976] | x[3977];
     layer0_out[2778] <= x[7575];
     layer0_out[2779] <= x[6459];
     layer0_out[2780] <= x[2517];
     layer0_out[2781] <= x[2505] & x[2507];
     layer0_out[2782] <= x[8478] & ~x[8479];
     layer0_out[2783] <= x[8722] & x[8723];
     layer0_out[2784] <= ~x[1133] | x[1132];
     layer0_out[2785] <= x[2953] & ~x[2952];
     layer0_out[2786] <= x[1163] & x[1164];
     layer0_out[2787] <= x[7403] | x[7404];
     layer0_out[2788] <= ~x[7716];
     layer0_out[2789] <= ~x[8961] | x[8960];
     layer0_out[2790] <= x[6462];
     layer0_out[2791] <= 1'b1;
     layer0_out[2792] <= x[3792];
     layer0_out[2793] <= ~(x[6883] ^ x[6884]);
     layer0_out[2794] <= ~(x[1734] & x[1735]);
     layer0_out[2795] <= x[613] & x[615];
     layer0_out[2796] <= ~(x[8792] | x[8793]);
     layer0_out[2797] <= ~(x[368] & x[369]);
     layer0_out[2798] <= ~(x[8041] | x[8042]);
     layer0_out[2799] <= x[6983];
     layer0_out[2800] <= x[7719] | x[7720];
     layer0_out[2801] <= ~x[168] | x[167];
     layer0_out[2802] <= x[388];
     layer0_out[2803] <= ~(x[1666] & x[1668]);
     layer0_out[2804] <= ~(x[7659] | x[7660]);
     layer0_out[2805] <= ~(x[735] ^ x[736]);
     layer0_out[2806] <= x[5946] & x[5947];
     layer0_out[2807] <= x[2173] & x[2175];
     layer0_out[2808] <= x[5319] & x[5320];
     layer0_out[2809] <= x[2129] & ~x[2127];
     layer0_out[2810] <= x[1623] ^ x[1624];
     layer0_out[2811] <= ~(x[1866] ^ x[1867]);
     layer0_out[2812] <= ~(x[7562] | x[7563]);
     layer0_out[2813] <= x[1449] & x[1450];
     layer0_out[2814] <= ~x[9205];
     layer0_out[2815] <= ~x[5638];
     layer0_out[2816] <= 1'b1;
     layer0_out[2817] <= 1'b0;
     layer0_out[2818] <= ~(x[7551] ^ x[7552]);
     layer0_out[2819] <= x[1025] & x[1026];
     layer0_out[2820] <= ~x[3768];
     layer0_out[2821] <= 1'b1;
     layer0_out[2822] <= x[1079] & x[1081];
     layer0_out[2823] <= ~(x[1630] ^ x[1631]);
     layer0_out[2824] <= ~(x[1222] | x[1223]);
     layer0_out[2825] <= x[2260] & x[2262];
     layer0_out[2826] <= ~x[748];
     layer0_out[2827] <= ~(x[2231] & x[2233]);
     layer0_out[2828] <= x[1101];
     layer0_out[2829] <= x[5753] | x[5754];
     layer0_out[2830] <= ~x[7703];
     layer0_out[2831] <= x[396];
     layer0_out[2832] <= ~x[9133];
     layer0_out[2833] <= ~x[2683];
     layer0_out[2834] <= x[2072] & x[2073];
     layer0_out[2835] <= x[2235] & ~x[2234];
     layer0_out[2836] <= ~x[7714];
     layer0_out[2837] <= x[467] & x[469];
     layer0_out[2838] <= x[5261] & x[5262];
     layer0_out[2839] <= x[7744] ^ x[7745];
     layer0_out[2840] <= ~(x[1879] | x[1881]);
     layer0_out[2841] <= x[5416] & x[5417];
     layer0_out[2842] <= ~(x[5735] | x[5736]);
     layer0_out[2843] <= ~(x[97] & x[98]);
     layer0_out[2844] <= x[6587] | x[6588];
     layer0_out[2845] <= ~(x[2118] & x[2120]);
     layer0_out[2846] <= ~x[4162];
     layer0_out[2847] <= x[619];
     layer0_out[2848] <= x[5413] & x[5414];
     layer0_out[2849] <= x[2070] & x[2071];
     layer0_out[2850] <= ~(x[1962] & x[1963]);
     layer0_out[2851] <= x[6439] ^ x[6440];
     layer0_out[2852] <= x[840] & x[841];
     layer0_out[2853] <= x[2130] | x[2132];
     layer0_out[2854] <= ~(x[4855] | x[4856]);
     layer0_out[2855] <= ~(x[729] ^ x[730]);
     layer0_out[2856] <= x[5783] & ~x[5784];
     layer0_out[2857] <= x[3532] & x[3533];
     layer0_out[2858] <= ~x[3052] | x[3053];
     layer0_out[2859] <= ~x[9194];
     layer0_out[2860] <= ~x[4927];
     layer0_out[2861] <= ~x[1802];
     layer0_out[2862] <= ~(x[1897] & x[1899]);
     layer0_out[2863] <= ~(x[3845] | x[3846]);
     layer0_out[2864] <= 1'b0;
     layer0_out[2865] <= ~x[258];
     layer0_out[2866] <= x[2464];
     layer0_out[2867] <= ~(x[1524] & x[1525]);
     layer0_out[2868] <= 1'b1;
     layer0_out[2869] <= ~(x[3136] & x[3137]);
     layer0_out[2870] <= ~(x[6710] & x[6711]);
     layer0_out[2871] <= 1'b0;
     layer0_out[2872] <= ~x[3644];
     layer0_out[2873] <= ~(x[410] ^ x[411]);
     layer0_out[2874] <= x[6050] & x[6051];
     layer0_out[2875] <= ~(x[1292] & x[1294]);
     layer0_out[2876] <= 1'b0;
     layer0_out[2877] <= ~x[1529] | x[1528];
     layer0_out[2878] <= ~(x[4516] ^ x[4517]);
     layer0_out[2879] <= x[1984];
     layer0_out[2880] <= x[3104] ^ x[3105];
     layer0_out[2881] <= ~(x[1841] & x[1842]);
     layer0_out[2882] <= x[2538] & x[2540];
     layer0_out[2883] <= ~(x[9139] ^ x[9140]);
     layer0_out[2884] <= ~x[6832];
     layer0_out[2885] <= ~x[4063];
     layer0_out[2886] <= ~x[3415];
     layer0_out[2887] <= ~x[9163];
     layer0_out[2888] <= ~(x[8728] ^ x[8729]);
     layer0_out[2889] <= x[1657] & x[1659];
     layer0_out[2890] <= ~(x[1173] | x[1174]);
     layer0_out[2891] <= x[7480] & x[7481];
     layer0_out[2892] <= x[6024] | x[6025];
     layer0_out[2893] <= ~x[975];
     layer0_out[2894] <= ~(x[83] ^ x[85]);
     layer0_out[2895] <= x[2213] & x[2214];
     layer0_out[2896] <= x[2932] ^ x[2933];
     layer0_out[2897] <= x[2744];
     layer0_out[2898] <= ~(x[19] & x[20]);
     layer0_out[2899] <= x[1498] & x[1499];
     layer0_out[2900] <= x[1724] & x[1726];
     layer0_out[2901] <= ~(x[8339] & x[8340]);
     layer0_out[2902] <= x[785] & x[787];
     layer0_out[2903] <= x[2339];
     layer0_out[2904] <= 1'b0;
     layer0_out[2905] <= ~(x[5650] & x[5651]);
     layer0_out[2906] <= ~(x[1417] & x[1419]);
     layer0_out[2907] <= x[284];
     layer0_out[2908] <= ~(x[3255] | x[3256]);
     layer0_out[2909] <= x[4532];
     layer0_out[2910] <= ~(x[7955] | x[7956]);
     layer0_out[2911] <= x[8986] | x[8987];
     layer0_out[2912] <= x[3095] & x[3096];
     layer0_out[2913] <= 1'b0;
     layer0_out[2914] <= ~x[3275];
     layer0_out[2915] <= x[8811] | x[8812];
     layer0_out[2916] <= 1'b0;
     layer0_out[2917] <= ~(x[4351] ^ x[4352]);
     layer0_out[2918] <= ~x[2352] | x[2351];
     layer0_out[2919] <= ~(x[5130] & x[5131]);
     layer0_out[2920] <= x[1116] & ~x[1118];
     layer0_out[2921] <= x[5509];
     layer0_out[2922] <= ~(x[781] & x[782]);
     layer0_out[2923] <= x[2719] & x[2720];
     layer0_out[2924] <= x[3438];
     layer0_out[2925] <= ~(x[759] ^ x[760]);
     layer0_out[2926] <= ~x[2126];
     layer0_out[2927] <= x[2898] & x[2899];
     layer0_out[2928] <= ~(x[8394] & x[8395]);
     layer0_out[2929] <= x[3141];
     layer0_out[2930] <= x[324] | x[325];
     layer0_out[2931] <= ~(x[8734] | x[8735]);
     layer0_out[2932] <= x[7148] & ~x[7149];
     layer0_out[2933] <= ~(x[7352] ^ x[7353]);
     layer0_out[2934] <= x[7268] & ~x[7269];
     layer0_out[2935] <= ~(x[3745] ^ x[3746]);
     layer0_out[2936] <= ~(x[7027] ^ x[7028]);
     layer0_out[2937] <= ~x[819] | x[818];
     layer0_out[2938] <= x[4539] & x[4540];
     layer0_out[2939] <= x[3556] & x[3557];
     layer0_out[2940] <= 1'b1;
     layer0_out[2941] <= x[2581] & x[2582];
     layer0_out[2942] <= ~(x[4460] & x[4461]);
     layer0_out[2943] <= x[6756] & ~x[6757];
     layer0_out[2944] <= x[1522] & x[1524];
     layer0_out[2945] <= x[7105] ^ x[7106];
     layer0_out[2946] <= x[142] & x[144];
     layer0_out[2947] <= ~(x[9110] & x[9111]);
     layer0_out[2948] <= x[8418];
     layer0_out[2949] <= x[6055] & ~x[6056];
     layer0_out[2950] <= x[9] & ~x[8];
     layer0_out[2951] <= x[3265] ^ x[3266];
     layer0_out[2952] <= x[854] & x[855];
     layer0_out[2953] <= 1'b0;
     layer0_out[2954] <= x[1744] & x[1746];
     layer0_out[2955] <= x[1394] & x[1395];
     layer0_out[2956] <= x[2131] & x[2132];
     layer0_out[2957] <= ~(x[3000] & x[3001]);
     layer0_out[2958] <= x[4593];
     layer0_out[2959] <= ~x[7882] | x[7881];
     layer0_out[2960] <= x[8172] & ~x[8171];
     layer0_out[2961] <= ~(x[7566] & x[7567]);
     layer0_out[2962] <= x[201] | x[203];
     layer0_out[2963] <= x[8266] & x[8267];
     layer0_out[2964] <= ~(x[1666] ^ x[1667]);
     layer0_out[2965] <= ~(x[5159] & x[5160]);
     layer0_out[2966] <= ~x[351];
     layer0_out[2967] <= x[4588];
     layer0_out[2968] <= ~x[510];
     layer0_out[2969] <= ~(x[7205] ^ x[7206]);
     layer0_out[2970] <= x[2092] & x[2093];
     layer0_out[2971] <= 1'b0;
     layer0_out[2972] <= x[3797];
     layer0_out[2973] <= x[6088];
     layer0_out[2974] <= ~(x[232] ^ x[234]);
     layer0_out[2975] <= ~(x[4108] & x[4109]);
     layer0_out[2976] <= ~(x[6448] | x[6449]);
     layer0_out[2977] <= x[156];
     layer0_out[2978] <= ~x[8509];
     layer0_out[2979] <= x[8752] | x[8753];
     layer0_out[2980] <= x[5097] & x[5098];
     layer0_out[2981] <= x[1680] & x[1682];
     layer0_out[2982] <= ~(x[2223] & x[2224]);
     layer0_out[2983] <= x[1190];
     layer0_out[2984] <= x[8914] | x[8915];
     layer0_out[2985] <= ~(x[181] | x[182]);
     layer0_out[2986] <= x[3796];
     layer0_out[2987] <= ~(x[2010] & x[2012]);
     layer0_out[2988] <= x[8289] | x[8290];
     layer0_out[2989] <= x[940] ^ x[942];
     layer0_out[2990] <= 1'b0;
     layer0_out[2991] <= ~(x[731] & x[733]);
     layer0_out[2992] <= ~(x[190] | x[191]);
     layer0_out[2993] <= 1'b0;
     layer0_out[2994] <= x[3362];
     layer0_out[2995] <= x[2897] & x[2898];
     layer0_out[2996] <= x[2566] | x[2568];
     layer0_out[2997] <= x[2679] & x[2681];
     layer0_out[2998] <= ~(x[1914] & x[1916]);
     layer0_out[2999] <= ~(x[4647] | x[4648]);
     layer0_out[3000] <= ~(x[2746] ^ x[2748]);
     layer0_out[3001] <= ~(x[756] | x[757]);
     layer0_out[3002] <= ~x[1954];
     layer0_out[3003] <= x[8002] | x[8003];
     layer0_out[3004] <= x[6821] & x[6822];
     layer0_out[3005] <= x[4832];
     layer0_out[3006] <= ~(x[8105] | x[8106]);
     layer0_out[3007] <= ~x[8702];
     layer0_out[3008] <= x[7958] | x[7959];
     layer0_out[3009] <= ~(x[518] ^ x[520]);
     layer0_out[3010] <= ~x[342];
     layer0_out[3011] <= ~(x[2636] ^ x[2637]);
     layer0_out[3012] <= ~(x[872] | x[874]);
     layer0_out[3013] <= x[333] | x[334];
     layer0_out[3014] <= ~(x[8304] | x[8305]);
     layer0_out[3015] <= x[1151] & x[1152];
     layer0_out[3016] <= x[820] | x[822];
     layer0_out[3017] <= 1'b0;
     layer0_out[3018] <= ~(x[7244] & x[7245]);
     layer0_out[3019] <= ~(x[951] & x[952]);
     layer0_out[3020] <= x[647] | x[648];
     layer0_out[3021] <= ~x[6243] | x[6244];
     layer0_out[3022] <= ~(x[3900] | x[3901]);
     layer0_out[3023] <= ~x[251] | x[250];
     layer0_out[3024] <= x[1527] & x[1528];
     layer0_out[3025] <= x[2108] & x[2109];
     layer0_out[3026] <= ~x[8930];
     layer0_out[3027] <= x[3607] ^ x[3608];
     layer0_out[3028] <= ~(x[5845] & x[5846]);
     layer0_out[3029] <= ~(x[1610] | x[1611]);
     layer0_out[3030] <= 1'b0;
     layer0_out[3031] <= x[4706] & x[4707];
     layer0_out[3032] <= ~(x[8683] & x[8684]);
     layer0_out[3033] <= ~x[4428];
     layer0_out[3034] <= ~(x[4326] ^ x[4327]);
     layer0_out[3035] <= x[3503] & x[3504];
     layer0_out[3036] <= x[7091] | x[7092];
     layer0_out[3037] <= x[4514];
     layer0_out[3038] <= ~(x[1215] ^ x[1217]);
     layer0_out[3039] <= ~x[8961];
     layer0_out[3040] <= ~x[36] | x[34];
     layer0_out[3041] <= ~(x[2030] & x[2031]);
     layer0_out[3042] <= x[88];
     layer0_out[3043] <= x[789] & x[790];
     layer0_out[3044] <= x[1178] & x[1180];
     layer0_out[3045] <= ~(x[9027] ^ x[9028]);
     layer0_out[3046] <= ~x[114];
     layer0_out[3047] <= x[3380] ^ x[3381];
     layer0_out[3048] <= ~(x[2296] & x[2298]);
     layer0_out[3049] <= x[3182] & x[3183];
     layer0_out[3050] <= ~(x[8747] | x[8748]);
     layer0_out[3051] <= x[7278];
     layer0_out[3052] <= x[2610];
     layer0_out[3053] <= ~(x[1894] | x[1895]);
     layer0_out[3054] <= x[500];
     layer0_out[3055] <= x[6110] & ~x[6111];
     layer0_out[3056] <= ~(x[6335] ^ x[6336]);
     layer0_out[3057] <= x[8429] | x[8430];
     layer0_out[3058] <= 1'b1;
     layer0_out[3059] <= 1'b0;
     layer0_out[3060] <= x[2312] & x[2314];
     layer0_out[3061] <= x[8981] & x[8982];
     layer0_out[3062] <= ~(x[1455] & x[1457]);
     layer0_out[3063] <= ~(x[1909] & x[1911]);
     layer0_out[3064] <= x[6238];
     layer0_out[3065] <= x[700] & ~x[702];
     layer0_out[3066] <= ~(x[5530] & x[5531]);
     layer0_out[3067] <= ~(x[2227] & x[2228]);
     layer0_out[3068] <= ~(x[1667] & x[1669]);
     layer0_out[3069] <= ~(x[2527] & x[2529]);
     layer0_out[3070] <= ~x[7472] | x[7471];
     layer0_out[3071] <= ~(x[459] & x[461]);
     layer0_out[3072] <= x[2608] ^ x[2609];
     layer0_out[3073] <= ~x[8843] | x[8842];
     layer0_out[3074] <= x[395] ^ x[396];
     layer0_out[3075] <= ~(x[4000] | x[4001]);
     layer0_out[3076] <= ~x[4942];
     layer0_out[3077] <= ~(x[1532] & x[1534]);
     layer0_out[3078] <= x[2236] ^ x[2237];
     layer0_out[3079] <= ~x[1465] | x[1466];
     layer0_out[3080] <= x[7927] | x[7928];
     layer0_out[3081] <= x[3281];
     layer0_out[3082] <= ~(x[2499] & x[2500]);
     layer0_out[3083] <= ~(x[5709] & x[5710]);
     layer0_out[3084] <= x[7059] & x[7060];
     layer0_out[3085] <= ~x[2527] | x[2525];
     layer0_out[3086] <= x[2099] & x[2101];
     layer0_out[3087] <= x[1249];
     layer0_out[3088] <= ~(x[5651] & x[5652]);
     layer0_out[3089] <= x[2098] & x[2100];
     layer0_out[3090] <= x[2660] ^ x[2662];
     layer0_out[3091] <= x[2975] & x[2976];
     layer0_out[3092] <= x[1284] & x[1285];
     layer0_out[3093] <= x[1294] & x[1295];
     layer0_out[3094] <= x[5306] & x[5307];
     layer0_out[3095] <= ~(x[1435] | x[1436]);
     layer0_out[3096] <= ~x[4106];
     layer0_out[3097] <= x[2153];
     layer0_out[3098] <= ~(x[1250] ^ x[1251]);
     layer0_out[3099] <= ~(x[1234] | x[1235]);
     layer0_out[3100] <= ~x[2991] | x[2990];
     layer0_out[3101] <= x[6280];
     layer0_out[3102] <= x[8354];
     layer0_out[3103] <= x[3228] & ~x[3229];
     layer0_out[3104] <= ~x[6389];
     layer0_out[3105] <= x[948] | x[949];
     layer0_out[3106] <= ~x[770];
     layer0_out[3107] <= ~x[2397];
     layer0_out[3108] <= ~(x[1031] & x[1033]);
     layer0_out[3109] <= x[3457] | x[3458];
     layer0_out[3110] <= ~x[1902];
     layer0_out[3111] <= x[7171] | x[7172];
     layer0_out[3112] <= x[6687] & x[6688];
     layer0_out[3113] <= ~x[5840] | x[5841];
     layer0_out[3114] <= x[5391] & x[5392];
     layer0_out[3115] <= x[6712];
     layer0_out[3116] <= 1'b0;
     layer0_out[3117] <= x[1292] ^ x[1293];
     layer0_out[3118] <= x[1673] & x[1674];
     layer0_out[3119] <= x[9145];
     layer0_out[3120] <= ~(x[5235] & x[5236]);
     layer0_out[3121] <= 1'b0;
     layer0_out[3122] <= x[1518] & x[1520];
     layer0_out[3123] <= ~x[8557];
     layer0_out[3124] <= x[3784] | x[3785];
     layer0_out[3125] <= x[8669] & x[8670];
     layer0_out[3126] <= ~(x[2238] & x[2239]);
     layer0_out[3127] <= x[4133] & x[4134];
     layer0_out[3128] <= x[6121] | x[6122];
     layer0_out[3129] <= x[8660] | x[8661];
     layer0_out[3130] <= 1'b1;
     layer0_out[3131] <= ~(x[4857] & x[4858]);
     layer0_out[3132] <= x[6963] & ~x[6962];
     layer0_out[3133] <= x[7188] ^ x[7189];
     layer0_out[3134] <= ~(x[2917] & x[2918]);
     layer0_out[3135] <= ~x[141] | x[139];
     layer0_out[3136] <= x[1487];
     layer0_out[3137] <= x[2635] & x[2637];
     layer0_out[3138] <= x[108] ^ x[109];
     layer0_out[3139] <= 1'b0;
     layer0_out[3140] <= x[2696] ^ x[2697];
     layer0_out[3141] <= x[6000] & x[6001];
     layer0_out[3142] <= ~(x[194] ^ x[196]);
     layer0_out[3143] <= x[1114] & x[1115];
     layer0_out[3144] <= x[1401];
     layer0_out[3145] <= ~x[1976];
     layer0_out[3146] <= x[1940] & x[1942];
     layer0_out[3147] <= 1'b1;
     layer0_out[3148] <= ~(x[452] | x[453]);
     layer0_out[3149] <= ~(x[7079] | x[7080]);
     layer0_out[3150] <= ~(x[158] & x[160]);
     layer0_out[3151] <= 1'b0;
     layer0_out[3152] <= x[9057];
     layer0_out[3153] <= ~(x[2369] | x[2371]);
     layer0_out[3154] <= x[1087];
     layer0_out[3155] <= x[1989] & x[1991];
     layer0_out[3156] <= x[2021] & x[2022];
     layer0_out[3157] <= x[7826];
     layer0_out[3158] <= x[2643];
     layer0_out[3159] <= x[3393] & ~x[3392];
     layer0_out[3160] <= ~x[7400];
     layer0_out[3161] <= x[409] ^ x[410];
     layer0_out[3162] <= x[1678] & x[1679];
     layer0_out[3163] <= ~x[4199] | x[4200];
     layer0_out[3164] <= 1'b1;
     layer0_out[3165] <= x[1030] & x[1032];
     layer0_out[3166] <= x[2023] & x[2024];
     layer0_out[3167] <= x[1755] | x[1757];
     layer0_out[3168] <= x[3606] & x[3607];
     layer0_out[3169] <= x[170] ^ x[171];
     layer0_out[3170] <= 1'b1;
     layer0_out[3171] <= x[1794] & x[1796];
     layer0_out[3172] <= x[8012] & x[8013];
     layer0_out[3173] <= ~(x[1239] | x[1240]);
     layer0_out[3174] <= ~x[1588];
     layer0_out[3175] <= ~(x[3036] & x[3037]);
     layer0_out[3176] <= ~x[1600] | x[1599];
     layer0_out[3177] <= ~(x[1779] | x[1780]);
     layer0_out[3178] <= x[1439] | x[1441];
     layer0_out[3179] <= ~(x[1651] | x[1652]);
     layer0_out[3180] <= ~(x[3219] & x[3220]);
     layer0_out[3181] <= x[1667] & x[1668];
     layer0_out[3182] <= ~(x[681] | x[682]);
     layer0_out[3183] <= x[9150] & x[9151];
     layer0_out[3184] <= 1'b0;
     layer0_out[3185] <= ~(x[2889] | x[2890]);
     layer0_out[3186] <= x[3152] | x[3153];
     layer0_out[3187] <= x[8883] & x[8884];
     layer0_out[3188] <= x[2549] & x[2551];
     layer0_out[3189] <= x[4640] ^ x[4641];
     layer0_out[3190] <= ~(x[1361] & x[1362]);
     layer0_out[3191] <= ~(x[3958] | x[3959]);
     layer0_out[3192] <= ~x[1836] | x[1835];
     layer0_out[3193] <= ~(x[4465] & x[4466]);
     layer0_out[3194] <= ~(x[1144] ^ x[1146]);
     layer0_out[3195] <= x[8056] ^ x[8057];
     layer0_out[3196] <= ~(x[3480] | x[3481]);
     layer0_out[3197] <= ~x[8840] | x[8841];
     layer0_out[3198] <= x[2317] ^ x[2319];
     layer0_out[3199] <= ~(x[293] & x[295]);
     layer0_out[3200] <= ~(x[370] & x[372]);
     layer0_out[3201] <= 1'b0;
     layer0_out[3202] <= x[1324] & x[1326];
     layer0_out[3203] <= ~(x[1101] & x[1103]);
     layer0_out[3204] <= ~(x[1538] | x[1539]);
     layer0_out[3205] <= ~(x[4645] & x[4646]);
     layer0_out[3206] <= x[3499] & ~x[3498];
     layer0_out[3207] <= x[1997] | x[1999];
     layer0_out[3208] <= 1'b0;
     layer0_out[3209] <= x[3260] | x[3261];
     layer0_out[3210] <= ~x[7832] | x[7833];
     layer0_out[3211] <= x[2673] & x[2674];
     layer0_out[3212] <= 1'b0;
     layer0_out[3213] <= x[5063] & x[5064];
     layer0_out[3214] <= ~x[4668];
     layer0_out[3215] <= ~(x[7707] ^ x[7708]);
     layer0_out[3216] <= ~(x[7153] | x[7154]);
     layer0_out[3217] <= ~x[4365] | x[4366];
     layer0_out[3218] <= ~x[8705] | x[8706];
     layer0_out[3219] <= x[6903] | x[6904];
     layer0_out[3220] <= x[8898] & x[8899];
     layer0_out[3221] <= ~x[1313];
     layer0_out[3222] <= ~(x[532] & x[534]);
     layer0_out[3223] <= x[3810];
     layer0_out[3224] <= x[1392] ^ x[1393];
     layer0_out[3225] <= x[1252] ^ x[1254];
     layer0_out[3226] <= x[3700] | x[3701];
     layer0_out[3227] <= ~x[6796];
     layer0_out[3228] <= ~x[826];
     layer0_out[3229] <= ~(x[6391] ^ x[6392]);
     layer0_out[3230] <= x[4481] & x[4482];
     layer0_out[3231] <= x[5271] & x[5272];
     layer0_out[3232] <= ~(x[7734] | x[7735]);
     layer0_out[3233] <= ~(x[3963] ^ x[3964]);
     layer0_out[3234] <= ~(x[3941] | x[3942]);
     layer0_out[3235] <= ~x[945] | x[946];
     layer0_out[3236] <= ~(x[1763] & x[1765]);
     layer0_out[3237] <= ~(x[2028] | x[2029]);
     layer0_out[3238] <= x[5479] & x[5480];
     layer0_out[3239] <= x[5189];
     layer0_out[3240] <= x[6066] & ~x[6065];
     layer0_out[3241] <= x[7764];
     layer0_out[3242] <= x[896];
     layer0_out[3243] <= x[7282];
     layer0_out[3244] <= x[7709] | x[7710];
     layer0_out[3245] <= ~x[1695];
     layer0_out[3246] <= x[1858];
     layer0_out[3247] <= ~x[143];
     layer0_out[3248] <= x[457];
     layer0_out[3249] <= ~x[8466];
     layer0_out[3250] <= ~(x[1323] ^ x[1325]);
     layer0_out[3251] <= ~(x[4041] | x[4042]);
     layer0_out[3252] <= ~(x[965] & x[966]);
     layer0_out[3253] <= 1'b0;
     layer0_out[3254] <= ~(x[8217] & x[8218]);
     layer0_out[3255] <= 1'b0;
     layer0_out[3256] <= ~(x[1533] ^ x[1534]);
     layer0_out[3257] <= x[3856] ^ x[3857];
     layer0_out[3258] <= ~(x[5618] | x[5619]);
     layer0_out[3259] <= x[9088] & x[9089];
     layer0_out[3260] <= x[9001] ^ x[9002];
     layer0_out[3261] <= x[5234] & x[5235];
     layer0_out[3262] <= ~(x[5032] ^ x[5033]);
     layer0_out[3263] <= x[5187] | x[5188];
     layer0_out[3264] <= x[9117] | x[9118];
     layer0_out[3265] <= ~x[3916];
     layer0_out[3266] <= ~(x[3279] | x[3280]);
     layer0_out[3267] <= x[6590] | x[6591];
     layer0_out[3268] <= x[7374] & x[7375];
     layer0_out[3269] <= x[1810] | x[1811];
     layer0_out[3270] <= x[2726] & x[2728];
     layer0_out[3271] <= x[8790];
     layer0_out[3272] <= ~x[8048];
     layer0_out[3273] <= ~(x[6104] & x[6105]);
     layer0_out[3274] <= ~x[53] | x[55];
     layer0_out[3275] <= ~(x[367] & x[368]);
     layer0_out[3276] <= ~(x[3880] ^ x[3881]);
     layer0_out[3277] <= ~(x[5164] & x[5165]);
     layer0_out[3278] <= x[5524] & x[5525];
     layer0_out[3279] <= x[1961];
     layer0_out[3280] <= ~(x[2746] ^ x[2747]);
     layer0_out[3281] <= x[1919];
     layer0_out[3282] <= x[4868] & x[4869];
     layer0_out[3283] <= ~(x[2753] | x[2754]);
     layer0_out[3284] <= ~x[1490];
     layer0_out[3285] <= ~x[1615];
     layer0_out[3286] <= ~(x[3254] ^ x[3255]);
     layer0_out[3287] <= ~x[1260] | x[1259];
     layer0_out[3288] <= ~(x[1637] & x[1638]);
     layer0_out[3289] <= ~(x[1855] & x[1856]);
     layer0_out[3290] <= ~x[833];
     layer0_out[3291] <= x[7814] ^ x[7815];
     layer0_out[3292] <= x[1262] & x[1263];
     layer0_out[3293] <= ~(x[1634] & x[1635]);
     layer0_out[3294] <= 1'b0;
     layer0_out[3295] <= x[2589] | x[2591];
     layer0_out[3296] <= x[2079] & x[2081];
     layer0_out[3297] <= ~x[4723] | x[4722];
     layer0_out[3298] <= ~x[1251];
     layer0_out[3299] <= ~(x[7404] ^ x[7405]);
     layer0_out[3300] <= ~(x[3954] & x[3955]);
     layer0_out[3301] <= x[1308] & x[1310];
     layer0_out[3302] <= x[8098];
     layer0_out[3303] <= ~x[600];
     layer0_out[3304] <= ~x[2308];
     layer0_out[3305] <= ~(x[1066] ^ x[1068]);
     layer0_out[3306] <= ~(x[2215] & x[2216]);
     layer0_out[3307] <= ~(x[1084] & x[1086]);
     layer0_out[3308] <= ~(x[2599] & x[2601]);
     layer0_out[3309] <= ~(x[1616] | x[1617]);
     layer0_out[3310] <= x[2945];
     layer0_out[3311] <= ~(x[8628] | x[8629]);
     layer0_out[3312] <= x[1193];
     layer0_out[3313] <= x[6830] & x[6831];
     layer0_out[3314] <= ~x[6325] | x[6324];
     layer0_out[3315] <= x[3990];
     layer0_out[3316] <= ~(x[463] & x[465]);
     layer0_out[3317] <= ~(x[904] | x[905]);
     layer0_out[3318] <= ~(x[1135] ^ x[1137]);
     layer0_out[3319] <= ~x[6302];
     layer0_out[3320] <= ~(x[973] ^ x[974]);
     layer0_out[3321] <= ~x[1691];
     layer0_out[3322] <= x[3796] | x[3797];
     layer0_out[3323] <= ~(x[4441] & x[4442]);
     layer0_out[3324] <= ~(x[94] & x[95]);
     layer0_out[3325] <= x[3120];
     layer0_out[3326] <= ~x[1575];
     layer0_out[3327] <= ~(x[8462] & x[8463]);
     layer0_out[3328] <= x[837] & x[838];
     layer0_out[3329] <= ~x[7242];
     layer0_out[3330] <= ~(x[1359] & x[1361]);
     layer0_out[3331] <= ~(x[2103] & x[2104]);
     layer0_out[3332] <= 1'b1;
     layer0_out[3333] <= ~(x[4946] & x[4947]);
     layer0_out[3334] <= 1'b0;
     layer0_out[3335] <= x[6350] | x[6351];
     layer0_out[3336] <= x[8232];
     layer0_out[3337] <= ~(x[2004] | x[2005]);
     layer0_out[3338] <= x[8844] & ~x[8843];
     layer0_out[3339] <= x[6337] | x[6338];
     layer0_out[3340] <= ~x[7545];
     layer0_out[3341] <= x[7350] & ~x[7351];
     layer0_out[3342] <= x[984];
     layer0_out[3343] <= x[2243] & x[2244];
     layer0_out[3344] <= x[1381] | x[1382];
     layer0_out[3345] <= ~(x[998] & x[1000]);
     layer0_out[3346] <= 1'b1;
     layer0_out[3347] <= x[6550] | x[6551];
     layer0_out[3348] <= x[2057] & x[2059];
     layer0_out[3349] <= x[2468] ^ x[2469];
     layer0_out[3350] <= ~x[7330] | x[7329];
     layer0_out[3351] <= ~(x[2374] & x[2375]);
     layer0_out[3352] <= ~(x[7899] | x[7900]);
     layer0_out[3353] <= x[573] ^ x[575];
     layer0_out[3354] <= x[1165];
     layer0_out[3355] <= ~x[2524];
     layer0_out[3356] <= x[303] | x[305];
     layer0_out[3357] <= 1'b0;
     layer0_out[3358] <= x[1928];
     layer0_out[3359] <= 1'b1;
     layer0_out[3360] <= ~(x[4293] & x[4294]);
     layer0_out[3361] <= ~(x[3862] | x[3863]);
     layer0_out[3362] <= x[1551] & x[1553];
     layer0_out[3363] <= ~(x[2585] & x[2587]);
     layer0_out[3364] <= 1'b1;
     layer0_out[3365] <= ~(x[7086] & x[7087]);
     layer0_out[3366] <= ~(x[1544] | x[1546]);
     layer0_out[3367] <= x[1078] ^ x[1080];
     layer0_out[3368] <= ~x[4291];
     layer0_out[3369] <= ~(x[4260] ^ x[4261]);
     layer0_out[3370] <= ~(x[8033] | x[8034]);
     layer0_out[3371] <= ~(x[1523] & x[1525]);
     layer0_out[3372] <= ~(x[8797] ^ x[8798]);
     layer0_out[3373] <= ~(x[4194] | x[4195]);
     layer0_out[3374] <= ~(x[2455] & x[2456]);
     layer0_out[3375] <= ~(x[400] | x[402]);
     layer0_out[3376] <= ~x[3511];
     layer0_out[3377] <= 1'b1;
     layer0_out[3378] <= x[444] & x[445];
     layer0_out[3379] <= x[5546];
     layer0_out[3380] <= ~(x[3877] | x[3878]);
     layer0_out[3381] <= 1'b0;
     layer0_out[3382] <= ~x[4184];
     layer0_out[3383] <= x[2020] & x[2022];
     layer0_out[3384] <= x[6851] & ~x[6850];
     layer0_out[3385] <= x[5427];
     layer0_out[3386] <= x[8983] | x[8984];
     layer0_out[3387] <= ~(x[2338] & x[2340]);
     layer0_out[3388] <= ~(x[2303] & x[2304]);
     layer0_out[3389] <= x[7756] | x[7757];
     layer0_out[3390] <= ~(x[2111] & x[2113]);
     layer0_out[3391] <= x[8783] | x[8784];
     layer0_out[3392] <= ~x[130];
     layer0_out[3393] <= x[8250] | x[8251];
     layer0_out[3394] <= x[3139] & x[3140];
     layer0_out[3395] <= 1'b1;
     layer0_out[3396] <= x[3861] | x[3862];
     layer0_out[3397] <= x[5031] & x[5032];
     layer0_out[3398] <= ~x[6818] | x[6817];
     layer0_out[3399] <= ~(x[746] | x[747]);
     layer0_out[3400] <= ~x[1493];
     layer0_out[3401] <= ~x[974];
     layer0_out[3402] <= x[388] ^ x[390];
     layer0_out[3403] <= ~(x[671] | x[672]);
     layer0_out[3404] <= ~x[5293];
     layer0_out[3405] <= ~(x[1992] & x[1993]);
     layer0_out[3406] <= x[3523];
     layer0_out[3407] <= ~(x[2164] & x[2166]);
     layer0_out[3408] <= x[2078];
     layer0_out[3409] <= x[345] ^ x[347];
     layer0_out[3410] <= ~x[474];
     layer0_out[3411] <= x[1054] & x[1056];
     layer0_out[3412] <= ~x[2116];
     layer0_out[3413] <= ~(x[910] | x[911]);
     layer0_out[3414] <= x[8698];
     layer0_out[3415] <= ~(x[737] | x[738]);
     layer0_out[3416] <= ~x[8326] | x[8327];
     layer0_out[3417] <= ~(x[5091] | x[5092]);
     layer0_out[3418] <= ~(x[8877] ^ x[8878]);
     layer0_out[3419] <= ~(x[615] ^ x[616]);
     layer0_out[3420] <= ~x[3804] | x[3803];
     layer0_out[3421] <= ~(x[6824] & x[6825]);
     layer0_out[3422] <= ~(x[3044] ^ x[3045]);
     layer0_out[3423] <= ~x[21] | x[22];
     layer0_out[3424] <= x[3172] & ~x[3171];
     layer0_out[3425] <= x[3833] & x[3834];
     layer0_out[3426] <= x[7214];
     layer0_out[3427] <= ~(x[2584] | x[2585]);
     layer0_out[3428] <= x[8563] | x[8564];
     layer0_out[3429] <= x[543] & x[544];
     layer0_out[3430] <= x[7558] ^ x[7559];
     layer0_out[3431] <= x[2799] & x[2800];
     layer0_out[3432] <= ~(x[7739] ^ x[7740]);
     layer0_out[3433] <= x[1604] & x[1606];
     layer0_out[3434] <= x[3163] ^ x[3164];
     layer0_out[3435] <= x[787] | x[789];
     layer0_out[3436] <= ~(x[72] | x[73]);
     layer0_out[3437] <= x[7522];
     layer0_out[3438] <= ~(x[2059] & x[2061]);
     layer0_out[3439] <= x[6271] ^ x[6272];
     layer0_out[3440] <= ~(x[4137] | x[4138]);
     layer0_out[3441] <= ~(x[320] & x[321]);
     layer0_out[3442] <= ~(x[5404] & x[5405]);
     layer0_out[3443] <= ~x[2392];
     layer0_out[3444] <= ~x[6700];
     layer0_out[3445] <= x[5695] | x[5696];
     layer0_out[3446] <= ~(x[1652] | x[1654]);
     layer0_out[3447] <= x[2590] | x[2591];
     layer0_out[3448] <= ~(x[3476] | x[3477]);
     layer0_out[3449] <= x[2485] & x[2486];
     layer0_out[3450] <= x[2319] & x[2321];
     layer0_out[3451] <= x[2440] & x[2442];
     layer0_out[3452] <= ~(x[2754] & x[2755]);
     layer0_out[3453] <= x[8822] | x[8823];
     layer0_out[3454] <= x[670];
     layer0_out[3455] <= x[154] & x[155];
     layer0_out[3456] <= x[3016] & x[3017];
     layer0_out[3457] <= x[7338] ^ x[7339];
     layer0_out[3458] <= ~(x[6683] ^ x[6684]);
     layer0_out[3459] <= x[4518] & x[4519];
     layer0_out[3460] <= x[4274] & x[4275];
     layer0_out[3461] <= ~(x[1413] ^ x[1414]);
     layer0_out[3462] <= x[4989];
     layer0_out[3463] <= x[421];
     layer0_out[3464] <= ~x[6494];
     layer0_out[3465] <= x[1675];
     layer0_out[3466] <= ~(x[976] | x[978]);
     layer0_out[3467] <= ~(x[6150] ^ x[6151]);
     layer0_out[3468] <= x[1423] ^ x[1425];
     layer0_out[3469] <= ~(x[4164] & x[4165]);
     layer0_out[3470] <= x[6162] ^ x[6163];
     layer0_out[3471] <= ~(x[4185] & x[4186]);
     layer0_out[3472] <= ~(x[340] | x[341]);
     layer0_out[3473] <= ~(x[4312] | x[4313]);
     layer0_out[3474] <= x[5100] & ~x[5101];
     layer0_out[3475] <= ~(x[4345] & x[4346]);
     layer0_out[3476] <= x[2038] & x[2039];
     layer0_out[3477] <= ~(x[1428] & x[1429]);
     layer0_out[3478] <= 1'b1;
     layer0_out[3479] <= x[7255] ^ x[7256];
     layer0_out[3480] <= x[1751] & x[1752];
     layer0_out[3481] <= ~(x[8122] | x[8123]);
     layer0_out[3482] <= ~(x[4467] ^ x[4468]);
     layer0_out[3483] <= x[176] ^ x[177];
     layer0_out[3484] <= ~x[2622] | x[2620];
     layer0_out[3485] <= x[6908] ^ x[6909];
     layer0_out[3486] <= x[2054] & x[2055];
     layer0_out[3487] <= x[5949] & x[5950];
     layer0_out[3488] <= ~(x[422] & x[424]);
     layer0_out[3489] <= ~(x[6579] | x[6580]);
     layer0_out[3490] <= ~(x[198] ^ x[200]);
     layer0_out[3491] <= ~x[6430] | x[6431];
     layer0_out[3492] <= x[8454] | x[8455];
     layer0_out[3493] <= ~(x[3876] ^ x[3877]);
     layer0_out[3494] <= x[2121] & x[2122];
     layer0_out[3495] <= ~(x[8096] & x[8097]);
     layer0_out[3496] <= x[536] ^ x[537];
     layer0_out[3497] <= ~x[3978];
     layer0_out[3498] <= ~x[2653];
     layer0_out[3499] <= x[4396] & x[4397];
     layer0_out[3500] <= x[4662];
     layer0_out[3501] <= ~(x[3001] & x[3002]);
     layer0_out[3502] <= ~x[5009];
     layer0_out[3503] <= x[5158];
     layer0_out[3504] <= ~x[3873] | x[3872];
     layer0_out[3505] <= ~(x[8766] | x[8767]);
     layer0_out[3506] <= ~(x[5431] & x[5432]);
     layer0_out[3507] <= ~(x[684] ^ x[685]);
     layer0_out[3508] <= x[180];
     layer0_out[3509] <= x[2421] ^ x[2423];
     layer0_out[3510] <= ~(x[687] ^ x[688]);
     layer0_out[3511] <= ~(x[7536] | x[7537]);
     layer0_out[3512] <= ~x[4953];
     layer0_out[3513] <= ~(x[3135] & x[3136]);
     layer0_out[3514] <= ~x[5991];
     layer0_out[3515] <= x[5244] & x[5245];
     layer0_out[3516] <= x[3006] & x[3007];
     layer0_out[3517] <= x[5557] & x[5558];
     layer0_out[3518] <= ~(x[4802] ^ x[4803]);
     layer0_out[3519] <= ~(x[280] ^ x[282]);
     layer0_out[3520] <= x[5982];
     layer0_out[3521] <= ~(x[2694] | x[2696]);
     layer0_out[3522] <= x[6373] & ~x[6374];
     layer0_out[3523] <= ~(x[1811] & x[1812]);
     layer0_out[3524] <= ~x[38];
     layer0_out[3525] <= x[1944] & x[1946];
     layer0_out[3526] <= x[5198] & x[5199];
     layer0_out[3527] <= ~x[1319];
     layer0_out[3528] <= x[255] & x[256];
     layer0_out[3529] <= x[6218] & ~x[6219];
     layer0_out[3530] <= ~x[7323] | x[7324];
     layer0_out[3531] <= x[9000] & x[9001];
     layer0_out[3532] <= 1'b0;
     layer0_out[3533] <= x[331] & ~x[330];
     layer0_out[3534] <= x[3509] & ~x[3510];
     layer0_out[3535] <= x[4265] & x[4266];
     layer0_out[3536] <= ~x[1208];
     layer0_out[3537] <= x[3722] | x[3723];
     layer0_out[3538] <= x[6007] & x[6008];
     layer0_out[3539] <= ~(x[7457] ^ x[7458]);
     layer0_out[3540] <= ~(x[5787] & x[5788]);
     layer0_out[3541] <= ~(x[4092] & x[4093]);
     layer0_out[3542] <= x[1813];
     layer0_out[3543] <= x[1119] & x[1121];
     layer0_out[3544] <= x[8142] ^ x[8143];
     layer0_out[3545] <= 1'b1;
     layer0_out[3546] <= ~(x[6338] | x[6339]);
     layer0_out[3547] <= x[8920] & x[8921];
     layer0_out[3548] <= ~(x[940] & x[941]);
     layer0_out[3549] <= 1'b1;
     layer0_out[3550] <= x[877] | x[878];
     layer0_out[3551] <= ~(x[5935] & x[5936]);
     layer0_out[3552] <= x[5097] & ~x[5096];
     layer0_out[3553] <= 1'b1;
     layer0_out[3554] <= ~(x[1149] & x[1150]);
     layer0_out[3555] <= ~(x[1183] ^ x[1184]);
     layer0_out[3556] <= x[2531] | x[2532];
     layer0_out[3557] <= ~(x[8409] & x[8410]);
     layer0_out[3558] <= ~(x[2837] & x[2838]);
     layer0_out[3559] <= x[2879] & ~x[2878];
     layer0_out[3560] <= x[1340];
     layer0_out[3561] <= x[3063];
     layer0_out[3562] <= ~(x[5305] & x[5306]);
     layer0_out[3563] <= x[3592];
     layer0_out[3564] <= x[5733] & x[5734];
     layer0_out[3565] <= x[3720] | x[3721];
     layer0_out[3566] <= x[1961] | x[1963];
     layer0_out[3567] <= x[511] & x[512];
     layer0_out[3568] <= ~x[230] | x[231];
     layer0_out[3569] <= x[5030] | x[5031];
     layer0_out[3570] <= x[1211] & x[1213];
     layer0_out[3571] <= ~(x[786] & x[788]);
     layer0_out[3572] <= x[108] & ~x[107];
     layer0_out[3573] <= x[2349] ^ x[2351];
     layer0_out[3574] <= ~x[8207];
     layer0_out[3575] <= x[2143] & x[2145];
     layer0_out[3576] <= x[3869];
     layer0_out[3577] <= x[3434];
     layer0_out[3578] <= x[4474] & x[4475];
     layer0_out[3579] <= ~x[8212];
     layer0_out[3580] <= ~x[2900] | x[2901];
     layer0_out[3581] <= x[8278] ^ x[8279];
     layer0_out[3582] <= x[1554] | x[1555];
     layer0_out[3583] <= ~x[1501] | x[1502];
     layer0_out[3584] <= ~(x[2438] & x[2440]);
     layer0_out[3585] <= 1'b0;
     layer0_out[3586] <= ~(x[8713] | x[8714]);
     layer0_out[3587] <= 1'b1;
     layer0_out[3588] <= x[2992] & ~x[2991];
     layer0_out[3589] <= 1'b1;
     layer0_out[3590] <= ~(x[651] ^ x[653]);
     layer0_out[3591] <= x[1352] & x[1354];
     layer0_out[3592] <= ~(x[3494] | x[3495]);
     layer0_out[3593] <= 1'b0;
     layer0_out[3594] <= x[395];
     layer0_out[3595] <= ~x[551];
     layer0_out[3596] <= ~(x[4242] & x[4243]);
     layer0_out[3597] <= ~(x[2321] & x[2322]);
     layer0_out[3598] <= ~(x[1272] & x[1274]);
     layer0_out[3599] <= x[897];
     layer0_out[3600] <= x[5377] | x[5378];
     layer0_out[3601] <= x[6792];
     layer0_out[3602] <= 1'b1;
     layer0_out[3603] <= x[6031] & x[6032];
     layer0_out[3604] <= ~(x[2739] & x[2741]);
     layer0_out[3605] <= ~x[8226];
     layer0_out[3606] <= x[1762] ^ x[1763];
     layer0_out[3607] <= ~x[6140];
     layer0_out[3608] <= x[1397] | x[1398];
     layer0_out[3609] <= ~x[1665];
     layer0_out[3610] <= ~x[5956];
     layer0_out[3611] <= x[1552];
     layer0_out[3612] <= x[5679];
     layer0_out[3613] <= ~(x[2300] & x[2301]);
     layer0_out[3614] <= ~(x[1210] | x[1212]);
     layer0_out[3615] <= x[1781] & x[1782];
     layer0_out[3616] <= x[1037];
     layer0_out[3617] <= ~x[5601];
     layer0_out[3618] <= ~x[3889] | x[3888];
     layer0_out[3619] <= ~x[3340];
     layer0_out[3620] <= x[7056] & x[7057];
     layer0_out[3621] <= x[7379] | x[7380];
     layer0_out[3622] <= x[3973] | x[3974];
     layer0_out[3623] <= ~(x[6185] | x[6186]);
     layer0_out[3624] <= x[302] ^ x[303];
     layer0_out[3625] <= ~x[3209];
     layer0_out[3626] <= ~x[6044];
     layer0_out[3627] <= x[2049];
     layer0_out[3628] <= ~x[2416] | x[2414];
     layer0_out[3629] <= ~(x[1319] & x[1320]);
     layer0_out[3630] <= x[94] | x[96];
     layer0_out[3631] <= 1'b1;
     layer0_out[3632] <= ~(x[2503] | x[2504]);
     layer0_out[3633] <= x[7208] | x[7209];
     layer0_out[3634] <= x[7977] & x[7978];
     layer0_out[3635] <= ~(x[1120] | x[1122]);
     layer0_out[3636] <= ~x[3529];
     layer0_out[3637] <= ~(x[881] | x[883]);
     layer0_out[3638] <= x[5747] & x[5748];
     layer0_out[3639] <= x[337] | x[339];
     layer0_out[3640] <= ~(x[718] & x[719]);
     layer0_out[3641] <= x[1342];
     layer0_out[3642] <= x[1776] | x[1778];
     layer0_out[3643] <= x[2533];
     layer0_out[3644] <= ~x[4990];
     layer0_out[3645] <= x[669] & ~x[671];
     layer0_out[3646] <= x[949] & ~x[951];
     layer0_out[3647] <= 1'b1;
     layer0_out[3648] <= 1'b1;
     layer0_out[3649] <= x[5578] | x[5579];
     layer0_out[3650] <= ~x[2134] | x[2135];
     layer0_out[3651] <= x[7889] & x[7890];
     layer0_out[3652] <= x[226] | x[227];
     layer0_out[3653] <= x[6310] | x[6311];
     layer0_out[3654] <= x[1096] & x[1097];
     layer0_out[3655] <= x[3018] ^ x[3019];
     layer0_out[3656] <= ~(x[6534] | x[6535]);
     layer0_out[3657] <= x[873] & x[875];
     layer0_out[3658] <= x[8100] & ~x[8099];
     layer0_out[3659] <= ~(x[2353] ^ x[2355]);
     layer0_out[3660] <= ~(x[2608] & x[2610]);
     layer0_out[3661] <= x[8203] | x[8204];
     layer0_out[3662] <= ~x[1190] | x[1191];
     layer0_out[3663] <= ~x[323];
     layer0_out[3664] <= x[888];
     layer0_out[3665] <= ~(x[5489] & x[5490]);
     layer0_out[3666] <= ~x[7595];
     layer0_out[3667] <= x[908] & x[910];
     layer0_out[3668] <= ~(x[1859] & x[1860]);
     layer0_out[3669] <= ~(x[7448] | x[7449]);
     layer0_out[3670] <= ~(x[4462] & x[4463]);
     layer0_out[3671] <= ~(x[391] ^ x[392]);
     layer0_out[3672] <= ~(x[1972] | x[1974]);
     layer0_out[3673] <= x[3307] | x[3308];
     layer0_out[3674] <= ~x[8819] | x[8820];
     layer0_out[3675] <= ~(x[1622] | x[1624]);
     layer0_out[3676] <= x[7287] | x[7288];
     layer0_out[3677] <= ~(x[3623] & x[3624]);
     layer0_out[3678] <= ~x[1772];
     layer0_out[3679] <= x[6210];
     layer0_out[3680] <= ~(x[632] ^ x[633]);
     layer0_out[3681] <= x[5587] | x[5588];
     layer0_out[3682] <= ~(x[6030] ^ x[6031]);
     layer0_out[3683] <= x[2161] & x[2162];
     layer0_out[3684] <= x[3322] | x[3323];
     layer0_out[3685] <= ~x[199] | x[200];
     layer0_out[3686] <= 1'b0;
     layer0_out[3687] <= x[7134];
     layer0_out[3688] <= ~x[4801] | x[4802];
     layer0_out[3689] <= 1'b1;
     layer0_out[3690] <= ~(x[8951] & x[8952]);
     layer0_out[3691] <= x[8751] | x[8752];
     layer0_out[3692] <= x[4357] ^ x[4358];
     layer0_out[3693] <= ~(x[576] ^ x[577]);
     layer0_out[3694] <= x[8397] & x[8398];
     layer0_out[3695] <= ~(x[4979] ^ x[4980]);
     layer0_out[3696] <= ~(x[6206] ^ x[6207]);
     layer0_out[3697] <= ~(x[7664] & x[7665]);
     layer0_out[3698] <= x[4376] & x[4377];
     layer0_out[3699] <= ~x[2031];
     layer0_out[3700] <= ~x[7087];
     layer0_out[3701] <= x[1600] | x[1601];
     layer0_out[3702] <= ~x[9124];
     layer0_out[3703] <= x[1719];
     layer0_out[3704] <= ~(x[6109] & x[6110]);
     layer0_out[3705] <= x[1211] ^ x[1212];
     layer0_out[3706] <= ~(x[4817] & x[4818]);
     layer0_out[3707] <= x[3908];
     layer0_out[3708] <= x[4778] | x[4779];
     layer0_out[3709] <= x[2763] | x[2765];
     layer0_out[3710] <= ~(x[7295] & x[7296]);
     layer0_out[3711] <= ~(x[6699] & x[6700]);
     layer0_out[3712] <= 1'b0;
     layer0_out[3713] <= ~(x[6813] ^ x[6814]);
     layer0_out[3714] <= x[6559] & ~x[6558];
     layer0_out[3715] <= ~x[3384];
     layer0_out[3716] <= x[2152] ^ x[2154];
     layer0_out[3717] <= ~x[1117] | x[1119];
     layer0_out[3718] <= x[2286] & ~x[2288];
     layer0_out[3719] <= x[4653];
     layer0_out[3720] <= ~(x[7386] & x[7387]);
     layer0_out[3721] <= x[629] | x[631];
     layer0_out[3722] <= 1'b0;
     layer0_out[3723] <= x[3264] ^ x[3265];
     layer0_out[3724] <= ~x[5276];
     layer0_out[3725] <= ~x[415];
     layer0_out[3726] <= 1'b1;
     layer0_out[3727] <= ~(x[2782] & x[2784]);
     layer0_out[3728] <= x[5288] & x[5289];
     layer0_out[3729] <= x[2191] & x[2192];
     layer0_out[3730] <= x[2479] & x[2481];
     layer0_out[3731] <= ~x[7894] | x[7895];
     layer0_out[3732] <= 1'b0;
     layer0_out[3733] <= 1'b1;
     layer0_out[3734] <= ~(x[7849] | x[7850]);
     layer0_out[3735] <= ~(x[1224] & x[1226]);
     layer0_out[3736] <= x[3525] | x[3526];
     layer0_out[3737] <= x[2403] ^ x[2405];
     layer0_out[3738] <= x[1088] & x[1090];
     layer0_out[3739] <= x[3236] & ~x[3235];
     layer0_out[3740] <= x[2400] & x[2401];
     layer0_out[3741] <= ~x[569] | x[571];
     layer0_out[3742] <= x[8355] & x[8356];
     layer0_out[3743] <= 1'b1;
     layer0_out[3744] <= x[9162] & x[9163];
     layer0_out[3745] <= ~x[6947] | x[6946];
     layer0_out[3746] <= 1'b1;
     layer0_out[3747] <= x[1887] & x[1888];
     layer0_out[3748] <= x[3076] ^ x[3077];
     layer0_out[3749] <= x[817] ^ x[819];
     layer0_out[3750] <= 1'b1;
     layer0_out[3751] <= ~(x[1894] ^ x[1896]);
     layer0_out[3752] <= ~x[267] | x[268];
     layer0_out[3753] <= x[1004] | x[1005];
     layer0_out[3754] <= x[8529] | x[8530];
     layer0_out[3755] <= ~(x[5689] | x[5690]);
     layer0_out[3756] <= ~(x[2026] & x[2027]);
     layer0_out[3757] <= 1'b0;
     layer0_out[3758] <= ~(x[2772] & x[2773]);
     layer0_out[3759] <= ~x[1151] | x[1149];
     layer0_out[3760] <= ~x[1150];
     layer0_out[3761] <= x[6143];
     layer0_out[3762] <= 1'b0;
     layer0_out[3763] <= x[5109] & ~x[5110];
     layer0_out[3764] <= x[2467] & x[2468];
     layer0_out[3765] <= x[2703] & x[2704];
     layer0_out[3766] <= x[952] & x[954];
     layer0_out[3767] <= ~(x[6604] & x[6605]);
     layer0_out[3768] <= x[5592] & x[5593];
     layer0_out[3769] <= x[2196] | x[2197];
     layer0_out[3770] <= ~(x[7531] | x[7532]);
     layer0_out[3771] <= ~(x[5659] & x[5660]);
     layer0_out[3772] <= x[2057] & x[2058];
     layer0_out[3773] <= 1'b1;
     layer0_out[3774] <= x[410] ^ x[412];
     layer0_out[3775] <= ~x[894];
     layer0_out[3776] <= ~(x[5337] & x[5338]);
     layer0_out[3777] <= x[36] & x[38];
     layer0_out[3778] <= ~x[885];
     layer0_out[3779] <= ~(x[3501] ^ x[3502]);
     layer0_out[3780] <= x[8296] & x[8297];
     layer0_out[3781] <= ~(x[2384] & x[2386]);
     layer0_out[3782] <= x[3660] & x[3661];
     layer0_out[3783] <= ~x[7565];
     layer0_out[3784] <= ~(x[1750] & x[1752]);
     layer0_out[3785] <= x[4094] | x[4095];
     layer0_out[3786] <= ~x[8760] | x[8761];
     layer0_out[3787] <= ~(x[2181] | x[2183]);
     layer0_out[3788] <= ~(x[4210] & x[4211]);
     layer0_out[3789] <= x[1151] & x[1153];
     layer0_out[3790] <= ~x[3427] | x[3428];
     layer0_out[3791] <= x[9119] ^ x[9120];
     layer0_out[3792] <= x[4035] | x[4036];
     layer0_out[3793] <= x[593] & x[595];
     layer0_out[3794] <= ~(x[8923] & x[8924]);
     layer0_out[3795] <= x[8803];
     layer0_out[3796] <= ~(x[2085] | x[2086]);
     layer0_out[3797] <= 1'b0;
     layer0_out[3798] <= ~(x[639] & x[640]);
     layer0_out[3799] <= ~x[8628];
     layer0_out[3800] <= ~(x[2324] & x[2326]);
     layer0_out[3801] <= x[1445] & x[1447];
     layer0_out[3802] <= ~(x[1698] & x[1699]);
     layer0_out[3803] <= ~x[598] | x[597];
     layer0_out[3804] <= ~x[5203];
     layer0_out[3805] <= ~(x[4853] | x[4854]);
     layer0_out[3806] <= x[9057] | x[9058];
     layer0_out[3807] <= x[4087] & x[4088];
     layer0_out[3808] <= x[474] & ~x[472];
     layer0_out[3809] <= 1'b1;
     layer0_out[3810] <= x[3773];
     layer0_out[3811] <= ~x[127] | x[129];
     layer0_out[3812] <= ~x[2221] | x[2223];
     layer0_out[3813] <= ~(x[1516] & x[1517]);
     layer0_out[3814] <= x[2487] ^ x[2488];
     layer0_out[3815] <= ~(x[8477] | x[8478]);
     layer0_out[3816] <= ~x[5556];
     layer0_out[3817] <= x[628];
     layer0_out[3818] <= ~(x[8972] & x[8973]);
     layer0_out[3819] <= ~(x[5051] & x[5052]);
     layer0_out[3820] <= x[1747] | x[1749];
     layer0_out[3821] <= ~(x[9039] & x[9040]);
     layer0_out[3822] <= 1'b0;
     layer0_out[3823] <= x[1315] ^ x[1317];
     layer0_out[3824] <= x[2019] & x[2021];
     layer0_out[3825] <= ~x[7933] | x[7934];
     layer0_out[3826] <= x[1082];
     layer0_out[3827] <= ~x[7363] | x[7362];
     layer0_out[3828] <= ~(x[2611] & x[2612]);
     layer0_out[3829] <= x[7538];
     layer0_out[3830] <= ~x[6729];
     layer0_out[3831] <= ~(x[638] ^ x[640]);
     layer0_out[3832] <= ~(x[1928] & x[1929]);
     layer0_out[3833] <= ~(x[3364] & x[3365]);
     layer0_out[3834] <= ~(x[1030] & x[1031]);
     layer0_out[3835] <= ~(x[1342] & x[1344]);
     layer0_out[3836] <= ~(x[4042] | x[4043]);
     layer0_out[3837] <= x[6548] & ~x[6549];
     layer0_out[3838] <= ~(x[4823] | x[4824]);
     layer0_out[3839] <= ~(x[3706] & x[3707]);
     layer0_out[3840] <= 1'b1;
     layer0_out[3841] <= ~(x[3292] | x[3293]);
     layer0_out[3842] <= ~(x[5002] & x[5003]);
     layer0_out[3843] <= x[7237];
     layer0_out[3844] <= ~(x[4294] ^ x[4295]);
     layer0_out[3845] <= x[5660] | x[5661];
     layer0_out[3846] <= x[9147];
     layer0_out[3847] <= x[5599];
     layer0_out[3848] <= x[3281] & x[3282];
     layer0_out[3849] <= ~x[3289];
     layer0_out[3850] <= ~(x[4781] ^ x[4782]);
     layer0_out[3851] <= ~(x[827] | x[828]);
     layer0_out[3852] <= x[5267] & x[5268];
     layer0_out[3853] <= x[6690] ^ x[6691];
     layer0_out[3854] <= ~(x[675] ^ x[677]);
     layer0_out[3855] <= ~(x[6464] | x[6465]);
     layer0_out[3856] <= ~(x[2652] & x[2653]);
     layer0_out[3857] <= x[649] | x[651];
     layer0_out[3858] <= x[8390] | x[8391];
     layer0_out[3859] <= ~(x[6003] & x[6004]);
     layer0_out[3860] <= x[126];
     layer0_out[3861] <= x[2598] & x[2599];
     layer0_out[3862] <= ~(x[1548] & x[1550]);
     layer0_out[3863] <= x[5444];
     layer0_out[3864] <= 1'b0;
     layer0_out[3865] <= ~(x[2836] & x[2837]);
     layer0_out[3866] <= ~(x[1572] & x[1574]);
     layer0_out[3867] <= ~(x[737] & x[739]);
     layer0_out[3868] <= ~x[6251];
     layer0_out[3869] <= ~(x[1258] & x[1259]);
     layer0_out[3870] <= ~x[2748] | x[2750];
     layer0_out[3871] <= x[4504] & x[4505];
     layer0_out[3872] <= ~(x[4634] & x[4635]);
     layer0_out[3873] <= ~(x[8949] | x[8950]);
     layer0_out[3874] <= ~(x[2807] & x[2808]);
     layer0_out[3875] <= ~x[2513];
     layer0_out[3876] <= x[4454];
     layer0_out[3877] <= x[2204] & x[2205];
     layer0_out[3878] <= x[613] & x[614];
     layer0_out[3879] <= ~x[200];
     layer0_out[3880] <= x[719] ^ x[721];
     layer0_out[3881] <= 1'b1;
     layer0_out[3882] <= ~x[8333];
     layer0_out[3883] <= ~x[4015];
     layer0_out[3884] <= x[7639] ^ x[7640];
     layer0_out[3885] <= ~(x[8620] | x[8621]);
     layer0_out[3886] <= ~(x[4670] ^ x[4671]);
     layer0_out[3887] <= x[2874] & x[2875];
     layer0_out[3888] <= x[1407] ^ x[1409];
     layer0_out[3889] <= ~x[6316] | x[6317];
     layer0_out[3890] <= ~(x[6555] | x[6556]);
     layer0_out[3891] <= ~(x[5336] & x[5337]);
     layer0_out[3892] <= ~(x[2023] & x[2025]);
     layer0_out[3893] <= ~(x[2823] & x[2824]);
     layer0_out[3894] <= ~x[8464];
     layer0_out[3895] <= 1'b1;
     layer0_out[3896] <= ~(x[5801] & x[5802]);
     layer0_out[3897] <= ~(x[7373] & x[7374]);
     layer0_out[3898] <= x[4405] & x[4406];
     layer0_out[3899] <= x[2062];
     layer0_out[3900] <= 1'b1;
     layer0_out[3901] <= ~(x[942] | x[943]);
     layer0_out[3902] <= 1'b0;
     layer0_out[3903] <= ~x[2299];
     layer0_out[3904] <= ~x[293] | x[291];
     layer0_out[3905] <= ~(x[3923] & x[3924]);
     layer0_out[3906] <= ~(x[937] | x[939]);
     layer0_out[3907] <= ~(x[2257] & x[2258]);
     layer0_out[3908] <= ~(x[3965] ^ x[3966]);
     layer0_out[3909] <= ~(x[274] | x[275]);
     layer0_out[3910] <= ~x[2536];
     layer0_out[3911] <= x[6922] | x[6923];
     layer0_out[3912] <= ~(x[2478] & x[2480]);
     layer0_out[3913] <= x[3939] ^ x[3940];
     layer0_out[3914] <= x[3789] & x[3790];
     layer0_out[3915] <= x[7846] | x[7847];
     layer0_out[3916] <= x[5834] & x[5835];
     layer0_out[3917] <= ~x[5604];
     layer0_out[3918] <= ~(x[2344] & x[2345]);
     layer0_out[3919] <= x[6562] | x[6563];
     layer0_out[3920] <= ~x[6537];
     layer0_out[3921] <= x[5185] & x[5186];
     layer0_out[3922] <= x[1576] & ~x[1577];
     layer0_out[3923] <= x[1648] ^ x[1649];
     layer0_out[3924] <= x[5540];
     layer0_out[3925] <= ~x[2054] | x[2052];
     layer0_out[3926] <= ~(x[7250] | x[7251]);
     layer0_out[3927] <= ~x[1121] | x[1123];
     layer0_out[3928] <= x[654] & x[656];
     layer0_out[3929] <= ~(x[2721] | x[2723]);
     layer0_out[3930] <= ~(x[674] ^ x[676]);
     layer0_out[3931] <= x[1484] & ~x[1485];
     layer0_out[3932] <= ~x[206];
     layer0_out[3933] <= ~x[8794] | x[8795];
     layer0_out[3934] <= ~(x[459] & x[460]);
     layer0_out[3935] <= ~(x[6070] & x[6071]);
     layer0_out[3936] <= ~x[9084] | x[9083];
     layer0_out[3937] <= ~(x[6208] & x[6209]);
     layer0_out[3938] <= x[5620] & ~x[5619];
     layer0_out[3939] <= ~(x[391] | x[393]);
     layer0_out[3940] <= ~(x[5243] & x[5244]);
     layer0_out[3941] <= 1'b0;
     layer0_out[3942] <= ~(x[5795] & x[5796]);
     layer0_out[3943] <= x[470] | x[472];
     layer0_out[3944] <= x[6295];
     layer0_out[3945] <= ~(x[5373] & x[5374]);
     layer0_out[3946] <= ~x[434];
     layer0_out[3947] <= x[3580] | x[3581];
     layer0_out[3948] <= x[8973] | x[8974];
     layer0_out[3949] <= x[5701];
     layer0_out[3950] <= ~(x[2382] ^ x[2384]);
     layer0_out[3951] <= x[3082];
     layer0_out[3952] <= 1'b0;
     layer0_out[3953] <= x[361] ^ x[362];
     layer0_out[3954] <= x[72] & x[74];
     layer0_out[3955] <= x[2304] & x[2306];
     layer0_out[3956] <= ~(x[2852] & x[2853]);
     layer0_out[3957] <= x[1938] & x[1940];
     layer0_out[3958] <= x[834] & ~x[835];
     layer0_out[3959] <= ~(x[1341] ^ x[1343]);
     layer0_out[3960] <= ~(x[2605] & x[2607]);
     layer0_out[3961] <= x[8382];
     layer0_out[3962] <= x[2063] & x[2065];
     layer0_out[3963] <= x[3603] & x[3604];
     layer0_out[3964] <= x[955];
     layer0_out[3965] <= ~x[1832];
     layer0_out[3966] <= x[1068];
     layer0_out[3967] <= x[2332] & x[2334];
     layer0_out[3968] <= x[473] & ~x[471];
     layer0_out[3969] <= 1'b0;
     layer0_out[3970] <= ~(x[2832] & x[2833]);
     layer0_out[3971] <= ~x[3835];
     layer0_out[3972] <= x[1741] ^ x[1743];
     layer0_out[3973] <= x[4245] | x[4246];
     layer0_out[3974] <= ~(x[2232] & x[2233]);
     layer0_out[3975] <= ~(x[9092] ^ x[9093]);
     layer0_out[3976] <= ~x[1521];
     layer0_out[3977] <= ~x[8231];
     layer0_out[3978] <= ~(x[3033] | x[3034]);
     layer0_out[3979] <= x[241] & x[242];
     layer0_out[3980] <= x[8648] | x[8649];
     layer0_out[3981] <= ~x[6576];
     layer0_out[3982] <= ~(x[1041] & x[1042]);
     layer0_out[3983] <= x[3426];
     layer0_out[3984] <= x[1461];
     layer0_out[3985] <= ~(x[8812] | x[8813]);
     layer0_out[3986] <= x[3519] | x[3520];
     layer0_out[3987] <= 1'b0;
     layer0_out[3988] <= x[596] & x[597];
     layer0_out[3989] <= ~(x[2026] & x[2028]);
     layer0_out[3990] <= ~x[2430];
     layer0_out[3991] <= x[4411] ^ x[4412];
     layer0_out[3992] <= ~(x[7115] | x[7116]);
     layer0_out[3993] <= ~x[8500] | x[8499];
     layer0_out[3994] <= x[2655] | x[2656];
     layer0_out[3995] <= 1'b0;
     layer0_out[3996] <= ~x[5927];
     layer0_out[3997] <= ~x[1298];
     layer0_out[3998] <= x[6940];
     layer0_out[3999] <= x[383] ^ x[384];
     layer0_out[4000] <= x[3060] ^ x[3061];
     layer0_out[4001] <= ~(x[9102] & x[9103]);
     layer0_out[4002] <= ~x[405];
     layer0_out[4003] <= x[8525] | x[8526];
     layer0_out[4004] <= ~(x[498] & x[500]);
     layer0_out[4005] <= x[1279] & x[1280];
     layer0_out[4006] <= x[1447] & x[1448];
     layer0_out[4007] <= ~(x[133] & x[134]);
     layer0_out[4008] <= x[8852] & x[8853];
     layer0_out[4009] <= 1'b0;
     layer0_out[4010] <= ~(x[2114] & x[2116]);
     layer0_out[4011] <= x[5299] & x[5300];
     layer0_out[4012] <= ~x[7428] | x[7429];
     layer0_out[4013] <= x[956] ^ x[957];
     layer0_out[4014] <= ~(x[5671] & x[5672]);
     layer0_out[4015] <= 1'b1;
     layer0_out[4016] <= x[4834] & x[4835];
     layer0_out[4017] <= ~(x[401] ^ x[403]);
     layer0_out[4018] <= ~x[7771] | x[7772];
     layer0_out[4019] <= 1'b0;
     layer0_out[4020] <= ~x[8203];
     layer0_out[4021] <= ~(x[4699] & x[4700]);
     layer0_out[4022] <= ~x[193] | x[195];
     layer0_out[4023] <= ~x[2910];
     layer0_out[4024] <= x[6987] ^ x[6988];
     layer0_out[4025] <= x[409];
     layer0_out[4026] <= ~(x[231] & x[233]);
     layer0_out[4027] <= x[9026] | x[9027];
     layer0_out[4028] <= ~(x[8724] | x[8725]);
     layer0_out[4029] <= x[810] & x[812];
     layer0_out[4030] <= x[1952];
     layer0_out[4031] <= x[6526];
     layer0_out[4032] <= 1'b0;
     layer0_out[4033] <= ~x[7896];
     layer0_out[4034] <= x[3818] | x[3819];
     layer0_out[4035] <= x[1285] ^ x[1287];
     layer0_out[4036] <= x[8988] ^ x[8989];
     layer0_out[4037] <= ~(x[3676] & x[3677]);
     layer0_out[4038] <= x[3455] & ~x[3454];
     layer0_out[4039] <= ~(x[1393] & x[1395]);
     layer0_out[4040] <= ~(x[6895] | x[6896]);
     layer0_out[4041] <= 1'b1;
     layer0_out[4042] <= ~(x[1328] & x[1329]);
     layer0_out[4043] <= 1'b1;
     layer0_out[4044] <= x[4625] & x[4626];
     layer0_out[4045] <= x[5205] & x[5206];
     layer0_out[4046] <= 1'b0;
     layer0_out[4047] <= ~x[4933];
     layer0_out[4048] <= x[2224] & x[2226];
     layer0_out[4049] <= ~(x[209] & x[210]);
     layer0_out[4050] <= ~(x[1873] & x[1874]);
     layer0_out[4051] <= ~(x[1713] & x[1714]);
     layer0_out[4052] <= 1'b0;
     layer0_out[4053] <= ~(x[846] & x[847]);
     layer0_out[4054] <= x[2744] ^ x[2745];
     layer0_out[4055] <= x[2530] | x[2531];
     layer0_out[4056] <= x[4826] | x[4827];
     layer0_out[4057] <= ~(x[3864] | x[3865]);
     layer0_out[4058] <= ~(x[5326] & x[5327]);
     layer0_out[4059] <= x[2075] & x[2076];
     layer0_out[4060] <= x[5520] | x[5521];
     layer0_out[4061] <= ~x[1946];
     layer0_out[4062] <= x[3764] | x[3765];
     layer0_out[4063] <= x[2258] ^ x[2260];
     layer0_out[4064] <= x[1880] & x[1882];
     layer0_out[4065] <= 1'b0;
     layer0_out[4066] <= x[1455] & x[1456];
     layer0_out[4067] <= ~x[8222];
     layer0_out[4068] <= ~(x[6641] & x[6642]);
     layer0_out[4069] <= x[1078] & x[1079];
     layer0_out[4070] <= x[6225] | x[6226];
     layer0_out[4071] <= x[906];
     layer0_out[4072] <= x[1422] & x[1423];
     layer0_out[4073] <= ~x[5050] | x[5051];
     layer0_out[4074] <= ~(x[4985] | x[4986]);
     layer0_out[4075] <= x[22] & ~x[20];
     layer0_out[4076] <= ~(x[3950] | x[3951]);
     layer0_out[4077] <= ~(x[3038] & x[3039]);
     layer0_out[4078] <= ~(x[3719] & x[3720]);
     layer0_out[4079] <= ~(x[3198] & x[3199]);
     layer0_out[4080] <= ~(x[7964] | x[7965]);
     layer0_out[4081] <= ~x[2201];
     layer0_out[4082] <= ~(x[2217] & x[2219]);
     layer0_out[4083] <= x[2508] & x[2510];
     layer0_out[4084] <= x[2087] & ~x[2086];
     layer0_out[4085] <= ~(x[7251] | x[7252]);
     layer0_out[4086] <= x[6260];
     layer0_out[4087] <= x[9178] | x[9179];
     layer0_out[4088] <= x[912] | x[913];
     layer0_out[4089] <= ~(x[7096] | x[7097]);
     layer0_out[4090] <= x[9175] | x[9176];
     layer0_out[4091] <= ~(x[3690] | x[3691]);
     layer0_out[4092] <= ~x[2168];
     layer0_out[4093] <= ~(x[1156] | x[1157]);
     layer0_out[4094] <= ~(x[6797] | x[6798]);
     layer0_out[4095] <= x[3339] & ~x[3338];
     layer0_out[4096] <= x[242] & ~x[240];
     layer0_out[4097] <= ~x[7410];
     layer0_out[4098] <= x[792] & ~x[791];
     layer0_out[4099] <= x[5065];
     layer0_out[4100] <= x[3118] | x[3119];
     layer0_out[4101] <= x[2411] & ~x[2410];
     layer0_out[4102] <= ~(x[5974] & x[5975]);
     layer0_out[4103] <= ~(x[6352] & x[6353]);
     layer0_out[4104] <= x[259] & ~x[260];
     layer0_out[4105] <= x[5304] & x[5305];
     layer0_out[4106] <= x[4076] & x[4077];
     layer0_out[4107] <= ~(x[3312] ^ x[3313]);
     layer0_out[4108] <= x[7136];
     layer0_out[4109] <= ~x[2274];
     layer0_out[4110] <= ~(x[466] & x[467]);
     layer0_out[4111] <= ~x[8876];
     layer0_out[4112] <= x[5121] & x[5122];
     layer0_out[4113] <= x[1010] & ~x[1012];
     layer0_out[4114] <= x[1858] & x[1860];
     layer0_out[4115] <= ~x[371];
     layer0_out[4116] <= ~(x[3756] & x[3757]);
     layer0_out[4117] <= 1'b1;
     layer0_out[4118] <= ~x[1950];
     layer0_out[4119] <= x[103] & x[104];
     layer0_out[4120] <= x[868] & x[869];
     layer0_out[4121] <= ~(x[1070] & x[1072]);
     layer0_out[4122] <= x[1187] & x[1188];
     layer0_out[4123] <= x[7827] | x[7828];
     layer0_out[4124] <= x[5123] & x[5124];
     layer0_out[4125] <= x[1858] | x[1859];
     layer0_out[4126] <= ~(x[725] & x[726]);
     layer0_out[4127] <= ~x[800];
     layer0_out[4128] <= ~(x[1661] ^ x[1663]);
     layer0_out[4129] <= x[9032];
     layer0_out[4130] <= ~x[2699];
     layer0_out[4131] <= x[838] & x[840];
     layer0_out[4132] <= ~(x[2351] & x[2353]);
     layer0_out[4133] <= ~(x[2244] & x[2245]);
     layer0_out[4134] <= x[5083] ^ x[5084];
     layer0_out[4135] <= x[2500] & x[2501];
     layer0_out[4136] <= x[1436] & x[1437];
     layer0_out[4137] <= ~x[6530] | x[6529];
     layer0_out[4138] <= ~x[238];
     layer0_out[4139] <= x[5108] & x[5109];
     layer0_out[4140] <= x[2440] & x[2441];
     layer0_out[4141] <= x[1869] & x[1870];
     layer0_out[4142] <= ~x[2312];
     layer0_out[4143] <= x[9022] & x[9023];
     layer0_out[4144] <= ~(x[8917] & x[8918]);
     layer0_out[4145] <= 1'b1;
     layer0_out[4146] <= ~(x[5223] & x[5224]);
     layer0_out[4147] <= x[735];
     layer0_out[4148] <= x[8316] & x[8317];
     layer0_out[4149] <= ~x[6265];
     layer0_out[4150] <= x[1239] & x[1241];
     layer0_out[4151] <= x[2390] & x[2392];
     layer0_out[4152] <= x[2036] & ~x[2034];
     layer0_out[4153] <= x[657] & x[659];
     layer0_out[4154] <= ~(x[22] ^ x[23]);
     layer0_out[4155] <= ~(x[5189] & x[5190]);
     layer0_out[4156] <= ~x[1181];
     layer0_out[4157] <= ~(x[8779] | x[8780]);
     layer0_out[4158] <= ~(x[6144] | x[6145]);
     layer0_out[4159] <= ~x[35];
     layer0_out[4160] <= x[2123] & ~x[2121];
     layer0_out[4161] <= ~(x[2535] ^ x[2537]);
     layer0_out[4162] <= x[6067] ^ x[6068];
     layer0_out[4163] <= x[8086] & ~x[8085];
     layer0_out[4164] <= x[2356] | x[2358];
     layer0_out[4165] <= 1'b0;
     layer0_out[4166] <= ~x[8245];
     layer0_out[4167] <= x[2016];
     layer0_out[4168] <= x[1614] & x[1615];
     layer0_out[4169] <= ~(x[2674] & x[2676]);
     layer0_out[4170] <= x[2451] & x[2453];
     layer0_out[4171] <= ~(x[704] ^ x[706]);
     layer0_out[4172] <= ~x[5353] | x[5354];
     layer0_out[4173] <= x[713] | x[714];
     layer0_out[4174] <= ~x[8392] | x[8393];
     layer0_out[4175] <= x[1935];
     layer0_out[4176] <= x[6981] & x[6982];
     layer0_out[4177] <= ~(x[1369] & x[1370]);
     layer0_out[4178] <= ~x[490] | x[488];
     layer0_out[4179] <= x[6719];
     layer0_out[4180] <= ~(x[5081] & x[5082]);
     layer0_out[4181] <= x[5352] & x[5353];
     layer0_out[4182] <= 1'b1;
     layer0_out[4183] <= x[3473] & x[3474];
     layer0_out[4184] <= ~x[1176] | x[1174];
     layer0_out[4185] <= x[8480] | x[8481];
     layer0_out[4186] <= ~x[2826] | x[2825];
     layer0_out[4187] <= ~x[267];
     layer0_out[4188] <= ~(x[1706] & x[1707]);
     layer0_out[4189] <= ~(x[7504] | x[7505]);
     layer0_out[4190] <= ~(x[8455] | x[8456]);
     layer0_out[4191] <= ~(x[8767] ^ x[8768]);
     layer0_out[4192] <= ~(x[2326] & x[2328]);
     layer0_out[4193] <= x[5019] | x[5020];
     layer0_out[4194] <= ~x[6254];
     layer0_out[4195] <= x[7755];
     layer0_out[4196] <= ~(x[6737] & x[6738]);
     layer0_out[4197] <= x[9029] & x[9030];
     layer0_out[4198] <= ~(x[8608] & x[8609]);
     layer0_out[4199] <= x[1633] | x[1634];
     layer0_out[4200] <= x[1868] & x[1869];
     layer0_out[4201] <= x[4354] ^ x[4355];
     layer0_out[4202] <= x[2543] & x[2545];
     layer0_out[4203] <= ~(x[3030] ^ x[3031]);
     layer0_out[4204] <= x[438] & ~x[440];
     layer0_out[4205] <= 1'b1;
     layer0_out[4206] <= 1'b0;
     layer0_out[4207] <= ~(x[3090] | x[3091]);
     layer0_out[4208] <= ~x[8953];
     layer0_out[4209] <= ~(x[7870] | x[7871]);
     layer0_out[4210] <= ~(x[7336] ^ x[7337]);
     layer0_out[4211] <= ~(x[7112] & x[7113]);
     layer0_out[4212] <= x[1908] | x[1909];
     layer0_out[4213] <= x[1856] | x[1857];
     layer0_out[4214] <= 1'b1;
     layer0_out[4215] <= x[2269] & x[2270];
     layer0_out[4216] <= ~(x[8241] ^ x[8242]);
     layer0_out[4217] <= x[4872] ^ x[4873];
     layer0_out[4218] <= ~x[3728];
     layer0_out[4219] <= x[1225] & x[1227];
     layer0_out[4220] <= x[3373] | x[3374];
     layer0_out[4221] <= x[9049] ^ x[9050];
     layer0_out[4222] <= ~x[1549] | x[1551];
     layer0_out[4223] <= x[9198] & x[9199];
     layer0_out[4224] <= x[4758] & x[4759];
     layer0_out[4225] <= x[5049] | x[5050];
     layer0_out[4226] <= x[8582] & x[8583];
     layer0_out[4227] <= ~(x[2754] & x[2756]);
     layer0_out[4228] <= x[3709] & x[3710];
     layer0_out[4229] <= ~(x[695] ^ x[697]);
     layer0_out[4230] <= x[8469];
     layer0_out[4231] <= x[2146] & ~x[2145];
     layer0_out[4232] <= x[3621] | x[3622];
     layer0_out[4233] <= x[31] & x[32];
     layer0_out[4234] <= x[102] ^ x[103];
     layer0_out[4235] <= x[4450] & ~x[4449];
     layer0_out[4236] <= ~(x[5977] & x[5978]);
     layer0_out[4237] <= x[6168] | x[6169];
     layer0_out[4238] <= ~(x[4779] & x[4780]);
     layer0_out[4239] <= x[6805] & x[6806];
     layer0_out[4240] <= x[3670] & x[3671];
     layer0_out[4241] <= 1'b1;
     layer0_out[4242] <= ~x[3778];
     layer0_out[4243] <= ~(x[4013] | x[4014]);
     layer0_out[4244] <= x[7070];
     layer0_out[4245] <= ~(x[749] ^ x[751]);
     layer0_out[4246] <= ~(x[741] & x[743]);
     layer0_out[4247] <= x[4258] & x[4259];
     layer0_out[4248] <= ~(x[7463] ^ x[7464]);
     layer0_out[4249] <= ~(x[217] & x[219]);
     layer0_out[4250] <= ~(x[6947] & x[6948]);
     layer0_out[4251] <= ~(x[5874] ^ x[5875]);
     layer0_out[4252] <= x[1494];
     layer0_out[4253] <= x[6870] & x[6871];
     layer0_out[4254] <= 1'b1;
     layer0_out[4255] <= ~(x[7962] & x[7963]);
     layer0_out[4256] <= x[4885] | x[4886];
     layer0_out[4257] <= 1'b1;
     layer0_out[4258] <= x[339];
     layer0_out[4259] <= x[2246];
     layer0_out[4260] <= x[2112] & x[2114];
     layer0_out[4261] <= x[2070];
     layer0_out[4262] <= x[172] & x[173];
     layer0_out[4263] <= x[821] & x[822];
     layer0_out[4264] <= ~x[1429] | x[1430];
     layer0_out[4265] <= ~x[2406];
     layer0_out[4266] <= ~x[6080];
     layer0_out[4267] <= ~(x[820] & x[821]);
     layer0_out[4268] <= x[6615] ^ x[6616];
     layer0_out[4269] <= x[3465] & x[3466];
     layer0_out[4270] <= x[5316] & x[5317];
     layer0_out[4271] <= x[1459];
     layer0_out[4272] <= ~x[4439];
     layer0_out[4273] <= ~(x[759] & x[761]);
     layer0_out[4274] <= x[879] & x[881];
     layer0_out[4275] <= x[2363] & ~x[2364];
     layer0_out[4276] <= ~(x[3624] | x[3625]);
     layer0_out[4277] <= x[245] ^ x[246];
     layer0_out[4278] <= ~x[7236];
     layer0_out[4279] <= ~(x[1013] | x[1015]);
     layer0_out[4280] <= x[4267] & x[4268];
     layer0_out[4281] <= x[2445] ^ x[2447];
     layer0_out[4282] <= ~(x[7553] ^ x[7554]);
     layer0_out[4283] <= x[6200] | x[6201];
     layer0_out[4284] <= ~x[7364];
     layer0_out[4285] <= x[8255] & x[8256];
     layer0_out[4286] <= x[4310] ^ x[4311];
     layer0_out[4287] <= x[9063];
     layer0_out[4288] <= x[4902] | x[4903];
     layer0_out[4289] <= ~x[7356];
     layer0_out[4290] <= x[640] ^ x[642];
     layer0_out[4291] <= x[1663] & x[1665];
     layer0_out[4292] <= x[2498] & x[2500];
     layer0_out[4293] <= x[7760] & x[7761];
     layer0_out[4294] <= x[7381];
     layer0_out[4295] <= ~x[2156];
     layer0_out[4296] <= x[1708] & x[1710];
     layer0_out[4297] <= ~(x[641] ^ x[642]);
     layer0_out[4298] <= ~x[4169] | x[4170];
     layer0_out[4299] <= ~(x[5364] | x[5365]);
     layer0_out[4300] <= x[2294];
     layer0_out[4301] <= ~(x[2037] & x[2039]);
     layer0_out[4302] <= x[186] & ~x[187];
     layer0_out[4303] <= x[86] & x[87];
     layer0_out[4304] <= ~(x[1947] & x[1949]);
     layer0_out[4305] <= x[7072];
     layer0_out[4306] <= ~x[8030];
     layer0_out[4307] <= ~x[550];
     layer0_out[4308] <= ~(x[2307] ^ x[2309]);
     layer0_out[4309] <= ~x[6116] | x[6115];
     layer0_out[4310] <= ~x[3961] | x[3962];
     layer0_out[4311] <= ~x[7019];
     layer0_out[4312] <= ~(x[6415] ^ x[6416]);
     layer0_out[4313] <= ~(x[8511] ^ x[8512]);
     layer0_out[4314] <= x[370] & x[371];
     layer0_out[4315] <= x[98] & x[99];
     layer0_out[4316] <= ~(x[5375] | x[5376]);
     layer0_out[4317] <= ~(x[7579] | x[7580]);
     layer0_out[4318] <= 1'b1;
     layer0_out[4319] <= x[2295] ^ x[2297];
     layer0_out[4320] <= ~(x[8549] | x[8550]);
     layer0_out[4321] <= ~(x[8437] & x[8438]);
     layer0_out[4322] <= ~x[5623];
     layer0_out[4323] <= x[1217] ^ x[1218];
     layer0_out[4324] <= ~x[6487];
     layer0_out[4325] <= ~x[8965];
     layer0_out[4326] <= ~(x[2633] ^ x[2634]);
     layer0_out[4327] <= ~x[6954] | x[6953];
     layer0_out[4328] <= x[1473] & x[1475];
     layer0_out[4329] <= x[7021] ^ x[7022];
     layer0_out[4330] <= x[4452];
     layer0_out[4331] <= ~(x[246] | x[248]);
     layer0_out[4332] <= ~(x[6123] ^ x[6124]);
     layer0_out[4333] <= ~(x[1058] | x[1059]);
     layer0_out[4334] <= x[2062] & x[2063];
     layer0_out[4335] <= 1'b0;
     layer0_out[4336] <= ~(x[2929] & x[2930]);
     layer0_out[4337] <= x[3705] & ~x[3704];
     layer0_out[4338] <= ~(x[1532] & x[1533]);
     layer0_out[4339] <= x[1115];
     layer0_out[4340] <= ~(x[1408] & x[1410]);
     layer0_out[4341] <= x[8909] | x[8910];
     layer0_out[4342] <= x[8189];
     layer0_out[4343] <= x[811] & ~x[813];
     layer0_out[4344] <= ~(x[6086] & x[6087]);
     layer0_out[4345] <= x[1967] ^ x[1969];
     layer0_out[4346] <= ~(x[9035] ^ x[9036]);
     layer0_out[4347] <= ~(x[4784] ^ x[4785]);
     layer0_out[4348] <= ~(x[3573] ^ x[3574]);
     layer0_out[4349] <= x[1449] & ~x[1448];
     layer0_out[4350] <= x[344] & x[346];
     layer0_out[4351] <= ~(x[1228] & x[1230]);
     layer0_out[4352] <= ~(x[2728] & x[2729]);
     layer0_out[4353] <= 1'b0;
     layer0_out[4354] <= ~(x[6733] ^ x[6734]);
     layer0_out[4355] <= ~x[4402] | x[4403];
     layer0_out[4356] <= ~x[15] | x[13];
     layer0_out[4357] <= ~x[1820] | x[1821];
     layer0_out[4358] <= x[2141] & x[2143];
     layer0_out[4359] <= x[782] ^ x[784];
     layer0_out[4360] <= x[1651] | x[1653];
     layer0_out[4361] <= 1'b0;
     layer0_out[4362] <= ~(x[547] | x[548]);
     layer0_out[4363] <= ~(x[3582] ^ x[3583]);
     layer0_out[4364] <= ~x[8788] | x[8789];
     layer0_out[4365] <= ~(x[6845] & x[6846]);
     layer0_out[4366] <= x[1221];
     layer0_out[4367] <= x[3115] & ~x[3116];
     layer0_out[4368] <= x[1550] & x[1552];
     layer0_out[4369] <= x[2646] & ~x[2644];
     layer0_out[4370] <= ~x[2458];
     layer0_out[4371] <= ~(x[5963] & x[5964]);
     layer0_out[4372] <= 1'b0;
     layer0_out[4373] <= x[5003] | x[5004];
     layer0_out[4374] <= 1'b1;
     layer0_out[4375] <= x[1365] & x[1367];
     layer0_out[4376] <= ~x[1696];
     layer0_out[4377] <= ~x[8837];
     layer0_out[4378] <= x[3436] | x[3437];
     layer0_out[4379] <= 1'b1;
     layer0_out[4380] <= x[2998] | x[2999];
     layer0_out[4381] <= ~x[2188];
     layer0_out[4382] <= ~(x[2164] & x[2165]);
     layer0_out[4383] <= x[8244] & x[8245];
     layer0_out[4384] <= ~(x[3353] | x[3354]);
     layer0_out[4385] <= ~(x[1790] & x[1791]);
     layer0_out[4386] <= ~(x[3565] | x[3566]);
     layer0_out[4387] <= x[1530] | x[1531];
     layer0_out[4388] <= x[3293];
     layer0_out[4389] <= x[8254];
     layer0_out[4390] <= x[8238] | x[8239];
     layer0_out[4391] <= ~x[7367];
     layer0_out[4392] <= ~x[7381];
     layer0_out[4393] <= ~(x[2259] & x[2260]);
     layer0_out[4394] <= x[936] | x[937];
     layer0_out[4395] <= 1'b0;
     layer0_out[4396] <= ~(x[1185] & x[1187]);
     layer0_out[4397] <= ~(x[521] | x[522]);
     layer0_out[4398] <= ~(x[4140] | x[4141]);
     layer0_out[4399] <= ~(x[934] | x[936]);
     layer0_out[4400] <= ~(x[5494] & x[5495]);
     layer0_out[4401] <= x[8726] & ~x[8727];
     layer0_out[4402] <= x[8708] & x[8709];
     layer0_out[4403] <= ~(x[8140] & x[8141]);
     layer0_out[4404] <= ~x[9079];
     layer0_out[4405] <= x[796] | x[798];
     layer0_out[4406] <= x[740] ^ x[741];
     layer0_out[4407] <= ~x[2160];
     layer0_out[4408] <= 1'b0;
     layer0_out[4409] <= ~(x[2516] & x[2518]);
     layer0_out[4410] <= x[6344] | x[6345];
     layer0_out[4411] <= ~x[2292] | x[2290];
     layer0_out[4412] <= x[1718];
     layer0_out[4413] <= ~(x[2150] & x[2151]);
     layer0_out[4414] <= ~(x[5467] & x[5468]);
     layer0_out[4415] <= x[6385] ^ x[6386];
     layer0_out[4416] <= ~x[42] | x[43];
     layer0_out[4417] <= x[776] ^ x[778];
     layer0_out[4418] <= 1'b0;
     layer0_out[4419] <= x[5383] & x[5384];
     layer0_out[4420] <= x[221] & x[223];
     layer0_out[4421] <= ~(x[1113] | x[1114]);
     layer0_out[4422] <= ~(x[7489] | x[7490]);
     layer0_out[4423] <= 1'b1;
     layer0_out[4424] <= ~x[7562];
     layer0_out[4425] <= x[7908] & ~x[7909];
     layer0_out[4426] <= x[3329];
     layer0_out[4427] <= ~(x[3105] | x[3106]);
     layer0_out[4428] <= x[6554];
     layer0_out[4429] <= ~(x[3665] | x[3666]);
     layer0_out[4430] <= x[7994] & x[7995];
     layer0_out[4431] <= ~(x[7289] | x[7290]);
     layer0_out[4432] <= 1'b1;
     layer0_out[4433] <= ~(x[6074] & x[6075]);
     layer0_out[4434] <= x[8169] & ~x[8168];
     layer0_out[4435] <= x[765] | x[767];
     layer0_out[4436] <= x[653] | x[654];
     layer0_out[4437] <= x[8186] | x[8187];
     layer0_out[4438] <= ~(x[755] ^ x[757]);
     layer0_out[4439] <= ~x[2940] | x[2939];
     layer0_out[4440] <= ~(x[6479] | x[6480]);
     layer0_out[4441] <= ~(x[2818] & x[2819]);
     layer0_out[4442] <= ~(x[4935] & x[4936]);
     layer0_out[4443] <= ~(x[430] & x[431]);
     layer0_out[4444] <= ~(x[622] & x[623]);
     layer0_out[4445] <= ~(x[7308] | x[7309]);
     layer0_out[4446] <= ~(x[3499] | x[3500]);
     layer0_out[4447] <= ~x[2231];
     layer0_out[4448] <= ~(x[4932] ^ x[4933]);
     layer0_out[4449] <= x[7451];
     layer0_out[4450] <= x[2281] & x[2282];
     layer0_out[4451] <= ~(x[1668] & x[1670]);
     layer0_out[4452] <= x[8754];
     layer0_out[4453] <= ~x[1893];
     layer0_out[4454] <= ~x[6874] | x[6875];
     layer0_out[4455] <= x[3654] ^ x[3655];
     layer0_out[4456] <= x[7033] ^ x[7034];
     layer0_out[4457] <= x[2082] & x[2084];
     layer0_out[4458] <= x[5286] & x[5287];
     layer0_out[4459] <= x[6828] | x[6829];
     layer0_out[4460] <= ~(x[2784] | x[2786]);
     layer0_out[4461] <= x[9190] ^ x[9191];
     layer0_out[4462] <= x[3290] | x[3291];
     layer0_out[4463] <= 1'b1;
     layer0_out[4464] <= x[3244] & x[3245];
     layer0_out[4465] <= x[919] | x[921];
     layer0_out[4466] <= ~(x[33] & x[35]);
     layer0_out[4467] <= ~(x[1380] ^ x[1381]);
     layer0_out[4468] <= ~(x[8165] & x[8166]);
     layer0_out[4469] <= x[4355] ^ x[4356];
     layer0_out[4470] <= x[7217] ^ x[7218];
     layer0_out[4471] <= ~x[6375];
     layer0_out[4472] <= x[7765] | x[7766];
     layer0_out[4473] <= x[8317] & x[8318];
     layer0_out[4474] <= x[553] & x[554];
     layer0_out[4475] <= x[4582] & ~x[4583];
     layer0_out[4476] <= ~(x[703] & x[705]);
     layer0_out[4477] <= x[768];
     layer0_out[4478] <= x[2659] & x[2661];
     layer0_out[4479] <= x[9017];
     layer0_out[4480] <= x[765];
     layer0_out[4481] <= x[4404] | x[4405];
     layer0_out[4482] <= ~x[7161] | x[7160];
     layer0_out[4483] <= x[1646] & x[1648];
     layer0_out[4484] <= ~(x[7140] & x[7141]);
     layer0_out[4485] <= x[5154] & x[5155];
     layer0_out[4486] <= ~(x[7272] ^ x[7273]);
     layer0_out[4487] <= x[929];
     layer0_out[4488] <= x[7869] & ~x[7868];
     layer0_out[4489] <= x[1288] | x[1289];
     layer0_out[4490] <= x[5190] & x[5191];
     layer0_out[4491] <= x[5129] & x[5130];
     layer0_out[4492] <= x[6792] | x[6793];
     layer0_out[4493] <= ~(x[1686] & x[1687]);
     layer0_out[4494] <= x[1994] ^ x[1996];
     layer0_out[4495] <= x[570] ^ x[571];
     layer0_out[4496] <= x[2405] ^ x[2406];
     layer0_out[4497] <= x[8101] & x[8102];
     layer0_out[4498] <= x[6970] ^ x[6971];
     layer0_out[4499] <= ~x[4188];
     layer0_out[4500] <= x[4211] | x[4212];
     layer0_out[4501] <= ~(x[2526] & x[2527]);
     layer0_out[4502] <= x[2736] & x[2738];
     layer0_out[4503] <= ~x[601] | x[600];
     layer0_out[4504] <= ~(x[2321] & x[2323]);
     layer0_out[4505] <= x[2173];
     layer0_out[4506] <= ~(x[4317] | x[4318]);
     layer0_out[4507] <= x[7930];
     layer0_out[4508] <= x[2739] | x[2740];
     layer0_out[4509] <= ~(x[693] | x[695]);
     layer0_out[4510] <= x[589] & x[590];
     layer0_out[4511] <= ~(x[327] | x[329]);
     layer0_out[4512] <= x[2639] ^ x[2640];
     layer0_out[4513] <= ~x[4002];
     layer0_out[4514] <= x[5805] & x[5806];
     layer0_out[4515] <= ~x[1130] | x[1129];
     layer0_out[4516] <= 1'b0;
     layer0_out[4517] <= ~(x[8458] | x[8459]);
     layer0_out[4518] <= ~x[4520];
     layer0_out[4519] <= ~(x[1729] ^ x[1731]);
     layer0_out[4520] <= ~(x[2154] | x[2156]);
     layer0_out[4521] <= ~(x[7201] & x[7202]);
     layer0_out[4522] <= x[2630] ^ x[2631];
     layer0_out[4523] <= x[6841] ^ x[6842];
     layer0_out[4524] <= 1'b1;
     layer0_out[4525] <= x[6056] & x[6057];
     layer0_out[4526] <= ~(x[719] & x[720]);
     layer0_out[4527] <= ~x[4027] | x[4026];
     layer0_out[4528] <= ~x[4992];
     layer0_out[4529] <= x[1135];
     layer0_out[4530] <= x[2948];
     layer0_out[4531] <= x[4390] & x[4391];
     layer0_out[4532] <= ~(x[1364] & x[1366]);
     layer0_out[4533] <= ~x[581];
     layer0_out[4534] <= ~(x[8447] & x[8448]);
     layer0_out[4535] <= x[7524];
     layer0_out[4536] <= 1'b1;
     layer0_out[4537] <= ~(x[8674] | x[8675]);
     layer0_out[4538] <= ~(x[593] ^ x[594]);
     layer0_out[4539] <= x[4429] | x[4430];
     layer0_out[4540] <= x[2771] & x[2773];
     layer0_out[4541] <= 1'b0;
     layer0_out[4542] <= ~(x[7685] ^ x[7686]);
     layer0_out[4543] <= x[4533] ^ x[4534];
     layer0_out[4544] <= ~(x[1658] & x[1659]);
     layer0_out[4545] <= x[8536];
     layer0_out[4546] <= ~x[8979];
     layer0_out[4547] <= x[6108] & x[6109];
     layer0_out[4548] <= x[433] & x[435];
     layer0_out[4549] <= ~(x[1964] | x[1966]);
     layer0_out[4550] <= x[3821] & x[3822];
     layer0_out[4551] <= x[886];
     layer0_out[4552] <= ~(x[8893] | x[8894]);
     layer0_out[4553] <= ~(x[2408] & x[2410]);
     layer0_out[4554] <= ~(x[3072] ^ x[3073]);
     layer0_out[4555] <= x[2770] ^ x[2771];
     layer0_out[4556] <= ~(x[3840] | x[3841]);
     layer0_out[4557] <= x[5665] & x[5666];
     layer0_out[4558] <= ~x[1892];
     layer0_out[4559] <= x[3765] ^ x[3766];
     layer0_out[4560] <= x[5726] & x[5727];
     layer0_out[4561] <= ~x[365] | x[363];
     layer0_out[4562] <= ~x[2698];
     layer0_out[4563] <= ~(x[4852] | x[4853]);
     layer0_out[4564] <= ~(x[2229] ^ x[2231]);
     layer0_out[4565] <= x[1559] ^ x[1560];
     layer0_out[4566] <= x[479] | x[481];
     layer0_out[4567] <= x[816] & x[818];
     layer0_out[4568] <= x[346];
     layer0_out[4569] <= 1'b0;
     layer0_out[4570] <= x[6334] | x[6335];
     layer0_out[4571] <= ~(x[7108] ^ x[7109]);
     layer0_out[4572] <= ~x[1746] | x[1748];
     layer0_out[4573] <= ~(x[1903] | x[1905]);
     layer0_out[4574] <= x[8717];
     layer0_out[4575] <= x[1485];
     layer0_out[4576] <= 1'b1;
     layer0_out[4577] <= ~x[550] | x[552];
     layer0_out[4578] <= 1'b0;
     layer0_out[4579] <= ~(x[4201] & x[4202]);
     layer0_out[4580] <= x[5062] | x[5063];
     layer0_out[4581] <= ~(x[1274] ^ x[1276]);
     layer0_out[4582] <= ~(x[9168] & x[9169]);
     layer0_out[4583] <= 1'b1;
     layer0_out[4584] <= ~(x[3153] ^ x[3154]);
     layer0_out[4585] <= ~(x[6659] ^ x[6660]);
     layer0_out[4586] <= ~x[448] | x[449];
     layer0_out[4587] <= x[1263] & ~x[1265];
     layer0_out[4588] <= ~(x[314] ^ x[316]);
     layer0_out[4589] <= x[8589] | x[8590];
     layer0_out[4590] <= x[802] | x[804];
     layer0_out[4591] <= 1'b1;
     layer0_out[4592] <= ~x[132] | x[133];
     layer0_out[4593] <= ~(x[857] & x[858]);
     layer0_out[4594] <= x[2807] & ~x[2806];
     layer0_out[4595] <= x[7388] | x[7389];
     layer0_out[4596] <= x[408] & ~x[410];
     layer0_out[4597] <= ~(x[801] ^ x[802]);
     layer0_out[4598] <= x[6873] & ~x[6872];
     layer0_out[4599] <= ~(x[2110] & x[2111]);
     layer0_out[4600] <= x[5972] ^ x[5973];
     layer0_out[4601] <= x[2637] & x[2639];
     layer0_out[4602] <= ~(x[8148] ^ x[8149]);
     layer0_out[4603] <= ~x[507];
     layer0_out[4604] <= x[6040] ^ x[6041];
     layer0_out[4605] <= x[3934] | x[3935];
     layer0_out[4606] <= x[4383] & x[4384];
     layer0_out[4607] <= x[4511] & x[4512];
     layer0_out[4608] <= x[4857];
     layer0_out[4609] <= ~(x[476] ^ x[477]);
     layer0_out[4610] <= x[631] ^ x[633];
     layer0_out[4611] <= 1'b0;
     layer0_out[4612] <= ~(x[3884] | x[3885]);
     layer0_out[4613] <= x[3972] | x[3973];
     layer0_out[4614] <= x[5865];
     layer0_out[4615] <= x[3086];
     layer0_out[4616] <= x[8102] | x[8103];
     layer0_out[4617] <= ~(x[8436] ^ x[8437]);
     layer0_out[4618] <= ~(x[4692] | x[4693]);
     layer0_out[4619] <= ~(x[1121] & x[1122]);
     layer0_out[4620] <= ~(x[1635] & x[1636]);
     layer0_out[4621] <= x[6890] ^ x[6891];
     layer0_out[4622] <= x[225] & x[226];
     layer0_out[4623] <= x[8885] ^ x[8886];
     layer0_out[4624] <= 1'b1;
     layer0_out[4625] <= x[2099] & x[2100];
     layer0_out[4626] <= 1'b0;
     layer0_out[4627] <= ~(x[536] & x[538]);
     layer0_out[4628] <= x[7378] | x[7379];
     layer0_out[4629] <= x[4043] | x[4044];
     layer0_out[4630] <= x[1207] ^ x[1209];
     layer0_out[4631] <= ~(x[3715] & x[3716]);
     layer0_out[4632] <= x[1365] & x[1366];
     layer0_out[4633] <= x[1282] & ~x[1280];
     layer0_out[4634] <= ~(x[5478] ^ x[5479]);
     layer0_out[4635] <= x[1116] ^ x[1117];
     layer0_out[4636] <= ~x[2738];
     layer0_out[4637] <= ~(x[7740] ^ x[7741]);
     layer0_out[4638] <= ~(x[1727] & x[1728]);
     layer0_out[4639] <= x[8252] & x[8253];
     layer0_out[4640] <= ~(x[286] | x[288]);
     layer0_out[4641] <= x[7075] ^ x[7076];
     layer0_out[4642] <= ~(x[1579] ^ x[1581]);
     layer0_out[4643] <= ~(x[2647] & x[2649]);
     layer0_out[4644] <= x[1883] & x[1884];
     layer0_out[4645] <= ~(x[8558] | x[8559]);
     layer0_out[4646] <= x[1244] & x[1245];
     layer0_out[4647] <= ~(x[1608] | x[1610]);
     layer0_out[4648] <= 1'b0;
     layer0_out[4649] <= ~(x[1969] & x[1970]);
     layer0_out[4650] <= ~(x[268] | x[270]);
     layer0_out[4651] <= ~(x[109] & x[111]);
     layer0_out[4652] <= ~(x[2389] & x[2390]);
     layer0_out[4653] <= x[945] & x[947];
     layer0_out[4654] <= ~x[6742];
     layer0_out[4655] <= x[8479] ^ x[8480];
     layer0_out[4656] <= x[6809] & x[6810];
     layer0_out[4657] <= x[4727] & x[4728];
     layer0_out[4658] <= ~(x[4125] & x[4126]);
     layer0_out[4659] <= ~x[8270];
     layer0_out[4660] <= ~x[2108];
     layer0_out[4661] <= 1'b1;
     layer0_out[4662] <= ~(x[2510] & x[2512]);
     layer0_out[4663] <= x[5072] & ~x[5071];
     layer0_out[4664] <= x[7159] ^ x[7160];
     layer0_out[4665] <= ~x[4152];
     layer0_out[4666] <= 1'b0;
     layer0_out[4667] <= x[6831];
     layer0_out[4668] <= x[732] ^ x[733];
     layer0_out[4669] <= ~(x[8232] & x[8233]);
     layer0_out[4670] <= x[5161] & x[5162];
     layer0_out[4671] <= x[5542] ^ x[5543];
     layer0_out[4672] <= ~(x[1787] ^ x[1789]);
     layer0_out[4673] <= 1'b0;
     layer0_out[4674] <= x[3913] | x[3914];
     layer0_out[4675] <= ~(x[7883] ^ x[7884]);
     layer0_out[4676] <= ~(x[1754] & x[1755]);
     layer0_out[4677] <= x[1588];
     layer0_out[4678] <= ~x[6350] | x[6349];
     layer0_out[4679] <= x[5671];
     layer0_out[4680] <= x[624] | x[626];
     layer0_out[4681] <= ~(x[406] | x[408]);
     layer0_out[4682] <= ~(x[8927] | x[8928]);
     layer0_out[4683] <= x[7984] | x[7985];
     layer0_out[4684] <= x[5289] & x[5290];
     layer0_out[4685] <= ~(x[2274] & x[2275]);
     layer0_out[4686] <= x[3874] ^ x[3875];
     layer0_out[4687] <= ~(x[1842] & x[1843]);
     layer0_out[4688] <= ~(x[4082] & x[4083]);
     layer0_out[4689] <= x[7196] ^ x[7197];
     layer0_out[4690] <= x[2517] & x[2518];
     layer0_out[4691] <= ~(x[3193] | x[3194]);
     layer0_out[4692] <= x[3134] ^ x[3135];
     layer0_out[4693] <= x[1980] & x[1982];
     layer0_out[4694] <= ~(x[716] | x[717]);
     layer0_out[4695] <= 1'b1;
     layer0_out[4696] <= ~(x[4432] & x[4433]);
     layer0_out[4697] <= x[8995] | x[8996];
     layer0_out[4698] <= x[5355] | x[5356];
     layer0_out[4699] <= x[5026] | x[5027];
     layer0_out[4700] <= ~(x[920] ^ x[922]);
     layer0_out[4701] <= ~(x[3147] & x[3148]);
     layer0_out[4702] <= x[1036];
     layer0_out[4703] <= ~(x[2635] & x[2636]);
     layer0_out[4704] <= x[7602] | x[7603];
     layer0_out[4705] <= x[9140];
     layer0_out[4706] <= ~(x[6105] & x[6106]);
     layer0_out[4707] <= 1'b1;
     layer0_out[4708] <= x[297] & ~x[298];
     layer0_out[4709] <= x[179] ^ x[180];
     layer0_out[4710] <= x[2673];
     layer0_out[4711] <= ~(x[95] | x[96]);
     layer0_out[4712] <= x[5432] & x[5433];
     layer0_out[4713] <= x[5422] | x[5423];
     layer0_out[4714] <= ~x[1937];
     layer0_out[4715] <= ~(x[4251] & x[4252]);
     layer0_out[4716] <= ~(x[119] | x[120]);
     layer0_out[4717] <= ~(x[6626] | x[6627]);
     layer0_out[4718] <= x[2426] | x[2428];
     layer0_out[4719] <= ~x[752];
     layer0_out[4720] <= x[1296] & x[1298];
     layer0_out[4721] <= ~(x[1378] ^ x[1380]);
     layer0_out[4722] <= ~x[8325];
     layer0_out[4723] <= ~(x[7197] & x[7198]);
     layer0_out[4724] <= 1'b1;
     layer0_out[4725] <= x[7997] | x[7998];
     layer0_out[4726] <= x[3173] & ~x[3172];
     layer0_out[4727] <= ~(x[6878] | x[6879]);
     layer0_out[4728] <= x[7952] | x[7953];
     layer0_out[4729] <= ~x[7769] | x[7770];
     layer0_out[4730] <= x[6226] ^ x[6227];
     layer0_out[4731] <= ~x[2125] | x[2123];
     layer0_out[4732] <= ~(x[9152] & x[9153]);
     layer0_out[4733] <= x[3522] ^ x[3523];
     layer0_out[4734] <= ~x[254];
     layer0_out[4735] <= ~(x[1339] & x[1341]);
     layer0_out[4736] <= ~(x[707] & x[708]);
     layer0_out[4737] <= ~(x[2210] & x[2212]);
     layer0_out[4738] <= ~(x[4119] & x[4120]);
     layer0_out[4739] <= x[3518];
     layer0_out[4740] <= x[497] & x[498];
     layer0_out[4741] <= 1'b0;
     layer0_out[4742] <= x[650] ^ x[651];
     layer0_out[4743] <= ~x[2098] | x[2099];
     layer0_out[4744] <= x[265] ^ x[266];
     layer0_out[4745] <= ~(x[853] & x[854]);
     layer0_out[4746] <= x[2399] ^ x[2401];
     layer0_out[4747] <= ~(x[7300] ^ x[7301]);
     layer0_out[4748] <= x[1584] & x[1586];
     layer0_out[4749] <= x[477] & ~x[475];
     layer0_out[4750] <= ~(x[1653] & x[1654]);
     layer0_out[4751] <= ~(x[8134] ^ x[8135]);
     layer0_out[4752] <= ~x[579];
     layer0_out[4753] <= x[6553] & ~x[6554];
     layer0_out[4754] <= ~x[2010];
     layer0_out[4755] <= ~(x[6958] | x[6959]);
     layer0_out[4756] <= 1'b0;
     layer0_out[4757] <= ~(x[5919] | x[5920]);
     layer0_out[4758] <= 1'b1;
     layer0_out[4759] <= ~(x[2778] & x[2779]);
     layer0_out[4760] <= 1'b1;
     layer0_out[4761] <= x[2496] ^ x[2498];
     layer0_out[4762] <= x[823] & x[825];
     layer0_out[4763] <= 1'b0;
     layer0_out[4764] <= x[7688] ^ x[7689];
     layer0_out[4765] <= 1'b1;
     layer0_out[4766] <= ~(x[7465] & x[7466]);
     layer0_out[4767] <= ~(x[4673] | x[4674]);
     layer0_out[4768] <= ~(x[3825] | x[3826]);
     layer0_out[4769] <= x[5000];
     layer0_out[4770] <= ~x[6157];
     layer0_out[4771] <= x[2625] | x[2627];
     layer0_out[4772] <= ~x[2857] | x[2856];
     layer0_out[4773] <= x[228] & ~x[230];
     layer0_out[4774] <= ~(x[1553] & x[1554]);
     layer0_out[4775] <= 1'b1;
     layer0_out[4776] <= x[8749] | x[8750];
     layer0_out[4777] <= x[2196] & x[2198];
     layer0_out[4778] <= x[568] ^ x[570];
     layer0_out[4779] <= x[2262] & x[2264];
     layer0_out[4780] <= ~(x[9155] | x[9156]);
     layer0_out[4781] <= x[922] | x[923];
     layer0_out[4782] <= ~(x[1113] & x[1115]);
     layer0_out[4783] <= x[4269] & x[4270];
     layer0_out[4784] <= ~x[312];
     layer0_out[4785] <= ~(x[8312] | x[8313]);
     layer0_out[4786] <= ~(x[5958] ^ x[5959]);
     layer0_out[4787] <= x[2882];
     layer0_out[4788] <= ~(x[6594] | x[6595]);
     layer0_out[4789] <= ~(x[3791] & x[3792]);
     layer0_out[4790] <= ~(x[1669] & x[1671]);
     layer0_out[4791] <= x[2650] ^ x[2651];
     layer0_out[4792] <= x[5126] & x[5127];
     layer0_out[4793] <= x[5351] & x[5352];
     layer0_out[4794] <= x[991] | x[992];
     layer0_out[4795] <= ~(x[2059] & x[2060]);
     layer0_out[4796] <= x[5440];
     layer0_out[4797] <= ~x[1553];
     layer0_out[4798] <= x[1195] & x[1197];
     layer0_out[4799] <= ~(x[2370] & x[2371]);
     layer0_out[4800] <= x[2621];
     layer0_out[4801] <= x[3234] | x[3235];
     layer0_out[4802] <= ~x[1207] | x[1208];
     layer0_out[4803] <= 1'b1;
     layer0_out[4804] <= x[4263] & x[4264];
     layer0_out[4805] <= ~(x[4115] & x[4116]);
     layer0_out[4806] <= x[1986];
     layer0_out[4807] <= x[9004] | x[9005];
     layer0_out[4808] <= ~x[2000] | x[1999];
     layer0_out[4809] <= ~(x[1613] | x[1614]);
     layer0_out[4810] <= ~(x[2676] & x[2677]);
     layer0_out[4811] <= ~x[2499] | x[2497];
     layer0_out[4812] <= ~(x[742] ^ x[744]);
     layer0_out[4813] <= ~(x[5155] & x[5156]);
     layer0_out[4814] <= ~(x[8596] | x[8597]);
     layer0_out[4815] <= x[5341] | x[5342];
     layer0_out[4816] <= x[1289] & x[1291];
     layer0_out[4817] <= ~(x[437] | x[439]);
     layer0_out[4818] <= ~x[2150];
     layer0_out[4819] <= ~x[3732] | x[3733];
     layer0_out[4820] <= x[7122] | x[7123];
     layer0_out[4821] <= ~(x[5264] & x[5265]);
     layer0_out[4822] <= 1'b1;
     layer0_out[4823] <= x[6592] | x[6593];
     layer0_out[4824] <= ~x[570] | x[569];
     layer0_out[4825] <= x[1683] ^ x[1685];
     layer0_out[4826] <= 1'b1;
     layer0_out[4827] <= x[2911] & x[2912];
     layer0_out[4828] <= x[5278] & x[5279];
     layer0_out[4829] <= ~(x[6975] | x[6976]);
     layer0_out[4830] <= x[6028];
     layer0_out[4831] <= x[7867] & x[7868];
     layer0_out[4832] <= ~(x[825] & x[826]);
     layer0_out[4833] <= ~(x[961] & x[962]);
     layer0_out[4834] <= ~(x[1110] | x[1111]);
     layer0_out[4835] <= x[543] & ~x[541];
     layer0_out[4836] <= x[1301] & ~x[1302];
     layer0_out[4837] <= x[8552] & x[8553];
     layer0_out[4838] <= ~(x[7836] | x[7837]);
     layer0_out[4839] <= ~(x[4170] & x[4171]);
     layer0_out[4840] <= ~(x[2567] | x[2568]);
     layer0_out[4841] <= ~x[8976] | x[8975];
     layer0_out[4842] <= ~(x[1196] ^ x[1198]);
     layer0_out[4843] <= 1'b1;
     layer0_out[4844] <= x[8389] & x[8390];
     layer0_out[4845] <= ~(x[7410] ^ x[7411]);
     layer0_out[4846] <= x[5236] & x[5237];
     layer0_out[4847] <= ~x[1143] | x[1142];
     layer0_out[4848] <= x[5541] & x[5542];
     layer0_out[4849] <= x[3439] | x[3440];
     layer0_out[4850] <= ~x[4798];
     layer0_out[4851] <= ~(x[1679] & x[1681]);
     layer0_out[4852] <= ~(x[3370] & x[3371]);
     layer0_out[4853] <= ~(x[8079] ^ x[8080]);
     layer0_out[4854] <= x[4887] | x[4888];
     layer0_out[4855] <= ~x[4626];
     layer0_out[4856] <= ~x[925] | x[923];
     layer0_out[4857] <= x[4631] & ~x[4632];
     layer0_out[4858] <= x[12] ^ x[13];
     layer0_out[4859] <= x[2018] & x[2020];
     layer0_out[4860] <= ~(x[1466] & x[1467]);
     layer0_out[4861] <= ~(x[1247] & x[1249]);
     layer0_out[4862] <= x[2292] & x[2293];
     layer0_out[4863] <= x[8048] & ~x[8049];
     layer0_out[4864] <= x[3273];
     layer0_out[4865] <= x[7376] & ~x[7375];
     layer0_out[4866] <= x[7632] | x[7633];
     layer0_out[4867] <= x[1173] & x[1175];
     layer0_out[4868] <= ~(x[9179] | x[9180]);
     layer0_out[4869] <= ~(x[3689] | x[3690]);
     layer0_out[4870] <= x[2685] & x[2686];
     layer0_out[4871] <= x[4882] & x[4883];
     layer0_out[4872] <= x[2439] & x[2440];
     layer0_out[4873] <= ~x[1904] | x[1903];
     layer0_out[4874] <= x[3599];
     layer0_out[4875] <= x[6580] | x[6581];
     layer0_out[4876] <= x[6026];
     layer0_out[4877] <= x[4910] | x[4911];
     layer0_out[4878] <= ~(x[6019] | x[6020]);
     layer0_out[4879] <= ~(x[6498] | x[6499]);
     layer0_out[4880] <= ~(x[1968] | x[1969]);
     layer0_out[4881] <= ~(x[8536] ^ x[8537]);
     layer0_out[4882] <= x[3481] ^ x[3482];
     layer0_out[4883] <= ~x[1647] | x[1648];
     layer0_out[4884] <= x[7154] | x[7155];
     layer0_out[4885] <= x[3020] & x[3021];
     layer0_out[4886] <= x[2737] & x[2739];
     layer0_out[4887] <= ~(x[1309] & x[1311]);
     layer0_out[4888] <= ~(x[560] & x[562]);
     layer0_out[4889] <= x[6893] & x[6894];
     layer0_out[4890] <= ~x[1855] | x[1853];
     layer0_out[4891] <= ~(x[1406] ^ x[1408]);
     layer0_out[4892] <= ~(x[2208] | x[2210]);
     layer0_out[4893] <= x[1372] & x[1373];
     layer0_out[4894] <= x[9093] | x[9094];
     layer0_out[4895] <= ~x[7535];
     layer0_out[4896] <= x[6135] & x[6136];
     layer0_out[4897] <= ~x[2570] | x[2571];
     layer0_out[4898] <= 1'b1;
     layer0_out[4899] <= x[5424];
     layer0_out[4900] <= ~(x[2383] & x[2384]);
     layer0_out[4901] <= x[4349];
     layer0_out[4902] <= ~(x[4827] & x[4828]);
     layer0_out[4903] <= x[628] & x[630];
     layer0_out[4904] <= x[4508] & ~x[4509];
     layer0_out[4905] <= x[6954] | x[6955];
     layer0_out[4906] <= x[191] & x[193];
     layer0_out[4907] <= ~(x[7337] | x[7338]);
     layer0_out[4908] <= ~(x[4870] | x[4871]);
     layer0_out[4909] <= 1'b0;
     layer0_out[4910] <= ~(x[9031] ^ x[9032]);
     layer0_out[4911] <= x[4721] | x[4722];
     layer0_out[4912] <= 1'b1;
     layer0_out[4913] <= ~x[6734];
     layer0_out[4914] <= x[5772] & x[5773];
     layer0_out[4915] <= x[6111] & x[6112];
     layer0_out[4916] <= x[4372];
     layer0_out[4917] <= x[3699] & x[3700];
     layer0_out[4918] <= ~x[6214] | x[6213];
     layer0_out[4919] <= x[1670] & x[1671];
     layer0_out[4920] <= ~x[7931];
     layer0_out[4921] <= ~(x[1718] & x[1720]);
     layer0_out[4922] <= x[3553] ^ x[3554];
     layer0_out[4923] <= x[5918];
     layer0_out[4924] <= ~x[1162];
     layer0_out[4925] <= ~x[183] | x[185];
     layer0_out[4926] <= ~(x[603] | x[605]);
     layer0_out[4927] <= ~(x[6927] | x[6928]);
     layer0_out[4928] <= x[1716];
     layer0_out[4929] <= x[2113] & x[2115];
     layer0_out[4930] <= 1'b1;
     layer0_out[4931] <= x[4096];
     layer0_out[4932] <= x[8021] | x[8022];
     layer0_out[4933] <= ~(x[1914] & x[1915]);
     layer0_out[4934] <= 1'b1;
     layer0_out[4935] <= ~x[4009];
     layer0_out[4936] <= ~x[317] | x[315];
     layer0_out[4937] <= ~(x[1261] & x[1262]);
     layer0_out[4938] <= ~(x[875] & x[877]);
     layer0_out[4939] <= 1'b0;
     layer0_out[4940] <= x[7292] & x[7293];
     layer0_out[4941] <= x[1470] ^ x[1472];
     layer0_out[4942] <= ~(x[4491] ^ x[4492]);
     layer0_out[4943] <= ~x[5294];
     layer0_out[4944] <= x[8438] | x[8439];
     layer0_out[4945] <= ~(x[1793] & x[1794]);
     layer0_out[4946] <= ~(x[2652] & x[2654]);
     layer0_out[4947] <= ~x[870];
     layer0_out[4948] <= x[638] | x[639];
     layer0_out[4949] <= 1'b0;
     layer0_out[4950] <= ~(x[1973] & x[1974]);
     layer0_out[4951] <= x[4234] & ~x[4235];
     layer0_out[4952] <= ~(x[795] | x[797]);
     layer0_out[4953] <= ~(x[4118] | x[4119]);
     layer0_out[4954] <= ~(x[5832] & x[5833]);
     layer0_out[4955] <= ~x[6665] | x[6666];
     layer0_out[4956] <= ~(x[6426] | x[6427]);
     layer0_out[4957] <= ~x[1560];
     layer0_out[4958] <= ~(x[1674] | x[1675]);
     layer0_out[4959] <= x[1221] & x[1222];
     layer0_out[4960] <= x[3483] | x[3484];
     layer0_out[4961] <= x[9045];
     layer0_out[4962] <= ~x[3161];
     layer0_out[4963] <= ~(x[1922] | x[1923]);
     layer0_out[4964] <= ~x[1191] | x[1189];
     layer0_out[4965] <= ~x[1960];
     layer0_out[4966] <= ~(x[1629] ^ x[1630]);
     layer0_out[4967] <= x[8180] & ~x[8181];
     layer0_out[4968] <= ~(x[320] | x[322]);
     layer0_out[4969] <= ~(x[5425] & x[5426]);
     layer0_out[4970] <= ~(x[7367] & x[7368]);
     layer0_out[4971] <= x[6782] & ~x[6783];
     layer0_out[4972] <= ~x[8341];
     layer0_out[4973] <= ~(x[4956] | x[4957]);
     layer0_out[4974] <= x[169] | x[170];
     layer0_out[4975] <= x[8955] & ~x[8956];
     layer0_out[4976] <= ~(x[4612] & x[4613]);
     layer0_out[4977] <= x[1828];
     layer0_out[4978] <= x[8039] | x[8040];
     layer0_out[4979] <= x[2781] & x[2783];
     layer0_out[4980] <= ~x[3067] | x[3068];
     layer0_out[4981] <= ~x[5708];
     layer0_out[4982] <= x[8243];
     layer0_out[4983] <= ~x[8162];
     layer0_out[4984] <= ~(x[5021] ^ x[5022]);
     layer0_out[4985] <= ~(x[2093] | x[2095]);
     layer0_out[4986] <= ~x[336];
     layer0_out[4987] <= ~(x[2348] & x[2350]);
     layer0_out[4988] <= ~(x[2338] & x[2339]);
     layer0_out[4989] <= x[947] & x[948];
     layer0_out[4990] <= 1'b0;
     layer0_out[4991] <= x[8647] | x[8648];
     layer0_out[4992] <= x[256] ^ x[258];
     layer0_out[4993] <= x[6362] | x[6363];
     layer0_out[4994] <= x[4045] | x[4046];
     layer0_out[4995] <= x[1754] & x[1756];
     layer0_out[4996] <= x[2718];
     layer0_out[4997] <= x[3781] | x[3782];
     layer0_out[4998] <= ~x[46] | x[45];
     layer0_out[4999] <= ~(x[4795] & x[4796]);
     layer0_out[5000] <= x[1940];
     layer0_out[5001] <= ~(x[8320] | x[8321]);
     layer0_out[5002] <= x[2950] & x[2951];
     layer0_out[5003] <= ~x[8730];
     layer0_out[5004] <= x[4812] | x[4813];
     layer0_out[5005] <= x[4433] & x[4434];
     layer0_out[5006] <= x[5338];
     layer0_out[5007] <= ~x[8201];
     layer0_out[5008] <= ~(x[2509] & x[2511]);
     layer0_out[5009] <= ~(x[3653] & x[3654]);
     layer0_out[5010] <= 1'b0;
     layer0_out[5011] <= x[5701] | x[5702];
     layer0_out[5012] <= x[121] ^ x[122];
     layer0_out[5013] <= 1'b0;
     layer0_out[5014] <= ~x[5582];
     layer0_out[5015] <= x[862] & x[863];
     layer0_out[5016] <= ~(x[1477] & x[1478]);
     layer0_out[5017] <= ~(x[6508] | x[6509]);
     layer0_out[5018] <= x[213] & ~x[212];
     layer0_out[5019] <= x[202];
     layer0_out[5020] <= x[1911] & ~x[1913];
     layer0_out[5021] <= x[1860] | x[1861];
     layer0_out[5022] <= ~(x[2007] | x[2009]);
     layer0_out[5023] <= x[5644] | x[5645];
     layer0_out[5024] <= 1'b1;
     layer0_out[5025] <= ~(x[81] | x[82]);
     layer0_out[5026] <= ~(x[7987] | x[7988]);
     layer0_out[5027] <= x[1977] & ~x[1976];
     layer0_out[5028] <= x[4298] & x[4299];
     layer0_out[5029] <= x[635] & x[637];
     layer0_out[5030] <= ~x[3181];
     layer0_out[5031] <= ~x[2099];
     layer0_out[5032] <= x[2918] & x[2919];
     layer0_out[5033] <= x[3335] | x[3336];
     layer0_out[5034] <= 1'b1;
     layer0_out[5035] <= x[2639] & x[2641];
     layer0_out[5036] <= x[7038] & x[7039];
     layer0_out[5037] <= x[2665] & ~x[2666];
     layer0_out[5038] <= ~x[6123];
     layer0_out[5039] <= x[5053] ^ x[5054];
     layer0_out[5040] <= ~(x[2471] & x[2472]);
     layer0_out[5041] <= x[3145] & x[3146];
     layer0_out[5042] <= ~(x[711] & x[712]);
     layer0_out[5043] <= x[2710] & x[2712];
     layer0_out[5044] <= ~(x[2910] | x[2911]);
     layer0_out[5045] <= x[4175] & x[4176];
     layer0_out[5046] <= ~(x[1348] & x[1349]);
     layer0_out[5047] <= ~(x[5472] & x[5473]);
     layer0_out[5048] <= ~(x[788] | x[790]);
     layer0_out[5049] <= ~x[3396] | x[3395];
     layer0_out[5050] <= ~(x[5423] | x[5424]);
     layer0_out[5051] <= ~(x[9043] | x[9044]);
     layer0_out[5052] <= ~x[2381] | x[2383];
     layer0_out[5053] <= ~x[6778];
     layer0_out[5054] <= x[4862] & x[4863];
     layer0_out[5055] <= x[5153];
     layer0_out[5056] <= x[1456] ^ x[1457];
     layer0_out[5057] <= x[2398];
     layer0_out[5058] <= ~(x[2755] & x[2756]);
     layer0_out[5059] <= x[4380] & x[4381];
     layer0_out[5060] <= ~(x[2140] & x[2142]);
     layer0_out[5061] <= x[6861] & x[6862];
     layer0_out[5062] <= x[6934];
     layer0_out[5063] <= x[5493] & x[5494];
     layer0_out[5064] <= 1'b1;
     layer0_out[5065] <= x[842] | x[844];
     layer0_out[5066] <= 1'b1;
     layer0_out[5067] <= x[3823] & x[3824];
     layer0_out[5068] <= x[6702] | x[6703];
     layer0_out[5069] <= 1'b0;
     layer0_out[5070] <= x[433] | x[434];
     layer0_out[5071] <= ~x[1267];
     layer0_out[5072] <= x[4982] | x[4983];
     layer0_out[5073] <= x[4957] & x[4958];
     layer0_out[5074] <= x[1532] & ~x[1530];
     layer0_out[5075] <= ~(x[2001] | x[2002]);
     layer0_out[5076] <= ~(x[1980] ^ x[1981]);
     layer0_out[5077] <= x[8832] | x[8833];
     layer0_out[5078] <= x[2043] & x[2045];
     layer0_out[5079] <= x[4666] & x[4667];
     layer0_out[5080] <= x[7848];
     layer0_out[5081] <= ~(x[1363] & x[1365]);
     layer0_out[5082] <= x[6680] & x[6681];
     layer0_out[5083] <= ~(x[285] & x[287]);
     layer0_out[5084] <= x[1641] & x[1642];
     layer0_out[5085] <= x[2548] ^ x[2550];
     layer0_out[5086] <= x[8078] & x[8079];
     layer0_out[5087] <= x[6839];
     layer0_out[5088] <= x[2425] & x[2427];
     layer0_out[5089] <= 1'b1;
     layer0_out[5090] <= ~(x[5767] | x[5768]);
     layer0_out[5091] <= x[5142] & x[5143];
     layer0_out[5092] <= x[2038] | x[2040];
     layer0_out[5093] <= x[500];
     layer0_out[5094] <= ~(x[6006] | x[6007]);
     layer0_out[5095] <= ~(x[1333] ^ x[1335]);
     layer0_out[5096] <= ~(x[1907] | x[1909]);
     layer0_out[5097] <= 1'b1;
     layer0_out[5098] <= ~(x[4947] | x[4948]);
     layer0_out[5099] <= 1'b0;
     layer0_out[5100] <= ~x[7225];
     layer0_out[5101] <= x[3937] & x[3938];
     layer0_out[5102] <= x[6880] | x[6881];
     layer0_out[5103] <= x[1846] & x[1847];
     layer0_out[5104] <= x[8967];
     layer0_out[5105] <= x[6640] | x[6641];
     layer0_out[5106] <= ~(x[4577] | x[4578]);
     layer0_out[5107] <= ~(x[1139] | x[1140]);
     layer0_out[5108] <= x[8550] | x[8551];
     layer0_out[5109] <= ~x[5200];
     layer0_out[5110] <= ~(x[979] | x[980]);
     layer0_out[5111] <= x[7384];
     layer0_out[5112] <= x[971] ^ x[973];
     layer0_out[5113] <= x[6212] | x[6213];
     layer0_out[5114] <= x[209] & ~x[211];
     layer0_out[5115] <= ~(x[3340] ^ x[3341]);
     layer0_out[5116] <= x[8849];
     layer0_out[5117] <= x[1344] & x[1346];
     layer0_out[5118] <= x[4604] & x[4605];
     layer0_out[5119] <= x[2666] & x[2668];
     layer0_out[5120] <= x[4747] | x[4748];
     layer0_out[5121] <= x[425] & ~x[423];
     layer0_out[5122] <= ~(x[6395] | x[6396]);
     layer0_out[5123] <= x[5125] & x[5126];
     layer0_out[5124] <= x[51] & ~x[53];
     layer0_out[5125] <= x[4466] & x[4467];
     layer0_out[5126] <= ~(x[2749] | x[2751]);
     layer0_out[5127] <= x[1299] & x[1300];
     layer0_out[5128] <= x[480] | x[481];
     layer0_out[5129] <= x[1311] & x[1312];
     layer0_out[5130] <= ~x[7377] | x[7376];
     layer0_out[5131] <= x[2252];
     layer0_out[5132] <= x[1836] & x[1837];
     layer0_out[5133] <= ~(x[6645] | x[6646]);
     layer0_out[5134] <= x[6956];
     layer0_out[5135] <= x[2723] ^ x[2725];
     layer0_out[5136] <= x[5900] & x[5901];
     layer0_out[5137] <= ~(x[738] ^ x[740]);
     layer0_out[5138] <= x[1439];
     layer0_out[5139] <= x[6021] & x[6022];
     layer0_out[5140] <= x[8383];
     layer0_out[5141] <= ~(x[430] & x[432]);
     layer0_out[5142] <= ~x[885];
     layer0_out[5143] <= ~(x[2001] | x[2003]);
     layer0_out[5144] <= ~(x[9013] | x[9014]);
     layer0_out[5145] <= x[1913] & x[1915];
     layer0_out[5146] <= x[6851] ^ x[6852];
     layer0_out[5147] <= x[3822] & x[3823];
     layer0_out[5148] <= x[1636] & x[1637];
     layer0_out[5149] <= ~(x[7625] ^ x[7626]);
     layer0_out[5150] <= ~(x[794] ^ x[796]);
     layer0_out[5151] <= x[7250];
     layer0_out[5152] <= x[5117] & x[5118];
     layer0_out[5153] <= x[2202] & x[2203];
     layer0_out[5154] <= ~(x[3124] ^ x[3125]);
     layer0_out[5155] <= x[8053] & ~x[8052];
     layer0_out[5156] <= x[7834] & ~x[7833];
     layer0_out[5157] <= ~x[2620] | x[2621];
     layer0_out[5158] <= ~(x[2482] & x[2483]);
     layer0_out[5159] <= x[4440] ^ x[4441];
     layer0_out[5160] <= x[939] ^ x[940];
     layer0_out[5161] <= x[839];
     layer0_out[5162] <= x[7877];
     layer0_out[5163] <= x[4515] ^ x[4516];
     layer0_out[5164] <= x[2554];
     layer0_out[5165] <= x[5936] | x[5937];
     layer0_out[5166] <= 1'b1;
     layer0_out[5167] <= ~(x[5720] & x[5721]);
     layer0_out[5168] <= ~x[712];
     layer0_out[5169] <= x[683] | x[684];
     layer0_out[5170] <= ~x[635];
     layer0_out[5171] <= x[184] ^ x[185];
     layer0_out[5172] <= ~(x[5692] | x[5693]);
     layer0_out[5173] <= x[1995];
     layer0_out[5174] <= ~(x[480] ^ x[482]);
     layer0_out[5175] <= x[953] ^ x[955];
     layer0_out[5176] <= x[1310] | x[1312];
     layer0_out[5177] <= ~(x[1792] & x[1793]);
     layer0_out[5178] <= ~(x[6957] ^ x[6958]);
     layer0_out[5179] <= ~(x[2169] & x[2170]);
     layer0_out[5180] <= ~(x[3761] ^ x[3762]);
     layer0_out[5181] <= x[6274] ^ x[6275];
     layer0_out[5182] <= x[3213] | x[3214];
     layer0_out[5183] <= 1'b1;
     layer0_out[5184] <= x[1815] & x[1817];
     layer0_out[5185] <= ~(x[190] | x[192]);
     layer0_out[5186] <= ~x[8957];
     layer0_out[5187] <= ~(x[7252] & x[7253]);
     layer0_out[5188] <= x[3630];
     layer0_out[5189] <= ~x[3698];
     layer0_out[5190] <= ~(x[5517] | x[5518]);
     layer0_out[5191] <= x[5564];
     layer0_out[5192] <= ~(x[358] | x[360]);
     layer0_out[5193] <= ~x[8544];
     layer0_out[5194] <= ~(x[2883] ^ x[2884]);
     layer0_out[5195] <= x[7904] | x[7905];
     layer0_out[5196] <= x[159] & x[160];
     layer0_out[5197] <= 1'b1;
     layer0_out[5198] <= ~(x[1025] ^ x[1027]);
     layer0_out[5199] <= ~(x[512] ^ x[513]);
     layer0_out[5200] <= x[542];
     layer0_out[5201] <= ~(x[7253] ^ x[7254]);
     layer0_out[5202] <= ~(x[2423] & x[2425]);
     layer0_out[5203] <= x[9058] & x[9059];
     layer0_out[5204] <= x[2514] & x[2515];
     layer0_out[5205] <= ~(x[8997] | x[8998]);
     layer0_out[5206] <= ~x[4085] | x[4084];
     layer0_out[5207] <= ~x[4489];
     layer0_out[5208] <= ~x[1187];
     layer0_out[5209] <= ~(x[3981] | x[3982]);
     layer0_out[5210] <= x[129] | x[131];
     layer0_out[5211] <= x[4159] & x[4160];
     layer0_out[5212] <= x[7507];
     layer0_out[5213] <= x[7793] | x[7794];
     layer0_out[5214] <= x[8284] & x[8285];
     layer0_out[5215] <= x[4760];
     layer0_out[5216] <= ~x[3221];
     layer0_out[5217] <= x[8218] | x[8219];
     layer0_out[5218] <= ~(x[90] & x[92]);
     layer0_out[5219] <= ~x[8604];
     layer0_out[5220] <= ~(x[8757] | x[8758]);
     layer0_out[5221] <= ~(x[5134] & x[5135]);
     layer0_out[5222] <= x[1062] & x[1063];
     layer0_out[5223] <= x[8410] & x[8411];
     layer0_out[5224] <= ~(x[6258] | x[6259]);
     layer0_out[5225] <= x[1497] ^ x[1499];
     layer0_out[5226] <= x[6764];
     layer0_out[5227] <= ~(x[5575] & x[5576]);
     layer0_out[5228] <= ~x[3216];
     layer0_out[5229] <= ~(x[386] ^ x[388]);
     layer0_out[5230] <= ~x[4927];
     layer0_out[5231] <= ~(x[469] ^ x[470]);
     layer0_out[5232] <= x[1002] & x[1004];
     layer0_out[5233] <= ~(x[1120] & x[1121]);
     layer0_out[5234] <= x[2100] & x[2101];
     layer0_out[5235] <= ~(x[9200] & x[9201]);
     layer0_out[5236] <= x[1787] | x[1788];
     layer0_out[5237] <= x[1664] ^ x[1666];
     layer0_out[5238] <= x[14];
     layer0_out[5239] <= ~x[638];
     layer0_out[5240] <= x[6066] & x[6067];
     layer0_out[5241] <= ~(x[2708] | x[2709]);
     layer0_out[5242] <= x[1397] & x[1399];
     layer0_out[5243] <= x[7398] & ~x[7399];
     layer0_out[5244] <= ~(x[1897] & x[1898]);
     layer0_out[5245] <= x[1929] & x[1930];
     layer0_out[5246] <= x[720] & x[722];
     layer0_out[5247] <= ~(x[2267] & x[2268]);
     layer0_out[5248] <= ~x[7628] | x[7629];
     layer0_out[5249] <= ~x[579] | x[581];
     layer0_out[5250] <= x[1625];
     layer0_out[5251] <= x[5491];
     layer0_out[5252] <= x[6901];
     layer0_out[5253] <= ~(x[162] | x[164]);
     layer0_out[5254] <= ~(x[9103] | x[9104]);
     layer0_out[5255] <= ~(x[6408] & x[6409]);
     layer0_out[5256] <= x[5280] ^ x[5281];
     layer0_out[5257] <= ~(x[6450] | x[6451]);
     layer0_out[5258] <= x[7230];
     layer0_out[5259] <= ~(x[7168] & x[7169]);
     layer0_out[5260] <= ~(x[5826] | x[5827]);
     layer0_out[5261] <= ~(x[1445] & x[1446]);
     layer0_out[5262] <= ~(x[1392] & x[1394]);
     layer0_out[5263] <= ~(x[3029] & x[3030]);
     layer0_out[5264] <= x[5240] & x[5241];
     layer0_out[5265] <= ~(x[3] | x[5]);
     layer0_out[5266] <= ~(x[6790] & x[6791]);
     layer0_out[5267] <= ~(x[5120] & x[5121]);
     layer0_out[5268] <= 1'b0;
     layer0_out[5269] <= x[5888] | x[5889];
     layer0_out[5270] <= ~(x[815] & x[816]);
     layer0_out[5271] <= x[918] | x[919];
     layer0_out[5272] <= ~x[7449];
     layer0_out[5273] <= ~(x[1580] & x[1581]);
     layer0_out[5274] <= x[9212] & ~x[9213];
     layer0_out[5275] <= x[4679] & ~x[4680];
     layer0_out[5276] <= ~(x[4816] | x[4817]);
     layer0_out[5277] <= 1'b1;
     layer0_out[5278] <= ~(x[6711] | x[6712]);
     layer0_out[5279] <= ~(x[505] & x[506]);
     layer0_out[5280] <= ~x[993];
     layer0_out[5281] <= ~(x[2707] | x[2708]);
     layer0_out[5282] <= ~(x[8977] | x[8978]);
     layer0_out[5283] <= ~x[7504];
     layer0_out[5284] <= x[3855] & x[3856];
     layer0_out[5285] <= ~x[1950];
     layer0_out[5286] <= ~(x[8954] | x[8955]);
     layer0_out[5287] <= x[207] & x[208];
     layer0_out[5288] <= ~(x[2429] | x[2430]);
     layer0_out[5289] <= ~x[4753];
     layer0_out[5290] <= x[2394] | x[2395];
     layer0_out[5291] <= ~(x[3317] ^ x[3318]);
     layer0_out[5292] <= x[2366] & x[2367];
     layer0_out[5293] <= 1'b1;
     layer0_out[5294] <= x[9075] | x[9076];
     layer0_out[5295] <= ~(x[6775] ^ x[6776]);
     layer0_out[5296] <= x[884] & ~x[886];
     layer0_out[5297] <= x[438] | x[439];
     layer0_out[5298] <= x[5862] | x[5863];
     layer0_out[5299] <= x[641] ^ x[643];
     layer0_out[5300] <= x[1426] & x[1428];
     layer0_out[5301] <= x[2078] & x[2079];
     layer0_out[5302] <= x[8935];
     layer0_out[5303] <= ~(x[7993] ^ x[7994]);
     layer0_out[5304] <= x[1786] & x[1787];
     layer0_out[5305] <= x[8089] | x[8090];
     layer0_out[5306] <= x[7184];
     layer0_out[5307] <= x[839] & x[840];
     layer0_out[5308] <= ~x[3472];
     layer0_out[5309] <= x[5419] | x[5420];
     layer0_out[5310] <= ~x[8046] | x[8045];
     layer0_out[5311] <= x[4361] | x[4362];
     layer0_out[5312] <= ~x[6683];
     layer0_out[5313] <= x[2949] | x[2950];
     layer0_out[5314] <= ~(x[1075] ^ x[1076]);
     layer0_out[5315] <= ~x[7032] | x[7031];
     layer0_out[5316] <= ~x[8652] | x[8651];
     layer0_out[5317] <= 1'b1;
     layer0_out[5318] <= x[411] & x[413];
     layer0_out[5319] <= x[125] & x[127];
     layer0_out[5320] <= x[4190] ^ x[4191];
     layer0_out[5321] <= x[8381] | x[8382];
     layer0_out[5322] <= ~(x[4331] & x[4332]);
     layer0_out[5323] <= ~x[3993];
     layer0_out[5324] <= ~(x[1690] & x[1692]);
     layer0_out[5325] <= ~(x[1216] | x[1217]);
     layer0_out[5326] <= ~(x[1098] & x[1100]);
     layer0_out[5327] <= ~x[3093];
     layer0_out[5328] <= x[1431];
     layer0_out[5329] <= ~(x[2699] ^ x[2701]);
     layer0_out[5330] <= x[1796] ^ x[1797];
     layer0_out[5331] <= x[5054] & x[5055];
     layer0_out[5332] <= ~x[6886];
     layer0_out[5333] <= x[3755] & x[3756];
     layer0_out[5334] <= ~x[7961];
     layer0_out[5335] <= 1'b0;
     layer0_out[5336] <= ~(x[7747] & x[7748]);
     layer0_out[5337] <= ~(x[635] ^ x[636]);
     layer0_out[5338] <= ~(x[4152] ^ x[4153]);
     layer0_out[5339] <= x[1821] ^ x[1822];
     layer0_out[5340] <= x[1327];
     layer0_out[5341] <= x[663] & x[664];
     layer0_out[5342] <= x[4027] | x[4028];
     layer0_out[5343] <= x[4875] | x[4876];
     layer0_out[5344] <= x[1042] & x[1044];
     layer0_out[5345] <= ~(x[1936] & x[1937]);
     layer0_out[5346] <= x[8636] & x[8637];
     layer0_out[5347] <= 1'b1;
     layer0_out[5348] <= ~(x[1443] & x[1445]);
     layer0_out[5349] <= 1'b1;
     layer0_out[5350] <= x[5473];
     layer0_out[5351] <= x[3860] ^ x[3861];
     layer0_out[5352] <= ~(x[4033] | x[4034]);
     layer0_out[5353] <= x[3040] & x[3041];
     layer0_out[5354] <= x[4395] & x[4396];
     layer0_out[5355] <= ~(x[959] | x[961]);
     layer0_out[5356] <= ~(x[2997] ^ x[2998]);
     layer0_out[5357] <= x[1755] & x[1756];
     layer0_out[5358] <= ~(x[614] ^ x[616]);
     layer0_out[5359] <= ~(x[7939] & x[7940]);
     layer0_out[5360] <= ~(x[497] & x[499]);
     layer0_out[5361] <= 1'b0;
     layer0_out[5362] <= ~x[2820];
     layer0_out[5363] <= ~(x[1241] & x[1243]);
     layer0_out[5364] <= ~x[8093] | x[8092];
     layer0_out[5365] <= 1'b1;
     layer0_out[5366] <= ~(x[2050] & x[2052]);
     layer0_out[5367] <= x[5968] & x[5969];
     layer0_out[5368] <= 1'b1;
     layer0_out[5369] <= x[7850] & x[7851];
     layer0_out[5370] <= ~x[1753];
     layer0_out[5371] <= x[7674] & ~x[7675];
     layer0_out[5372] <= x[8169] | x[8170];
     layer0_out[5373] <= x[883] | x[884];
     layer0_out[5374] <= x[3178] ^ x[3179];
     layer0_out[5375] <= ~(x[1117] & x[1118]);
     layer0_out[5376] <= ~(x[2465] ^ x[2466]);
     layer0_out[5377] <= x[1140] & x[1141];
     layer0_out[5378] <= ~x[2925];
     layer0_out[5379] <= ~(x[5318] | x[5319]);
     layer0_out[5380] <= ~x[3383];
     layer0_out[5381] <= x[599] & ~x[597];
     layer0_out[5382] <= ~(x[2628] & x[2630]);
     layer0_out[5383] <= x[4203] & x[4204];
     layer0_out[5384] <= 1'b1;
     layer0_out[5385] <= x[5168] & x[5169];
     layer0_out[5386] <= x[1780] & x[1782];
     layer0_out[5387] <= 1'b0;
     layer0_out[5388] <= x[1746] & x[1747];
     layer0_out[5389] <= ~x[207] | x[206];
     layer0_out[5390] <= x[8688] | x[8689];
     layer0_out[5391] <= x[2855] & ~x[2856];
     layer0_out[5392] <= ~x[1876];
     layer0_out[5393] <= x[7766];
     layer0_out[5394] <= x[2429];
     layer0_out[5395] <= ~(x[664] ^ x[666]);
     layer0_out[5396] <= ~(x[3455] | x[3456]);
     layer0_out[5397] <= x[1515];
     layer0_out[5398] <= x[5285] | x[5286];
     layer0_out[5399] <= ~(x[5314] | x[5315]);
     layer0_out[5400] <= ~(x[5438] & x[5439]);
     layer0_out[5401] <= ~(x[1566] ^ x[1567]);
     layer0_out[5402] <= x[3837];
     layer0_out[5403] <= ~x[7264];
     layer0_out[5404] <= x[376] & x[377];
     layer0_out[5405] <= ~(x[6246] | x[6247]);
     layer0_out[5406] <= ~(x[2528] | x[2530]);
     layer0_out[5407] <= ~x[5987] | x[5986];
     layer0_out[5408] <= ~(x[4510] & x[4511]);
     layer0_out[5409] <= ~x[7300];
     layer0_out[5410] <= x[7591] | x[7592];
     layer0_out[5411] <= ~(x[6616] & x[6617]);
     layer0_out[5412] <= ~(x[7472] | x[7473]);
     layer0_out[5413] <= ~(x[1959] | x[1960]);
     layer0_out[5414] <= x[2977] | x[2978];
     layer0_out[5415] <= x[8184] | x[8185];
     layer0_out[5416] <= x[5621] & x[5622];
     layer0_out[5417] <= ~x[6279];
     layer0_out[5418] <= 1'b1;
     layer0_out[5419] <= ~x[1986];
     layer0_out[5420] <= ~(x[743] | x[744]);
     layer0_out[5421] <= ~(x[30] | x[32]);
     layer0_out[5422] <= ~(x[6858] ^ x[6859]);
     layer0_out[5423] <= ~(x[6421] | x[6422]);
     layer0_out[5424] <= 1'b0;
     layer0_out[5425] <= ~x[181] | x[183];
     layer0_out[5426] <= x[914];
     layer0_out[5427] <= x[2640] & x[2641];
     layer0_out[5428] <= x[6888] | x[6889];
     layer0_out[5429] <= ~(x[7157] & x[7158]);
     layer0_out[5430] <= ~(x[7145] & x[7146]);
     layer0_out[5431] <= ~(x[1130] ^ x[1132]);
     layer0_out[5432] <= ~(x[3361] | x[3362]);
     layer0_out[5433] <= x[8258] | x[8259];
     layer0_out[5434] <= ~(x[4831] & x[4832]);
     layer0_out[5435] <= ~x[2361] | x[2359];
     layer0_out[5436] <= ~(x[8630] | x[8631]);
     layer0_out[5437] <= 1'b0;
     layer0_out[5438] <= ~x[4566] | x[4567];
     layer0_out[5439] <= x[6884] ^ x[6885];
     layer0_out[5440] <= 1'b0;
     layer0_out[5441] <= x[2582] ^ x[2584];
     layer0_out[5442] <= ~x[4564] | x[4563];
     layer0_out[5443] <= ~(x[9141] | x[9142]);
     layer0_out[5444] <= ~x[5172];
     layer0_out[5445] <= x[5202] | x[5203];
     layer0_out[5446] <= ~x[8188];
     layer0_out[5447] <= ~x[8965];
     layer0_out[5448] <= x[2019] & x[2020];
     layer0_out[5449] <= x[632] & ~x[631];
     layer0_out[5450] <= x[2784];
     layer0_out[5451] <= x[6196] | x[6197];
     layer0_out[5452] <= ~(x[2752] | x[2754]);
     layer0_out[5453] <= x[577] & x[579];
     layer0_out[5454] <= ~(x[1640] & x[1641]);
     layer0_out[5455] <= x[8691];
     layer0_out[5456] <= ~(x[1875] | x[1876]);
     layer0_out[5457] <= ~x[3865];
     layer0_out[5458] <= x[1502] & x[1504];
     layer0_out[5459] <= x[8641];
     layer0_out[5460] <= x[51] ^ x[52];
     layer0_out[5461] <= ~(x[5106] ^ x[5107]);
     layer0_out[5462] <= 1'b1;
     layer0_out[5463] <= 1'b0;
     layer0_out[5464] <= x[512] & ~x[510];
     layer0_out[5465] <= ~(x[2683] | x[2685]);
     layer0_out[5466] <= ~x[4358] | x[4359];
     layer0_out[5467] <= x[5997] & x[5998];
     layer0_out[5468] <= 1'b0;
     layer0_out[5469] <= x[6786] & x[6787];
     layer0_out[5470] <= x[8673] ^ x[8674];
     layer0_out[5471] <= x[571] & ~x[573];
     layer0_out[5472] <= ~x[2459];
     layer0_out[5473] <= ~(x[334] & x[336]);
     layer0_out[5474] <= ~(x[972] | x[973]);
     layer0_out[5475] <= 1'b1;
     layer0_out[5476] <= ~(x[8539] & x[8540]);
     layer0_out[5477] <= ~(x[745] & x[747]);
     layer0_out[5478] <= x[2797] & x[2798];
     layer0_out[5479] <= x[5841] & x[5842];
     layer0_out[5480] <= ~x[4593] | x[4592];
     layer0_out[5481] <= x[1242];
     layer0_out[5482] <= ~(x[1727] & x[1729]);
     layer0_out[5483] <= ~(x[5697] | x[5698]);
     layer0_out[5484] <= ~(x[2512] & x[2514]);
     layer0_out[5485] <= x[2379] & x[2380];
     layer0_out[5486] <= x[8503] & x[8504];
     layer0_out[5487] <= ~x[1302];
     layer0_out[5488] <= x[2074] | x[2075];
     layer0_out[5489] <= x[1006] | x[1007];
     layer0_out[5490] <= x[7944] | x[7945];
     layer0_out[5491] <= ~x[6758];
     layer0_out[5492] <= ~(x[8044] | x[8045]);
     layer0_out[5493] <= x[2611] ^ x[2613];
     layer0_out[5494] <= x[171] | x[172];
     layer0_out[5495] <= x[4486] & x[4487];
     layer0_out[5496] <= ~x[2019] | x[2018];
     layer0_out[5497] <= ~(x[5163] & x[5164]);
     layer0_out[5498] <= ~(x[1815] | x[1816]);
     layer0_out[5499] <= ~x[3327] | x[3326];
     layer0_out[5500] <= ~(x[6180] | x[6181]);
     layer0_out[5501] <= x[3077];
     layer0_out[5502] <= x[5507] & x[5508];
     layer0_out[5503] <= ~x[7611] | x[7610];
     layer0_out[5504] <= x[1329] & x[1330];
     layer0_out[5505] <= ~x[2733] | x[2735];
     layer0_out[5506] <= ~(x[2094] & x[2096]);
     layer0_out[5507] <= ~(x[855] & x[857]);
     layer0_out[5508] <= ~(x[2871] & x[2872]);
     layer0_out[5509] <= x[750];
     layer0_out[5510] <= ~(x[812] & x[813]);
     layer0_out[5511] <= 1'b0;
     layer0_out[5512] <= ~(x[3944] | x[3945]);
     layer0_out[5513] <= 1'b1;
     layer0_out[5514] <= x[4453] & ~x[4454];
     layer0_out[5515] <= x[3738];
     layer0_out[5516] <= ~x[1919];
     layer0_out[5517] <= ~(x[7724] | x[7725]);
     layer0_out[5518] <= ~x[261];
     layer0_out[5519] <= ~x[6443] | x[6442];
     layer0_out[5520] <= ~x[6343] | x[6344];
     layer0_out[5521] <= ~(x[2268] & x[2270]);
     layer0_out[5522] <= x[4973] | x[4974];
     layer0_out[5523] <= x[2973];
     layer0_out[5524] <= ~(x[5272] & x[5273]);
     layer0_out[5525] <= ~x[6085] | x[6084];
     layer0_out[5526] <= ~(x[4085] | x[4086]);
     layer0_out[5527] <= x[2358] & x[2359];
     layer0_out[5528] <= x[5947] & ~x[5948];
     layer0_out[5529] <= ~x[1248];
     layer0_out[5530] <= ~x[2221];
     layer0_out[5531] <= ~x[6457];
     layer0_out[5532] <= ~x[2920];
     layer0_out[5533] <= ~(x[6301] | x[6302]);
     layer0_out[5534] <= x[4830] | x[4831];
     layer0_out[5535] <= ~(x[1596] ^ x[1598]);
     layer0_out[5536] <= x[2741] ^ x[2743];
     layer0_out[5537] <= x[7885] | x[7886];
     layer0_out[5538] <= ~(x[2643] & x[2644]);
     layer0_out[5539] <= x[9072];
     layer0_out[5540] <= x[900];
     layer0_out[5541] <= ~(x[2114] & x[2115]);
     layer0_out[5542] <= 1'b0;
     layer0_out[5543] <= ~(x[4553] ^ x[4554]);
     layer0_out[5544] <= x[346];
     layer0_out[5545] <= x[4209] ^ x[4210];
     layer0_out[5546] <= x[662] | x[664];
     layer0_out[5547] <= ~x[6878];
     layer0_out[5548] <= ~(x[5859] ^ x[5860]);
     layer0_out[5549] <= ~(x[6020] ^ x[6021]);
     layer0_out[5550] <= x[4324] | x[4325];
     layer0_out[5551] <= ~(x[2762] & x[2764]);
     layer0_out[5552] <= x[6911] & x[6912];
     layer0_out[5553] <= x[663] | x[665];
     layer0_out[5554] <= ~x[7737];
     layer0_out[5555] <= ~(x[8887] | x[8888]);
     layer0_out[5556] <= x[1688];
     layer0_out[5557] <= ~x[3769];
     layer0_out[5558] <= x[5884] | x[5885];
     layer0_out[5559] <= ~x[1424];
     layer0_out[5560] <= x[8258];
     layer0_out[5561] <= ~(x[6726] & x[6727]);
     layer0_out[5562] <= x[8739] ^ x[8740];
     layer0_out[5563] <= x[7712] ^ x[7713];
     layer0_out[5564] <= ~x[7517];
     layer0_out[5565] <= ~(x[6843] ^ x[6844]);
     layer0_out[5566] <= x[5393] & x[5394];
     layer0_out[5567] <= ~x[775] | x[777];
     layer0_out[5568] <= ~(x[2041] & x[2043]);
     layer0_out[5569] <= ~(x[1937] & x[1939]);
     layer0_out[5570] <= x[1073];
     layer0_out[5571] <= x[3847] & ~x[3848];
     layer0_out[5572] <= ~(x[5486] | x[5487]);
     layer0_out[5573] <= ~(x[7780] | x[7781]);
     layer0_out[5574] <= ~(x[1061] | x[1062]);
     layer0_out[5575] <= ~(x[17] & x[18]);
     layer0_out[5576] <= ~(x[735] & x[737]);
     layer0_out[5577] <= ~(x[2996] | x[2997]);
     layer0_out[5578] <= x[5250];
     layer0_out[5579] <= x[2445] ^ x[2446];
     layer0_out[5580] <= x[754] & x[755];
     layer0_out[5581] <= ~x[8668] | x[8669];
     layer0_out[5582] <= ~(x[911] | x[912]);
     layer0_out[5583] <= ~x[2341] | x[2340];
     layer0_out[5584] <= x[740] & x[742];
     layer0_out[5585] <= ~x[2264] | x[2263];
     layer0_out[5586] <= ~(x[7071] | x[7072]);
     layer0_out[5587] <= ~(x[2600] & x[2601]);
     layer0_out[5588] <= 1'b0;
     layer0_out[5589] <= x[8054] & x[8055];
     layer0_out[5590] <= x[6633] | x[6634];
     layer0_out[5591] <= 1'b1;
     layer0_out[5592] <= ~x[1421];
     layer0_out[5593] <= ~x[7918];
     layer0_out[5594] <= x[4686] | x[4687];
     layer0_out[5595] <= x[529] | x[530];
     layer0_out[5596] <= ~(x[9133] ^ x[9134]);
     layer0_out[5597] <= x[2408] & x[2409];
     layer0_out[5598] <= ~x[1988] | x[1989];
     layer0_out[5599] <= ~(x[3948] | x[3949]);
     layer0_out[5600] <= x[5313] & x[5314];
     layer0_out[5601] <= 1'b0;
     layer0_out[5602] <= x[2724] & x[2725];
     layer0_out[5603] <= 1'b0;
     layer0_out[5604] <= x[3935] ^ x[3936];
     layer0_out[5605] <= 1'b0;
     layer0_out[5606] <= 1'b1;
     layer0_out[5607] <= x[1417] | x[1418];
     layer0_out[5608] <= ~(x[1843] & x[1844]);
     layer0_out[5609] <= x[2033] & x[2035];
     layer0_out[5610] <= x[2505] ^ x[2506];
     layer0_out[5611] <= ~(x[4810] ^ x[4811]);
     layer0_out[5612] <= x[76] ^ x[77];
     layer0_out[5613] <= x[2956] & x[2957];
     layer0_out[5614] <= x[4250] ^ x[4251];
     layer0_out[5615] <= ~x[7098];
     layer0_out[5616] <= ~(x[3804] & x[3805]);
     layer0_out[5617] <= x[5916] & x[5917];
     layer0_out[5618] <= ~(x[1138] | x[1140]);
     layer0_out[5619] <= ~(x[6835] ^ x[6836]);
     layer0_out[5620] <= x[6900] ^ x[6901];
     layer0_out[5621] <= x[3315] & x[3316];
     layer0_out[5622] <= x[549] | x[551];
     layer0_out[5623] <= x[180] & ~x[181];
     layer0_out[5624] <= x[3429];
     layer0_out[5625] <= x[9183] | x[9184];
     layer0_out[5626] <= x[5211] & x[5212];
     layer0_out[5627] <= ~(x[3863] ^ x[3864]);
     layer0_out[5628] <= x[8403] & x[8404];
     layer0_out[5629] <= x[8908] | x[8909];
     layer0_out[5630] <= x[744] & x[745];
     layer0_out[5631] <= ~(x[4876] & x[4877]);
     layer0_out[5632] <= ~(x[7797] | x[7798]);
     layer0_out[5633] <= ~(x[5186] & x[5187]);
     layer0_out[5634] <= x[1148] & ~x[1146];
     layer0_out[5635] <= x[5470] & x[5471];
     layer0_out[5636] <= ~(x[108] ^ x[110]);
     layer0_out[5637] <= x[749] ^ x[750];
     layer0_out[5638] <= ~(x[245] & x[247]);
     layer0_out[5639] <= ~x[3547];
     layer0_out[5640] <= 1'b1;
     layer0_out[5641] <= 1'b0;
     layer0_out[5642] <= ~(x[2703] ^ x[2705]);
     layer0_out[5643] <= 1'b1;
     layer0_out[5644] <= ~x[3788];
     layer0_out[5645] <= x[1851] & x[1852];
     layer0_out[5646] <= x[7864] ^ x[7865];
     layer0_out[5647] <= ~(x[5929] & x[5930]);
     layer0_out[5648] <= x[133] & x[135];
     layer0_out[5649] <= ~(x[6380] | x[6381]);
     layer0_out[5650] <= ~(x[4016] & x[4017]);
     layer0_out[5651] <= x[7988] ^ x[7989];
     layer0_out[5652] <= x[8470] | x[8471];
     layer0_out[5653] <= x[4480] ^ x[4481];
     layer0_out[5654] <= ~x[2684];
     layer0_out[5655] <= ~(x[6992] | x[6993]);
     layer0_out[5656] <= ~(x[3559] & x[3560]);
     layer0_out[5657] <= 1'b0;
     layer0_out[5658] <= ~(x[4630] & x[4631]);
     layer0_out[5659] <= x[8867];
     layer0_out[5660] <= x[6405];
     layer0_out[5661] <= x[5037] | x[5038];
     layer0_out[5662] <= 1'b0;
     layer0_out[5663] <= x[8959] ^ x[8960];
     layer0_out[5664] <= 1'b1;
     layer0_out[5665] <= ~(x[3045] & x[3046]);
     layer0_out[5666] <= x[351] & x[352];
     layer0_out[5667] <= x[2251] & x[2252];
     layer0_out[5668] <= 1'b1;
     layer0_out[5669] <= ~(x[8494] | x[8495]);
     layer0_out[5670] <= x[8734];
     layer0_out[5671] <= ~(x[4259] & x[4260]);
     layer0_out[5672] <= ~x[6899];
     layer0_out[5673] <= ~(x[7434] | x[7435]);
     layer0_out[5674] <= ~(x[1132] & x[1134]);
     layer0_out[5675] <= ~(x[1233] & x[1235]);
     layer0_out[5676] <= x[1852] & x[1853];
     layer0_out[5677] <= x[5094] & x[5095];
     layer0_out[5678] <= ~(x[7601] ^ x[7602]);
     layer0_out[5679] <= x[6480] | x[6481];
     layer0_out[5680] <= x[988] | x[989];
     layer0_out[5681] <= ~x[6979];
     layer0_out[5682] <= 1'b0;
     layer0_out[5683] <= ~(x[2173] & x[2174]);
     layer0_out[5684] <= ~x[3900] | x[3899];
     layer0_out[5685] <= ~x[2179];
     layer0_out[5686] <= x[5941] ^ x[5942];
     layer0_out[5687] <= x[1249] & x[1250];
     layer0_out[5688] <= ~(x[5370] & x[5371]);
     layer0_out[5689] <= ~x[4572];
     layer0_out[5690] <= ~(x[110] & x[112]);
     layer0_out[5691] <= ~(x[1421] & x[1422]);
     layer0_out[5692] <= ~(x[5487] | x[5488]);
     layer0_out[5693] <= ~x[4525] | x[4524];
     layer0_out[5694] <= x[3738] & x[3739];
     layer0_out[5695] <= x[2053];
     layer0_out[5696] <= x[5739] & x[5740];
     layer0_out[5697] <= x[7398];
     layer0_out[5698] <= ~(x[3319] & x[3320]);
     layer0_out[5699] <= x[5807];
     layer0_out[5700] <= x[4171] & x[4172];
     layer0_out[5701] <= x[9055] & x[9056];
     layer0_out[5702] <= ~(x[3942] | x[3943]);
     layer0_out[5703] <= x[1619] & ~x[1618];
     layer0_out[5704] <= ~(x[7900] | x[7901]);
     layer0_out[5705] <= 1'b1;
     layer0_out[5706] <= ~x[1996];
     layer0_out[5707] <= x[6815] | x[6816];
     layer0_out[5708] <= ~(x[976] ^ x[977]);
     layer0_out[5709] <= ~(x[5282] ^ x[5283]);
     layer0_out[5710] <= x[2467] ^ x[2469];
     layer0_out[5711] <= x[491] & ~x[490];
     layer0_out[5712] <= x[1338] & x[1339];
     layer0_out[5713] <= ~(x[1930] ^ x[1931]);
     layer0_out[5714] <= ~x[907];
     layer0_out[5715] <= 1'b1;
     layer0_out[5716] <= x[2718];
     layer0_out[5717] <= ~(x[4864] | x[4865]);
     layer0_out[5718] <= ~x[6591] | x[6592];
     layer0_out[5719] <= x[4599];
     layer0_out[5720] <= x[5209];
     layer0_out[5721] <= ~x[9175];
     layer0_out[5722] <= x[3194];
     layer0_out[5723] <= ~(x[3601] ^ x[3602]);
     layer0_out[5724] <= ~x[5399];
     layer0_out[5725] <= ~(x[6964] | x[6965]);
     layer0_out[5726] <= x[583];
     layer0_out[5727] <= x[847] | x[848];
     layer0_out[5728] <= ~(x[440] & x[441]);
     layer0_out[5729] <= ~(x[8157] & x[8158]);
     layer0_out[5730] <= x[1040] ^ x[1042];
     layer0_out[5731] <= x[5148] & x[5149];
     layer0_out[5732] <= ~(x[5617] & x[5618]);
     layer0_out[5733] <= x[5627] & x[5628];
     layer0_out[5734] <= x[8285] | x[8286];
     layer0_out[5735] <= x[1144] ^ x[1145];
     layer0_out[5736] <= x[2477] & x[2478];
     layer0_out[5737] <= x[5277] & x[5278];
     layer0_out[5738] <= ~(x[6194] | x[6195]);
     layer0_out[5739] <= ~x[601];
     layer0_out[5740] <= x[1438] & x[1440];
     layer0_out[5741] <= x[2115];
     layer0_out[5742] <= 1'b0;
     layer0_out[5743] <= ~x[5087] | x[5086];
     layer0_out[5744] <= ~x[633];
     layer0_out[5745] <= x[6612];
     layer0_out[5746] <= ~x[403];
     layer0_out[5747] <= ~(x[1299] & x[1301]);
     layer0_out[5748] <= x[8605] & x[8606];
     layer0_out[5749] <= 1'b1;
     layer0_out[5750] <= ~(x[445] ^ x[446]);
     layer0_out[5751] <= ~x[276];
     layer0_out[5752] <= ~x[7066];
     layer0_out[5753] <= ~x[4312];
     layer0_out[5754] <= ~(x[8598] & x[8599]);
     layer0_out[5755] <= x[6976] | x[6977];
     layer0_out[5756] <= ~(x[2470] & x[2472]);
     layer0_out[5757] <= x[2278] ^ x[2280];
     layer0_out[5758] <= ~x[7697];
     layer0_out[5759] <= ~x[7885] | x[7884];
     layer0_out[5760] <= x[6152] | x[6153];
     layer0_out[5761] <= x[7371] | x[7372];
     layer0_out[5762] <= x[8530] | x[8531];
     layer0_out[5763] <= ~(x[7158] | x[7159]);
     layer0_out[5764] <= ~(x[6755] | x[6756]);
     layer0_out[5765] <= ~(x[5829] & x[5830]);
     layer0_out[5766] <= x[2381];
     layer0_out[5767] <= ~(x[6491] | x[6492]);
     layer0_out[5768] <= x[3744] | x[3745];
     layer0_out[5769] <= ~x[727] | x[725];
     layer0_out[5770] <= x[1201] ^ x[1203];
     layer0_out[5771] <= x[6518] | x[6519];
     layer0_out[5772] <= x[2558];
     layer0_out[5773] <= x[1000];
     layer0_out[5774] <= x[1863] & x[1864];
     layer0_out[5775] <= ~x[1111] | x[1113];
     layer0_out[5776] <= ~(x[642] ^ x[643]);
     layer0_out[5777] <= x[7000] ^ x[7001];
     layer0_out[5778] <= ~(x[2303] & x[2305]);
     layer0_out[5779] <= x[3314];
     layer0_out[5780] <= ~(x[6119] & x[6120]);
     layer0_out[5781] <= x[1731] & x[1733];
     layer0_out[5782] <= ~(x[715] | x[717]);
     layer0_out[5783] <= x[2914];
     layer0_out[5784] <= 1'b1;
     layer0_out[5785] <= x[604] | x[605];
     layer0_out[5786] <= x[8996];
     layer0_out[5787] <= ~(x[7934] | x[7935]);
     layer0_out[5788] <= ~(x[7238] | x[7239]);
     layer0_out[5789] <= x[2404];
     layer0_out[5790] <= ~(x[2064] | x[2065]);
     layer0_out[5791] <= ~(x[836] & x[837]);
     layer0_out[5792] <= ~(x[1243] | x[1245]);
     layer0_out[5793] <= ~(x[3953] ^ x[3954]);
     layer0_out[5794] <= ~(x[605] | x[606]);
     layer0_out[5795] <= x[6820] ^ x[6821];
     layer0_out[5796] <= x[2357] & x[2358];
     layer0_out[5797] <= 1'b1;
     layer0_out[5798] <= x[1395] & x[1396];
     layer0_out[5799] <= x[5029] | x[5030];
     layer0_out[5800] <= x[1777] | x[1778];
     layer0_out[5801] <= x[2796] & ~x[2795];
     layer0_out[5802] <= ~(x[6622] | x[6623]);
     layer0_out[5803] <= ~(x[354] | x[355]);
     layer0_out[5804] <= ~(x[2289] & x[2290]);
     layer0_out[5805] <= x[5620];
     layer0_out[5806] <= x[4128] & x[4129];
     layer0_out[5807] <= ~(x[2986] & x[2987]);
     layer0_out[5808] <= x[4937] ^ x[4938];
     layer0_out[5809] <= ~(x[3109] | x[3110]);
     layer0_out[5810] <= ~(x[2474] ^ x[2476]);
     layer0_out[5811] <= x[2093] | x[2094];
     layer0_out[5812] <= ~(x[4667] & x[4668]);
     layer0_out[5813] <= ~x[1880] | x[1878];
     layer0_out[5814] <= x[1705] & ~x[1707];
     layer0_out[5815] <= x[4805];
     layer0_out[5816] <= x[8971];
     layer0_out[5817] <= ~(x[1768] | x[1769]);
     layer0_out[5818] <= ~(x[2483] & x[2484]);
     layer0_out[5819] <= 1'b1;
     layer0_out[5820] <= x[917] ^ x[918];
     layer0_out[5821] <= ~x[929];
     layer0_out[5822] <= ~(x[6096] ^ x[6097]);
     layer0_out[5823] <= ~(x[1001] & x[1003]);
     layer0_out[5824] <= ~(x[1805] & x[1807]);
     layer0_out[5825] <= ~(x[971] | x[972]);
     layer0_out[5826] <= x[1577] | x[1578];
     layer0_out[5827] <= x[4071] & x[4072];
     layer0_out[5828] <= x[143] | x[145];
     layer0_out[5829] <= x[1391] & x[1392];
     layer0_out[5830] <= 1'b0;
     layer0_out[5831] <= 1'b0;
     layer0_out[5832] <= x[4881] & x[4882];
     layer0_out[5833] <= x[1581] & x[1583];
     layer0_out[5834] <= ~x[468];
     layer0_out[5835] <= x[1290] & x[1291];
     layer0_out[5836] <= ~x[8543] | x[8542];
     layer0_out[5837] <= x[9148] & ~x[9149];
     layer0_out[5838] <= x[731] | x[732];
     layer0_out[5839] <= ~(x[6224] | x[6225]);
     layer0_out[5840] <= ~(x[214] & x[215]);
     layer0_out[5841] <= x[1528] & x[1530];
     layer0_out[5842] <= ~(x[6017] ^ x[6018]);
     layer0_out[5843] <= ~(x[782] & x[783]);
     layer0_out[5844] <= x[1891] & ~x[1893];
     layer0_out[5845] <= x[7542];
     layer0_out[5846] <= ~x[4879];
     layer0_out[5847] <= x[4050];
     layer0_out[5848] <= ~(x[1179] | x[1180]);
     layer0_out[5849] <= 1'b1;
     layer0_out[5850] <= x[1003] | x[1005];
     layer0_out[5851] <= ~x[2696] | x[2695];
     layer0_out[5852] <= ~(x[3203] & x[3204]);
     layer0_out[5853] <= 1'b1;
     layer0_out[5854] <= ~(x[2833] & x[2834]);
     layer0_out[5855] <= ~(x[3504] & x[3505]);
     layer0_out[5856] <= x[7928] ^ x[7929];
     layer0_out[5857] <= ~x[1793];
     layer0_out[5858] <= x[6507] | x[6508];
     layer0_out[5859] <= x[5380] & x[5381];
     layer0_out[5860] <= ~(x[6513] ^ x[6514]);
     layer0_out[5861] <= ~(x[8624] & x[8625]);
     layer0_out[5862] <= x[2268] & x[2269];
     layer0_out[5863] <= ~x[2151];
     layer0_out[5864] <= x[5440] | x[5441];
     layer0_out[5865] <= ~x[8845] | x[8846];
     layer0_out[5866] <= ~x[4562] | x[4561];
     layer0_out[5867] <= ~(x[3391] | x[3392]);
     layer0_out[5868] <= x[706] & ~x[707];
     layer0_out[5869] <= x[1726] ^ x[1728];
     layer0_out[5870] <= x[7302] | x[7303];
     layer0_out[5871] <= ~x[7877];
     layer0_out[5872] <= ~(x[7980] | x[7981]);
     layer0_out[5873] <= ~(x[1991] & x[1993]);
     layer0_out[5874] <= x[6708] | x[6709];
     layer0_out[5875] <= x[5577] & x[5578];
     layer0_out[5876] <= ~x[1854];
     layer0_out[5877] <= x[2935] & x[2936];
     layer0_out[5878] <= ~x[900];
     layer0_out[5879] <= x[8] & ~x[10];
     layer0_out[5880] <= ~(x[5177] | x[5178]);
     layer0_out[5881] <= 1'b1;
     layer0_out[5882] <= 1'b1;
     layer0_out[5883] <= ~(x[522] & x[524]);
     layer0_out[5884] <= x[291] | x[292];
     layer0_out[5885] <= ~(x[1146] ^ x[1147]);
     layer0_out[5886] <= x[187] ^ x[189];
     layer0_out[5887] <= x[4238] & x[4239];
     layer0_out[5888] <= ~x[2228];
     layer0_out[5889] <= ~x[7494];
     layer0_out[5890] <= x[1300] & x[1301];
     layer0_out[5891] <= ~(x[6293] & x[6294]);
     layer0_out[5892] <= 1'b0;
     layer0_out[5893] <= x[880] | x[882];
     layer0_out[5894] <= ~(x[2765] & x[2767]);
     layer0_out[5895] <= x[2879] | x[2880];
     layer0_out[5896] <= ~(x[8555] & x[8556]);
     layer0_out[5897] <= x[1389] | x[1391];
     layer0_out[5898] <= x[3394] | x[3395];
     layer0_out[5899] <= ~(x[63] & x[64]);
     layer0_out[5900] <= ~(x[1871] & x[1873]);
     layer0_out[5901] <= ~x[823];
     layer0_out[5902] <= ~x[8552] | x[8551];
     layer0_out[5903] <= x[7546] | x[7547];
     layer0_out[5904] <= ~(x[1662] & x[1663]);
     layer0_out[5905] <= 1'b0;
     layer0_out[5906] <= x[8882] & ~x[8881];
     layer0_out[5907] <= x[2761] & x[2762];
     layer0_out[5908] <= 1'b0;
     layer0_out[5909] <= ~x[1828] | x[1827];
     layer0_out[5910] <= ~(x[2322] & x[2323]);
     layer0_out[5911] <= ~x[5960];
     layer0_out[5912] <= 1'b0;
     layer0_out[5913] <= x[1682] & x[1683];
     layer0_out[5914] <= x[4685] & x[4686];
     layer0_out[5915] <= x[8830] & ~x[8831];
     layer0_out[5916] <= x[847] ^ x[849];
     layer0_out[5917] <= ~x[9067];
     layer0_out[5918] <= x[8254] | x[8255];
     layer0_out[5919] <= ~(x[2569] ^ x[2570]);
     layer0_out[5920] <= x[2902] ^ x[2903];
     layer0_out[5921] <= ~(x[958] & x[960]);
     layer0_out[5922] <= 1'b1;
     layer0_out[5923] <= x[2144] & x[2146];
     layer0_out[5924] <= x[7775];
     layer0_out[5925] <= ~(x[9] ^ x[10]);
     layer0_out[5926] <= x[1267] & x[1269];
     layer0_out[5927] <= ~(x[1476] & x[1478]);
     layer0_out[5928] <= ~x[496] | x[495];
     layer0_out[5929] <= x[4615] & x[4616];
     layer0_out[5930] <= ~(x[4338] & x[4339]);
     layer0_out[5931] <= ~(x[6854] ^ x[6855]);
     layer0_out[5932] <= x[4643] & x[4644];
     layer0_out[5933] <= x[7037] & ~x[7038];
     layer0_out[5934] <= ~(x[6410] ^ x[6411]);
     layer0_out[5935] <= x[1752] | x[1753];
     layer0_out[5936] <= x[893] | x[894];
     layer0_out[5937] <= x[2419] & x[2421];
     layer0_out[5938] <= x[1311] & x[1313];
     layer0_out[5939] <= x[1955] | x[1957];
     layer0_out[5940] <= x[8947];
     layer0_out[5941] <= ~(x[2527] & x[2528]);
     layer0_out[5942] <= 1'b1;
     layer0_out[5943] <= x[5522];
     layer0_out[5944] <= x[1424] & x[1426];
     layer0_out[5945] <= ~(x[123] ^ x[125]);
     layer0_out[5946] <= x[1375] & x[1376];
     layer0_out[5947] <= ~x[7357] | x[7356];
     layer0_out[5948] <= ~x[1134];
     layer0_out[5949] <= ~(x[1091] & x[1092]);
     layer0_out[5950] <= ~x[7931];
     layer0_out[5951] <= x[5327] & x[5328];
     layer0_out[5952] <= 1'b1;
     layer0_out[5953] <= x[8528] | x[8529];
     layer0_out[5954] <= ~(x[3012] & x[3013]);
     layer0_out[5955] <= x[6599] | x[6600];
     layer0_out[5956] <= ~x[8721] | x[8722];
     layer0_out[5957] <= ~(x[656] | x[657]);
     layer0_out[5958] <= x[5760] & x[5761];
     layer0_out[5959] <= x[2081];
     layer0_out[5960] <= x[1716] & x[1717];
     layer0_out[5961] <= ~(x[5799] ^ x[5800]);
     layer0_out[5962] <= ~x[8444];
     layer0_out[5963] <= ~(x[1374] ^ x[1376]);
     layer0_out[5964] <= ~(x[1480] & x[1481]);
     layer0_out[5965] <= ~x[6517];
     layer0_out[5966] <= x[469] ^ x[471];
     layer0_out[5967] <= x[4052] | x[4053];
     layer0_out[5968] <= ~(x[5034] & x[5035]);
     layer0_out[5969] <= x[4060] & x[4061];
     layer0_out[5970] <= ~(x[7640] ^ x[7641]);
     layer0_out[5971] <= x[9153] & x[9154];
     layer0_out[5972] <= ~x[6383];
     layer0_out[5973] <= x[5042] & x[5043];
     layer0_out[5974] <= ~x[2333] | x[2331];
     layer0_out[5975] <= x[6816] ^ x[6817];
     layer0_out[5976] <= ~(x[1933] & x[1934]);
     layer0_out[5977] <= ~(x[64] & x[65]);
     layer0_out[5978] <= 1'b1;
     layer0_out[5979] <= ~(x[7360] ^ x[7361]);
     layer0_out[5980] <= ~(x[8365] | x[8366]);
     layer0_out[5981] <= x[1191];
     layer0_out[5982] <= x[1560];
     layer0_out[5983] <= ~(x[1942] | x[1944]);
     layer0_out[5984] <= 1'b1;
     layer0_out[5985] <= x[815] & x[817];
     layer0_out[5986] <= 1'b0;
     layer0_out[5987] <= ~(x[6062] & x[6063]);
     layer0_out[5988] <= ~x[1493] | x[1494];
     layer0_out[5989] <= x[4574] ^ x[4575];
     layer0_out[5990] <= ~x[6769] | x[6768];
     layer0_out[5991] <= ~x[323];
     layer0_out[5992] <= x[1732] & x[1734];
     layer0_out[5993] <= x[7496] & ~x[7495];
     layer0_out[5994] <= ~(x[566] ^ x[568]);
     layer0_out[5995] <= ~x[2270] | x[2271];
     layer0_out[5996] <= x[2617] & x[2618];
     layer0_out[5997] <= x[8075];
     layer0_out[5998] <= 1'b0;
     layer0_out[5999] <= x[1545] & ~x[1546];
     layer0_out[6000] <= ~x[203] | x[204];
     layer0_out[6001] <= x[2904] ^ x[2905];
     layer0_out[6002] <= ~x[5555];
     layer0_out[6003] <= x[8190] | x[8191];
     layer0_out[6004] <= x[5183];
     layer0_out[6005] <= ~(x[9161] & x[9162]);
     layer0_out[6006] <= ~x[7619];
     layer0_out[6007] <= ~(x[1238] & x[1239]);
     layer0_out[6008] <= x[1264] & x[1265];
     layer0_out[6009] <= 1'b0;
     layer0_out[6010] <= ~(x[1898] & x[1900]);
     layer0_out[6011] <= ~(x[8915] | x[8916]);
     layer0_out[6012] <= ~(x[8897] & x[8898]);
     layer0_out[6013] <= ~x[3591] | x[3592];
     layer0_out[6014] <= ~(x[1421] & x[1423]);
     layer0_out[6015] <= x[5599] ^ x[5600];
     layer0_out[6016] <= ~(x[6092] | x[6093]);
     layer0_out[6017] <= x[4382] & x[4383];
     layer0_out[6018] <= x[6409] | x[6410];
     layer0_out[6019] <= 1'b1;
     layer0_out[6020] <= ~(x[5093] ^ x[5094]);
     layer0_out[6021] <= ~x[2614] | x[2612];
     layer0_out[6022] <= x[525] & x[527];
     layer0_out[6023] <= ~x[1257];
     layer0_out[6024] <= x[2336];
     layer0_out[6025] <= x[471] & ~x[470];
     layer0_out[6026] <= x[1775] ^ x[1777];
     layer0_out[6027] <= x[4842];
     layer0_out[6028] <= ~x[6296] | x[6297];
     layer0_out[6029] <= ~x[5616];
     layer0_out[6030] <= 1'b0;
     layer0_out[6031] <= x[399] | x[401];
     layer0_out[6032] <= ~x[1927] | x[1925];
     layer0_out[6033] <= ~(x[5279] & x[5280]);
     layer0_out[6034] <= ~x[243];
     layer0_out[6035] <= ~x[5710];
     layer0_out[6036] <= ~(x[1184] & x[1185]);
     layer0_out[6037] <= ~x[6502] | x[6501];
     layer0_out[6038] <= x[3062] ^ x[3063];
     layer0_out[6039] <= ~(x[4341] | x[4342]);
     layer0_out[6040] <= ~(x[106] & x[108]);
     layer0_out[6041] <= ~(x[3378] & x[3379]);
     layer0_out[6042] <= x[1452] | x[1453];
     layer0_out[6043] <= x[5625] & x[5626];
     layer0_out[6044] <= x[78] & ~x[76];
     layer0_out[6045] <= ~(x[1485] ^ x[1486]);
     layer0_out[6046] <= ~(x[2375] ^ x[2377]);
     layer0_out[6047] <= ~x[6937];
     layer0_out[6048] <= ~(x[1849] & x[1851]);
     layer0_out[6049] <= 1'b1;
     layer0_out[6050] <= 1'b1;
     layer0_out[6051] <= ~x[8061];
     layer0_out[6052] <= ~x[5385];
     layer0_out[6053] <= x[8087] ^ x[8088];
     layer0_out[6054] <= ~(x[4286] ^ x[4287]);
     layer0_out[6055] <= ~x[4080];
     layer0_out[6056] <= x[4918] | x[4919];
     layer0_out[6057] <= ~(x[4939] | x[4940]);
     layer0_out[6058] <= x[4374] | x[4375];
     layer0_out[6059] <= ~(x[1495] & x[1496]);
     layer0_out[6060] <= ~(x[4687] & x[4688]);
     layer0_out[6061] <= x[9181];
     layer0_out[6062] <= x[7211] ^ x[7212];
     layer0_out[6063] <= x[4106] & x[4107];
     layer0_out[6064] <= x[6400];
     layer0_out[6065] <= ~(x[1981] | x[1982]);
     layer0_out[6066] <= x[5802] & x[5803];
     layer0_out[6067] <= ~(x[1504] | x[1506]);
     layer0_out[6068] <= ~(x[3257] | x[3258]);
     layer0_out[6069] <= x[7257] & x[7258];
     layer0_out[6070] <= ~(x[8611] | x[8612]);
     layer0_out[6071] <= x[1317] & x[1319];
     layer0_out[6072] <= x[7515] | x[7516];
     layer0_out[6073] <= ~x[4865];
     layer0_out[6074] <= ~(x[2382] & x[2383]);
     layer0_out[6075] <= x[2238] | x[2240];
     layer0_out[6076] <= ~x[2185];
     layer0_out[6077] <= x[8937];
     layer0_out[6078] <= ~x[8587];
     layer0_out[6079] <= x[3300] & ~x[3301];
     layer0_out[6080] <= x[858] & x[859];
     layer0_out[6081] <= ~(x[2039] ^ x[2040]);
     layer0_out[6082] <= ~(x[1965] | x[1967]);
     layer0_out[6083] <= ~(x[5748] & x[5749]);
     layer0_out[6084] <= ~(x[1839] | x[1840]);
     layer0_out[6085] <= ~(x[7219] | x[7220]);
     layer0_out[6086] <= x[2357] & ~x[2355];
     layer0_out[6087] <= ~x[234] | x[236];
     layer0_out[6088] <= ~(x[1540] & x[1541]);
     layer0_out[6089] <= x[4796] ^ x[4797];
     layer0_out[6090] <= ~(x[2908] & x[2909]);
     layer0_out[6091] <= ~(x[6750] ^ x[6751]);
     layer0_out[6092] <= x[2458] ^ x[2460];
     layer0_out[6093] <= 1'b0;
     layer0_out[6094] <= ~(x[2406] & x[2408]);
     layer0_out[6095] <= ~x[1840] | x[1841];
     layer0_out[6096] <= x[8684] | x[8685];
     layer0_out[6097] <= x[1779] | x[1781];
     layer0_out[6098] <= x[6443] | x[6444];
     layer0_out[6099] <= x[16] | x[18];
     layer0_out[6100] <= x[7118] ^ x[7119];
     layer0_out[6101] <= ~x[5058];
     layer0_out[6102] <= x[2012] & x[2013];
     layer0_out[6103] <= x[341] ^ x[342];
     layer0_out[6104] <= x[6232] ^ x[6233];
     layer0_out[6105] <= ~(x[2271] ^ x[2272]);
     layer0_out[6106] <= 1'b1;
     layer0_out[6107] <= ~(x[4202] ^ x[4203]);
     layer0_out[6108] <= ~(x[3785] ^ x[3786]);
     layer0_out[6109] <= x[530];
     layer0_out[6110] <= x[5595] & x[5596];
     layer0_out[6111] <= x[6051] | x[6052];
     layer0_out[6112] <= ~(x[4138] | x[4139]);
     layer0_out[6113] <= ~(x[1480] & x[1482]);
     layer0_out[6114] <= ~(x[4427] | x[4428]);
     layer0_out[6115] <= x[4731];
     layer0_out[6116] <= ~(x[3126] | x[3127]);
     layer0_out[6117] <= ~(x[3742] | x[3743]);
     layer0_out[6118] <= ~(x[3474] & x[3475]);
     layer0_out[6119] <= ~(x[3053] ^ x[3054]);
     layer0_out[6120] <= ~(x[2575] & x[2577]);
     layer0_out[6121] <= x[2543] & x[2544];
     layer0_out[6122] <= x[173] & x[175];
     layer0_out[6123] <= ~(x[5368] & x[5369]);
     layer0_out[6124] <= x[4044] | x[4045];
     layer0_out[6125] <= x[2109] & x[2111];
     layer0_out[6126] <= x[1414] & x[1416];
     layer0_out[6127] <= x[3121] & ~x[3122];
     layer0_out[6128] <= ~(x[2045] & x[2046]);
     layer0_out[6129] <= ~(x[4200] | x[4201]);
     layer0_out[6130] <= x[4703] & x[4704];
     layer0_out[6131] <= ~(x[8578] & x[8579]);
     layer0_out[6132] <= ~x[8866];
     layer0_out[6133] <= ~(x[5687] | x[5688]);
     layer0_out[6134] <= 1'b0;
     layer0_out[6135] <= ~(x[5191] | x[5192]);
     layer0_out[6136] <= x[4154] ^ x[4155];
     layer0_out[6137] <= x[6250] & ~x[6251];
     layer0_out[6138] <= x[919] & x[920];
     layer0_out[6139] <= x[2922] & x[2923];
     layer0_out[6140] <= x[589];
     layer0_out[6141] <= 1'b1;
     layer0_out[6142] <= ~(x[1670] & x[1672]);
     layer0_out[6143] <= ~(x[257] & x[258]);
     layer0_out[6144] <= ~x[4348] | x[4347];
     layer0_out[6145] <= x[7823] & ~x[7822];
     layer0_out[6146] <= x[4873] & x[4874];
     layer0_out[6147] <= 1'b1;
     layer0_out[6148] <= x[5891] & x[5892];
     layer0_out[6149] <= x[8727] | x[8728];
     layer0_out[6150] <= ~(x[42] & x[44]);
     layer0_out[6151] <= x[2926] & x[2927];
     layer0_out[6152] <= x[1491] & x[1492];
     layer0_out[6153] <= x[2705] & x[2707];
     layer0_out[6154] <= 1'b0;
     layer0_out[6155] <= ~(x[4622] & x[4623]);
     layer0_out[6156] <= 1'b1;
     layer0_out[6157] <= 1'b0;
     layer0_out[6158] <= x[2720] ^ x[2721];
     layer0_out[6159] <= x[2993] & x[2994];
     layer0_out[6160] <= x[5693] ^ x[5694];
     layer0_out[6161] <= x[5658];
     layer0_out[6162] <= ~x[8406];
     layer0_out[6163] <= x[1772];
     layer0_out[6164] <= ~(x[1298] & x[1299]);
     layer0_out[6165] <= ~x[3052] | x[3051];
     layer0_out[6166] <= ~(x[913] & x[915]);
     layer0_out[6167] <= 1'b0;
     layer0_out[6168] <= 1'b0;
     layer0_out[6169] <= ~(x[3089] & x[3090]);
     layer0_out[6170] <= ~(x[1918] & x[1920]);
     layer0_out[6171] <= x[8440] & x[8441];
     layer0_out[6172] <= x[2051];
     layer0_out[6173] <= x[1665] & x[1667];
     layer0_out[6174] <= ~(x[1118] & x[1120]);
     layer0_out[6175] <= ~(x[579] ^ x[580]);
     layer0_out[6176] <= x[2669] & x[2670];
     layer0_out[6177] <= x[249] & ~x[248];
     layer0_out[6178] <= ~x[1554];
     layer0_out[6179] <= x[3669] & ~x[3668];
     layer0_out[6180] <= ~(x[5691] | x[5692]);
     layer0_out[6181] <= x[2211] & x[2213];
     layer0_out[6182] <= ~x[8776] | x[8775];
     layer0_out[6183] <= ~(x[6191] | x[6192]);
     layer0_out[6184] <= ~(x[7054] | x[7055]);
     layer0_out[6185] <= x[799] & x[800];
     layer0_out[6186] <= x[2370] & ~x[2372];
     layer0_out[6187] <= ~(x[3321] ^ x[3322]);
     layer0_out[6188] <= x[390] & ~x[389];
     layer0_out[6189] <= ~(x[704] ^ x[705]);
     layer0_out[6190] <= x[620] | x[622];
     layer0_out[6191] <= x[213] & x[214];
     layer0_out[6192] <= 1'b0;
     layer0_out[6193] <= x[7020] ^ x[7021];
     layer0_out[6194] <= ~(x[5798] & x[5799]);
     layer0_out[6195] <= 1'b0;
     layer0_out[6196] <= x[3537] | x[3538];
     layer0_out[6197] <= x[5914] & x[5915];
     layer0_out[6198] <= ~(x[5135] & x[5136]);
     layer0_out[6199] <= 1'b0;
     layer0_out[6200] <= ~x[8263];
     layer0_out[6201] <= x[5629];
     layer0_out[6202] <= x[112] & ~x[113];
     layer0_out[6203] <= ~(x[689] & x[690]);
     layer0_out[6204] <= ~x[324] | x[326];
     layer0_out[6205] <= ~(x[7490] | x[7491]);
     layer0_out[6206] <= ~(x[6358] | x[6359]);
     layer0_out[6207] <= ~(x[1800] & x[1801]);
     layer0_out[6208] <= ~(x[675] ^ x[676]);
     layer0_out[6209] <= ~(x[2291] & x[2293]);
     layer0_out[6210] <= x[124];
     layer0_out[6211] <= x[2628] ^ x[2629];
     layer0_out[6212] <= ~x[2647];
     layer0_out[6213] <= x[2742];
     layer0_out[6214] <= x[5369] & x[5370];
     layer0_out[6215] <= x[9180];
     layer0_out[6216] <= x[5397] & x[5398];
     layer0_out[6217] <= x[2239] ^ x[2241];
     layer0_out[6218] <= x[1704] & x[1706];
     layer0_out[6219] <= ~x[7574];
     layer0_out[6220] <= x[6907] & x[6908];
     layer0_out[6221] <= ~(x[1163] | x[1165]);
     layer0_out[6222] <= ~(x[8484] | x[8485]);
     layer0_out[6223] <= x[590] & x[592];
     layer0_out[6224] <= x[1834] | x[1835];
     layer0_out[6225] <= ~(x[3994] & x[3995]);
     layer0_out[6226] <= x[2177] & x[2178];
     layer0_out[6227] <= ~x[5868];
     layer0_out[6228] <= x[2704] & x[2706];
     layer0_out[6229] <= ~(x[2992] | x[2993]);
     layer0_out[6230] <= x[115] | x[117];
     layer0_out[6231] <= ~(x[1699] & x[1700]);
     layer0_out[6232] <= ~(x[2760] & x[2761]);
     layer0_out[6233] <= ~(x[6113] | x[6114]);
     layer0_out[6234] <= ~(x[6952] | x[6953]);
     layer0_out[6235] <= x[1844];
     layer0_out[6236] <= x[8362] | x[8363];
     layer0_out[6237] <= ~(x[1650] & x[1652]);
     layer0_out[6238] <= ~x[1024];
     layer0_out[6239] <= ~(x[2951] & x[2952]);
     layer0_out[6240] <= ~(x[4996] | x[4997]);
     layer0_out[6241] <= ~(x[4006] | x[4007]);
     layer0_out[6242] <= ~(x[5844] & x[5845]);
     layer0_out[6243] <= x[1923] | x[1925];
     layer0_out[6244] <= x[7089] & x[7090];
     layer0_out[6245] <= x[1946];
     layer0_out[6246] <= ~(x[4254] ^ x[4255]);
     layer0_out[6247] <= x[1785] & x[1786];
     layer0_out[6248] <= x[2700] & x[2702];
     layer0_out[6249] <= ~(x[75] & x[77]);
     layer0_out[6250] <= x[347];
     layer0_out[6251] <= ~(x[8124] & x[8125]);
     layer0_out[6252] <= ~(x[2702] ^ x[2703]);
     layer0_out[6253] <= ~x[6022];
     layer0_out[6254] <= x[6608] ^ x[6609];
     layer0_out[6255] <= x[4772] & x[4773];
     layer0_out[6256] <= ~x[1648] | x[1650];
     layer0_out[6257] <= ~(x[2872] & x[2873]);
     layer0_out[6258] <= ~(x[3438] | x[3439]);
     layer0_out[6259] <= ~(x[8274] ^ x[8275]);
     layer0_out[6260] <= ~(x[4653] | x[4654]);
     layer0_out[6261] <= ~(x[6523] ^ x[6524]);
     layer0_out[6262] <= x[5813] & x[5814];
     layer0_out[6263] <= ~x[6309];
     layer0_out[6264] <= ~(x[1781] & x[1783]);
     layer0_out[6265] <= ~x[1244] | x[1242];
     layer0_out[6266] <= ~x[8424];
     layer0_out[6267] <= ~(x[6033] & x[6034]);
     layer0_out[6268] <= ~(x[3977] | x[3978]);
     layer0_out[6269] <= x[1047];
     layer0_out[6270] <= x[6322];
     layer0_out[6271] <= ~x[6916] | x[6917];
     layer0_out[6272] <= ~(x[5041] | x[5042]);
     layer0_out[6273] <= ~(x[4627] & x[4628]);
     layer0_out[6274] <= x[3618] | x[3619];
     layer0_out[6275] <= ~x[4410];
     layer0_out[6276] <= x[534] | x[535];
     layer0_out[6277] <= x[1586] & x[1588];
     layer0_out[6278] <= ~x[1019] | x[1018];
     layer0_out[6279] <= x[2153] & ~x[2154];
     layer0_out[6280] <= x[360] ^ x[361];
     layer0_out[6281] <= ~(x[1500] & x[1501]);
     layer0_out[6282] <= ~x[9080];
     layer0_out[6283] <= ~(x[4591] ^ x[4592]);
     layer0_out[6284] <= ~(x[6445] | x[6446]);
     layer0_out[6285] <= 1'b1;
     layer0_out[6286] <= ~(x[2376] & x[2377]);
     layer0_out[6287] <= x[2166] & x[2168];
     layer0_out[6288] <= ~(x[2779] | x[2780]);
     layer0_out[6289] <= x[4770] | x[4771];
     layer0_out[6290] <= ~(x[1806] | x[1807]);
     layer0_out[6291] <= x[7580] ^ x[7581];
     layer0_out[6292] <= x[610];
     layer0_out[6293] <= x[8875];
     layer0_out[6294] <= x[3707];
     layer0_out[6295] <= x[4388] & x[4389];
     layer0_out[6296] <= ~(x[4040] | x[4041]);
     layer0_out[6297] <= x[7606];
     layer0_out[6298] <= 1'b0;
     layer0_out[6299] <= x[2799];
     layer0_out[6300] <= x[905] | x[907];
     layer0_out[6301] <= x[5583];
     layer0_out[6302] <= ~(x[2854] | x[2855]);
     layer0_out[6303] <= x[5920] | x[5921];
     layer0_out[6304] <= ~(x[5339] | x[5340]);
     layer0_out[6305] <= ~(x[787] ^ x[788]);
     layer0_out[6306] <= x[4758] & ~x[4757];
     layer0_out[6307] <= x[724];
     layer0_out[6308] <= x[1050] | x[1051];
     layer0_out[6309] <= ~(x[9214] | x[9215]);
     layer0_out[6310] <= x[2633] ^ x[2635];
     layer0_out[6311] <= x[5549] ^ x[5550];
     layer0_out[6312] <= x[8833] & x[8834];
     layer0_out[6313] <= ~(x[2851] & x[2852]);
     layer0_out[6314] <= x[6826];
     layer0_out[6315] <= ~(x[2155] & x[2157]);
     layer0_out[6316] <= x[4966] & ~x[4965];
     layer0_out[6317] <= x[3633];
     layer0_out[6318] <= ~x[538];
     layer0_out[6319] <= ~(x[7880] & x[7881]);
     layer0_out[6320] <= x[6848] & ~x[6849];
     layer0_out[6321] <= x[1285];
     layer0_out[6322] <= ~x[2970];
     layer0_out[6323] <= 1'b1;
     layer0_out[6324] <= ~(x[7125] & x[7126]);
     layer0_out[6325] <= ~(x[5764] & x[5765]);
     layer0_out[6326] <= x[5989] & x[5990];
     layer0_out[6327] <= x[5360] & x[5361];
     layer0_out[6328] <= ~x[7694];
     layer0_out[6329] <= ~x[322];
     layer0_out[6330] <= x[4548];
     layer0_out[6331] <= x[4115];
     layer0_out[6332] <= 1'b0;
     layer0_out[6333] <= ~(x[3217] & x[3218]);
     layer0_out[6334] <= ~x[134];
     layer0_out[6335] <= x[2138] & x[2140];
     layer0_out[6336] <= x[6923] ^ x[6924];
     layer0_out[6337] <= x[4950] | x[4951];
     layer0_out[6338] <= 1'b0;
     layer0_out[6339] <= ~x[2170];
     layer0_out[6340] <= ~x[944];
     layer0_out[6341] <= ~x[1551] | x[1550];
     layer0_out[6342] <= x[7938] ^ x[7939];
     layer0_out[6343] <= x[5786] & x[5787];
     layer0_out[6344] <= x[1795] | x[1796];
     layer0_out[6345] <= x[3512] & x[3513];
     layer0_out[6346] <= ~(x[3956] | x[3957]);
     layer0_out[6347] <= x[5046] | x[5047];
     layer0_out[6348] <= x[4866] & x[4867];
     layer0_out[6349] <= ~x[797];
     layer0_out[6350] <= x[2280] & x[2281];
     layer0_out[6351] <= ~(x[6789] | x[6790]);
     layer0_out[6352] <= 1'b0;
     layer0_out[6353] <= ~x[5520];
     layer0_out[6354] <= x[2405] & x[2407];
     layer0_out[6355] <= x[7016] | x[7017];
     layer0_out[6356] <= x[7648] ^ x[7649];
     layer0_out[6357] <= ~(x[557] | x[559]);
     layer0_out[6358] <= x[938] & x[940];
     layer0_out[6359] <= 1'b1;
     layer0_out[6360] <= ~(x[8755] | x[8756]);
     layer0_out[6361] <= ~x[8368] | x[8367];
     layer0_out[6362] <= ~(x[788] & x[789]);
     layer0_out[6363] <= ~(x[4913] & x[4914]);
     layer0_out[6364] <= x[7317] | x[7318];
     layer0_out[6365] <= ~(x[1627] ^ x[1629]);
     layer0_out[6366] <= ~x[3682];
     layer0_out[6367] <= x[2228];
     layer0_out[6368] <= x[415] ^ x[416];
     layer0_out[6369] <= x[4740] | x[4741];
     layer0_out[6370] <= ~x[1296] | x[1294];
     layer0_out[6371] <= x[8112] & x[8113];
     layer0_out[6372] <= x[5463] & x[5464];
     layer0_out[6373] <= x[2736] & ~x[2734];
     layer0_out[6374] <= x[8118] ^ x[8119];
     layer0_out[6375] <= x[2580] & x[2581];
     layer0_out[6376] <= 1'b0;
     layer0_out[6377] <= ~(x[4150] & x[4151]);
     layer0_out[6378] <= ~x[8220];
     layer0_out[6379] <= ~(x[491] | x[492]);
     layer0_out[6380] <= ~x[66];
     layer0_out[6381] <= ~x[1093] | x[1095];
     layer0_out[6382] <= x[7143] | x[7144];
     layer0_out[6383] <= x[312] & x[314];
     layer0_out[6384] <= ~(x[5501] ^ x[5502]);
     layer0_out[6385] <= ~(x[2613] ^ x[2614]);
     layer0_out[6386] <= ~(x[548] ^ x[550]);
     layer0_out[6387] <= ~(x[6879] ^ x[6880]);
     layer0_out[6388] <= ~x[1387];
     layer0_out[6389] <= ~(x[1509] | x[1511]);
     layer0_out[6390] <= ~x[1509];
     layer0_out[6391] <= x[8701];
     layer0_out[6392] <= ~(x[1633] & x[1635]);
     layer0_out[6393] <= x[7548] ^ x[7549];
     layer0_out[6394] <= ~x[2925];
     layer0_out[6395] <= x[6666] ^ x[6667];
     layer0_out[6396] <= x[1291] & x[1293];
     layer0_out[6397] <= x[5847] ^ x[5848];
     layer0_out[6398] <= ~(x[4505] | x[4506]);
     layer0_out[6399] <= x[1106] & x[1107];
     layer0_out[6400] <= 1'b0;
     layer0_out[6401] <= ~(x[2994] ^ x[2995]);
     layer0_out[6402] <= x[6272] | x[6273];
     layer0_out[6403] <= x[217] | x[218];
     layer0_out[6404] <= ~(x[4768] ^ x[4769]);
     layer0_out[6405] <= ~(x[2725] ^ x[2727]);
     layer0_out[6406] <= ~(x[2392] & x[2394]);
     layer0_out[6407] <= x[3725] | x[3726];
     layer0_out[6408] <= ~(x[501] & x[502]);
     layer0_out[6409] <= 1'b0;
     layer0_out[6410] <= x[1749] | x[1751];
     layer0_out[6411] <= x[608] ^ x[609];
     layer0_out[6412] <= x[5147] & x[5148];
     layer0_out[6413] <= ~x[1916];
     layer0_out[6414] <= x[9143];
     layer0_out[6415] <= ~x[277];
     layer0_out[6416] <= ~(x[1256] & x[1258]);
     layer0_out[6417] <= ~(x[1269] & x[1271]);
     layer0_out[6418] <= ~(x[2676] & x[2678]);
     layer0_out[6419] <= x[3333];
     layer0_out[6420] <= ~x[3429];
     layer0_out[6421] <= x[1205] & x[1207];
     layer0_out[6422] <= ~(x[4083] | x[4084]);
     layer0_out[6423] <= ~(x[3042] & x[3043]);
     layer0_out[6424] <= x[3082] & ~x[3083];
     layer0_out[6425] <= ~(x[3802] & x[3803]);
     layer0_out[6426] <= x[5329] & x[5330];
     layer0_out[6427] <= ~x[666] | x[665];
     layer0_out[6428] <= x[9043];
     layer0_out[6429] <= ~(x[6532] | x[6533]);
     layer0_out[6430] <= x[503] ^ x[504];
     layer0_out[6431] <= ~(x[8189] ^ x[8190]);
     layer0_out[6432] <= x[4005];
     layer0_out[6433] <= ~x[7436] | x[7437];
     layer0_out[6434] <= ~x[937];
     layer0_out[6435] <= ~(x[7703] ^ x[7704]);
     layer0_out[6436] <= ~x[7460];
     layer0_out[6437] <= ~x[5614];
     layer0_out[6438] <= ~x[4117];
     layer0_out[6439] <= ~(x[8293] & x[8294]);
     layer0_out[6440] <= x[7918] | x[7919];
     layer0_out[6441] <= ~x[5062];
     layer0_out[6442] <= x[7596] | x[7597];
     layer0_out[6443] <= ~(x[4700] & x[4701]);
     layer0_out[6444] <= ~(x[1675] & x[1676]);
     layer0_out[6445] <= x[5219] & ~x[5220];
     layer0_out[6446] <= ~(x[4217] & x[4218]);
     layer0_out[6447] <= x[147] ^ x[148];
     layer0_out[6448] <= ~x[7705];
     layer0_out[6449] <= x[1888];
     layer0_out[6450] <= 1'b0;
     layer0_out[6451] <= ~x[1164] | x[1165];
     layer0_out[6452] <= x[1849];
     layer0_out[6453] <= x[578] ^ x[580];
     layer0_out[6454] <= ~(x[623] & x[625]);
     layer0_out[6455] <= x[3757] ^ x[3758];
     layer0_out[6456] <= x[720] ^ x[721];
     layer0_out[6457] <= ~x[7314];
     layer0_out[6458] <= x[5323] & x[5324];
     layer0_out[6459] <= x[1457] & x[1458];
     layer0_out[6460] <= x[3590];
     layer0_out[6461] <= ~(x[7144] | x[7145]);
     layer0_out[6462] <= 1'b0;
     layer0_out[6463] <= x[1265] & x[1266];
     layer0_out[6464] <= ~x[1177];
     layer0_out[6465] <= ~(x[2333] & x[2334]);
     layer0_out[6466] <= x[8360];
     layer0_out[6467] <= ~(x[2563] & x[2564]);
     layer0_out[6468] <= ~(x[730] ^ x[731]);
     layer0_out[6469] <= ~(x[8663] ^ x[8664]);
     layer0_out[6470] <= ~(x[4614] & x[4615]);
     layer0_out[6471] <= x[4270];
     layer0_out[6472] <= 1'b0;
     layer0_out[6473] <= ~(x[3943] | x[3944]);
     layer0_out[6474] <= ~(x[7290] ^ x[7291]);
     layer0_out[6475] <= x[2452] & x[2454];
     layer0_out[6476] <= ~(x[1107] | x[1109]);
     layer0_out[6477] <= x[2005];
     layer0_out[6478] <= x[7775] | x[7776];
     layer0_out[6479] <= ~(x[7618] & x[7619]);
     layer0_out[6480] <= ~(x[451] | x[452]);
     layer0_out[6481] <= ~x[222] | x[223];
     layer0_out[6482] <= ~(x[527] & x[528]);
     layer0_out[6483] <= ~(x[1654] ^ x[1656]);
     layer0_out[6484] <= ~(x[7207] | x[7208]);
     layer0_out[6485] <= x[1710] & x[1711];
     layer0_out[6486] <= x[7972];
     layer0_out[6487] <= x[7285] | x[7286];
     layer0_out[6488] <= x[1962] | x[1964];
     layer0_out[6489] <= x[5915] ^ x[5916];
     layer0_out[6490] <= x[7121] & ~x[7120];
     layer0_out[6491] <= ~x[1];
     layer0_out[6492] <= x[6061] & x[6062];
     layer0_out[6493] <= ~(x[1690] & x[1691]);
     layer0_out[6494] <= ~(x[705] | x[707]);
     layer0_out[6495] <= ~(x[762] & x[764]);
     layer0_out[6496] <= 1'b1;
     layer0_out[6497] <= ~(x[8892] & x[8893]);
     layer0_out[6498] <= ~(x[5610] & x[5611]);
     layer0_out[6499] <= ~x[1447];
     layer0_out[6500] <= x[3313] | x[3314];
     layer0_out[6501] <= ~x[1036] | x[1037];
     layer0_out[6502] <= x[2735] & ~x[2734];
     layer0_out[6503] <= ~(x[8617] | x[8618]);
     layer0_out[6504] <= x[4102] | x[4103];
     layer0_out[6505] <= x[705] ^ x[706];
     layer0_out[6506] <= ~x[9207];
     layer0_out[6507] <= x[1540] & x[1542];
     layer0_out[6508] <= x[5016] | x[5017];
     layer0_out[6509] <= ~(x[8768] ^ x[8769]);
     layer0_out[6510] <= ~x[8569];
     layer0_out[6511] <= ~x[5438];
     layer0_out[6512] <= x[90] & x[91];
     layer0_out[6513] <= ~(x[32] & x[33]);
     layer0_out[6514] <= x[2511];
     layer0_out[6515] <= x[1127] & x[1128];
     layer0_out[6516] <= ~x[3924];
     layer0_out[6517] <= ~x[6941];
     layer0_out[6518] <= x[7879] | x[7880];
     layer0_out[6519] <= x[5873];
     layer0_out[6520] <= x[3269] | x[3270];
     layer0_out[6521] <= ~(x[656] ^ x[658]);
     layer0_out[6522] <= ~x[114];
     layer0_out[6523] <= ~(x[3487] | x[3488]);
     layer0_out[6524] <= x[6227] ^ x[6228];
     layer0_out[6525] <= ~(x[1643] ^ x[1645]);
     layer0_out[6526] <= x[8310] & x[8311];
     layer0_out[6527] <= 1'b1;
     layer0_out[6528] <= x[6419];
     layer0_out[6529] <= x[124] | x[126];
     layer0_out[6530] <= ~(x[2225] & x[2226]);
     layer0_out[6531] <= x[762] & x[763];
     layer0_out[6532] <= ~(x[1551] ^ x[1552]);
     layer0_out[6533] <= ~(x[97] & x[99]);
     layer0_out[6534] <= x[3727];
     layer0_out[6535] <= x[5045] ^ x[5046];
     layer0_out[6536] <= x[1564];
     layer0_out[6537] <= x[304] & x[306];
     layer0_out[6538] <= 1'b0;
     layer0_out[6539] <= x[1208] ^ x[1209];
     layer0_out[6540] <= ~(x[2328] & x[2330]);
     layer0_out[6541] <= x[1486] ^ x[1487];
     layer0_out[6542] <= x[1254] & x[1255];
     layer0_out[6543] <= ~(x[7084] & x[7085]);
     layer0_out[6544] <= x[8571] | x[8572];
     layer0_out[6545] <= ~x[8449];
     layer0_out[6546] <= ~x[4613];
     layer0_out[6547] <= ~(x[2239] | x[2240]);
     layer0_out[6548] <= ~(x[2082] | x[2083]);
     layer0_out[6549] <= x[1810] & x[1812];
     layer0_out[6550] <= ~x[976];
     layer0_out[6551] <= ~(x[2767] ^ x[2768]);
     layer0_out[6552] <= x[5102] & x[5103];
     layer0_out[6553] <= ~(x[8229] | x[8230]);
     layer0_out[6554] <= ~(x[33] | x[34]);
     layer0_out[6555] <= x[1827] | x[1829];
     layer0_out[6556] <= x[6400] ^ x[6401];
     layer0_out[6557] <= x[1860] & x[1862];
     layer0_out[6558] <= x[9159];
     layer0_out[6559] <= x[7858] | x[7859];
     layer0_out[6560] <= ~(x[1356] & x[1357]);
     layer0_out[6561] <= ~(x[1057] ^ x[1059]);
     layer0_out[6562] <= ~x[88];
     layer0_out[6563] <= ~(x[4436] & x[4437]);
     layer0_out[6564] <= x[7028] & x[7029];
     layer0_out[6565] <= ~(x[1739] | x[1740]);
     layer0_out[6566] <= x[1362] & x[1363];
     layer0_out[6567] <= ~(x[5414] & x[5415]);
     layer0_out[6568] <= x[242];
     layer0_out[6569] <= ~(x[736] | x[737]);
     layer0_out[6570] <= 1'b1;
     layer0_out[6571] <= 1'b0;
     layer0_out[6572] <= x[498] & x[499];
     layer0_out[6573] <= x[1200] & ~x[1202];
     layer0_out[6574] <= x[520] & x[522];
     layer0_out[6575] <= ~(x[1703] & x[1705]);
     layer0_out[6576] <= x[2421];
     layer0_out[6577] <= x[5827] & x[5828];
     layer0_out[6578] <= x[5434] & x[5435];
     layer0_out[6579] <= x[5956] & x[5957];
     layer0_out[6580] <= ~(x[3918] | x[3919]);
     layer0_out[6581] <= x[1437];
     layer0_out[6582] <= ~(x[1957] & x[1958]);
     layer0_out[6583] <= ~(x[1926] | x[1927]);
     layer0_out[6584] <= ~(x[7324] | x[7325]);
     layer0_out[6585] <= ~(x[998] ^ x[999]);
     layer0_out[6586] <= ~(x[4555] & x[4556]);
     layer0_out[6587] <= ~(x[3983] & x[3984]);
     layer0_out[6588] <= x[7265];
     layer0_out[6589] <= ~(x[3212] | x[3213]);
     layer0_out[6590] <= ~x[8204];
     layer0_out[6591] <= x[2714] ^ x[2715];
     layer0_out[6592] <= x[3813] ^ x[3814];
     layer0_out[6593] <= x[7830] | x[7831];
     layer0_out[6594] <= x[2360] ^ x[2362];
     layer0_out[6595] <= x[1426] & x[1427];
     layer0_out[6596] <= x[1059] & x[1060];
     layer0_out[6597] <= ~x[7910];
     layer0_out[6598] <= x[140] & ~x[139];
     layer0_out[6599] <= ~x[1975];
     layer0_out[6600] <= ~(x[500] | x[501]);
     layer0_out[6601] <= ~(x[141] & x[143]);
     layer0_out[6602] <= x[1039] & x[1041];
     layer0_out[6603] <= ~(x[1913] & x[1914]);
     layer0_out[6604] <= x[7327];
     layer0_out[6605] <= 1'b0;
     layer0_out[6606] <= ~(x[974] ^ x[975]);
     layer0_out[6607] <= ~x[205];
     layer0_out[6608] <= ~(x[210] | x[211]);
     layer0_out[6609] <= ~x[5481];
     layer0_out[6610] <= 1'b1;
     layer0_out[6611] <= x[6114] & x[6115];
     layer0_out[6612] <= ~x[3316];
     layer0_out[6613] <= ~(x[1893] ^ x[1895]);
     layer0_out[6614] <= x[3688] & ~x[3689];
     layer0_out[6615] <= x[90];
     layer0_out[6616] <= ~x[1117];
     layer0_out[6617] <= x[1429] ^ x[1431];
     layer0_out[6618] <= ~(x[1357] & x[1358]);
     layer0_out[6619] <= x[7731];
     layer0_out[6620] <= x[603] ^ x[604];
     layer0_out[6621] <= x[5632] ^ x[5633];
     layer0_out[6622] <= ~(x[809] | x[810]);
     layer0_out[6623] <= x[7496] & x[7497];
     layer0_out[6624] <= ~(x[302] & x[304]);
     layer0_out[6625] <= ~x[2530];
     layer0_out[6626] <= x[760] | x[762];
     layer0_out[6627] <= ~x[5458];
     layer0_out[6628] <= x[662] & ~x[663];
     layer0_out[6629] <= x[1194] & x[1196];
     layer0_out[6630] <= ~(x[1671] | x[1673]);
     layer0_out[6631] <= ~(x[1479] | x[1481]);
     layer0_out[6632] <= x[6614] & x[6615];
     layer0_out[6633] <= x[2094] & x[2095];
     layer0_out[6634] <= ~(x[2345] & x[2346]);
     layer0_out[6635] <= 1'b0;
     layer0_out[6636] <= ~(x[755] & x[756]);
     layer0_out[6637] <= x[891];
     layer0_out[6638] <= x[1745] | x[1747];
     layer0_out[6639] <= x[1089] & x[1090];
     layer0_out[6640] <= 1'b0;
     layer0_out[6641] <= ~(x[3520] ^ x[3521]);
     layer0_out[6642] <= ~(x[1927] | x[1928]);
     layer0_out[6643] <= x[3007] & x[3008];
     layer0_out[6644] <= x[5607] & x[5608];
     layer0_out[6645] <= 1'b0;
     layer0_out[6646] <= ~(x[5741] | x[5742]);
     layer0_out[6647] <= 1'b1;
     layer0_out[6648] <= x[1583] & x[1584];
     layer0_out[6649] <= x[1490] & x[1492];
     layer0_out[6650] <= x[6621] ^ x[6622];
     layer0_out[6651] <= ~(x[4755] | x[4756]);
     layer0_out[6652] <= 1'b1;
     layer0_out[6653] <= x[1982] & x[1984];
     layer0_out[6654] <= ~(x[7227] | x[7228]);
     layer0_out[6655] <= ~(x[7111] & x[7112]);
     layer0_out[6656] <= x[2540] & x[2541];
     layer0_out[6657] <= ~x[2471] | x[2469];
     layer0_out[6658] <= ~(x[5165] | x[5166]);
     layer0_out[6659] <= ~(x[4086] & x[4087]);
     layer0_out[6660] <= x[144] & ~x[143];
     layer0_out[6661] <= x[6131] & x[6132];
     layer0_out[6662] <= x[75] & ~x[73];
     layer0_out[6663] <= x[5967] & x[5968];
     layer0_out[6664] <= x[1479] ^ x[1480];
     layer0_out[6665] <= ~x[4623];
     layer0_out[6666] <= x[7418] & x[7419];
     layer0_out[6667] <= ~(x[6770] | x[6771]);
     layer0_out[6668] <= 1'b1;
     layer0_out[6669] <= ~(x[5221] & x[5222]);
     layer0_out[6670] <= x[188] | x[190];
     layer0_out[6671] <= ~(x[7179] & x[7180]);
     layer0_out[6672] <= x[4552] & x[4553];
     layer0_out[6673] <= 1'b0;
     layer0_out[6674] <= x[8199] | x[8200];
     layer0_out[6675] <= x[8283] | x[8284];
     layer0_out[6676] <= ~(x[2448] & x[2450]);
     layer0_out[6677] <= ~(x[4220] & x[4221]);
     layer0_out[6678] <= x[369];
     layer0_out[6679] <= ~(x[7458] | x[7459]);
     layer0_out[6680] <= ~(x[2293] & x[2295]);
     layer0_out[6681] <= ~x[3003];
     layer0_out[6682] <= x[8151] | x[8152];
     layer0_out[6683] <= x[2302] & x[2304];
     layer0_out[6684] <= ~(x[677] ^ x[678]);
     layer0_out[6685] <= ~(x[8824] | x[8825]);
     layer0_out[6686] <= ~(x[8703] & x[8704]);
     layer0_out[6687] <= 1'b0;
     layer0_out[6688] <= 1'b0;
     layer0_out[6689] <= x[2776] ^ x[2778];
     layer0_out[6690] <= ~(x[8433] ^ x[8434]);
     layer0_out[6691] <= ~(x[481] | x[482]);
     layer0_out[6692] <= x[5759];
     layer0_out[6693] <= x[3647] & x[3648];
     layer0_out[6694] <= ~(x[8008] | x[8009]);
     layer0_out[6695] <= x[7746];
     layer0_out[6696] <= x[406];
     layer0_out[6697] <= ~(x[4384] | x[4385]);
     layer0_out[6698] <= ~x[6054];
     layer0_out[6699] <= x[8723] | x[8724];
     layer0_out[6700] <= x[353] & x[355];
     layer0_out[6701] <= ~x[6278];
     layer0_out[6702] <= x[373];
     layer0_out[6703] <= x[7435] & x[7436];
     layer0_out[6704] <= ~x[2106];
     layer0_out[6705] <= x[7035] | x[7036];
     layer0_out[6706] <= ~(x[2175] & x[2177]);
     layer0_out[6707] <= ~(x[6545] & x[6546]);
     layer0_out[6708] <= x[1376] & x[1378];
     layer0_out[6709] <= x[4458] & x[4459];
     layer0_out[6710] <= ~x[4881];
     layer0_out[6711] <= x[7910];
     layer0_out[6712] <= ~x[3169];
     layer0_out[6713] <= ~(x[1737] & x[1738]);
     layer0_out[6714] <= x[2161] & x[2163];
     layer0_out[6715] <= x[1488] & x[1490];
     layer0_out[6716] <= x[3562] & ~x[3561];
     layer0_out[6717] <= x[8329] | x[8330];
     layer0_out[6718] <= x[3406];
     layer0_out[6719] <= x[1605];
     layer0_out[6720] <= x[1590] | x[1592];
     layer0_out[6721] <= x[6939] | x[6940];
     layer0_out[6722] <= 1'b0;
     layer0_out[6723] <= x[849] & x[850];
     layer0_out[6724] <= x[3536];
     layer0_out[6725] <= ~(x[6290] | x[6291]);
     layer0_out[6726] <= ~x[7204];
     layer0_out[6727] <= 1'b1;
     layer0_out[6728] <= ~(x[5846] & x[5847]);
     layer0_out[6729] <= x[4707] & x[4708];
     layer0_out[6730] <= ~x[9026] | x[9025];
     layer0_out[6731] <= x[7690] | x[7691];
     layer0_out[6732] <= x[6650] & ~x[6651];
     layer0_out[6733] <= ~(x[1037] & x[1038]);
     layer0_out[6734] <= ~(x[1943] & x[1945]);
     layer0_out[6735] <= x[3597] | x[3598];
     layer0_out[6736] <= x[5234] & ~x[5233];
     layer0_out[6737] <= ~(x[978] | x[979]);
     layer0_out[6738] <= ~(x[1536] & x[1537]);
     layer0_out[6739] <= ~(x[2188] & x[2190]);
     layer0_out[6740] <= x[7857] | x[7858];
     layer0_out[6741] <= ~x[2510];
     layer0_out[6742] <= 1'b0;
     layer0_out[6743] <= x[8476] ^ x[8477];
     layer0_out[6744] <= ~(x[5415] & x[5416]);
     layer0_out[6745] <= ~(x[3555] ^ x[3556]);
     layer0_out[6746] <= ~x[4741];
     layer0_out[6747] <= ~x[270] | x[271];
     layer0_out[6748] <= x[2654] ^ x[2655];
     layer0_out[6749] <= x[826] | x[828];
     layer0_out[6750] <= ~(x[1731] | x[1732]);
     layer0_out[6751] <= ~(x[8745] | x[8746]);
     layer0_out[6752] <= x[210] & x[212];
     layer0_out[6753] <= x[416] & x[418];
     layer0_out[6754] <= ~(x[7187] | x[7188]);
     layer0_out[6755] <= x[1099] & x[1101];
     layer0_out[6756] <= x[5811] & x[5812];
     layer0_out[6757] <= ~(x[8619] | x[8620]);
     layer0_out[6758] <= x[8268];
     layer0_out[6759] <= x[4743] & ~x[4742];
     layer0_out[6760] <= x[4182] | x[4183];
     layer0_out[6761] <= ~x[1159] | x[1160];
     layer0_out[6762] <= x[2195] & x[2196];
     layer0_out[6763] <= x[5315] & x[5316];
     layer0_out[6764] <= x[517] & x[519];
     layer0_out[6765] <= ~(x[1175] ^ x[1177]);
     layer0_out[6766] <= ~(x[3766] | x[3767]);
     layer0_out[6767] <= ~(x[2210] | x[2211]);
     layer0_out[6768] <= x[1357] & x[1359];
     layer0_out[6769] <= x[2248] & x[2250];
     layer0_out[6770] <= x[8831] & ~x[8832];
     layer0_out[6771] <= ~(x[6905] | x[6906]);
     layer0_out[6772] <= x[6408];
     layer0_out[6773] <= ~(x[7990] & x[7991]);
     layer0_out[6774] <= x[7905] & x[7906];
     layer0_out[6775] <= ~(x[764] ^ x[766]);
     layer0_out[6776] <= x[2808] | x[2809];
     layer0_out[6777] <= x[4847] & x[4848];
     layer0_out[6778] <= ~(x[1236] & x[1238]);
     layer0_out[6779] <= x[3004];
     layer0_out[6780] <= x[7921] & x[7922];
     layer0_out[6781] <= ~x[3998] | x[3997];
     layer0_out[6782] <= x[9208] | x[9209];
     layer0_out[6783] <= ~(x[4444] & x[4445]);
     layer0_out[6784] <= x[1054] & x[1055];
     layer0_out[6785] <= x[2728] & x[2730];
     layer0_out[6786] <= x[7560];
     layer0_out[6787] <= ~x[4737];
     layer0_out[6788] <= x[8153] & x[8154];
     layer0_out[6789] <= x[0] | x[2];
     layer0_out[6790] <= ~x[5639];
     layer0_out[6791] <= 1'b0;
     layer0_out[6792] <= 1'b1;
     layer0_out[6793] <= ~(x[1797] & x[1798]);
     layer0_out[6794] <= x[709] & x[711];
     layer0_out[6795] <= x[1634] & x[1636];
     layer0_out[6796] <= x[7996];
     layer0_out[6797] <= ~(x[7924] & x[7925]);
     layer0_out[6798] <= x[7948] | x[7949];
     layer0_out[6799] <= ~x[9077];
     layer0_out[6800] <= ~x[5834];
     layer0_out[6801] <= ~(x[6010] ^ x[6011]);
     layer0_out[6802] <= ~x[2373] | x[2374];
     layer0_out[6803] <= x[1883] & x[1885];
     layer0_out[6804] <= 1'b1;
     layer0_out[6805] <= x[3146] | x[3147];
     layer0_out[6806] <= x[5292] & x[5293];
     layer0_out[6807] <= ~(x[5249] & x[5250]);
     layer0_out[6808] <= x[4113] & ~x[4112];
     layer0_out[6809] <= x[590] ^ x[591];
     layer0_out[6810] <= 1'b0;
     layer0_out[6811] <= x[7359] ^ x[7360];
     layer0_out[6812] <= x[7221] | x[7222];
     layer0_out[6813] <= x[6721];
     layer0_out[6814] <= x[2921];
     layer0_out[6815] <= ~(x[1709] & x[1711]);
     layer0_out[6816] <= x[3696] | x[3697];
     layer0_out[6817] <= x[1872];
     layer0_out[6818] <= x[1364] & ~x[1363];
     layer0_out[6819] <= ~x[801] | x[803];
     layer0_out[6820] <= x[5896] & x[5897];
     layer0_out[6821] <= ~(x[326] | x[327]);
     layer0_out[6822] <= x[2655] & x[2657];
     layer0_out[6823] <= x[54] ^ x[56];
     layer0_out[6824] <= ~(x[5464] | x[5465]);
     layer0_out[6825] <= x[7631] | x[7632];
     layer0_out[6826] <= ~(x[7838] ^ x[7839]);
     layer0_out[6827] <= ~(x[1326] ^ x[1327]);
     layer0_out[6828] <= ~(x[8170] & x[8171]);
     layer0_out[6829] <= ~(x[1560] & x[1561]);
     layer0_out[6830] <= ~x[6920] | x[6919];
     layer0_out[6831] <= x[5925] & x[5926];
     layer0_out[6832] <= x[4261] | x[4262];
     layer0_out[6833] <= ~x[8986];
     layer0_out[6834] <= ~(x[2202] | x[2204]);
     layer0_out[6835] <= ~x[58];
     layer0_out[6836] <= ~x[3190];
     layer0_out[6837] <= ~x[7683];
     layer0_out[6838] <= ~x[800];
     layer0_out[6839] <= x[7350] & ~x[7349];
     layer0_out[6840] <= x[9007] | x[9008];
     layer0_out[6841] <= ~(x[1884] | x[1886]);
     layer0_out[6842] <= ~(x[1449] & x[1451]);
     layer0_out[6843] <= x[980] | x[981];
     layer0_out[6844] <= x[8566] ^ x[8567];
     layer0_out[6845] <= ~(x[775] & x[776]);
     layer0_out[6846] <= x[5854] & x[5855];
     layer0_out[6847] <= ~x[8373];
     layer0_out[6848] <= ~x[1846];
     layer0_out[6849] <= x[993];
     layer0_out[6850] <= 1'b1;
     layer0_out[6851] <= x[2579] & x[2581];
     layer0_out[6852] <= ~(x[451] | x[453]);
     layer0_out[6853] <= x[4497] & ~x[4498];
     layer0_out[6854] <= ~x[2042];
     layer0_out[6855] <= ~(x[1728] & x[1730]);
     layer0_out[6856] <= x[3148] & x[3149];
     layer0_out[6857] <= x[2241] & x[2243];
     layer0_out[6858] <= ~(x[6577] & x[6578]);
     layer0_out[6859] <= ~(x[3401] | x[3402]);
     layer0_out[6860] <= ~x[225] | x[224];
     layer0_out[6861] <= x[2218] & ~x[2216];
     layer0_out[6862] <= x[1303] & x[1304];
     layer0_out[6863] <= ~x[7708];
     layer0_out[6864] <= x[3188] | x[3189];
     layer0_out[6865] <= x[6779];
     layer0_out[6866] <= x[6619] ^ x[6620];
     layer0_out[6867] <= x[5429];
     layer0_out[6868] <= ~(x[6365] ^ x[6366]);
     layer0_out[6869] <= ~(x[1107] & x[1108]);
     layer0_out[6870] <= x[5716] & x[5717];
     layer0_out[6871] <= x[2489] ^ x[2491];
     layer0_out[6872] <= ~(x[8375] | x[8376]);
     layer0_out[6873] <= ~x[5930];
     layer0_out[6874] <= 1'b0;
     layer0_out[6875] <= x[6547] | x[6548];
     layer0_out[6876] <= 1'b1;
     layer0_out[6877] <= x[879];
     layer0_out[6878] <= ~(x[727] | x[728]);
     layer0_out[6879] <= x[82] & x[83];
     layer0_out[6880] <= x[8595] | x[8596];
     layer0_out[6881] <= x[7945] | x[7946];
     layer0_out[6882] <= ~(x[5633] & x[5634]);
     layer0_out[6883] <= ~x[11] | x[12];
     layer0_out[6884] <= ~(x[6379] | x[6380]);
     layer0_out[6885] <= ~(x[7882] ^ x[7883]);
     layer0_out[6886] <= ~(x[2495] ^ x[2497]);
     layer0_out[6887] <= x[5048] & x[5049];
     layer0_out[6888] <= ~(x[5297] & x[5298]);
     layer0_out[6889] <= x[4538] ^ x[4539];
     layer0_out[6890] <= x[3107] | x[3108];
     layer0_out[6891] <= ~(x[6053] | x[6054]);
     layer0_out[6892] <= ~(x[232] | x[233]);
     layer0_out[6893] <= ~(x[5980] & x[5981]);
     layer0_out[6894] <= 1'b0;
     layer0_out[6895] <= ~x[236];
     layer0_out[6896] <= ~(x[1992] & x[1994]);
     layer0_out[6897] <= ~x[4784];
     layer0_out[6898] <= ~x[3628] | x[3629];
     layer0_out[6899] <= x[387] & x[389];
     layer0_out[6900] <= x[7804];
     layer0_out[6901] <= ~(x[8971] | x[8972]);
     layer0_out[6902] <= x[344] & ~x[345];
     layer0_out[6903] <= x[4166] & x[4167];
     layer0_out[6904] <= ~(x[3832] | x[3833]);
     layer0_out[6905] <= 1'b1;
     layer0_out[6906] <= x[285];
     layer0_out[6907] <= x[1579];
     layer0_out[6908] <= ~x[8685];
     layer0_out[6909] <= ~(x[4414] | x[4415]);
     layer0_out[6910] <= 1'b0;
     layer0_out[6911] <= x[8654] | x[8655];
     layer0_out[6912] <= ~(x[2669] ^ x[2671]);
     layer0_out[6913] <= ~x[5564];
     layer0_out[6914] <= ~(x[2684] & x[2686]);
     layer0_out[6915] <= x[2522] | x[2524];
     layer0_out[6916] <= x[1597] & x[1598];
     layer0_out[6917] <= ~x[3979];
     layer0_out[6918] <= x[49] & x[51];
     layer0_out[6919] <= x[2999] & x[3000];
     layer0_out[6920] <= x[1367] & x[1368];
     layer0_out[6921] <= x[4143];
     layer0_out[6922] <= x[2948] & x[2949];
     layer0_out[6923] <= x[2767] & ~x[2766];
     layer0_out[6924] <= ~x[6283];
     layer0_out[6925] <= ~(x[6593] | x[6594]);
     layer0_out[6926] <= ~x[1291] | x[1292];
     layer0_out[6927] <= ~(x[1157] | x[1158]);
     layer0_out[6928] <= x[4320] & x[4321];
     layer0_out[6929] <= ~(x[4301] | x[4302]);
     layer0_out[6930] <= ~(x[882] | x[884]);
     layer0_out[6931] <= x[2521] ^ x[2523];
     layer0_out[6932] <= 1'b1;
     layer0_out[6933] <= x[4417] & x[4418];
     layer0_out[6934] <= ~x[7954];
     layer0_out[6935] <= ~(x[3914] | x[3915]);
     layer0_out[6936] <= ~(x[4271] | x[4272]);
     layer0_out[6937] <= x[4237] | x[4238];
     layer0_out[6938] <= ~x[1453];
     layer0_out[6939] <= x[157] & ~x[158];
     layer0_out[6940] <= ~(x[2282] | x[2284]);
     layer0_out[6941] <= ~(x[2962] | x[2963]);
     layer0_out[6942] <= x[2749];
     layer0_out[6943] <= x[2662] | x[2663];
     layer0_out[6944] <= ~x[3968];
     layer0_out[6945] <= 1'b0;
     layer0_out[6946] <= ~(x[1483] & x[1484]);
     layer0_out[6947] <= x[557];
     layer0_out[6948] <= 1'b1;
     layer0_out[6949] <= x[491] ^ x[493];
     layer0_out[6950] <= x[3483];
     layer0_out[6951] <= 1'b1;
     layer0_out[6952] <= ~x[3784];
     layer0_out[6953] <= x[2299];
     layer0_out[6954] <= ~(x[1569] | x[1570]);
     layer0_out[6955] <= x[4070] ^ x[4071];
     layer0_out[6956] <= ~x[6842] | x[6843];
     layer0_out[6957] <= ~(x[1180] & x[1181]);
     layer0_out[6958] <= x[8670] ^ x[8671];
     layer0_out[6959] <= ~(x[7761] & x[7762]);
     layer0_out[6960] <= x[8673] & ~x[8672];
     layer0_out[6961] <= x[5441] & x[5442];
     layer0_out[6962] <= x[1391] & x[1393];
     layer0_out[6963] <= x[1568] ^ x[1570];
     layer0_out[6964] <= 1'b0;
     layer0_out[6965] <= ~(x[5238] ^ x[5239]);
     layer0_out[6966] <= ~(x[1359] & x[1360]);
     layer0_out[6967] <= x[812];
     layer0_out[6968] <= x[1793] & x[1795];
     layer0_out[6969] <= ~x[362] | x[363];
     layer0_out[6970] <= x[1496] | x[1498];
     layer0_out[6971] <= ~x[1390] | x[1392];
     layer0_out[6972] <= 1'b1;
     layer0_out[6973] <= x[283] ^ x[285];
     layer0_out[6974] <= x[559] & ~x[561];
     layer0_out[6975] <= x[1104];
     layer0_out[6976] <= ~x[557];
     layer0_out[6977] <= ~(x[5886] & x[5887]);
     layer0_out[6978] <= x[3551] & x[3552];
     layer0_out[6979] <= x[4632] ^ x[4633];
     layer0_out[6980] <= ~(x[2711] & x[2713]);
     layer0_out[6981] <= ~(x[7818] | x[7819]);
     layer0_out[6982] <= x[2848] | x[2849];
     layer0_out[6983] <= ~(x[7455] | x[7456]);
     layer0_out[6984] <= x[4255] ^ x[4256];
     layer0_out[6985] <= ~(x[581] | x[582]);
     layer0_out[6986] <= x[1895] & x[1896];
     layer0_out[6987] <= ~x[4551];
     layer0_out[6988] <= ~(x[7076] ^ x[7077]);
     layer0_out[6989] <= ~(x[2107] & x[2108]);
     layer0_out[6990] <= ~(x[2323] & x[2324]);
     layer0_out[6991] <= ~(x[2742] & x[2743]);
     layer0_out[6992] <= ~(x[2434] ^ x[2436]);
     layer0_out[6993] <= ~(x[1698] & x[1700]);
     layer0_out[6994] <= ~(x[4099] | x[4100]);
     layer0_out[6995] <= x[8981] & ~x[8980];
     layer0_out[6996] <= x[5743] & x[5744];
     layer0_out[6997] <= x[1775] & x[1776];
     layer0_out[6998] <= x[742] & x[743];
     layer0_out[6999] <= x[7751] & ~x[7750];
     layer0_out[7000] <= ~x[6458] | x[6457];
     layer0_out[7001] <= x[729] & x[731];
     layer0_out[7002] <= ~(x[7358] ^ x[7359]);
     layer0_out[7003] <= ~x[7979];
     layer0_out[7004] <= x[8548] | x[8549];
     layer0_out[7005] <= ~(x[5085] & x[5086]);
     layer0_out[7006] <= ~(x[2008] ^ x[2009]);
     layer0_out[7007] <= ~x[8103] | x[8104];
     layer0_out[7008] <= ~x[3841] | x[3842];
     layer0_out[7009] <= ~(x[7193] | x[7194]);
     layer0_out[7010] <= x[1035] & x[1037];
     layer0_out[7011] <= x[6244] & ~x[6245];
     layer0_out[7012] <= ~(x[918] & x[920]);
     layer0_out[7013] <= x[3851] | x[3852];
     layer0_out[7014] <= ~x[3287] | x[3288];
     layer0_out[7015] <= x[170] | x[172];
     layer0_out[7016] <= ~(x[1412] | x[1413]);
     layer0_out[7017] <= x[5828] & x[5829];
     layer0_out[7018] <= x[6729] & ~x[6730];
     layer0_out[7019] <= ~(x[3693] | x[3694]);
     layer0_out[7020] <= ~x[9112];
     layer0_out[7021] <= x[20] & ~x[21];
     layer0_out[7022] <= x[5877] & x[5878];
     layer0_out[7023] <= ~(x[4178] & x[4179]);
     layer0_out[7024] <= 1'b1;
     layer0_out[7025] <= x[1077] & x[1079];
     layer0_out[7026] <= x[2240] & x[2241];
     layer0_out[7027] <= x[80];
     layer0_out[7028] <= ~(x[8123] & x[8124]);
     layer0_out[7029] <= x[4031] ^ x[4032];
     layer0_out[7030] <= 1'b0;
     layer0_out[7031] <= ~(x[4936] | x[4937]);
     layer0_out[7032] <= 1'b1;
     layer0_out[7033] <= x[7842] & ~x[7843];
     layer0_out[7034] <= ~(x[3790] | x[3791]);
     layer0_out[7035] <= x[4472] & ~x[4473];
     layer0_out[7036] <= x[1427] & x[1428];
     layer0_out[7037] <= x[1286] & x[1288];
     layer0_out[7038] <= ~x[5613];
     layer0_out[7039] <= 1'b0;
     layer0_out[7040] <= x[621];
     layer0_out[7041] <= x[2022];
     layer0_out[7042] <= ~(x[679] | x[680]);
     layer0_out[7043] <= x[7382] & x[7383];
     layer0_out[7044] <= x[1347] | x[1349];
     layer0_out[7045] <= x[5124] & x[5125];
     layer0_out[7046] <= ~(x[2718] & x[2719]);
     layer0_out[7047] <= ~x[1020] | x[1019];
     layer0_out[7048] <= x[2232] & x[2234];
     layer0_out[7049] <= x[674] & ~x[673];
     layer0_out[7050] <= ~(x[3358] | x[3359]);
     layer0_out[7051] <= x[414];
     layer0_out[7052] <= x[9081] | x[9082];
     layer0_out[7053] <= ~x[80];
     layer0_out[7054] <= ~(x[5077] | x[5078]);
     layer0_out[7055] <= ~x[8842];
     layer0_out[7056] <= ~(x[8370] & x[8371]);
     layer0_out[7057] <= x[418] | x[419];
     layer0_out[7058] <= 1'b1;
     layer0_out[7059] <= ~(x[322] & x[323]);
     layer0_out[7060] <= ~(x[2687] ^ x[2689]);
     layer0_out[7061] <= x[5079] ^ x[5080];
     layer0_out[7062] <= x[1029] & x[1031];
     layer0_out[7063] <= ~(x[1410] | x[1412]);
     layer0_out[7064] <= ~(x[5141] & x[5142]);
     layer0_out[7065] <= ~x[3932] | x[3931];
     layer0_out[7066] <= ~(x[3014] & x[3015]);
     layer0_out[7067] <= ~(x[4556] | x[4557]);
     layer0_out[7068] <= ~(x[1506] & x[1508]);
     layer0_out[7069] <= x[573] | x[574];
     layer0_out[7070] <= ~x[364];
     layer0_out[7071] <= ~(x[6259] & x[6260]);
     layer0_out[7072] <= 1'b0;
     layer0_out[7073] <= x[424];
     layer0_out[7074] <= ~x[1219];
     layer0_out[7075] <= ~(x[1555] | x[1557]);
     layer0_out[7076] <= ~x[7220];
     layer0_out[7077] <= x[2149] ^ x[2150];
     layer0_out[7078] <= x[2618] ^ x[2620];
     layer0_out[7079] <= ~(x[6794] | x[6795]);
     layer0_out[7080] <= x[7645] | x[7646];
     layer0_out[7081] <= x[8547] | x[8548];
     layer0_out[7082] <= x[4897] & x[4898];
     layer0_out[7083] <= ~(x[953] | x[954]);
     layer0_out[7084] <= ~(x[269] | x[271]);
     layer0_out[7085] <= x[5664] | x[5665];
     layer0_out[7086] <= ~x[3325] | x[3326];
     layer0_out[7087] <= ~x[2706];
     layer0_out[7088] <= x[7637] | x[7638];
     layer0_out[7089] <= 1'b0;
     layer0_out[7090] <= x[8308] & x[8309];
     layer0_out[7091] <= x[3270] & x[3271];
     layer0_out[7092] <= ~(x[1119] & x[1120]);
     layer0_out[7093] <= x[6606];
     layer0_out[7094] <= 1'b1;
     layer0_out[7095] <= ~(x[8400] ^ x[8401]);
     layer0_out[7096] <= 1'b1;
     layer0_out[7097] <= ~x[1335];
     layer0_out[7098] <= ~(x[1388] & x[1390]);
     layer0_out[7099] <= x[524];
     layer0_out[7100] <= ~(x[8459] | x[8460]);
     layer0_out[7101] <= x[4891];
     layer0_out[7102] <= x[1462];
     layer0_out[7103] <= x[2071] & ~x[2072];
     layer0_out[7104] <= x[2847] ^ x[2848];
     layer0_out[7105] <= x[9000];
     layer0_out[7106] <= x[5177];
     layer0_out[7107] <= ~(x[7981] | x[7982]);
     layer0_out[7108] <= x[7344] | x[7345];
     layer0_out[7109] <= x[1040];
     layer0_out[7110] <= ~(x[4694] & x[4695]);
     layer0_out[7111] <= x[58] & x[59];
     layer0_out[7112] <= ~(x[3492] & x[3493]);
     layer0_out[7113] <= ~(x[6470] | x[6471]);
     layer0_out[7114] <= x[6651] & x[6652];
     layer0_out[7115] <= x[3909] & x[3910];
     layer0_out[7116] <= ~(x[7919] | x[7920]);
     layer0_out[7117] <= ~(x[3011] | x[3012]);
     layer0_out[7118] <= x[4509] | x[4510];
     layer0_out[7119] <= ~(x[8517] ^ x[8518]);
     layer0_out[7120] <= x[3212] & ~x[3211];
     layer0_out[7121] <= x[1672] | x[1673];
     layer0_out[7122] <= ~x[881];
     layer0_out[7123] <= x[1979] & x[1981];
     layer0_out[7124] <= ~(x[4296] & x[4297]);
     layer0_out[7125] <= 1'b0;
     layer0_out[7126] <= x[2783] & x[2785];
     layer0_out[7127] <= 1'b1;
     layer0_out[7128] <= 1'b0;
     layer0_out[7129] <= x[338] & x[340];
     layer0_out[7130] <= ~(x[4447] ^ x[4448]);
     layer0_out[7131] <= x[6342] | x[6343];
     layer0_out[7132] <= x[726] | x[728];
     layer0_out[7133] <= 1'b1;
     layer0_out[7134] <= x[561] & x[562];
     layer0_out[7135] <= x[606] & x[608];
     layer0_out[7136] <= x[2965] & x[2966];
     layer0_out[7137] <= ~(x[8679] ^ x[8680]);
     layer0_out[7138] <= x[736] | x[738];
     layer0_out[7139] <= ~(x[2588] | x[2589]);
     layer0_out[7140] <= x[1797] & x[1799];
     layer0_out[7141] <= ~(x[1607] & x[1609]);
     layer0_out[7142] <= ~x[8386];
     layer0_out[7143] <= x[7795] & x[7796];
     layer0_out[7144] <= x[2411] & x[2413];
     layer0_out[7145] <= ~(x[1167] & x[1169]);
     layer0_out[7146] <= ~(x[3472] ^ x[3473]);
     layer0_out[7147] <= x[1123] & x[1125];
     layer0_out[7148] <= ~(x[8846] | x[8847]);
     layer0_out[7149] <= x[1505] & x[1507];
     layer0_out[7150] <= x[3078];
     layer0_out[7151] <= ~(x[1585] & x[1587]);
     layer0_out[7152] <= ~x[8025] | x[8024];
     layer0_out[7153] <= x[8901] | x[8902];
     layer0_out[7154] <= ~(x[7469] & x[7470]);
     layer0_out[7155] <= ~(x[1270] & x[1272]);
     layer0_out[7156] <= ~(x[4372] & x[4373]);
     layer0_out[7157] <= ~(x[5088] ^ x[5089]);
     layer0_out[7158] <= x[163] & ~x[164];
     layer0_out[7159] <= ~x[4822] | x[4823];
     layer0_out[7160] <= ~(x[4678] & x[4679]);
     layer0_out[7161] <= x[1612];
     layer0_out[7162] <= 1'b0;
     layer0_out[7163] <= x[849] | x[851];
     layer0_out[7164] <= x[6083] & x[6084];
     layer0_out[7165] <= ~x[7908] | x[7907];
     layer0_out[7166] <= ~(x[5897] & x[5898]);
     layer0_out[7167] <= ~(x[5661] & x[5662]);
     layer0_out[7168] <= ~(x[6510] | x[6511]);
     layer0_out[7169] <= x[317] | x[319];
     layer0_out[7170] <= x[760] | x[761];
     layer0_out[7171] <= x[5537];
     layer0_out[7172] <= ~(x[2958] ^ x[2959]);
     layer0_out[7173] <= 1'b0;
     layer0_out[7174] <= x[4386] & x[4387];
     layer0_out[7175] <= ~(x[1360] & x[1362]);
     layer0_out[7176] <= x[3475] ^ x[3476];
     layer0_out[7177] <= ~(x[6490] & x[6491]);
     layer0_out[7178] <= x[2777] ^ x[2779];
     layer0_out[7179] <= x[3511];
     layer0_out[7180] <= ~(x[5703] ^ x[5704]);
     layer0_out[7181] <= x[2775] & x[2776];
     layer0_out[7182] <= x[153] ^ x[154];
     layer0_out[7183] <= x[941];
     layer0_out[7184] <= ~x[3693];
     layer0_out[7185] <= x[5815];
     layer0_out[7186] <= x[8136] ^ x[8137];
     layer0_out[7187] <= x[3009];
     layer0_out[7188] <= ~(x[1044] | x[1045]);
     layer0_out[7189] <= ~x[5076] | x[5077];
     layer0_out[7190] <= ~(x[1638] ^ x[1639]);
     layer0_out[7191] <= ~x[6974];
     layer0_out[7192] <= x[3116] & x[3117];
     layer0_out[7193] <= x[2891] ^ x[2892];
     layer0_out[7194] <= x[6397];
     layer0_out[7195] <= x[1011] & ~x[1013];
     layer0_out[7196] <= ~(x[1517] & x[1519]);
     layer0_out[7197] <= ~x[4145];
     layer0_out[7198] <= x[8679];
     layer0_out[7199] <= ~x[7840];
     layer0_out[7200] <= ~(x[6694] | x[6695]);
     layer0_out[7201] <= x[9045];
     layer0_out[7202] <= ~x[767];
     layer0_out[7203] <= x[3431] | x[3432];
     layer0_out[7204] <= ~x[7798];
     layer0_out[7205] <= x[152] & ~x[154];
     layer0_out[7206] <= x[466] | x[468];
     layer0_out[7207] <= ~(x[6537] | x[6538]);
     layer0_out[7208] <= x[8873] | x[8874];
     layer0_out[7209] <= x[6751] ^ x[6752];
     layer0_out[7210] <= x[4861] & x[4862];
     layer0_out[7211] <= ~(x[8094] & x[8095]);
     layer0_out[7212] <= ~(x[1902] & x[1904]);
     layer0_out[7213] <= ~(x[179] ^ x[181]);
     layer0_out[7214] <= ~(x[2532] ^ x[2534]);
     layer0_out[7215] <= x[1476] & x[1477];
     layer0_out[7216] <= x[2553] & x[2554];
     layer0_out[7217] <= x[6252] | x[6253];
     layer0_out[7218] <= ~(x[8050] ^ x[8051]);
     layer0_out[7219] <= ~(x[2805] ^ x[2806]);
     layer0_out[7220] <= ~x[8247] | x[8248];
     layer0_out[7221] <= ~(x[828] | x[830]);
     layer0_out[7222] <= x[4223] | x[4224];
     layer0_out[7223] <= ~(x[7057] & x[7058]);
     layer0_out[7224] <= ~(x[4998] ^ x[4999]);
     layer0_out[7225] <= ~(x[8813] ^ x[8814]);
     layer0_out[7226] <= ~(x[1215] & x[1216]);
     layer0_out[7227] <= ~x[5877];
     layer0_out[7228] <= x[5944] & x[5945];
     layer0_out[7229] <= ~x[1619];
     layer0_out[7230] <= x[6239] | x[6240];
     layer0_out[7231] <= x[2868] | x[2869];
     layer0_out[7232] <= x[5006] | x[5007];
     layer0_out[7233] <= ~x[305];
     layer0_out[7234] <= x[1017] | x[1018];
     layer0_out[7235] <= x[2753];
     layer0_out[7236] <= x[9191];
     layer0_out[7237] <= x[7246] ^ x[7247];
     layer0_out[7238] <= x[632];
     layer0_out[7239] <= ~(x[6926] | x[6927]);
     layer0_out[7240] <= x[6037] & ~x[6036];
     layer0_out[7241] <= ~(x[5490] & x[5491]);
     layer0_out[7242] <= 1'b1;
     layer0_out[7243] <= x[2013] & x[2015];
     layer0_out[7244] <= x[7407] | x[7408];
     layer0_out[7245] <= ~x[4906] | x[4905];
     layer0_out[7246] <= x[2016] & x[2018];
     layer0_out[7247] <= x[3025] | x[3026];
     layer0_out[7248] <= x[2192] & x[2193];
     layer0_out[7249] <= ~(x[2857] ^ x[2858]);
     layer0_out[7250] <= ~(x[6521] | x[6522]);
     layer0_out[7251] <= x[7590];
     layer0_out[7252] <= x[5284] & x[5285];
     layer0_out[7253] <= x[2761] ^ x[2763];
     layer0_out[7254] <= ~(x[6787] & x[6788]);
     layer0_out[7255] <= ~(x[2086] & x[2088]);
     layer0_out[7256] <= ~(x[1102] & x[1103]);
     layer0_out[7257] <= x[5678] & x[5679];
     layer0_out[7258] <= ~(x[8652] | x[8653]);
     layer0_out[7259] <= 1'b1;
     layer0_out[7260] <= ~x[7395];
     layer0_out[7261] <= ~(x[2051] & x[2053]);
     layer0_out[7262] <= x[38] ^ x[40];
     layer0_out[7263] <= ~x[3215];
     layer0_out[7264] <= x[4842];
     layer0_out[7265] <= ~(x[5881] & x[5882]);
     layer0_out[7266] <= x[2607] & x[2609];
     layer0_out[7267] <= 1'b0;
     layer0_out[7268] <= x[4709] & x[4710];
     layer0_out[7269] <= x[7805] ^ x[7806];
     layer0_out[7270] <= 1'b0;
     layer0_out[7271] <= x[188];
     layer0_out[7272] <= x[8110] | x[8111];
     layer0_out[7273] <= ~(x[6994] | x[6995]);
     layer0_out[7274] <= x[843] ^ x[845];
     layer0_out[7275] <= x[2447] ^ x[2448];
     layer0_out[7276] <= x[3470] | x[3471];
     layer0_out[7277] <= x[1340] ^ x[1342];
     layer0_out[7278] <= x[8501];
     layer0_out[7279] <= ~x[394];
     layer0_out[7280] <= x[1428] ^ x[1430];
     layer0_out[7281] <= ~(x[3159] | x[3160]);
     layer0_out[7282] <= x[9169] | x[9170];
     layer0_out[7283] <= ~x[7861];
     layer0_out[7284] <= ~x[6485];
     layer0_out[7285] <= x[7789] | x[7790];
     layer0_out[7286] <= x[1751];
     layer0_out[7287] <= 1'b0;
     layer0_out[7288] <= ~(x[4609] | x[4610]);
     layer0_out[7289] <= x[2185] & x[2187];
     layer0_out[7290] <= x[1190] & x[1192];
     layer0_out[7291] <= 1'b1;
     layer0_out[7292] <= ~x[7997] | x[7996];
     layer0_out[7293] <= x[2750] ^ x[2751];
     layer0_out[7294] <= x[5255] | x[5256];
     layer0_out[7295] <= x[4903] ^ x[4904];
     layer0_out[7296] <= x[308] & ~x[310];
     layer0_out[7297] <= x[840] | x[842];
     layer0_out[7298] <= ~(x[8502] | x[8503]);
     layer0_out[7299] <= x[7425] & ~x[7426];
     layer0_out[7300] <= x[1153] & x[1155];
     layer0_out[7301] <= ~x[7670];
     layer0_out[7302] <= x[4639];
     layer0_out[7303] <= x[616];
     layer0_out[7304] <= ~(x[2565] & x[2566]);
     layer0_out[7305] <= x[723];
     layer0_out[7306] <= x[4649] ^ x[4650];
     layer0_out[7307] <= x[6693];
     layer0_out[7308] <= ~x[23];
     layer0_out[7309] <= x[1420] & x[1422];
     layer0_out[7310] <= x[4469] | x[4470];
     layer0_out[7311] <= ~x[9185];
     layer0_out[7312] <= ~(x[5789] & x[5790]);
     layer0_out[7313] <= 1'b1;
     layer0_out[7314] <= ~(x[800] | x[802]);
     layer0_out[7315] <= ~(x[7248] | x[7249]);
     layer0_out[7316] <= ~(x[3195] | x[3196]);
     layer0_out[7317] <= x[6042] & x[6043];
     layer0_out[7318] <= ~(x[4034] | x[4035]);
     layer0_out[7319] <= ~x[2616] | x[2617];
     layer0_out[7320] <= ~(x[2241] & x[2242]);
     layer0_out[7321] <= x[3410] | x[3411];
     layer0_out[7322] <= ~x[8756] | x[8757];
     layer0_out[7323] <= x[31] | x[33];
     layer0_out[7324] <= x[1862] | x[1863];
     layer0_out[7325] <= x[2223];
     layer0_out[7326] <= ~x[646];
     layer0_out[7327] <= x[2020] & x[2021];
     layer0_out[7328] <= x[2614] & x[2615];
     layer0_out[7329] <= x[6220];
     layer0_out[7330] <= ~x[6353];
     layer0_out[7331] <= x[6849] & ~x[6850];
     layer0_out[7332] <= x[9061] | x[9062];
     layer0_out[7333] <= ~(x[1021] & x[1022]);
     layer0_out[7334] <= ~x[3223];
     layer0_out[7335] <= x[1537];
     layer0_out[7336] <= x[2740] & x[2742];
     layer0_out[7337] <= ~x[1979];
     layer0_out[7338] <= ~(x[9051] ^ x[9052]);
     layer0_out[7339] <= ~x[3854];
     layer0_out[7340] <= ~x[1977] | x[1979];
     layer0_out[7341] <= ~x[3787] | x[3786];
     layer0_out[7342] <= x[4124] | x[4125];
     layer0_out[7343] <= x[8694] | x[8695];
     layer0_out[7344] <= 1'b1;
     layer0_out[7345] <= ~x[1453];
     layer0_out[7346] <= x[7273];
     layer0_out[7347] <= x[2206] & x[2207];
     layer0_out[7348] <= 1'b0;
     layer0_out[7349] <= ~x[3347];
     layer0_out[7350] <= x[4285] & x[4286];
     layer0_out[7351] <= ~(x[9156] | x[9157]);
     layer0_out[7352] <= ~(x[1386] & x[1387]);
     layer0_out[7353] <= ~(x[7450] & x[7451]);
     layer0_out[7354] <= 1'b0;
     layer0_out[7355] <= ~(x[4944] ^ x[4945]);
     layer0_out[7356] <= 1'b0;
     layer0_out[7357] <= ~x[988];
     layer0_out[7358] <= ~x[3529];
     layer0_out[7359] <= ~(x[4205] & x[4206]);
     layer0_out[7360] <= x[881] | x[882];
     layer0_out[7361] <= x[1262] & x[1264];
     layer0_out[7362] <= x[1243];
     layer0_out[7363] <= x[1416] & x[1418];
     layer0_out[7364] <= x[8213] & x[8214];
     layer0_out[7365] <= ~(x[8910] | x[8911]);
     layer0_out[7366] <= ~(x[7543] ^ x[7544]);
     layer0_out[7367] <= x[5151] & x[5152];
     layer0_out[7368] <= x[3805] & x[3806];
     layer0_out[7369] <= x[863] ^ x[865];
     layer0_out[7370] <= x[9109] & x[9110];
     layer0_out[7371] <= x[711] | x[713];
     layer0_out[7372] <= 1'b1;
     layer0_out[7373] <= ~(x[4221] & x[4222]);
     layer0_out[7374] <= ~(x[46] | x[47]);
     layer0_out[7375] <= ~x[3627];
     layer0_out[7376] <= x[2648] & ~x[2650];
     layer0_out[7377] <= ~(x[4300] & x[4301]);
     layer0_out[7378] <= x[6052] & x[6053];
     layer0_out[7379] <= x[6552];
     layer0_out[7380] <= ~(x[8179] & x[8180]);
     layer0_out[7381] <= x[786] & x[787];
     layer0_out[7382] <= ~(x[2136] ^ x[2138]);
     layer0_out[7383] <= x[7124] & x[7125];
     layer0_out[7384] <= ~(x[4160] | x[4161]);
     layer0_out[7385] <= ~x[596];
     layer0_out[7386] <= x[6516] | x[6517];
     layer0_out[7387] <= x[4030];
     layer0_out[7388] <= x[796] | x[797];
     layer0_out[7389] <= x[9078] & ~x[9077];
     layer0_out[7390] <= x[2781] ^ x[2782];
     layer0_out[7391] <= ~(x[1324] & x[1325]);
     layer0_out[7392] <= ~x[626];
     layer0_out[7393] <= ~(x[196] | x[198]);
     layer0_out[7394] <= ~(x[4749] | x[4750]);
     layer0_out[7395] <= x[3882] | x[3883];
     layer0_out[7396] <= x[1567] & x[1569];
     layer0_out[7397] <= ~(x[2253] & x[2254]);
     layer0_out[7398] <= x[2410] & x[2412];
     layer0_out[7399] <= ~(x[7267] | x[7268]);
     layer0_out[7400] <= ~(x[8637] ^ x[8638]);
     layer0_out[7401] <= x[7848] & ~x[7849];
     layer0_out[7402] <= x[5657] & x[5658];
     layer0_out[7403] <= x[1177];
     layer0_out[7404] <= x[5820] & x[5821];
     layer0_out[7405] <= ~(x[1174] | x[1175]);
     layer0_out[7406] <= x[4675] & ~x[4676];
     layer0_out[7407] <= x[6437] | x[6438];
     layer0_out[7408] <= x[3661] & x[3662];
     layer0_out[7409] <= ~(x[2473] | x[2475]);
     layer0_out[7410] <= ~(x[1042] ^ x[1043]);
     layer0_out[7411] <= x[2546] & x[2548];
     layer0_out[7412] <= x[7142] & ~x[7141];
     layer0_out[7413] <= 1'b0;
     layer0_out[7414] <= ~(x[6139] | x[6140]);
     layer0_out[7415] <= ~(x[2487] & x[2489]);
     layer0_out[7416] <= ~x[6291] | x[6292];
     layer0_out[7417] <= ~x[5782];
     layer0_out[7418] <= 1'b0;
     layer0_out[7419] <= x[7698];
     layer0_out[7420] <= x[3143];
     layer0_out[7421] <= ~x[682];
     layer0_out[7422] <= x[1127] | x[1129];
     layer0_out[7423] <= x[7421] & x[7422];
     layer0_out[7424] <= ~(x[4891] & x[4892]);
     layer0_out[7425] <= ~(x[6008] & x[6009]);
     layer0_out[7426] <= 1'b1;
     layer0_out[7427] <= x[724] & x[726];
     layer0_out[7428] <= ~(x[2521] & x[2522]);
     layer0_out[7429] <= x[4423] ^ x[4424];
     layer0_out[7430] <= ~x[4652] | x[4651];
     layer0_out[7431] <= x[272] & x[274];
     layer0_out[7432] <= ~(x[864] & x[865]);
     layer0_out[7433] <= ~(x[843] | x[844]);
     layer0_out[7434] <= ~(x[8276] ^ x[8277]);
     layer0_out[7435] <= ~(x[7347] ^ x[7348]);
     layer0_out[7436] <= ~x[2065];
     layer0_out[7437] <= x[316] & ~x[315];
     layer0_out[7438] <= x[531] | x[532];
     layer0_out[7439] <= ~(x[1133] & x[1134]);
     layer0_out[7440] <= ~(x[1097] & x[1098]);
     layer0_out[7441] <= ~(x[2128] & x[2129]);
     layer0_out[7442] <= 1'b1;
     layer0_out[7443] <= x[4601] & x[4602];
     layer0_out[7444] <= x[2269];
     layer0_out[7445] <= ~x[5597];
     layer0_out[7446] <= x[855];
     layer0_out[7447] <= x[5825];
     layer0_out[7448] <= x[7298] & x[7299];
     layer0_out[7449] <= x[7135] | x[7136];
     layer0_out[7450] <= x[860] ^ x[862];
     layer0_out[7451] <= ~x[4736];
     layer0_out[7452] <= x[233] & x[235];
     layer0_out[7453] <= ~(x[2831] & x[2832]);
     layer0_out[7454] <= ~(x[2609] & x[2610]);
     layer0_out[7455] <= ~x[1368] | x[1366];
     layer0_out[7456] <= ~(x[1691] & x[1693]);
     layer0_out[7457] <= x[3875] ^ x[3876];
     layer0_out[7458] <= x[5855] ^ x[5856];
     layer0_out[7459] <= x[5911] & x[5912];
     layer0_out[7460] <= x[1034] & x[1036];
     layer0_out[7461] <= x[1329];
     layer0_out[7462] <= x[8839];
     layer0_out[7463] <= ~x[2170];
     layer0_out[7464] <= ~(x[3739] | x[3740]);
     layer0_out[7465] <= x[1649];
     layer0_out[7466] <= ~(x[5907] | x[5908]);
     layer0_out[7467] <= 1'b1;
     layer0_out[7468] <= ~(x[4153] | x[4154]);
     layer0_out[7469] <= x[8393] & x[8394];
     layer0_out[7470] <= x[64] | x[66];
     layer0_out[7471] <= ~(x[4559] | x[4560]);
     layer0_out[7472] <= x[2515] & x[2517];
     layer0_out[7473] <= ~(x[7213] ^ x[7214]);
     layer0_out[7474] <= ~x[456];
     layer0_out[7475] <= x[3070] | x[3071];
     layer0_out[7476] <= x[3382] ^ x[3383];
     layer0_out[7477] <= ~(x[2377] ^ x[2379]);
     layer0_out[7478] <= x[5391];
     layer0_out[7479] <= ~(x[9106] & x[9107]);
     layer0_out[7480] <= x[1906] | x[1908];
     layer0_out[7481] <= ~(x[4392] | x[4393]);
     layer0_out[7482] <= x[3748] & x[3749];
     layer0_out[7483] <= x[1825];
     layer0_out[7484] <= ~(x[1799] & x[1800]);
     layer0_out[7485] <= 1'b0;
     layer0_out[7486] <= x[2601] & x[2602];
     layer0_out[7487] <= x[1235] ^ x[1236];
     layer0_out[7488] <= ~x[1230];
     layer0_out[7489] <= ~x[2624];
     layer0_out[7490] <= x[4701] & x[4702];
     layer0_out[7491] <= ~x[957];
     layer0_out[7492] <= ~(x[8419] ^ x[8420]);
     layer0_out[7493] <= x[848] & x[850];
     layer0_out[7494] <= ~(x[5879] & x[5880]);
     layer0_out[7495] <= ~(x[2204] & x[2206]);
     layer0_out[7496] <= ~(x[2757] & x[2758]);
     layer0_out[7497] <= x[1368] | x[1370];
     layer0_out[7498] <= ~(x[5765] ^ x[5766]);
     layer0_out[7499] <= 1'b0;
     layer0_out[7500] <= ~(x[2569] ^ x[2571]);
     layer0_out[7501] <= ~(x[1930] & x[1932]);
     layer0_out[7502] <= ~(x[2420] & x[2421]);
     layer0_out[7503] <= x[1582] & x[1583];
     layer0_out[7504] <= ~(x[1627] & x[1628]);
     layer0_out[7505] <= ~x[7767] | x[7768];
     layer0_out[7506] <= ~x[7477];
     layer0_out[7507] <= x[1036] | x[1038];
     layer0_out[7508] <= ~(x[586] | x[587]);
     layer0_out[7509] <= ~(x[5540] & x[5541]);
     layer0_out[7510] <= ~(x[2449] & x[2450]);
     layer0_out[7511] <= x[7673];
     layer0_out[7512] <= ~x[4226];
     layer0_out[7513] <= ~(x[9020] | x[9021]);
     layer0_out[7514] <= x[5883] & x[5884];
     layer0_out[7515] <= ~(x[8127] & x[8128]);
     layer0_out[7516] <= ~(x[7170] ^ x[7171]);
     layer0_out[7517] <= 1'b1;
     layer0_out[7518] <= ~(x[3088] | x[3089]);
     layer0_out[7519] <= x[798] & x[799];
     layer0_out[7520] <= x[7539] & ~x[7538];
     layer0_out[7521] <= ~x[780];
     layer0_out[7522] <= x[8687] | x[8688];
     layer0_out[7523] <= x[3557] & ~x[3558];
     layer0_out[7524] <= ~x[868];
     layer0_out[7525] <= 1'b1;
     layer0_out[7526] <= ~(x[3141] | x[3142]);
     layer0_out[7527] <= x[4791];
     layer0_out[7528] <= x[2363];
     layer0_out[7529] <= ~(x[1726] ^ x[1727]);
     layer0_out[7530] <= x[5857] & x[5858];
     layer0_out[7531] <= ~(x[7452] & x[7453]);
     layer0_out[7532] <= ~(x[1525] & x[1527]);
     layer0_out[7533] <= ~(x[1298] & x[1300]);
     layer0_out[7534] <= ~(x[8046] & x[8047]);
     layer0_out[7535] <= ~x[7973];
     layer0_out[7536] <= x[3885] | x[3886];
     layer0_out[7537] <= x[5973] & x[5974];
     layer0_out[7538] <= x[6219] | x[6220];
     layer0_out[7539] <= ~x[637] | x[636];
     layer0_out[7540] <= ~(x[2358] ^ x[2360]);
     layer0_out[7541] <= ~x[2080];
     layer0_out[7542] <= ~(x[6175] ^ x[6176]);
     layer0_out[7543] <= ~x[590];
     layer0_out[7544] <= ~x[6697] | x[6696];
     layer0_out[7545] <= x[1837] & x[1839];
     layer0_out[7546] <= x[7794] ^ x[7795];
     layer0_out[7547] <= x[6925];
     layer0_out[7548] <= ~(x[2623] & x[2624]);
     layer0_out[7549] <= ~x[531];
     layer0_out[7550] <= x[1934] ^ x[1936];
     layer0_out[7551] <= x[5442] ^ x[5443];
     layer0_out[7552] <= ~x[4926] | x[4925];
     layer0_out[7553] <= x[1854] & ~x[1852];
     layer0_out[7554] <= ~(x[6481] | x[6482]);
     layer0_out[7555] <= x[2146] & x[2147];
     layer0_out[7556] <= ~(x[2325] & x[2327]);
     layer0_out[7557] <= x[1320] & x[1321];
     layer0_out[7558] <= ~(x[931] ^ x[932]);
     layer0_out[7559] <= x[6273];
     layer0_out[7560] <= x[352] | x[354];
     layer0_out[7561] <= 1'b0;
     layer0_out[7562] <= ~x[3100];
     layer0_out[7563] <= x[779] ^ x[780];
     layer0_out[7564] <= x[8125] & x[8126];
     layer0_out[7565] <= x[1375] ^ x[1377];
     layer0_out[7566] <= x[831] & x[832];
     layer0_out[7567] <= x[2590] | x[2592];
     layer0_out[7568] <= ~(x[4886] | x[4887]);
     layer0_out[7569] <= x[8848] | x[8849];
     layer0_out[7570] <= ~(x[5909] & x[5910]);
     layer0_out[7571] <= x[5652] & x[5653];
     layer0_out[7572] <= x[4655];
     layer0_out[7573] <= x[2475] & x[2477];
     layer0_out[7574] <= ~(x[8298] & x[8299]);
     layer0_out[7575] <= ~x[2603] | x[2602];
     layer0_out[7576] <= x[1779];
     layer0_out[7577] <= x[1847];
     layer0_out[7578] <= ~(x[2101] | x[2103]);
     layer0_out[7579] <= x[4471] & x[4472];
     layer0_out[7580] <= ~(x[1941] | x[1942]);
     layer0_out[7581] <= ~x[1271];
     layer0_out[7582] <= ~(x[1989] & x[1990]);
     layer0_out[7583] <= ~(x[8003] & x[8004]);
     layer0_out[7584] <= ~(x[797] | x[798]);
     layer0_out[7585] <= ~(x[2191] | x[2193]);
     layer0_out[7586] <= ~(x[7080] | x[7081]);
     layer0_out[7587] <= x[1188] ^ x[1189];
     layer0_out[7588] <= ~(x[4145] | x[4146]);
     layer0_out[7589] <= x[1315];
     layer0_out[7590] <= x[1191];
     layer0_out[7591] <= ~(x[1353] ^ x[1355]);
     layer0_out[7592] <= x[1732] & x[1733];
     layer0_out[7593] <= x[450];
     layer0_out[7594] <= ~x[1749];
     layer0_out[7595] <= ~x[2437] | x[2438];
     layer0_out[7596] <= x[1777] | x[1779];
     layer0_out[7597] <= x[574] | x[575];
     layer0_out[7598] <= x[8522] | x[8523];
     layer0_out[7599] <= x[5114] & ~x[5113];
     layer0_out[7600] <= ~(x[848] & x[849]);
     layer0_out[7601] <= ~x[8335];
     layer0_out[7602] <= x[4192] & ~x[4193];
     layer0_out[7603] <= x[3174] & x[3175];
     layer0_out[7604] <= ~x[2473];
     layer0_out[7605] <= ~(x[5600] & x[5601]);
     layer0_out[7606] <= ~x[1910];
     layer0_out[7607] <= x[1597] ^ x[1599];
     layer0_out[7608] <= ~(x[784] & x[785]);
     layer0_out[7609] <= x[3282] & x[3283];
     layer0_out[7610] <= ~x[5869];
     layer0_out[7611] <= x[3960] | x[3961];
     layer0_out[7612] <= ~(x[1674] ^ x[1676]);
     layer0_out[7613] <= x[4179] & x[4180];
     layer0_out[7614] <= x[6652] | x[6653];
     layer0_out[7615] <= x[1317] & x[1318];
     layer0_out[7616] <= x[6937] & x[6938];
     layer0_out[7617] <= ~(x[1639] & x[1641]);
     layer0_out[7618] <= x[1075] & x[1077];
     layer0_out[7619] <= ~(x[5663] | x[5664]);
     layer0_out[7620] <= 1'b1;
     layer0_out[7621] <= ~x[4190];
     layer0_out[7622] <= ~x[1889];
     layer0_out[7623] <= 1'b0;
     layer0_out[7624] <= x[1414] & ~x[1415];
     layer0_out[7625] <= ~(x[6569] | x[6570]);
     layer0_out[7626] <= x[1099];
     layer0_out[7627] <= x[1905] & x[1906];
     layer0_out[7628] <= x[7967] & ~x[7968];
     layer0_out[7629] <= ~(x[531] & x[533]);
     layer0_out[7630] <= ~(x[7078] | x[7079]);
     layer0_out[7631] <= x[4057];
     layer0_out[7632] <= ~(x[1227] & x[1229]);
     layer0_out[7633] <= x[9122] ^ x[9123];
     layer0_out[7634] <= ~(x[126] & x[128]);
     layer0_out[7635] <= ~x[2149] | x[2148];
     layer0_out[7636] <= ~x[1497];
     layer0_out[7637] <= x[6636] ^ x[6637];
     layer0_out[7638] <= ~x[1790];
     layer0_out[7639] <= ~x[6318];
     layer0_out[7640] <= ~(x[444] ^ x[446]);
     layer0_out[7641] <= ~(x[2327] & x[2328]);
     layer0_out[7642] <= x[2477];
     layer0_out[7643] <= ~(x[2490] | x[2491]);
     layer0_out[7644] <= ~(x[629] ^ x[630]);
     layer0_out[7645] <= x[2434] & ~x[2433];
     layer0_out[7646] <= x[5994] | x[5995];
     layer0_out[7647] <= ~(x[7937] | x[7938]);
     layer0_out[7648] <= x[1983] & x[1985];
     layer0_out[7649] <= x[6171];
     layer0_out[7650] <= ~x[3268];
     layer0_out[7651] <= x[220] ^ x[221];
     layer0_out[7652] <= ~x[7200];
     layer0_out[7653] <= x[5698] | x[5699];
     layer0_out[7654] <= ~x[2003];
     layer0_out[7655] <= x[5923] & x[5924];
     layer0_out[7656] <= x[4064] | x[4065];
     layer0_out[7657] <= x[7180] ^ x[7181];
     layer0_out[7658] <= x[1652] & x[1653];
     layer0_out[7659] <= ~x[6077];
     layer0_out[7660] <= x[8076] | x[8077];
     layer0_out[7661] <= ~x[4416];
     layer0_out[7662] <= ~(x[8200] | x[8201]);
     layer0_out[7663] <= x[2766] ^ x[2768];
     layer0_out[7664] <= ~(x[8500] ^ x[8501]);
     layer0_out[7665] <= x[1251] & ~x[1252];
     layer0_out[7666] <= x[4091] & x[4092];
     layer0_out[7667] <= ~x[8413];
     layer0_out[7668] <= x[744] | x[746];
     layer0_out[7669] <= x[356] & x[358];
     layer0_out[7670] <= x[8504];
     layer0_out[7671] <= ~(x[773] & x[774]);
     layer0_out[7672] <= x[6197];
     layer0_out[7673] <= x[3975] & ~x[3976];
     layer0_out[7674] <= x[8331] & x[8332];
     layer0_out[7675] <= ~(x[3183] | x[3184]);
     layer0_out[7676] <= x[4994] ^ x[4995];
     layer0_out[7677] <= ~(x[987] & x[989]);
     layer0_out[7678] <= x[6406] ^ x[6407];
     layer0_out[7679] <= ~x[3642] | x[3643];
     layer0_out[7680] <= x[2498] & x[2499];
     layer0_out[7681] <= ~(x[7680] ^ x[7681]);
     layer0_out[7682] <= ~(x[5730] ^ x[5731]);
     layer0_out[7683] <= x[1407] & x[1408];
     layer0_out[7684] <= x[67] & x[68];
     layer0_out[7685] <= ~(x[2399] & x[2400]);
     layer0_out[7686] <= x[5047] ^ x[5048];
     layer0_out[7687] <= ~x[6368];
     layer0_out[7688] <= ~x[4833];
     layer0_out[7689] <= 1'b1;
     layer0_out[7690] <= x[6497] | x[6498];
     layer0_out[7691] <= x[1083] | x[1084];
     layer0_out[7692] <= ~x[1066];
     layer0_out[7693] <= x[8130] & x[8131];
     layer0_out[7694] <= x[2450] & x[2451];
     layer0_out[7695] <= x[6287] ^ x[6288];
     layer0_out[7696] <= x[8064] | x[8065];
     layer0_out[7697] <= ~(x[3672] ^ x[3673]);
     layer0_out[7698] <= ~(x[9053] | x[9054]);
     layer0_out[7699] <= ~(x[6745] | x[6746]);
     layer0_out[7700] <= x[686];
     layer0_out[7701] <= ~(x[611] ^ x[613]);
     layer0_out[7702] <= ~(x[8635] | x[8636]);
     layer0_out[7703] <= ~(x[5602] & x[5603]);
     layer0_out[7704] <= ~(x[2002] | x[2003]);
     layer0_out[7705] <= x[1110];
     layer0_out[7706] <= ~(x[6746] ^ x[6747]);
     layer0_out[7707] <= x[509];
     layer0_out[7708] <= ~(x[6752] & x[6753]);
     layer0_out[7709] <= ~(x[2689] & x[2690]);
     layer0_out[7710] <= x[6826];
     layer0_out[7711] <= x[6669] & x[6670];
     layer0_out[7712] <= ~(x[642] & x[644]);
     layer0_out[7713] <= ~(x[887] & x[888]);
     layer0_out[7714] <= x[2697] & ~x[2695];
     layer0_out[7715] <= x[1293] & x[1295];
     layer0_out[7716] <= x[2632] & x[2634];
     layer0_out[7717] <= 1'b0;
     layer0_out[7718] <= x[5793] & x[5794];
     layer0_out[7719] <= x[7563] | x[7564];
     layer0_out[7720] <= x[1654] | x[1655];
     layer0_out[7721] <= x[2811];
     layer0_out[7722] <= x[4800] | x[4801];
     layer0_out[7723] <= ~(x[2100] & x[2102]);
     layer0_out[7724] <= x[6254] | x[6255];
     layer0_out[7725] <= x[1278] | x[1279];
     layer0_out[7726] <= x[6840] ^ x[6841];
     layer0_out[7727] <= x[8686] | x[8687];
     layer0_out[7728] <= x[2334] & x[2335];
     layer0_out[7729] <= 1'b1;
     layer0_out[7730] <= ~(x[1009] ^ x[1011]);
     layer0_out[7731] <= x[4997] | x[4998];
     layer0_out[7732] <= ~x[2618];
     layer0_out[7733] <= x[8880] | x[8881];
     layer0_out[7734] <= x[8587] ^ x[8588];
     layer0_out[7735] <= ~(x[48] & x[49]);
     layer0_out[7736] <= ~(x[2481] & x[2482]);
     layer0_out[7737] <= x[5450];
     layer0_out[7738] <= ~(x[1967] ^ x[1968]);
     layer0_out[7739] <= ~(x[8154] | x[8155]);
     layer0_out[7740] <= x[1473] & x[1474];
     layer0_out[7741] <= ~(x[1425] & x[1427]);
     layer0_out[7742] <= x[4954] | x[4955];
     layer0_out[7743] <= x[4545] ^ x[4546];
     layer0_out[7744] <= x[819];
     layer0_out[7745] <= x[1850] & x[1851];
     layer0_out[7746] <= x[6383] ^ x[6384];
     layer0_out[7747] <= x[8963] | x[8964];
     layer0_out[7748] <= x[5172] & x[5173];
     layer0_out[7749] <= ~x[1359] | x[1358];
     layer0_out[7750] <= x[5863] ^ x[5864];
     layer0_out[7751] <= x[2368];
     layer0_out[7752] <= ~(x[7612] | x[7613]);
     layer0_out[7753] <= x[8486];
     layer0_out[7754] <= ~(x[2656] | x[2657]);
     layer0_out[7755] <= 1'b1;
     layer0_out[7756] <= x[790] & x[791];
     layer0_out[7757] <= ~x[3807] | x[3806];
     layer0_out[7758] <= x[3839] ^ x[3840];
     layer0_out[7759] <= x[7202] & ~x[7203];
     layer0_out[7760] <= ~(x[331] & x[332]);
     layer0_out[7761] <= x[66] | x[68];
     layer0_out[7762] <= ~(x[7834] & x[7835]);
     layer0_out[7763] <= ~(x[2183] & x[2185]);
     layer0_out[7764] <= x[4077] & x[4078];
     layer0_out[7765] <= ~(x[4959] ^ x[4960]);
     layer0_out[7766] <= x[2076] & x[2078];
     layer0_out[7767] <= ~x[661];
     layer0_out[7768] <= x[4899] & x[4900];
     layer0_out[7769] <= x[473] ^ x[475];
     layer0_out[7770] <= ~(x[6124] & x[6125]);
     layer0_out[7771] <= x[4616] & x[4617];
     layer0_out[7772] <= x[2162] ^ x[2163];
     layer0_out[7773] <= x[8807] ^ x[8808];
     layer0_out[7774] <= ~(x[1169] & x[1170]);
     layer0_out[7775] <= ~(x[1984] | x[1985]);
     layer0_out[7776] <= ~x[6561];
     layer0_out[7777] <= x[3847];
     layer0_out[7778] <= ~(x[8545] & x[8546]);
     layer0_out[7779] <= x[4323] | x[4324];
     layer0_out[7780] <= ~(x[8680] | x[8681]);
     layer0_out[7781] <= x[4379] & x[4380];
     layer0_out[7782] <= 1'b0;
     layer0_out[7783] <= x[5156] & x[5157];
     layer0_out[7784] <= ~(x[4322] ^ x[4323]);
     layer0_out[7785] <= x[6930];
     layer0_out[7786] <= ~(x[5001] | x[5002]);
     layer0_out[7787] <= ~x[4628] | x[4629];
     layer0_out[7788] <= x[7646] | x[7647];
     layer0_out[7789] <= ~(x[659] & x[661]);
     layer0_out[7790] <= x[6789];
     layer0_out[7791] <= ~(x[6347] | x[6348]);
     layer0_out[7792] <= x[1433] | x[1434];
     layer0_out[7793] <= x[8036] & ~x[8037];
     layer0_out[7794] <= x[1943] ^ x[1944];
     layer0_out[7795] <= ~(x[7077] | x[7078]);
     layer0_out[7796] <= ~x[8991];
     layer0_out[7797] <= ~x[2549] | x[2548];
     layer0_out[7798] <= ~x[6155];
     layer0_out[7799] <= x[6495] | x[6496];
     layer0_out[7800] <= ~(x[8093] ^ x[8094]);
     layer0_out[7801] <= ~x[4309];
     layer0_out[7802] <= ~(x[553] | x[555]);
     layer0_out[7803] <= x[5705] & x[5706];
     layer0_out[7804] <= x[7873];
     layer0_out[7805] <= ~x[2871];
     layer0_out[7806] <= x[3430] ^ x[3431];
     layer0_out[7807] <= x[30] ^ x[31];
     layer0_out[7808] <= ~(x[5880] & x[5881]);
     layer0_out[7809] <= 1'b0;
     layer0_out[7810] <= x[6112] & x[6113];
     layer0_out[7811] <= x[2734] & ~x[2733];
     layer0_out[7812] <= ~x[4543] | x[4542];
     layer0_out[7813] <= x[7679] & x[7680];
     layer0_out[7814] <= x[8632] | x[8633];
     layer0_out[7815] <= ~(x[2526] | x[2528]);
     layer0_out[7816] <= x[4806] & x[4807];
     layer0_out[7817] <= ~(x[7978] ^ x[7979]);
     layer0_out[7818] <= x[1453] & x[1455];
     layer0_out[7819] <= x[7309];
     layer0_out[7820] <= ~(x[781] & x[783]);
     layer0_out[7821] <= 1'b0;
     layer0_out[7822] <= x[4233];
     layer0_out[7823] <= ~x[6590] | x[6589];
     layer0_out[7824] <= ~(x[622] ^ x[624]);
     layer0_out[7825] <= x[1932] ^ x[1933];
     layer0_out[7826] <= x[3225] | x[3226];
     layer0_out[7827] <= 1'b1;
     layer0_out[7828] <= ~(x[2942] & x[2943]);
     layer0_out[7829] <= ~(x[2568] & x[2570]);
     layer0_out[7830] <= x[1725] ^ x[1726];
     layer0_out[7831] <= x[7891] ^ x[7892];
     layer0_out[7832] <= ~(x[1763] & x[1764]);
     layer0_out[7833] <= x[2679] & x[2680];
     layer0_out[7834] <= ~(x[1804] | x[1806]);
     layer0_out[7835] <= x[1768] & x[1770];
     layer0_out[7836] <= ~x[7741];
     layer0_out[7837] <= ~(x[1009] & x[1010]);
     layer0_out[7838] <= x[693] | x[694];
     layer0_out[7839] <= ~(x[8718] | x[8719]);
     layer0_out[7840] <= ~x[6509];
     layer0_out[7841] <= x[5527] & x[5528];
     layer0_out[7842] <= ~x[8518] | x[8519];
     layer0_out[7843] <= x[2429] & ~x[2428];
     layer0_out[7844] <= 1'b0;
     layer0_out[7845] <= 1'b1;
     layer0_out[7846] <= x[1531] ^ x[1533];
     layer0_out[7847] <= x[7316];
     layer0_out[7848] <= ~(x[6688] & x[6689]);
     layer0_out[7849] <= x[1090];
     layer0_out[7850] <= ~(x[1468] & x[1469]);
     layer0_out[7851] <= x[5942] & x[5943];
     layer0_out[7852] <= x[696] & x[698];
     layer0_out[7853] <= ~(x[4107] & x[4108]);
     layer0_out[7854] <= ~(x[9136] ^ x[9137]);
     layer0_out[7855] <= x[2444] & x[2445];
     layer0_out[7856] <= 1'b1;
     layer0_out[7857] <= ~(x[6101] & x[6102]);
     layer0_out[7858] <= x[2559] ^ x[2561];
     layer0_out[7859] <= ~(x[3467] & x[3468]);
     layer0_out[7860] <= ~(x[6103] | x[6104]);
     layer0_out[7861] <= ~(x[5070] ^ x[5071]);
     layer0_out[7862] <= ~(x[3897] | x[3898]);
     layer0_out[7863] <= ~(x[2009] | x[2010]);
     layer0_out[7864] <= 1'b1;
     layer0_out[7865] <= x[5356] & x[5357];
     layer0_out[7866] <= x[7564] | x[7565];
     layer0_out[7867] <= x[16] & x[17];
     layer0_out[7868] <= x[7720] & x[7721];
     layer0_out[7869] <= ~(x[2651] ^ x[2653]);
     layer0_out[7870] <= ~(x[6256] | x[6257]);
     layer0_out[7871] <= x[6979];
     layer0_out[7872] <= ~(x[1570] & x[1571]);
     layer0_out[7873] <= 1'b0;
     layer0_out[7874] <= x[62] & x[63];
     layer0_out[7875] <= ~(x[6793] & x[6794]);
     layer0_out[7876] <= x[6744];
     layer0_out[7877] <= ~x[2752] | x[2751];
     layer0_out[7878] <= 1'b0;
     layer0_out[7879] <= ~(x[1618] & x[1620]);
     layer0_out[7880] <= ~x[5932] | x[5931];
     layer0_out[7881] <= ~(x[1816] | x[1817]);
     layer0_out[7882] <= ~(x[429] & x[431]);
     layer0_out[7883] <= x[905] & x[906];
     layer0_out[7884] <= x[962];
     layer0_out[7885] <= ~(x[685] & x[687]);
     layer0_out[7886] <= x[8856];
     layer0_out[7887] <= x[1647];
     layer0_out[7888] <= x[8619];
     layer0_out[7889] <= ~x[3634];
     layer0_out[7890] <= x[1231] | x[1233];
     layer0_out[7891] <= x[1749] ^ x[1750];
     layer0_out[7892] <= x[3533] & x[3534];
     layer0_out[7893] <= ~(x[2557] | x[2558]);
     layer0_out[7894] <= ~(x[3974] | x[3975]);
     layer0_out[7895] <= ~(x[6834] & x[6835]);
     layer0_out[7896] <= 1'b1;
     layer0_out[7897] <= ~x[5804];
     layer0_out[7898] <= ~(x[7483] & x[7484]);
     layer0_out[7899] <= x[4206] & x[4207];
     layer0_out[7900] <= ~(x[4401] | x[4402]);
     layer0_out[7901] <= x[5406] & x[5407];
     layer0_out[7902] <= x[6216] ^ x[6217];
     layer0_out[7903] <= ~(x[4208] & x[4209]);
     layer0_out[7904] <= ~(x[8520] | x[8521]);
     layer0_out[7905] <= x[7500] | x[7501];
     layer0_out[7906] <= x[2254] ^ x[2256];
     layer0_out[7907] <= x[1104] | x[1105];
     layer0_out[7908] <= x[652] | x[653];
     layer0_out[7909] <= ~(x[6942] | x[6943]);
     layer0_out[7910] <= ~(x[56] | x[57]);
     layer0_out[7911] <= ~(x[5068] & x[5069]);
     layer0_out[7912] <= x[8343] | x[8344];
     layer0_out[7913] <= x[3287] & ~x[3286];
     layer0_out[7914] <= x[1761] | x[1763];
     layer0_out[7915] <= x[980] | x[982];
     layer0_out[7916] <= ~(x[1978] & x[1979]);
     layer0_out[7917] <= ~(x[973] | x[975]);
     layer0_out[7918] <= x[515] & x[516];
     layer0_out[7919] <= ~x[1620];
     layer0_out[7920] <= ~(x[1735] | x[1737]);
     layer0_out[7921] <= x[8214] ^ x[8215];
     layer0_out[7922] <= x[6613];
     layer0_out[7923] <= x[391] & ~x[390];
     layer0_out[7924] <= ~(x[7985] | x[7986]);
     layer0_out[7925] <= 1'b0;
     layer0_out[7926] <= x[5514];
     layer0_out[7927] <= x[2041];
     layer0_out[7928] <= ~(x[5411] & x[5412]);
     layer0_out[7929] <= ~(x[1544] & x[1545]);
     layer0_out[7930] <= x[7776];
     layer0_out[7931] <= x[5713];
     layer0_out[7932] <= ~(x[1520] | x[1522]);
     layer0_out[7933] <= ~x[5641];
     layer0_out[7934] <= x[1232] & x[1234];
     layer0_out[7935] <= x[1048] ^ x[1049];
     layer0_out[7936] <= x[7957] | x[7958];
     layer0_out[7937] <= ~(x[8016] ^ x[8017]);
     layer0_out[7938] <= x[1136] & x[1137];
     layer0_out[7939] <= x[9068] & x[9069];
     layer0_out[7940] <= x[2735] & ~x[2737];
     layer0_out[7941] <= x[5447] & x[5448];
     layer0_out[7942] <= ~x[2294] | x[2292];
     layer0_out[7943] <= ~x[4859];
     layer0_out[7944] <= x[1947] & x[1948];
     layer0_out[7945] <= ~(x[6069] & x[6070]);
     layer0_out[7946] <= 1'b0;
     layer0_out[7947] <= x[4967] ^ x[4968];
     layer0_out[7948] <= ~x[5704] | x[5705];
     layer0_out[7949] <= x[5938];
     layer0_out[7950] <= x[2865] & x[2866];
     layer0_out[7951] <= x[7256] | x[7257];
     layer0_out[7952] <= x[887] & ~x[889];
     layer0_out[7953] <= x[7497] & x[7498];
     layer0_out[7954] <= x[1255] & x[1257];
     layer0_out[7955] <= ~(x[7721] ^ x[7722]);
     layer0_out[7956] <= ~(x[3711] ^ x[3712]);
     layer0_out[7957] <= x[9033] | x[9034];
     layer0_out[7958] <= ~(x[2756] ^ x[2757]);
     layer0_out[7959] <= ~(x[5152] & x[5153]);
     layer0_out[7960] <= ~x[6402];
     layer0_out[7961] <= x[1021] & x[1023];
     layer0_out[7962] <= x[1366] & x[1367];
     layer0_out[7963] <= ~(x[1321] & x[1323]);
     layer0_out[7964] <= ~(x[7417] | x[7418]);
     layer0_out[7965] <= ~x[518] | x[517];
     layer0_out[7966] <= ~x[411] | x[412];
     layer0_out[7967] <= x[970] | x[972];
     layer0_out[7968] <= x[7639];
     layer0_out[7969] <= x[5558] & x[5559];
     layer0_out[7970] <= x[7772] & x[7773];
     layer0_out[7971] <= ~(x[1823] & x[1824]);
     layer0_out[7972] <= ~x[7388];
     layer0_out[7973] <= ~(x[8580] | x[8581]);
     layer0_out[7974] <= ~(x[6235] | x[6236]);
     layer0_out[7975] <= x[7681] ^ x[7682];
     layer0_out[7976] <= ~x[593] | x[592];
     layer0_out[7977] <= ~x[7326];
     layer0_out[7978] <= ~(x[1513] & x[1514]);
     layer0_out[7979] <= ~(x[700] & x[701]);
     layer0_out[7980] <= ~(x[2169] & x[2171]);
     layer0_out[7981] <= ~(x[866] & x[867]);
     layer0_out[7982] <= x[8226];
     layer0_out[7983] <= x[3017] ^ x[3018];
     layer0_out[7984] <= ~(x[1519] & x[1521]);
     layer0_out[7985] <= x[8982] & x[8983];
     layer0_out[7986] <= x[2574] & x[2575];
     layer0_out[7987] <= x[6286] | x[6287];
     layer0_out[7988] <= ~(x[5921] & x[5922]);
     layer0_out[7989] <= x[1529] & x[1531];
     layer0_out[7990] <= x[689] ^ x[691];
     layer0_out[7991] <= x[8430] & x[8431];
     layer0_out[7992] <= x[5169];
     layer0_out[7993] <= x[8858] & x[8859];
     layer0_out[7994] <= ~(x[9034] | x[9035]);
     layer0_out[7995] <= ~x[8386];
     layer0_out[7996] <= x[5166] & x[5167];
     layer0_out[7997] <= ~(x[4660] | x[4661]);
     layer0_out[7998] <= ~(x[8233] | x[8234]);
     layer0_out[7999] <= ~x[8442];
     layer0_out[8000] <= x[2622] & x[2623];
     layer0_out[8001] <= x[1688] & ~x[1689];
     layer0_out[8002] <= ~x[8787];
     layer0_out[8003] <= x[3710] ^ x[3711];
     layer0_out[8004] <= ~x[483] | x[484];
     layer0_out[8005] <= ~(x[2769] & x[2771]);
     layer0_out[8006] <= 1'b1;
     layer0_out[8007] <= x[2105];
     layer0_out[8008] <= x[4127] ^ x[4128];
     layer0_out[8009] <= ~(x[8936] & x[8937]);
     layer0_out[8010] <= ~x[1612];
     layer0_out[8011] <= x[4292] & x[4293];
     layer0_out[8012] <= x[8246] | x[8247];
     layer0_out[8013] <= x[1762] ^ x[1764];
     layer0_out[8014] <= x[3911] | x[3912];
     layer0_out[8015] <= x[3770] & x[3771];
     layer0_out[8016] <= 1'b1;
     layer0_out[8017] <= x[2175] & x[2176];
     layer0_out[8018] <= ~(x[2741] & x[2742]);
     layer0_out[8019] <= ~x[476] | x[475];
     layer0_out[8020] <= ~(x[6796] | x[6797]);
     layer0_out[8021] <= x[2319] ^ x[2320];
     layer0_out[8022] <= x[1482] & x[1483];
     layer0_out[8023] <= ~(x[6308] & x[6309]);
     layer0_out[8024] <= x[7528] | x[7529];
     layer0_out[8025] <= x[3179] | x[3180];
     layer0_out[8026] <= ~(x[2395] ^ x[2396]);
     layer0_out[8027] <= ~x[349];
     layer0_out[8028] <= x[7569] | x[7570];
     layer0_out[8029] <= ~(x[6844] | x[6845]);
     layer0_out[8030] <= x[6381] | x[6382];
     layer0_out[8031] <= ~(x[1758] | x[1759]);
     layer0_out[8032] <= ~(x[1017] & x[1019]);
     layer0_out[8033] <= ~(x[2534] ^ x[2535]);
     layer0_out[8034] <= ~(x[886] | x[887]);
     layer0_out[8035] <= ~x[1696];
     layer0_out[8036] <= ~(x[5220] & x[5221]);
     layer0_out[8037] <= ~(x[3274] | x[3275]);
     layer0_out[8038] <= ~(x[6078] & x[6079]);
     layer0_out[8039] <= x[8182];
     layer0_out[8040] <= x[3299] | x[3300];
     layer0_out[8041] <= ~(x[2056] & x[2057]);
     layer0_out[8042] <= x[4224];
     layer0_out[8043] <= ~x[7572];
     layer0_out[8044] <= x[7540];
     layer0_out[8045] <= ~(x[2236] & x[2238]);
     layer0_out[8046] <= 1'b0;
     layer0_out[8047] <= ~(x[140] ^ x[142]);
     layer0_out[8048] <= 1'b1;
     layer0_out[8049] <= ~x[734] | x[732];
     layer0_out[8050] <= ~(x[501] ^ x[503]);
     layer0_out[8051] <= x[1304] & x[1306];
     layer0_out[8052] <= x[6497];
     layer0_out[8053] <= x[5588];
     layer0_out[8054] <= x[2842] ^ x[2843];
     layer0_out[8055] <= 1'b0;
     layer0_out[8056] <= ~x[1580];
     layer0_out[8057] <= x[8856] ^ x[8857];
     layer0_out[8058] <= x[6323] | x[6324];
     layer0_out[8059] <= ~x[5385];
     layer0_out[8060] <= x[1644] & x[1646];
     layer0_out[8061] <= x[2722];
     layer0_out[8062] <= x[9030];
     layer0_out[8063] <= 1'b0;
     layer0_out[8064] <= ~x[8063];
     layer0_out[8065] <= ~x[6010] | x[6009];
     layer0_out[8066] <= ~(x[2442] & x[2444]);
     layer0_out[8067] <= ~x[1513] | x[1512];
     layer0_out[8068] <= x[5197] & x[5198];
     layer0_out[8069] <= ~x[1529] | x[1527];
     layer0_out[8070] <= ~(x[7198] | x[7199]);
     layer0_out[8071] <= x[6257] ^ x[6258];
     layer0_out[8072] <= x[1222] & x[1224];
     layer0_out[8073] <= x[5837] & x[5838];
     layer0_out[8074] <= x[4098];
     layer0_out[8075] <= x[7788] & ~x[7789];
     layer0_out[8076] <= x[758] & x[760];
     layer0_out[8077] <= 1'b1;
     layer0_out[8078] <= x[2828] & x[2829];
     layer0_out[8079] <= x[1136] & x[1138];
     layer0_out[8080] <= x[977] | x[978];
     layer0_out[8081] <= ~(x[4231] & x[4232]);
     layer0_out[8082] <= x[2784] ^ x[2785];
     layer0_out[8083] <= ~(x[6543] | x[6544]);
     layer0_out[8084] <= ~(x[8744] | x[8745]);
     layer0_out[8085] <= ~(x[120] & x[121]);
     layer0_out[8086] <= x[5312] ^ x[5313];
     layer0_out[8087] <= x[3442] & ~x[3443];
     layer0_out[8088] <= x[2648] & x[2649];
     layer0_out[8089] <= ~(x[5727] ^ x[5728]);
     layer0_out[8090] <= x[1203] & x[1205];
     layer0_out[8091] <= x[6314] | x[6315];
     layer0_out[8092] <= x[5568] ^ x[5569];
     layer0_out[8093] <= ~(x[1012] | x[1014]);
     layer0_out[8094] <= ~(x[7729] ^ x[7730]);
     layer0_out[8095] <= 1'b1;
     layer0_out[8096] <= x[2055] & x[2057];
     layer0_out[8097] <= x[851] & x[852];
     layer0_out[8098] <= x[4919] | x[4920];
     layer0_out[8099] <= x[5593] ^ x[5594];
     layer0_out[8100] <= ~(x[1478] | x[1479]);
     layer0_out[8101] <= x[3776] & x[3777];
     layer0_out[8102] <= ~x[595];
     layer0_out[8103] <= x[1421];
     layer0_out[8104] <= x[805];
     layer0_out[8105] <= x[1689] | x[1690];
     layer0_out[8106] <= ~x[7314];
     layer0_out[8107] <= x[2525] | x[2526];
     layer0_out[8108] <= x[7780];
     layer0_out[8109] <= x[514] & ~x[516];
     layer0_out[8110] <= x[4589] & ~x[4588];
     layer0_out[8111] <= x[2533] ^ x[2535];
     layer0_out[8112] <= ~x[2502] | x[2501];
     layer0_out[8113] <= x[2104] | x[2106];
     layer0_out[8114] <= x[1369] & x[1371];
     layer0_out[8115] <= x[7667];
     layer0_out[8116] <= x[2869] ^ x[2870];
     layer0_out[8117] <= 1'b0;
     layer0_out[8118] <= ~x[6687];
     layer0_out[8119] <= ~x[4188];
     layer0_out[8120] <= ~(x[5069] | x[5070]);
     layer0_out[8121] <= ~(x[8626] | x[8627]);
     layer0_out[8122] <= ~(x[7550] | x[7551]);
     layer0_out[8123] <= ~(x[6875] & x[6876]);
     layer0_out[8124] <= ~(x[6023] ^ x[6024]);
     layer0_out[8125] <= ~(x[2619] & x[2621]);
     layer0_out[8126] <= ~(x[7521] | x[7522]);
     layer0_out[8127] <= 1'b1;
     layer0_out[8128] <= ~(x[149] & x[151]);
     layer0_out[8129] <= ~(x[7786] & x[7787]);
     layer0_out[8130] <= x[8616];
     layer0_out[8131] <= ~(x[4450] & x[4451]);
     layer0_out[8132] <= x[6117] & x[6118];
     layer0_out[8133] <= ~x[4220];
     layer0_out[8134] <= x[8449];
     layer0_out[8135] <= ~x[5952];
     layer0_out[8136] <= ~(x[5201] & x[5202]);
     layer0_out[8137] <= x[8074] ^ x[8075];
     layer0_out[8138] <= x[1512] & x[1514];
     layer0_out[8139] <= ~x[1150];
     layer0_out[8140] <= x[40] ^ x[41];
     layer0_out[8141] <= ~(x[6270] | x[6271]);
     layer0_out[8142] <= x[1398];
     layer0_out[8143] <= x[3057] | x[3058];
     layer0_out[8144] <= ~(x[5928] & x[5929]);
     layer0_out[8145] <= x[8748] | x[8749];
     layer0_out[8146] <= ~x[4475] | x[4476];
     layer0_out[8147] <= ~(x[5702] & x[5703]);
     layer0_out[8148] <= x[8629] | x[8630];
     layer0_out[8149] <= x[2015] & x[2016];
     layer0_out[8150] <= x[3157] | x[3158];
     layer0_out[8151] <= x[637] ^ x[639];
     layer0_out[8152] <= ~x[199] | x[198];
     layer0_out[8153] <= ~(x[3] & x[4]);
     layer0_out[8154] <= ~(x[92] & x[93]);
     layer0_out[8155] <= ~(x[908] | x[909]);
     layer0_out[8156] <= x[3925] | x[3926];
     layer0_out[8157] <= x[8967] & x[8968];
     layer0_out[8158] <= x[7340];
     layer0_out[8159] <= ~x[2529];
     layer0_out[8160] <= 1'b0;
     layer0_out[8161] <= ~(x[8770] ^ x[8771]);
     layer0_out[8162] <= x[1725] & x[1727];
     layer0_out[8163] <= 1'b1;
     layer0_out[8164] <= x[709] & x[710];
     layer0_out[8165] <= ~(x[1253] & x[1254]);
     layer0_out[8166] <= x[4212];
     layer0_out[8167] <= ~x[2466] | x[2467];
     layer0_out[8168] <= x[7723] | x[7724];
     layer0_out[8169] <= 1'b1;
     layer0_out[8170] <= ~x[428] | x[427];
     layer0_out[8171] <= x[9157] | x[9158];
     layer0_out[8172] <= ~x[1641] | x[1643];
     layer0_out[8173] <= x[7271] | x[7272];
     layer0_out[8174] <= x[9211];
     layer0_out[8175] <= 1'b1;
     layer0_out[8176] <= x[2561] | x[2562];
     layer0_out[8177] <= x[431] & ~x[433];
     layer0_out[8178] <= ~(x[969] ^ x[970]);
     layer0_out[8179] <= ~(x[5359] & x[5360]);
     layer0_out[8180] <= x[938] | x[939];
     layer0_out[8181] <= x[8610] ^ x[8611];
     layer0_out[8182] <= x[2547] & x[2549];
     layer0_out[8183] <= x[4394];
     layer0_out[8184] <= ~(x[7614] & x[7615]);
     layer0_out[8185] <= x[4651];
     layer0_out[8186] <= ~(x[1802] & x[1804]);
     layer0_out[8187] <= 1'b0;
     layer0_out[8188] <= x[676] ^ x[678];
     layer0_out[8189] <= x[727] ^ x[729];
     layer0_out[8190] <= x[2215] & ~x[2217];
     layer0_out[8191] <= x[2200] ^ x[2201];
     layer0_out[8192] <= ~x[1975];
     layer0_out[8193] <= ~(x[4023] | x[4024]);
     layer0_out[8194] <= x[2604] & x[2605];
     layer0_out[8195] <= ~(x[6029] & x[6030]);
     layer0_out[8196] <= x[8183] | x[8184];
     layer0_out[8197] <= x[1129] & x[1131];
     layer0_out[8198] <= ~x[484] | x[482];
     layer0_out[8199] <= ~(x[3563] | x[3564]);
     layer0_out[8200] <= ~(x[6420] | x[6421]);
     layer0_out[8201] <= x[2906] | x[2907];
     layer0_out[8202] <= ~(x[5894] ^ x[5895]);
     layer0_out[8203] <= x[103] & x[105];
     layer0_out[8204] <= ~(x[2346] ^ x[2347]);
     layer0_out[8205] <= ~(x[1165] ^ x[1167]);
     layer0_out[8206] <= ~(x[319] ^ x[320]);
     layer0_out[8207] <= x[6013] | x[6014];
     layer0_out[8208] <= x[7406] | x[7407];
     layer0_out[8209] <= 1'b1;
     layer0_out[8210] <= 1'b0;
     layer0_out[8211] <= 1'b1;
     layer0_out[8212] <= x[408];
     layer0_out[8213] <= ~(x[83] & x[84]);
     layer0_out[8214] <= ~x[7467];
     layer0_out[8215] <= x[1999];
     layer0_out[8216] <= ~(x[1312] & x[1314]);
     layer0_out[8217] <= ~x[1952] | x[1951];
     layer0_out[8218] <= x[3857] & x[3858];
     layer0_out[8219] <= 1'b1;
     layer0_out[8220] <= ~x[6263];
     layer0_out[8221] <= x[2347] & x[2348];
     layer0_out[8222] <= 1'b1;
     layer0_out[8223] <= x[2240] & x[2242];
     layer0_out[8224] <= x[671] & x[673];
     layer0_out[8225] <= x[1503];
     layer0_out[8226] <= ~(x[5215] | x[5216]);
     layer0_out[8227] <= ~x[4254] | x[4253];
     layer0_out[8228] <= ~(x[3740] ^ x[3741]);
     layer0_out[8229] <= ~x[2078];
     layer0_out[8230] <= ~(x[6170] ^ x[6171]);
     layer0_out[8231] <= x[3989] ^ x[3990];
     layer0_out[8232] <= ~(x[4451] & x[4452]);
     layer0_out[8233] <= x[3242] | x[3243];
     layer0_out[8234] <= x[627] | x[628];
     layer0_out[8235] <= ~x[6646];
     layer0_out[8236] <= ~(x[2545] & x[2546]);
     layer0_out[8237] <= 1'b1;
     layer0_out[8238] <= ~(x[2286] & x[2287]);
     layer0_out[8239] <= ~x[107];
     layer0_out[8240] <= ~(x[5324] & x[5325]);
     layer0_out[8241] <= x[8607] ^ x[8608];
     layer0_out[8242] <= ~x[2745];
     layer0_out[8243] <= x[741];
     layer0_out[8244] <= ~(x[4493] | x[4494]);
     layer0_out[8245] <= x[6193] & x[6194];
     layer0_out[8246] <= x[8737] & ~x[8738];
     layer0_out[8247] <= x[4369];
     layer0_out[8248] <= ~x[335];
     layer0_out[8249] <= ~(x[199] & x[201]);
     layer0_out[8250] <= ~x[7486];
     layer0_out[8251] <= ~x[2038];
     layer0_out[8252] <= 1'b1;
     layer0_out[8253] <= x[6631];
     layer0_out[8254] <= 1'b1;
     layer0_out[8255] <= x[1791] ^ x[1792];
     layer0_out[8256] <= x[7062] | x[7063];
     layer0_out[8257] <= x[8505];
     layer0_out[8258] <= ~x[8351];
     layer0_out[8259] <= ~x[2472];
     layer0_out[8260] <= ~(x[1628] & x[1629]);
     layer0_out[8261] <= x[2084] & x[2086];
     layer0_out[8262] <= x[6532] & ~x[6531];
     layer0_out[8263] <= 1'b0;
     layer0_out[8264] <= x[233] ^ x[234];
     layer0_out[8265] <= ~x[5309];
     layer0_out[8266] <= ~x[4730];
     layer0_out[8267] <= x[7492] | x[7493];
     layer0_out[8268] <= ~(x[890] | x[892]);
     layer0_out[8269] <= x[2750] & ~x[2749];
     layer0_out[8270] <= x[6897] | x[6898];
     layer0_out[8271] <= x[8194];
     layer0_out[8272] <= ~x[8578];
     layer0_out[8273] <= x[2297] & x[2299];
     layer0_out[8274] <= ~(x[5965] & x[5966]);
     layer0_out[8275] <= x[3071];
     layer0_out[8276] <= x[456] ^ x[458];
     layer0_out[8277] <= ~(x[7624] ^ x[7625]);
     layer0_out[8278] <= x[4776] ^ x[4777];
     layer0_out[8279] <= x[1106] & ~x[1105];
     layer0_out[8280] <= x[6560];
     layer0_out[8281] <= x[1135] & ~x[1133];
     layer0_out[8282] <= 1'b0;
     layer0_out[8283] <= 1'b1;
     layer0_out[8284] <= x[7456] | x[7457];
     layer0_out[8285] <= ~(x[6217] | x[6218]);
     layer0_out[8286] <= 1'b1;
     layer0_out[8287] <= ~(x[5345] | x[5346]);
     layer0_out[8288] <= x[3240] ^ x[3241];
     layer0_out[8289] <= ~(x[3055] & x[3056]);
     layer0_out[8290] <= x[6833] | x[6834];
     layer0_out[8291] <= x[1620] | x[1621];
     layer0_out[8292] <= ~(x[1747] & x[1748]);
     layer0_out[8293] <= x[344] & ~x[343];
     layer0_out[8294] <= ~(x[5200] | x[5201]);
     layer0_out[8295] <= x[1339] | x[1340];
     layer0_out[8296] <= ~x[4486];
     layer0_out[8297] <= x[400] ^ x[401];
     layer0_out[8298] <= x[4583] & x[4584];
     layer0_out[8299] <= x[7190] & x[7191];
     layer0_out[8300] <= x[3460] ^ x[3461];
     layer0_out[8301] <= x[5115] & ~x[5114];
     layer0_out[8302] <= ~(x[690] & x[691]);
     layer0_out[8303] <= ~(x[9112] | x[9113]);
     layer0_out[8304] <= ~(x[1966] ^ x[1967]);
     layer0_out[8305] <= ~(x[6478] | x[6479]);
     layer0_out[8306] <= ~(x[5335] & x[5336]);
     layer0_out[8307] <= ~x[4719] | x[4718];
     layer0_out[8308] <= ~(x[5792] & x[5793]);
     layer0_out[8309] <= x[7534] & ~x[7535];
     layer0_out[8310] <= ~(x[8294] & x[8295]);
     layer0_out[8311] <= x[3610] | x[3611];
     layer0_out[8312] <= x[1879] & x[1880];
     layer0_out[8313] <= ~x[253];
     layer0_out[8314] <= ~(x[7400] | x[7401]);
     layer0_out[8315] <= ~(x[7577] | x[7578]);
     layer0_out[8316] <= x[677] ^ x[679];
     layer0_out[8317] <= x[2080] & x[2082];
     layer0_out[8318] <= x[8088] ^ x[8089];
     layer0_out[8319] <= x[2596] | x[2598];
     layer0_out[8320] <= ~(x[6063] & x[6064]);
     layer0_out[8321] <= x[4305];
     layer0_out[8322] <= x[6393] & x[6394];
     layer0_out[8323] <= x[2320] | x[2321];
     layer0_out[8324] <= ~(x[2534] & x[2536]);
     layer0_out[8325] <= ~(x[5475] & x[5476]);
     layer0_out[8326] <= x[2450] & x[2452];
     layer0_out[8327] <= x[239] & x[240];
     layer0_out[8328] <= ~(x[8553] & x[8554]);
     layer0_out[8329] <= x[2349] | x[2350];
     layer0_out[8330] <= x[1506] ^ x[1507];
     layer0_out[8331] <= x[1954];
     layer0_out[8332] <= ~(x[254] & x[256]);
     layer0_out[8333] <= ~(x[1819] & x[1821]);
     layer0_out[8334] <= x[7412] ^ x[7413];
     layer0_out[8335] <= 1'b1;
     layer0_out[8336] <= x[8716] | x[8717];
     layer0_out[8337] <= x[7306] & x[7307];
     layer0_out[8338] <= x[502] | x[503];
     layer0_out[8339] <= 1'b1;
     layer0_out[8340] <= ~(x[3484] ^ x[3485]);
     layer0_out[8341] <= ~(x[2491] & x[2492]);
     layer0_out[8342] <= ~(x[2306] & x[2307]);
     layer0_out[8343] <= ~(x[8866] & x[8867]);
     layer0_out[8344] <= 1'b1;
     layer0_out[8345] <= x[5252] & x[5253];
     layer0_out[8346] <= ~x[102];
     layer0_out[8347] <= ~(x[1715] & x[1717]);
     layer0_out[8348] <= x[9160] & x[9161];
     layer0_out[8349] <= x[7333] | x[7334];
     layer0_out[8350] <= 1'b0;
     layer0_out[8351] <= ~(x[8557] | x[8558]);
     layer0_out[8352] <= ~(x[1329] ^ x[1331]);
     layer0_out[8353] <= ~x[793];
     layer0_out[8354] <= x[8932] ^ x[8933];
     layer0_out[8355] <= ~x[288] | x[290];
     layer0_out[8356] <= x[4750] & x[4751];
     layer0_out[8357] <= ~(x[9073] & x[9074]);
     layer0_out[8358] <= x[2434] & x[2435];
     layer0_out[8359] <= ~(x[1318] & x[1320]);
     layer0_out[8360] <= x[1800];
     layer0_out[8361] <= ~(x[1386] | x[1388]);
     layer0_out[8362] <= x[5643] & x[5644];
     layer0_out[8363] <= 1'b1;
     layer0_out[8364] <= ~(x[2572] & x[2573]);
     layer0_out[8365] <= x[7138] & x[7139];
     layer0_out[8366] <= ~(x[8221] | x[8222]);
     layer0_out[8367] <= ~(x[7920] & x[7921]);
     layer0_out[8368] <= ~(x[6248] | x[6249]);
     layer0_out[8369] <= 1'b0;
     layer0_out[8370] <= x[1593] | x[1595];
     layer0_out[8371] <= ~(x[8057] ^ x[8058]);
     layer0_out[8372] <= x[5333] & x[5334];
     layer0_out[8373] <= x[150] & x[151];
     layer0_out[8374] <= x[2151] & x[2152];
     layer0_out[8375] <= ~(x[219] ^ x[221]);
     layer0_out[8376] <= ~(x[6372] ^ x[6373]);
     layer0_out[8377] <= ~(x[5614] & x[5615]);
     layer0_out[8378] <= x[6503];
     layer0_out[8379] <= ~(x[7597] | x[7598]);
     layer0_out[8380] <= ~(x[1978] & x[1980]);
     layer0_out[8381] <= x[3763] & ~x[3764];
     layer0_out[8382] <= ~(x[6360] | x[6361]);
     layer0_out[8383] <= 1'b0;
     layer0_out[8384] <= 1'b1;
     layer0_out[8385] <= x[5298] & x[5299];
     layer0_out[8386] <= x[1733] & x[1734];
     layer0_out[8387] <= ~(x[906] & x[908]);
     layer0_out[8388] <= x[7727];
     layer0_out[8389] <= x[8814] | x[8815];
     layer0_out[8390] <= x[1448] & x[1450];
     layer0_out[8391] <= x[7312] | x[7313];
     layer0_out[8392] <= x[5738];
     layer0_out[8393] <= ~(x[8452] ^ x[8453]);
     layer0_out[8394] <= 1'b1;
     layer0_out[8395] <= x[1987];
     layer0_out[8396] <= x[4308] & x[4309];
     layer0_out[8397] <= x[2162] & x[2164];
     layer0_out[8398] <= x[2187] ^ x[2189];
     layer0_out[8399] <= x[2603] ^ x[2605];
     layer0_out[8400] <= ~(x[1285] ^ x[1286]);
     layer0_out[8401] <= x[7161] & ~x[7162];
     layer0_out[8402] <= x[1064] & ~x[1063];
     layer0_out[8403] <= x[7898] & ~x[7899];
     layer0_out[8404] <= ~(x[8750] | x[8751]);
     layer0_out[8405] <= ~(x[1886] & x[1888]);
     layer0_out[8406] <= ~x[2226] | x[2227];
     layer0_out[8407] <= ~x[7346];
     layer0_out[8408] <= ~(x[4367] | x[4368]);
     layer0_out[8409] <= 1'b1;
     layer0_out[8410] <= x[3968];
     layer0_out[8411] <= 1'b0;
     layer0_out[8412] <= 1'b1;
     layer0_out[8413] <= 1'b0;
     layer0_out[8414] <= ~(x[9108] ^ x[9109]);
     layer0_out[8415] <= x[572] & ~x[574];
     layer0_out[8416] <= x[18] ^ x[19];
     layer0_out[8417] <= x[1833];
     layer0_out[8418] <= ~(x[2899] & x[2900]);
     layer0_out[8419] <= x[5688] & ~x[5689];
     layer0_out[8420] <= ~(x[3538] | x[3539]);
     layer0_out[8421] <= x[472] | x[473];
     layer0_out[8422] <= x[8940] | x[8941];
     layer0_out[8423] <= x[680] | x[681];
     layer0_out[8424] <= ~x[4987] | x[4988];
     layer0_out[8425] <= x[2801] ^ x[2802];
     layer0_out[8426] <= x[3886] ^ x[3887];
     layer0_out[8427] <= x[2551] & x[2553];
     layer0_out[8428] <= x[1004] ^ x[1006];
     layer0_out[8429] <= x[8009] & ~x[8010];
     layer0_out[8430] <= ~x[4328];
     layer0_out[8431] <= ~x[6696] | x[6695];
     layer0_out[8432] <= x[7512] & ~x[7513];
     layer0_out[8433] <= x[4641] & x[4642];
     layer0_out[8434] <= x[1186];
     layer0_out[8435] <= x[1176];
     layer0_out[8436] <= x[1795];
     layer0_out[8437] <= x[3196] & x[3197];
     layer0_out[8438] <= x[6155] | x[6156];
     layer0_out[8439] <= ~x[8754];
     layer0_out[8440] <= x[6484] ^ x[6485];
     layer0_out[8441] <= x[121];
     layer0_out[8442] <= x[3655] | x[3656];
     layer0_out[8443] <= ~(x[676] & x[677]);
     layer0_out[8444] <= ~x[645] | x[644];
     layer0_out[8445] <= x[4637] & x[4638];
     layer0_out[8446] <= ~x[8249];
     layer0_out[8447] <= x[1899];
     layer0_out[8448] <= ~x[2026];
     layer0_out[8449] <= ~(x[790] & x[792]);
     layer0_out[8450] <= x[2747] ^ x[2749];
     layer0_out[8451] <= ~(x[4544] & x[4545]);
     layer0_out[8452] <= x[958];
     layer0_out[8453] <= ~(x[4117] | x[4118]);
     layer0_out[8454] <= 1'b1;
     layer0_out[8455] <= ~(x[5268] & x[5269]);
     layer0_out[8456] <= ~(x[2895] & x[2896]);
     layer0_out[8457] <= x[7657] & ~x[7658];
     layer0_out[8458] <= ~(x[4130] & x[4131]);
     layer0_out[8459] <= ~(x[15] | x[17]);
     layer0_out[8460] <= ~(x[263] ^ x[264]);
     layer0_out[8461] <= ~(x[6974] | x[6975]);
     layer0_out[8462] <= ~x[1270] | x[1268];
     layer0_out[8463] <= x[8224] | x[8225];
     layer0_out[8464] <= ~x[4648] | x[4649];
     layer0_out[8465] <= x[2787] & ~x[2788];
     layer0_out[8466] <= ~(x[225] | x[227]);
     layer0_out[8467] <= 1'b1;
     layer0_out[8468] <= ~(x[4840] ^ x[4841]);
     layer0_out[8469] <= x[3991] | x[3992];
     layer0_out[8470] <= ~(x[52] & x[53]);
     layer0_out[8471] <= x[7183] ^ x[7184];
     layer0_out[8472] <= x[1379] & ~x[1381];
     layer0_out[8473] <= x[8164] | x[8165];
     layer0_out[8474] <= ~x[9188];
     layer0_out[8475] <= ~(x[3986] | x[3987]);
     layer0_out[8476] <= ~x[8927];
     layer0_out[8477] <= ~(x[8354] | x[8355]);
     layer0_out[8478] <= ~(x[8784] | x[8785]);
     layer0_out[8479] <= x[4818] | x[4819];
     layer0_out[8480] <= ~(x[3921] | x[3922]);
     layer0_out[8481] <= x[7117];
     layer0_out[8482] <= ~(x[996] ^ x[997]);
     layer0_out[8483] <= ~(x[8943] & x[8944]);
     layer0_out[8484] <= x[9129] | x[9130];
     layer0_out[8485] <= ~(x[8906] | x[8907]);
     layer0_out[8486] <= 1'b1;
     layer0_out[8487] <= x[7916] | x[7917];
     layer0_out[8488] <= x[7320];
     layer0_out[8489] <= x[7871] & ~x[7872];
     layer0_out[8490] <= x[667] | x[669];
     layer0_out[8491] <= x[357];
     layer0_out[8492] <= x[2963] & ~x[2964];
     layer0_out[8493] <= 1'b0;
     layer0_out[8494] <= ~(x[8240] | x[8241]);
     layer0_out[8495] <= ~(x[7514] & x[7515]);
     layer0_out[8496] <= ~(x[7354] | x[7355]);
     layer0_out[8497] <= ~x[1389];
     layer0_out[8498] <= x[3586] | x[3587];
     layer0_out[8499] <= x[3622] | x[3623];
     layer0_out[8500] <= x[7672] & ~x[7671];
     layer0_out[8501] <= ~x[757];
     layer0_out[8502] <= x[2486] & x[2488];
     layer0_out[8503] <= x[2544] & x[2545];
     layer0_out[8504] <= ~x[7557] | x[7558];
     layer0_out[8505] <= ~x[5129];
     layer0_out[8506] <= ~(x[5759] | x[5760]);
     layer0_out[8507] <= ~(x[1085] ^ x[1087]);
     layer0_out[8508] <= ~(x[5722] & x[5723]);
     layer0_out[8509] <= 1'b1;
     layer0_out[8510] <= x[4352] | x[4353];
     layer0_out[8511] <= ~(x[1944] | x[1945]);
     layer0_out[8512] <= x[432] & x[433];
     layer0_out[8513] <= x[1050] ^ x[1052];
     layer0_out[8514] <= ~(x[7519] ^ x[7520]);
     layer0_out[8515] <= x[5838] & x[5839];
     layer0_out[8516] <= ~x[7029] | x[7030];
     layer0_out[8517] <= ~(x[1195] & x[1196]);
     layer0_out[8518] <= ~x[3393];
     layer0_out[8519] <= ~(x[515] | x[517]);
     layer0_out[8520] <= x[7270];
     layer0_out[8521] <= x[1548];
     layer0_out[8522] <= ~(x[1673] & x[1675]);
     layer0_out[8523] <= ~(x[351] | x[353]);
     layer0_out[8524] <= ~(x[9189] | x[9190]);
     layer0_out[8525] <= x[4459] & x[4460];
     layer0_out[8526] <= ~(x[474] & x[475]);
     layer0_out[8527] <= ~(x[118] & x[120]);
     layer0_out[8528] <= x[855] | x[856];
     layer0_out[8529] <= x[6199];
     layer0_out[8530] <= ~(x[9172] & x[9173]);
     layer0_out[8531] <= ~x[5739];
     layer0_out[8532] <= ~(x[60] ^ x[61]);
     layer0_out[8533] <= ~x[3291];
     layer0_out[8534] <= ~(x[1902] & x[1903]);
     layer0_out[8535] <= ~(x[2180] ^ x[2182]);
     layer0_out[8536] <= x[4143] | x[4144];
     layer0_out[8537] <= x[2624] ^ x[2625];
     layer0_out[8538] <= x[966];
     layer0_out[8539] <= ~(x[4762] & x[4763]);
     layer0_out[8540] <= x[7068];
     layer0_out[8541] <= ~(x[5649] | x[5650]);
     layer0_out[8542] <= x[6761] ^ x[6762];
     layer0_out[8543] <= ~(x[897] & x[899]);
     layer0_out[8544] <= ~(x[2636] & x[2638]);
     layer0_out[8545] <= x[7179];
     layer0_out[8546] <= x[5573];
     layer0_out[8547] <= x[85] ^ x[87];
     layer0_out[8548] <= x[4523] & x[4524];
     layer0_out[8549] <= x[2707] ^ x[2709];
     layer0_out[8550] <= ~x[7652];
     layer0_out[8551] <= x[7476] | x[7477];
     layer0_out[8552] <= ~(x[1446] ^ x[1448]);
     layer0_out[8553] <= ~(x[3838] | x[3839]);
     layer0_out[8554] <= ~x[2939] | x[2938];
     layer0_out[8555] <= x[6469] | x[6470];
     layer0_out[8556] <= ~(x[1481] ^ x[1483]);
     layer0_out[8557] <= ~x[2385];
     layer0_out[8558] <= x[8282] ^ x[8283];
     layer0_out[8559] <= x[1951];
     layer0_out[8560] <= x[1881] & x[1883];
     layer0_out[8561] <= 1'b0;
     layer0_out[8562] <= ~x[8439];
     layer0_out[8563] <= 1'b1;
     layer0_out[8564] <= x[9154] & x[9155];
     layer0_out[8565] <= x[7791] | x[7792];
     layer0_out[8566] <= ~(x[7865] ^ x[7866]);
     layer0_out[8567] <= 1'b0;
     layer0_out[8568] <= ~x[9174];
     layer0_out[8569] <= x[516] | x[518];
     layer0_out[8570] <= 1'b0;
     layer0_out[8571] <= x[4825] & x[4826];
     layer0_out[8572] <= ~(x[3229] | x[3230]);
     layer0_out[8573] <= ~(x[9040] | x[9041]);
     layer0_out[8574] <= x[1038] & x[1039];
     layer0_out[8575] <= ~x[395];
     layer0_out[8576] <= ~x[166] | x[168];
     layer0_out[8577] <= 1'b0;
     layer0_out[8578] <= ~(x[2233] & x[2234]);
     layer0_out[8579] <= ~x[1612] | x[1614];
     layer0_out[8580] <= x[3259] | x[3260];
     layer0_out[8581] <= x[7807];
     layer0_out[8582] <= ~(x[2112] & x[2113]);
     layer0_out[8583] <= ~(x[2123] & x[2124]);
     layer0_out[8584] <= ~(x[8191] ^ x[8192]);
     layer0_out[8585] <= x[6772];
     layer0_out[8586] <= ~(x[1601] & x[1603]);
     layer0_out[8587] <= x[6784] | x[6785];
     layer0_out[8588] <= ~x[8378];
     layer0_out[8589] <= ~x[7683];
     layer0_out[8590] <= ~(x[2482] & x[2484]);
     layer0_out[8591] <= ~x[7685] | x[7684];
     layer0_out[8592] <= ~(x[1261] & x[1263]);
     layer0_out[8593] <= ~(x[2243] & x[2245]);
     layer0_out[8594] <= x[6404] ^ x[6405];
     layer0_out[8595] <= x[2717] | x[2719];
     layer0_out[8596] <= ~x[3553] | x[3552];
     layer0_out[8597] <= ~(x[5861] & x[5862]);
     layer0_out[8598] <= ~(x[183] ^ x[184]);
     layer0_out[8599] <= ~x[4502];
     layer0_out[8600] <= ~(x[1958] & x[1960]);
     layer0_out[8601] <= x[67] & x[69];
     layer0_out[8602] <= x[4278] & x[4279];
     layer0_out[8603] <= ~x[4761];
     layer0_out[8604] <= ~x[4815];
     layer0_out[8605] <= ~(x[2464] & x[2465]);
     layer0_out[8606] <= ~(x[5913] | x[5914]);
     layer0_out[8607] <= x[1660] | x[1662];
     layer0_out[8608] <= ~(x[1890] & x[1892]);
     layer0_out[8609] <= x[1769];
     layer0_out[8610] <= x[2508];
     layer0_out[8611] <= ~x[79] | x[81];
     layer0_out[8612] <= 1'b0;
     layer0_out[8613] <= ~(x[4854] | x[4855]);
     layer0_out[8614] <= x[5174];
     layer0_out[8615] <= ~x[4242];
     layer0_out[8616] <= x[979];
     layer0_out[8617] <= x[2591] & x[2592];
     layer0_out[8618] <= x[8780] | x[8781];
     layer0_out[8619] <= x[9113] | x[9114];
     layer0_out[8620] <= ~(x[6307] | x[6308]);
     layer0_out[8621] <= ~(x[837] & x[839]);
     layer0_out[8622] <= x[1138] & x[1139];
     layer0_out[8623] <= x[3350] & ~x[3349];
     layer0_out[8624] <= ~x[8942] | x[8943];
     layer0_out[8625] <= ~(x[9008] | x[9009]);
     layer0_out[8626] <= ~(x[2843] & x[2844]);
     layer0_out[8627] <= x[806] & x[807];
     layer0_out[8628] <= ~(x[1451] & x[1452]);
     layer0_out[8629] <= ~(x[2726] & x[2727]);
     layer0_out[8630] <= x[495];
     layer0_out[8631] <= x[4850] & x[4851];
     layer0_out[8632] <= ~x[2201] | x[2199];
     layer0_out[8633] <= ~(x[1587] & x[1589]);
     layer0_out[8634] <= x[8205] | x[8206];
     layer0_out[8635] <= x[3249] ^ x[3250];
     layer0_out[8636] <= ~x[8115] | x[8114];
     layer0_out[8637] <= ~(x[3479] | x[3480]);
     layer0_out[8638] <= ~x[1211] | x[1210];
     layer0_out[8639] <= ~(x[2178] & x[2179]);
     layer0_out[8640] <= x[1516] & ~x[1515];
     layer0_out[8641] <= x[5966] | x[5967];
     layer0_out[8642] <= ~x[8070];
     layer0_out[8643] <= ~x[6707] | x[6706];
     layer0_out[8644] <= ~x[1065] | x[1066];
     layer0_out[8645] <= x[1353] & x[1354];
     layer0_out[8646] <= x[5547] & x[5548];
     layer0_out[8647] <= ~(x[1271] | x[1273]);
     layer0_out[8648] <= ~(x[5170] | x[5171]);
     layer0_out[8649] <= x[1900] & x[1901];
     layer0_out[8650] <= ~x[1010];
     layer0_out[8651] <= ~(x[2664] ^ x[2666]);
     layer0_out[8652] <= x[1345] ^ x[1346];
     layer0_out[8653] <= ~(x[4821] & x[4822]);
     layer0_out[8654] <= ~(x[6452] | x[6453]);
     layer0_out[8655] <= x[686] & x[688];
     layer0_out[8656] <= ~(x[4321] & x[4322]);
     layer0_out[8657] <= ~x[189];
     layer0_out[8658] <= x[8115] | x[8116];
     layer0_out[8659] <= ~x[8128];
     layer0_out[8660] <= ~(x[8889] & x[8890]);
     layer0_out[8661] <= x[1564] & x[1566];
     layer0_out[8662] <= ~(x[2322] ^ x[2324]);
     layer0_out[8663] <= x[4519] & x[4520];
     layer0_out[8664] <= ~x[6857];
     layer0_out[8665] <= ~x[1204] | x[1206];
     layer0_out[8666] <= x[750] & x[751];
     layer0_out[8667] <= ~x[1488];
     layer0_out[8668] <= x[9095];
     layer0_out[8669] <= ~(x[3798] | x[3799]);
     layer0_out[8670] <= ~x[2445] | x[2443];
     layer0_out[8671] <= ~(x[2678] & x[2680]);
     layer0_out[8672] <= x[398] & x[399];
     layer0_out[8673] <= x[2423] ^ x[2424];
     layer0_out[8674] <= x[2690] ^ x[2692];
     layer0_out[8675] <= 1'b0;
     layer0_out[8676] <= x[8277] | x[8278];
     layer0_out[8677] <= 1'b1;
     layer0_out[8678] <= x[877] | x[879];
     layer0_out[8679] <= x[771] ^ x[773];
     layer0_out[8680] <= ~x[398];
     layer0_out[8681] <= ~(x[3458] ^ x[3459]);
     layer0_out[8682] <= ~(x[8139] | x[8140]);
     layer0_out[8683] <= ~(x[2691] & x[2692]);
     layer0_out[8684] <= x[7866] & ~x[7867];
     layer0_out[8685] <= ~(x[5095] | x[5096]);
     layer0_out[8686] <= x[50] ^ x[52];
     layer0_out[8687] <= ~(x[4884] | x[4885]);
     layer0_out[8688] <= ~(x[1511] ^ x[1513]);
     layer0_out[8689] <= x[8369] & x[8370];
     layer0_out[8690] <= x[8493] ^ x[8494];
     layer0_out[8691] <= x[4736] ^ x[4737];
     layer0_out[8692] <= ~x[7046];
     layer0_out[8693] <= x[2046] | x[2047];
     layer0_out[8694] <= x[7343] & x[7344];
     layer0_out[8695] <= ~(x[2595] & x[2596]);
     layer0_out[8696] <= x[4056] & x[4057];
     layer0_out[8697] <= ~(x[2444] & x[2446]);
     layer0_out[8698] <= ~(x[6049] & x[6050]);
     layer0_out[8699] <= ~x[7611];
     layer0_out[8700] <= ~(x[7394] ^ x[7395]);
     layer0_out[8701] <= ~(x[844] | x[845]);
     layer0_out[8702] <= x[1331] & x[1333];
     layer0_out[8703] <= ~(x[1696] & x[1697]);
     layer0_out[8704] <= ~x[5935] | x[5934];
     layer0_out[8705] <= ~(x[2329] ^ x[2330]);
     layer0_out[8706] <= ~(x[906] | x[907]);
     layer0_out[8707] <= x[1692] ^ x[1694];
     layer0_out[8708] <= ~(x[9131] ^ x[9132]);
     layer0_out[8709] <= x[4753] & x[4754];
     layer0_out[8710] <= ~(x[3546] | x[3547]);
     layer0_out[8711] <= x[2745] | x[2747];
     layer0_out[8712] <= x[1157] & x[1159];
     layer0_out[8713] <= x[1226] & x[1228];
     layer0_out[8714] <= ~(x[1836] & x[1838]);
     layer0_out[8715] <= x[272];
     layer0_out[8716] <= ~x[245];
     layer0_out[8717] <= x[3828];
     layer0_out[8718] <= x[2485];
     layer0_out[8719] <= x[1154] | x[1155];
     layer0_out[8720] <= x[3288] | x[3289];
     layer0_out[8721] <= x[5677];
     layer0_out[8722] <= ~x[6823];
     layer0_out[8723] <= x[152];
     layer0_out[8724] <= ~(x[366] & x[367]);
     layer0_out[8725] <= ~x[1861];
     layer0_out[8726] <= ~(x[8451] & x[8452]);
     layer0_out[8727] <= ~(x[7167] ^ x[7168]);
     layer0_out[8728] <= ~(x[6950] | x[6951]);
     layer0_out[8729] <= x[2493] & x[2494];
     layer0_out[8730] <= ~(x[6458] ^ x[6459]);
     layer0_out[8731] <= ~x[1232];
     layer0_out[8732] <= ~x[5953];
     layer0_out[8733] <= x[3657] & ~x[3656];
     layer0_out[8734] <= x[6432] | x[6433];
     layer0_out[8735] <= x[2775] ^ x[2777];
     layer0_out[8736] <= x[412] | x[413];
     layer0_out[8737] <= x[84] & x[85];
     layer0_out[8738] <= ~(x[8567] ^ x[8568]);
     layer0_out[8739] <= ~(x[978] | x[980]);
     layer0_out[8740] <= x[7733] | x[7734];
     layer0_out[8741] <= ~x[5686];
     layer0_out[8742] <= ~(x[1171] ^ x[1173]);
     layer0_out[8743] <= ~(x[1557] & x[1558]);
     layer0_out[8744] <= 1'b1;
     layer0_out[8745] <= ~(x[2157] & x[2158]);
     layer0_out[8746] <= ~(x[3615] & x[3616]);
     layer0_out[8747] <= x[1248] & x[1249];
     layer0_out[8748] <= ~x[8665] | x[8664];
     layer0_out[8749] <= ~x[5875];
     layer0_out[8750] <= x[5643];
     layer0_out[8751] <= x[3750] | x[3751];
     layer0_out[8752] <= x[3464] | x[3465];
     layer0_out[8753] <= ~(x[5615] | x[5616]);
     layer0_out[8754] <= x[8720];
     layer0_out[8755] <= x[2593] & ~x[2594];
     layer0_out[8756] <= x[6767] & ~x[6768];
     layer0_out[8757] <= ~(x[1060] ^ x[1062]);
     layer0_out[8758] <= ~x[78] | x[79];
     layer0_out[8759] <= x[1966] & x[1968];
     layer0_out[8760] <= ~(x[7464] & x[7465]);
     layer0_out[8761] <= x[3130];
     layer0_out[8762] <= x[8904] & x[8905];
     layer0_out[8763] <= ~(x[7520] ^ x[7521]);
     layer0_out[8764] <= x[373];
     layer0_out[8765] <= x[7527];
     layer0_out[8766] <= x[2750] & x[2752];
     layer0_out[8767] <= x[6500] & x[6501];
     layer0_out[8768] <= ~(x[3646] | x[3647]);
     layer0_out[8769] <= x[6869] & ~x[6870];
     layer0_out[8770] <= x[8590] | x[8591];
     layer0_out[8771] <= x[4360] ^ x[4361];
     layer0_out[8772] <= ~(x[2587] & x[2588]);
     layer0_out[8773] <= ~(x[5007] | x[5008]);
     layer0_out[8774] <= x[437] | x[438];
     layer0_out[8775] <= ~x[2412] | x[2411];
     layer0_out[8776] <= ~(x[8347] & x[8348]);
     layer0_out[8777] <= x[6718];
     layer0_out[8778] <= ~x[3920];
     layer0_out[8779] <= x[960] | x[961];
     layer0_out[8780] <= 1'b0;
     layer0_out[8781] <= x[4805] & x[4806];
     layer0_out[8782] <= ~(x[8676] ^ x[8677]);
     layer0_out[8783] <= x[2793];
     layer0_out[8784] <= ~x[5732];
     layer0_out[8785] <= x[1281] ^ x[1282];
     layer0_out[8786] <= ~x[5971] | x[5970];
     layer0_out[8787] <= ~(x[4820] & x[4821]);
     layer0_out[8788] <= 1'b1;
     layer0_out[8789] <= ~(x[6961] ^ x[6962]);
     layer0_out[8790] <= ~(x[2629] ^ x[2631]);
     layer0_out[8791] <= 1'b1;
     layer0_out[8792] <= ~x[6542];
     layer0_out[8793] <= ~(x[4148] & x[4149]);
     layer0_out[8794] <= ~(x[4478] ^ x[4479]);
     layer0_out[8795] <= x[7013] & x[7014];
     layer0_out[8796] <= ~x[384] | x[386];
     layer0_out[8797] <= x[2504];
     layer0_out[8798] <= x[1015] ^ x[1016];
     layer0_out[8799] <= x[1314] & x[1316];
     layer0_out[8800] <= ~(x[6653] | x[6654]);
     layer0_out[8801] <= x[6027] & x[6028];
     layer0_out[8802] <= x[2627] ^ x[2629];
     layer0_out[8803] <= x[8198];
     layer0_out[8804] <= ~x[1469] | x[1467];
     layer0_out[8805] <= ~(x[1247] & x[1248]);
     layer0_out[8806] <= x[6436];
     layer0_out[8807] <= ~x[9139];
     layer0_out[8808] <= x[184] | x[186];
     layer0_out[8809] <= x[752];
     layer0_out[8810] <= x[2646] & x[2647];
     layer0_out[8811] <= 1'b1;
     layer0_out[8812] <= ~(x[1995] | x[1997]);
     layer0_out[8813] <= x[4564] ^ x[4565];
     layer0_out[8814] <= ~(x[2542] & x[2543]);
     layer0_out[8815] <= ~x[8879] | x[8878];
     layer0_out[8816] <= ~(x[2764] & x[2765]);
     layer0_out[8817] <= ~(x[2933] ^ x[2934]);
     layer0_out[8818] <= x[110];
     layer0_out[8819] <= ~(x[739] & x[740]);
     layer0_out[8820] <= ~x[369];
     layer0_out[8821] <= x[235];
     layer0_out[8822] <= x[3780] & x[3781];
     layer0_out[8823] <= x[3123] | x[3124];
     layer0_out[8824] <= ~(x[1605] & x[1606]);
     layer0_out[8825] <= x[61] & x[62];
     layer0_out[8826] <= x[990];
     layer0_out[8827] <= ~x[8121];
     layer0_out[8828] <= ~(x[2042] | x[2043]);
     layer0_out[8829] <= x[1925] | x[1926];
     layer0_out[8830] <= x[2056] & x[2058];
     layer0_out[8831] <= ~x[398];
     layer0_out[8832] <= ~(x[5910] ^ x[5911]);
     layer0_out[8833] <= x[5681] & x[5682];
     layer0_out[8834] <= ~(x[1901] & x[1902]);
     layer0_out[8835] <= ~(x[2017] & x[2019]);
     layer0_out[8836] <= ~x[8905];
     layer0_out[8837] <= ~(x[4761] & x[4762]);
     layer0_out[8838] <= x[8017] | x[8018];
     layer0_out[8839] <= ~(x[4037] ^ x[4038]);
     layer0_out[8840] <= ~x[1605];
     layer0_out[8841] <= x[1444] & ~x[1443];
     layer0_out[8842] <= ~(x[1032] & x[1033]);
     layer0_out[8843] <= x[6441] & ~x[6440];
     layer0_out[8844] <= x[2395] ^ x[2397];
     layer0_out[8845] <= x[1355] & x[1356];
     layer0_out[8846] <= ~(x[2002] | x[2004]);
     layer0_out[8847] <= 1'b0;
     layer0_out[8848] <= x[9184] | x[9185];
     layer0_out[8849] <= ~(x[1201] | x[1202]);
     layer0_out[8850] <= ~x[1917];
     layer0_out[8851] <= ~(x[3185] & x[3186]);
     layer0_out[8852] <= x[7004] ^ x[7005];
     layer0_out[8853] <= x[8944] & ~x[8945];
     layer0_out[8854] <= x[4387] ^ x[4388];
     layer0_out[8855] <= x[5014] & x[5015];
     layer0_out[8856] <= 1'b1;
     layer0_out[8857] <= ~x[2424] | x[2425];
     layer0_out[8858] <= ~(x[8710] | x[8711]);
     layer0_out[8859] <= x[4039] & x[4040];
     layer0_out[8860] <= x[1014] | x[1015];
     layer0_out[8861] <= ~x[1509];
     layer0_out[8862] <= ~(x[7008] & x[7009]);
     layer0_out[8863] <= ~x[3312] | x[3311];
     layer0_out[8864] <= x[1773] | x[1774];
     layer0_out[8865] <= ~(x[6376] | x[6377]);
     layer0_out[8866] <= ~(x[1485] | x[1487]);
     layer0_out[8867] <= x[874];
     layer0_out[8868] <= 1'b0;
     layer0_out[8869] <= ~x[2565];
     layer0_out[8870] <= ~(x[2266] ^ x[2268]);
     layer0_out[8871] <= ~(x[3253] | x[3254]);
     layer0_out[8872] <= ~(x[4446] ^ x[4447]);
     layer0_out[8873] <= ~(x[5246] & x[5247]);
     layer0_out[8874] <= ~x[5418];
     layer0_out[8875] <= 1'b0;
     layer0_out[8876] <= x[5646] & x[5647];
     layer0_out[8877] <= ~(x[4521] & x[4522]);
     layer0_out[8878] <= ~(x[2070] | x[2072]);
     layer0_out[8879] <= x[698] & x[699];
     layer0_out[8880] <= ~(x[1118] & x[1119]);
     layer0_out[8881] <= ~(x[2067] & x[2068]);
     layer0_out[8882] <= ~(x[5291] & x[5292]);
     layer0_out[8883] <= x[547] ^ x[549];
     layer0_out[8884] <= ~x[6331];
     layer0_out[8885] <= ~x[901];
     layer0_out[8886] <= 1'b0;
     layer0_out[8887] <= ~(x[5182] & x[5183]);
     layer0_out[8888] <= ~(x[587] ^ x[588]);
     layer0_out[8889] <= x[101] & x[102];
     layer0_out[8890] <= x[2586] & ~x[2585];
     layer0_out[8891] <= x[2669] & ~x[2667];
     layer0_out[8892] <= ~(x[6753] & x[6754]);
     layer0_out[8893] <= ~(x[4835] | x[4836]);
     layer0_out[8894] <= x[4698] & x[4699];
     layer0_out[8895] <= ~(x[6472] & x[6473]);
     layer0_out[8896] <= ~(x[6367] | x[6368]);
     layer0_out[8897] <= ~(x[494] & x[495]);
     layer0_out[8898] <= x[3381] | x[3382];
     layer0_out[8899] <= x[2675] | x[2676];
     layer0_out[8900] <= x[2394];
     layer0_out[8901] <= x[281] & x[282];
     layer0_out[8902] <= ~(x[3652] | x[3653]);
     layer0_out[8903] <= ~(x[3678] | x[3679]);
     layer0_out[8904] <= x[1289] & x[1290];
     layer0_out[8905] <= ~x[2295];
     layer0_out[8906] <= x[4529];
     layer0_out[8907] <= ~x[1190];
     layer0_out[8908] <= ~(x[5999] ^ x[6000]);
     layer0_out[8909] <= 1'b0;
     layer0_out[8910] <= x[1951] & x[1953];
     layer0_out[8911] <= x[7926];
     layer0_out[8912] <= ~(x[3747] & x[3748]);
     layer0_out[8913] <= x[4139];
     layer0_out[8914] <= ~(x[2335] | x[2336]);
     layer0_out[8915] <= 1'b1;
     layer0_out[8916] <= x[3449] | x[3450];
     layer0_out[8917] <= ~(x[2311] & x[2313]);
     layer0_out[8918] <= ~(x[4073] | x[4074]);
     layer0_out[8919] <= x[1622] & x[1623];
     layer0_out[8920] <= x[861];
     layer0_out[8921] <= ~(x[8847] | x[8848]);
     layer0_out[8922] <= 1'b0;
     layer0_out[8923] <= ~(x[5290] & x[5291]);
     layer0_out[8924] <= 1'b0;
     layer0_out[8925] <= ~(x[1844] & x[1846]);
     layer0_out[8926] <= ~(x[769] ^ x[771]);
     layer0_out[8927] <= x[2601] & x[2603];
     layer0_out[8928] <= x[4113] & ~x[4114];
     layer0_out[8929] <= ~(x[171] ^ x[173]);
     layer0_out[8930] <= ~(x[5745] | x[5746]);
     layer0_out[8931] <= ~x[1346];
     layer0_out[8932] <= ~(x[5058] & x[5059]);
     layer0_out[8933] <= ~x[3816];
     layer0_out[8934] <= ~x[4155] | x[4156];
     layer0_out[8935] <= x[1515] & x[1517];
     layer0_out[8936] <= ~(x[424] | x[425]);
     layer0_out[8937] <= x[5469] & x[5470];
     layer0_out[8938] <= 1'b0;
     layer0_out[8939] <= 1'b1;
     layer0_out[8940] <= x[1851] & x[1853];
     layer0_out[8941] <= ~(x[417] | x[418]);
     layer0_out[8942] <= x[3066];
     layer0_out[8943] <= x[8605];
     layer0_out[8944] <= ~(x[3550] & x[3551]);
     layer0_out[8945] <= ~x[2758];
     layer0_out[8946] <= ~(x[540] ^ x[542]);
     layer0_out[8947] <= x[1621];
     layer0_out[8948] <= x[3274];
     layer0_out[8949] <= x[2013] | x[2014];
     layer0_out[8950] <= x[8172];
     layer0_out[8951] <= x[238] | x[240];
     layer0_out[8952] <= ~(x[293] | x[294]);
     layer0_out[8953] <= ~(x[1984] & x[1986]);
     layer0_out[8954] <= ~(x[810] & x[811]);
     layer0_out[8955] <= 1'b0;
     layer0_out[8956] <= ~x[147];
     layer0_out[8957] <= 1'b1;
     layer0_out[8958] <= ~(x[2894] & x[2895]);
     layer0_out[8959] <= ~(x[2907] & x[2908]);
     layer0_out[8960] <= 1'b0;
     layer0_out[8961] <= ~(x[3167] ^ x[3168]);
     layer0_out[8962] <= x[6013];
     layer0_out[8963] <= ~(x[1737] & x[1739]);
     layer0_out[8964] <= x[496];
     layer0_out[8965] <= ~x[1593] | x[1594];
     layer0_out[8966] <= x[8228] ^ x[8229];
     layer0_out[8967] <= ~x[891] | x[893];
     layer0_out[8968] <= x[7989] & x[7990];
     layer0_out[8969] <= x[2502] & x[2503];
     layer0_out[8970] <= x[3571] ^ x[3572];
     layer0_out[8971] <= x[856] & x[857];
     layer0_out[8972] <= x[1572] & ~x[1573];
     layer0_out[8973] <= ~(x[6093] & x[6094]);
     layer0_out[8974] <= 1'b1;
     layer0_out[8975] <= x[697] ^ x[699];
     layer0_out[8976] <= x[1411] ^ x[1413];
     layer0_out[8977] <= ~x[4111];
     layer0_out[8978] <= ~x[595] | x[594];
     layer0_out[8979] <= x[1123] | x[1124];
     layer0_out[8980] <= ~(x[3367] ^ x[3368]);
     layer0_out[8981] <= x[749];
     layer0_out[8982] <= x[3144] ^ x[3145];
     layer0_out[8983] <= x[2418] & x[2420];
     layer0_out[8984] <= ~x[7613];
     layer0_out[8985] <= ~(x[428] & x[429]);
     layer0_out[8986] <= x[5348] & ~x[5349];
     layer0_out[8987] <= x[7603] | x[7604];
     layer0_out[8988] <= x[552] ^ x[553];
     layer0_out[8989] <= ~(x[8270] & x[8271]);
     layer0_out[8990] <= ~(x[284] | x[286]);
     layer0_out[8991] <= ~x[7817] | x[7816];
     layer0_out[8992] <= x[4872];
     layer0_out[8993] <= x[2287] & x[2289];
     layer0_out[8994] <= ~x[8844];
     layer0_out[8995] <= x[2446] & x[2447];
     layer0_out[8996] <= x[2494] & x[2495];
     layer0_out[8997] <= ~x[1168];
     layer0_out[8998] <= x[3895] ^ x[3896];
     layer0_out[8999] <= ~(x[5796] & x[5797]);
     layer0_out[9000] <= x[8037] ^ x[8038];
     layer0_out[9001] <= x[5699] ^ x[5700];
     layer0_out[9002] <= x[4517] & x[4518];
     layer0_out[9003] <= x[4252] & x[4253];
     layer0_out[9004] <= 1'b1;
     layer0_out[9005] <= ~x[4711];
     layer0_out[9006] <= x[336];
     layer0_out[9007] <= x[1227] & x[1228];
     layer0_out[9008] <= ~x[3817];
     layer0_out[9009] <= 1'b1;
     layer0_out[9010] <= ~(x[872] & x[873]);
     layer0_out[9011] <= x[7294];
     layer0_out[9012] <= ~x[504];
     layer0_out[9013] <= x[1193] & x[1194];
     layer0_out[9014] <= ~(x[5849] | x[5850]);
     layer0_out[9015] <= ~(x[6120] & x[6121]);
     layer0_out[9016] <= ~x[529] | x[531];
     layer0_out[9017] <= x[5735];
     layer0_out[9018] <= x[1897];
     layer0_out[9019] <= x[8863];
     layer0_out[9020] <= ~x[3596];
     layer0_out[9021] <= ~(x[7677] ^ x[7678]);
     layer0_out[9022] <= x[5719];
     layer0_out[9023] <= 1'b0;
     layer0_out[9024] <= x[5848] & x[5849];
     layer0_out[9025] <= x[2154];
     layer0_out[9026] <= ~(x[7567] | x[7568]);
     layer0_out[9027] <= ~x[1465];
     layer0_out[9028] <= ~(x[2357] & x[2359]);
     layer0_out[9029] <= ~x[5786];
     layer0_out[9030] <= x[362] ^ x[364];
     layer0_out[9031] <= x[1150] & x[1152];
     layer0_out[9032] <= x[3718] & ~x[3717];
     layer0_out[9033] <= ~(x[1511] ^ x[1512]);
     layer0_out[9034] <= x[5510] | x[5511];
     layer0_out[9035] <= x[836];
     layer0_out[9036] <= ~(x[261] & x[263]);
     layer0_out[9037] <= ~(x[7392] | x[7393]);
     layer0_out[9038] <= ~x[4249];
     layer0_out[9039] <= x[916] & ~x[918];
     layer0_out[9040] <= x[4334];
     layer0_out[9041] <= ~(x[3817] | x[3818]);
     layer0_out[9042] <= ~x[6];
     layer0_out[9043] <= ~x[2511];
     layer0_out[9044] <= ~x[4894];
     layer0_out[9045] <= x[7181] & x[7182];
     layer0_out[9046] <= x[9094] & x[9095];
     layer0_out[9047] <= x[2819] | x[2820];
     layer0_out[9048] <= ~(x[3266] | x[3267]);
     layer0_out[9049] <= ~(x[6447] ^ x[6448]);
     layer0_out[9050] <= x[970] & ~x[971];
     layer0_out[9051] <= x[2668] & x[2670];
     layer0_out[9052] <= ~x[1563];
     layer0_out[9053] <= ~(x[4952] ^ x[4953]);
     layer0_out[9054] <= ~(x[958] & x[959]);
     layer0_out[9055] <= x[6977] ^ x[6978];
     layer0_out[9056] <= x[2815] & x[2816];
     layer0_out[9057] <= 1'b0;
     layer0_out[9058] <= ~(x[2066] & x[2067]);
     layer0_out[9059] <= ~x[6720];
     layer0_out[9060] <= 1'b0;
     layer0_out[9061] <= ~x[592];
     layer0_out[9062] <= x[1911];
     layer0_out[9063] <= ~(x[7660] | x[7661]);
     layer0_out[9064] <= x[884] & x[885];
     layer0_out[9065] <= ~(x[5214] & x[5215]);
     layer0_out[9066] <= x[4534] | x[4535];
     layer0_out[9067] <= ~(x[2285] & x[2287]);
     layer0_out[9068] <= x[47] ^ x[49];
     layer0_out[9069] <= ~(x[2298] ^ x[2300]);
     layer0_out[9070] <= x[789] | x[791];
     layer0_out[9071] <= x[2574] | x[2576];
     layer0_out[9072] <= ~(x[1044] & x[1046]);
     layer0_out[9073] <= ~(x[1360] ^ x[1361]);
     layer0_out[9074] <= ~(x[5044] ^ x[5045]);
     layer0_out[9075] <= ~x[846];
     layer0_out[9076] <= ~(x[6522] ^ x[6523]);
     layer0_out[9077] <= ~x[4558];
     layer0_out[9078] <= x[5404];
     layer0_out[9079] <= ~(x[9205] | x[9206]);
     layer0_out[9080] <= x[443] & x[444];
     layer0_out[9081] <= ~(x[7479] & x[7480]);
     layer0_out[9082] <= ~(x[9009] | x[9010]);
     layer0_out[9083] <= x[8209] | x[8210];
     layer0_out[9084] <= 1'b1;
     layer0_out[9085] <= x[2393] ^ x[2395];
     layer0_out[9086] <= ~(x[2216] & x[2217]);
     layer0_out[9087] <= ~(x[4248] | x[4249]);
     layer0_out[9088] <= ~(x[5334] | x[5335]);
     layer0_out[9089] <= 1'b1;
     layer0_out[9090] <= ~(x[2305] & x[2306]);
     layer0_out[9091] <= x[5092] & x[5093];
     layer0_out[9092] <= ~(x[4100] & x[4101]);
     layer0_out[9093] <= x[1053] & x[1054];
     layer0_out[9094] <= ~x[459] | x[458];
     layer0_out[9095] <= ~(x[301] | x[303]);
     layer0_out[9096] <= ~x[3893] | x[3894];
     layer0_out[9097] <= x[8928];
     layer0_out[9098] <= x[2496] | x[2497];
     layer0_out[9099] <= x[4483];
     layer0_out[9100] <= ~x[5979] | x[5978];
     layer0_out[9101] <= x[25] & x[26];
     layer0_out[9102] <= ~(x[7746] | x[7747]);
     layer0_out[9103] <= x[8318];
     layer0_out[9104] <= x[7131] | x[7132];
     layer0_out[9105] <= ~(x[2637] & x[2638]);
     layer0_out[9106] <= x[2587] & x[2589];
     layer0_out[9107] <= x[3106] | x[3107];
     layer0_out[9108] <= ~(x[2277] & x[2279]);
     layer0_out[9109] <= x[765] ^ x[766];
     layer0_out[9110] <= ~(x[8359] ^ x[8360]);
     layer0_out[9111] <= ~(x[244] ^ x[245]);
     layer0_out[9112] <= x[5263] & x[5264];
     layer0_out[9113] <= x[1929] & x[1931];
     layer0_out[9114] <= x[5503] ^ x[5504];
     layer0_out[9115] <= x[5232] & x[5233];
     layer0_out[9116] <= x[2916] ^ x[2917];
     layer0_out[9117] <= x[2349];
     layer0_out[9118] <= x[4904];
     layer0_out[9119] <= x[793] ^ x[795];
     layer0_out[9120] <= 1'b1;
     layer0_out[9121] <= ~x[3507];
     layer0_out[9122] <= x[8133] | x[8134];
     layer0_out[9123] <= ~(x[8090] ^ x[8091]);
     layer0_out[9124] <= ~(x[1403] & x[1404]);
     layer0_out[9125] <= x[3187] ^ x[3188];
     layer0_out[9126] <= ~(x[1782] ^ x[1783]);
     layer0_out[9127] <= x[256];
     layer0_out[9128] <= x[8597] & x[8598];
     layer0_out[9129] <= x[2036] & x[2037];
     layer0_out[9130] <= x[4584] ^ x[4585];
     layer0_out[9131] <= ~x[2276];
     layer0_out[9132] <= x[5012] | x[5013];
     layer0_out[9133] <= ~(x[4512] & x[4513]);
     layer0_out[9134] <= x[7922];
     layer0_out[9135] <= ~x[6216] | x[6215];
     layer0_out[9136] <= ~x[3834];
     layer0_out[9137] <= x[5566];
     layer0_out[9138] <= x[1431] & x[1433];
     layer0_out[9139] <= x[4437] & x[4438];
     layer0_out[9140] <= x[8492] | x[8493];
     layer0_out[9141] <= 1'b0;
     layer0_out[9142] <= x[2581] ^ x[2583];
     layer0_out[9143] <= ~(x[4216] | x[4217]);
     layer0_out[9144] <= ~(x[751] & x[753]);
     layer0_out[9145] <= ~(x[7813] & x[7814]);
     layer0_out[9146] <= x[2130] | x[2131];
     layer0_out[9147] <= x[5585];
     layer0_out[9148] <= ~(x[5769] & x[5770]);
     layer0_out[9149] <= ~(x[2398] & x[2399]);
     layer0_out[9150] <= ~x[6268];
     layer0_out[9151] <= x[7083];
     layer0_out[9152] <= ~(x[5957] ^ x[5958]);
     layer0_out[9153] <= x[5892] & ~x[5893];
     layer0_out[9154] <= x[2006] | x[2007];
     layer0_out[9155] <= 1'b1;
     layer0_out[9156] <= ~(x[2186] & x[2187]);
     layer0_out[9157] <= x[1259] & x[1261];
     layer0_out[9158] <= ~(x[1452] ^ x[1454]);
     layer0_out[9159] <= x[299] & ~x[300];
     layer0_out[9160] <= ~(x[8303] & x[8304]);
     layer0_out[9161] <= 1'b1;
     layer0_out[9162] <= x[5253] & x[5254];
     layer0_out[9163] <= 1'b1;
     layer0_out[9164] <= x[2365] & ~x[2367];
     layer0_out[9165] <= x[964] | x[965];
     layer0_out[9166] <= x[1196] & x[1197];
     layer0_out[9167] <= ~(x[450] ^ x[452]);
     layer0_out[9168] <= ~(x[8481] | x[8482]);
     layer0_out[9169] <= x[5082] ^ x[5083];
     layer0_out[9170] <= ~(x[5579] & x[5580]);
     layer0_out[9171] <= x[3539] ^ x[3540];
     layer0_out[9172] <= ~x[8100] | x[8101];
     layer0_out[9173] <= x[6132] & x[6133];
     layer0_out[9174] <= x[8066] ^ x[8067];
     layer0_out[9175] <= x[614] | x[615];
     layer0_out[9176] <= ~x[2163];
     layer0_out[9177] <= ~(x[366] & x[368]);
     layer0_out[9178] <= ~(x[418] | x[420]);
     layer0_out[9179] <= 1'b1;
     layer0_out[9180] <= ~(x[6011] & x[6012]);
     layer0_out[9181] <= ~x[8647];
     layer0_out[9182] <= ~(x[9] ^ x[11]);
     layer0_out[9183] <= ~(x[1325] & x[1327]);
     layer0_out[9184] <= x[1635] & x[1637];
     layer0_out[9185] <= ~x[8399];
     layer0_out[9186] <= ~(x[306] & x[307]);
     layer0_out[9187] <= x[7015] & x[7016];
     layer0_out[9188] <= ~x[8027];
     layer0_out[9189] <= 1'b1;
     layer0_out[9190] <= x[1204] | x[1205];
     layer0_out[9191] <= x[1111] | x[1112];
     layer0_out[9192] <= ~(x[5371] & x[5372]);
     layer0_out[9193] <= x[2568] ^ x[2569];
     layer0_out[9194] <= 1'b0;
     layer0_out[9195] <= x[1526] | x[1528];
     layer0_out[9196] <= x[8301] ^ x[8302];
     layer0_out[9197] <= ~(x[4378] & x[4379]);
     layer0_out[9198] <= ~x[7024] | x[7025];
     layer0_out[9199] <= ~(x[9123] & x[9124]);
     layer0_out[9200] <= 1'b0;
     layer0_out[9201] <= ~(x[6463] | x[6464]);
     layer0_out[9202] <= x[2604] & x[2606];
     layer0_out[9203] <= ~(x[25] | x[27]);
     layer0_out[9204] <= ~x[3444] | x[3443];
     layer0_out[9205] <= ~(x[992] & x[993]);
     layer0_out[9206] <= ~(x[831] & x[833]);
     layer0_out[9207] <= x[307] & x[308];
     layer0_out[9208] <= ~x[1785] | x[1787];
     layer0_out[9209] <= x[429];
     layer0_out[9210] <= x[8272] & ~x[8271];
     layer0_out[9211] <= ~(x[4664] & x[4665]);
     layer0_out[9212] <= x[210];
     layer0_out[9213] <= ~(x[8159] | x[8160]);
     layer0_out[9214] <= x[1525] & x[1526];
     layer0_out[9215] <= x[1277] & x[1279];
     layer0_out[9216] <= ~x[1219];
     layer0_out[9217] <= x[2485];
     layer0_out[9218] <= ~(x[5629] & x[5630]);
     layer0_out[9219] <= ~x[2326];
     layer0_out[9220] <= ~(x[4851] | x[4852]);
     layer0_out[9221] <= x[967];
     layer0_out[9222] <= 1'b1;
     layer0_out[9223] <= x[2710] & ~x[2709];
     layer0_out[9224] <= x[5639] ^ x[5640];
     layer0_out[9225] <= x[4273];
     layer0_out[9226] <= ~(x[3536] ^ x[3537]);
     layer0_out[9227] <= x[8010] & x[8011];
     layer0_out[9228] <= ~(x[4272] & x[4273]);
     layer0_out[9229] <= x[3878] | x[3879];
     layer0_out[9230] <= 1'b0;
     layer0_out[9231] <= x[1804] ^ x[1805];
     layer0_out[9232] <= x[144] & x[146];
     layer0_out[9233] <= ~(x[2979] & x[2980]);
     layer0_out[9234] <= 1'b1;
     layer0_out[9235] <= x[930];
     layer0_out[9236] <= 1'b0;
     layer0_out[9237] <= x[318] | x[320];
     layer0_out[9238] <= ~(x[1957] & x[1959]);
     layer0_out[9239] <= 1'b1;
     layer0_out[9240] <= x[3920] | x[3921];
     layer0_out[9241] <= x[9128] | x[9129];
     layer0_out[9242] <= 1'b1;
     layer0_out[9243] <= x[680] & x[682];
     layer0_out[9244] <= ~x[2216] | x[2214];
     layer0_out[9245] <= ~(x[7286] | x[7287]);
     layer0_out[9246] <= x[8167] & ~x[8168];
     layer0_out[9247] <= x[6091] & x[6092];
     layer0_out[9248] <= ~(x[2474] ^ x[2475]);
     layer0_out[9249] <= x[404] ^ x[406];
     layer0_out[9250] <= ~x[8990];
     layer0_out[9251] <= ~(x[1659] | x[1661]);
     layer0_out[9252] <= x[4973];
     layer0_out[9253] <= x[3204] ^ x[3205];
     layer0_out[9254] <= x[1468] | x[1470];
     layer0_out[9255] <= x[5969] & x[5970];
     layer0_out[9256] <= x[2468] ^ x[2470];
     layer0_out[9257] <= ~x[5756] | x[5757];
     layer0_out[9258] <= ~x[4464];
     layer0_out[9259] <= ~x[1856];
     layer0_out[9260] <= x[615] ^ x[617];
     layer0_out[9261] <= 1'b1;
     layer0_out[9262] <= x[6713] | x[6714];
     layer0_out[9263] <= ~(x[6483] ^ x[6484]);
     layer0_out[9264] <= ~(x[5256] & x[5257]);
     layer0_out[9265] <= ~(x[572] ^ x[573]);
     layer0_out[9266] <= ~x[3197];
     layer0_out[9267] <= 1'b1;
     layer0_out[9268] <= x[2386] & x[2387];
     layer0_out[9269] <= x[5932] | x[5933];
     layer0_out[9270] <= x[1686] & x[1688];
     layer0_out[9271] <= ~(x[162] ^ x[163]);
     layer0_out[9272] <= x[1877] | x[1878];
     layer0_out[9273] <= x[6080];
     layer0_out[9274] <= ~(x[6098] & x[6099]);
     layer0_out[9275] <= x[2136] ^ x[2137];
     layer0_out[9276] <= ~x[3754];
     layer0_out[9277] <= ~(x[3701] & x[3702]);
     layer0_out[9278] <= x[7094] | x[7095];
     layer0_out[9279] <= x[6799] ^ x[6800];
     layer0_out[9280] <= x[1617] & x[1619];
     layer0_out[9281] <= x[3762] | x[3763];
     layer0_out[9282] <= ~(x[1430] ^ x[1431]);
     layer0_out[9283] <= ~(x[4961] ^ x[4962]);
     layer0_out[9284] <= x[3674];
     layer0_out[9285] <= x[2887];
     layer0_out[9286] <= x[3447] | x[3448];
     layer0_out[9287] <= ~(x[7742] & x[7743]);
     layer0_out[9288] <= x[486] & x[487];
     layer0_out[9289] <= ~(x[1287] & x[1288]);
     layer0_out[9290] <= ~x[2212];
     layer0_out[9291] <= ~x[3328] | x[3327];
     layer0_out[9292] <= ~(x[3664] | x[3665]);
     layer0_out[9293] <= ~(x[420] | x[422]);
     layer0_out[9294] <= ~(x[214] & x[216]);
     layer0_out[9295] <= ~(x[3716] ^ x[3717]);
     layer0_out[9296] <= x[3180] & ~x[3181];
     layer0_out[9297] <= x[5259] & x[5260];
     layer0_out[9298] <= 1'b0;
     layer0_out[9299] <= x[6073] | x[6074];
     layer0_out[9300] <= ~x[523] | x[521];
     layer0_out[9301] <= x[2544] & x[2546];
     layer0_out[9302] <= x[6442];
     layer0_out[9303] <= ~(x[41] & x[43]);
     layer0_out[9304] <= x[3627] & x[3628];
     layer0_out[9305] <= x[2944] & x[2945];
     layer0_out[9306] <= x[7629] | x[7630];
     layer0_out[9307] <= ~(x[5022] & x[5023]);
     layer0_out[9308] <= x[60] & x[62];
     layer0_out[9309] <= x[1427] & x[1429];
     layer0_out[9310] <= ~x[926] | x[924];
     layer0_out[9311] <= ~x[1566];
     layer0_out[9312] <= ~(x[2670] | x[2672]);
     layer0_out[9313] <= x[1798] | x[1799];
     layer0_out[9314] <= x[2288] | x[2290];
     layer0_out[9315] <= 1'b0;
     layer0_out[9316] <= x[467] & ~x[465];
     layer0_out[9317] <= x[933];
     layer0_out[9318] <= ~(x[4677] | x[4678]);
     layer0_out[9319] <= x[626] & x[627];
     layer0_out[9320] <= x[1305] & x[1307];
     layer0_out[9321] <= ~x[809];
     layer0_out[9322] <= 1'b1;
     layer0_out[9323] <= x[6624] | x[6625];
     layer0_out[9324] <= x[111];
     layer0_out[9325] <= 1'b1;
     layer0_out[9326] <= 1'b0;
     layer0_out[9327] <= ~(x[4540] & x[4541]);
     layer0_out[9328] <= x[903] | x[904];
     layer0_out[9329] <= ~x[1661];
     layer0_out[9330] <= x[1521];
     layer0_out[9331] <= ~x[2457];
     layer0_out[9332] <= ~(x[6620] | x[6621]);
     layer0_out[9333] <= x[733] | x[734];
     layer0_out[9334] <= ~(x[7182] | x[7183]);
     layer0_out[9335] <= x[2102] & x[2104];
     layer0_out[9336] <= ~(x[2657] | x[2658]);
     layer0_out[9337] <= x[29] | x[30];
     layer0_out[9338] <= ~(x[6476] | x[6477]);
     layer0_out[9339] <= ~(x[841] & x[842]);
     layer0_out[9340] <= 1'b0;
     layer0_out[9341] <= x[3562] | x[3563];
     layer0_out[9342] <= ~(x[58] & x[60]);
     layer0_out[9343] <= x[9090] | x[9091];
     layer0_out[9344] <= x[2301] & ~x[2303];
     layer0_out[9345] <= x[5906] & x[5907];
     layer0_out[9346] <= x[713] ^ x[715];
     layer0_out[9347] <= ~x[8274] | x[8273];
     layer0_out[9348] <= x[4537] & x[4538];
     layer0_out[9349] <= ~(x[1346] | x[1348]);
     layer0_out[9350] <= ~x[8602];
     layer0_out[9351] <= ~x[869] | x[871];
     layer0_out[9352] <= ~(x[8659] | x[8660]);
     layer0_out[9353] <= ~x[1305];
     layer0_out[9354] <= x[7105];
     layer0_out[9355] <= ~(x[4786] | x[4787]);
     layer0_out[9356] <= ~(x[2071] & x[2073]);
     layer0_out[9357] <= ~(x[1711] ^ x[1712]);
     layer0_out[9358] <= ~(x[57] & x[58]);
     layer0_out[9359] <= x[8514] ^ x[8515];
     layer0_out[9360] <= ~x[115];
     layer0_out[9361] <= ~x[7966];
     layer0_out[9362] <= x[6142];
     layer0_out[9363] <= x[1489] & x[1491];
     layer0_out[9364] <= ~(x[6137] ^ x[6138]);
     layer0_out[9365] <= ~(x[2134] | x[2136]);
     layer0_out[9366] <= ~(x[4288] | x[4289]);
     layer0_out[9367] <= x[1534] & x[1536];
     layer0_out[9368] <= x[168] & x[169];
     layer0_out[9369] <= 1'b1;
     layer0_out[9370] <= x[8028] ^ x[8029];
     layer0_out[9371] <= ~(x[1013] & x[1014]);
     layer0_out[9372] <= ~x[3420];
     layer0_out[9373] <= ~x[8911];
     layer0_out[9374] <= x[8572] ^ x[8573];
     layer0_out[9375] <= ~x[5431];
     layer0_out[9376] <= x[8388] & x[8389];
     layer0_out[9377] <= ~x[45] | x[43];
     layer0_out[9378] <= ~(x[5023] & x[5024]);
     layer0_out[9379] <= ~(x[8150] & x[8151]);
     layer0_out[9380] <= ~(x[6928] | x[6929]);
     layer0_out[9381] <= x[2720] | x[2722];
     layer0_out[9382] <= ~(x[5605] & x[5606]);
     layer0_out[9383] <= ~x[5589];
     layer0_out[9384] <= ~(x[696] & x[697]);
     layer0_out[9385] <= ~(x[2033] & x[2034]);
     layer0_out[9386] <= ~(x[5674] & x[5675]);
     layer0_out[9387] <= ~(x[2227] ^ x[2229]);
     layer0_out[9388] <= ~(x[3377] ^ x[3378]);
     layer0_out[9389] <= x[5089] | x[5090];
     layer0_out[9390] <= ~x[4067] | x[4068];
     layer0_out[9391] <= ~x[7453];
     layer0_out[9392] <= x[3414];
     layer0_out[9393] <= ~(x[3679] | x[3680]);
     layer0_out[9394] <= x[8223] | x[8224];
     layer0_out[9395] <= x[1895];
     layer0_out[9396] <= ~(x[1330] & x[1332]);
     layer0_out[9397] <= x[1632] & x[1634];
     layer0_out[9398] <= x[7554] | x[7555];
     layer0_out[9399] <= x[7239] & x[7240];
     layer0_out[9400] <= ~(x[8288] & x[8289]);
     layer0_out[9401] <= ~(x[8777] | x[8778]);
     layer0_out[9402] <= ~(x[1172] | x[1173]);
     layer0_out[9403] <= ~x[7093];
     layer0_out[9404] <= x[7924] & ~x[7923];
     layer0_out[9405] <= ~x[478] | x[480];
     layer0_out[9406] <= ~(x[721] ^ x[723]);
     layer0_out[9407] <= x[5560] | x[5561];
     layer0_out[9408] <= ~(x[298] & x[300]);
     layer0_out[9409] <= 1'b0;
     layer0_out[9410] <= ~(x[4282] ^ x[4283]);
     layer0_out[9411] <= ~(x[932] & x[933]);
     layer0_out[9412] <= ~(x[8006] ^ x[8007]);
     layer0_out[9413] <= x[3723] & x[3724];
     layer0_out[9414] <= x[2417] & x[2418];
     layer0_out[9415] <= x[8398] | x[8399];
     layer0_out[9416] <= 1'b0;
     layer0_out[9417] <= x[4879] | x[4880];
     layer0_out[9418] <= 1'b1;
     layer0_out[9419] <= ~x[1017];
     layer0_out[9420] <= x[778] | x[780];
     layer0_out[9421] <= ~(x[896] & x[897]);
     layer0_out[9422] <= x[119] & ~x[118];
     layer0_out[9423] <= ~x[1499];
     layer0_out[9424] <= 1'b1;
     layer0_out[9425] <= ~(x[278] | x[280]);
     layer0_out[9426] <= ~(x[4869] ^ x[4870]);
     layer0_out[9427] <= x[484] ^ x[486];
     layer0_out[9428] <= ~(x[2964] & x[2965]);
     layer0_out[9429] <= ~(x[6837] & x[6838]);
     layer0_out[9430] <= ~(x[8743] & x[8744]);
     layer0_out[9431] <= ~(x[1394] & x[1396]);
     layer0_out[9432] <= ~(x[3830] | x[3831]);
     layer0_out[9433] <= ~(x[5350] & x[5351]);
     layer0_out[9434] <= ~(x[9195] ^ x[9196]);
     layer0_out[9435] <= x[4008] ^ x[4009];
     layer0_out[9436] <= x[1606] & x[1608];
     layer0_out[9437] <= ~x[5635];
     layer0_out[9438] <= ~x[3149];
     layer0_out[9439] <= ~(x[39] | x[41]);
     layer0_out[9440] <= ~(x[303] ^ x[304]);
     layer0_out[9441] <= ~x[2302] | x[2301];
     layer0_out[9442] <= ~(x[1990] ^ x[1991]);
     layer0_out[9443] <= x[858] & x[860];
     layer0_out[9444] <= x[2774] | x[2775];
     layer0_out[9445] <= ~(x[1162] ^ x[1163]);
     layer0_out[9446] <= x[6424] | x[6425];
     layer0_out[9447] <= x[1723] & x[1724];
     layer0_out[9448] <= x[659] & x[660];
     layer0_out[9449] <= ~(x[694] & x[696]);
     layer0_out[9450] <= x[5055] & x[5056];
     layer0_out[9451] <= ~(x[248] ^ x[250]);
     layer0_out[9452] <= x[5810] & x[5811];
     layer0_out[9453] <= ~(x[1007] | x[1009]);
     layer0_out[9454] <= x[5666] & x[5667];
     layer0_out[9455] <= ~(x[1022] & x[1023]);
     layer0_out[9456] <= x[6868] ^ x[6869];
     layer0_out[9457] <= ~(x[926] ^ x[928]);
     layer0_out[9458] <= ~(x[1679] ^ x[1680]);
     layer0_out[9459] <= x[4654] | x[4655];
     layer0_out[9460] <= x[2792] & x[2793];
     layer0_out[9461] <= ~(x[3360] & x[3361]);
     layer0_out[9462] <= ~(x[644] & x[646]);
     layer0_out[9463] <= x[9115] ^ x[9116];
     layer0_out[9464] <= x[53];
     layer0_out[9465] <= ~x[1571] | x[1573];
     layer0_out[9466] <= x[2513] & x[2514];
     layer0_out[9467] <= x[2523];
     layer0_out[9468] <= x[7147] ^ x[7148];
     layer0_out[9469] <= x[5964];
     layer0_out[9470] <= x[1806] & x[1808];
     layer0_out[9471] <= x[3929];
     layer0_out[9472] <= ~x[7906];
     layer0_out[9473] <= x[443] | x[445];
     layer0_out[9474] <= ~(x[4291] ^ x[4292]);
     layer0_out[9475] <= x[6781];
     layer0_out[9476] <= ~(x[39] ^ x[40]);
     layer0_out[9477] <= ~x[1154] | x[1153];
     layer0_out[9478] <= ~x[3608] | x[3609];
     layer0_out[9479] <= ~(x[1183] & x[1185]);
     layer0_out[9480] <= x[172] & x[174];
     layer0_out[9481] <= x[7751] | x[7752];
     layer0_out[9482] <= ~(x[1405] & x[1406]);
     layer0_out[9483] <= ~(x[4888] & x[4889]);
     layer0_out[9484] <= ~x[6741];
     layer0_out[9485] <= x[1646] & ~x[1645];
     layer0_out[9486] <= ~(x[8696] & x[8697]);
     layer0_out[9487] <= ~(x[5] | x[6]);
     layer0_out[9488] <= x[2954] & x[2955];
     layer0_out[9489] <= ~(x[5332] & x[5333]);
     layer0_out[9490] <= x[1742] & x[1743];
     layer0_out[9491] <= ~(x[7943] ^ x[7944]);
     layer0_out[9492] <= ~(x[7647] & x[7648]);
     layer0_out[9493] <= ~(x[1589] | x[1590]);
     layer0_out[9494] <= x[4889];
     layer0_out[9495] <= ~(x[3521] & x[3522]);
     layer0_out[9496] <= x[7415] ^ x[7416];
     layer0_out[9497] <= x[2656] & x[2658];
     layer0_out[9498] <= ~x[8817];
     layer0_out[9499] <= x[8217];
     layer0_out[9500] <= ~x[8416];
     layer0_out[9501] <= ~(x[1748] ^ x[1750]);
     layer0_out[9502] <= x[2125] & x[2127];
     layer0_out[9503] <= ~(x[8177] ^ x[8178]);
     layer0_out[9504] <= ~(x[2035] | x[2036]);
     layer0_out[9505] <= x[3250] & x[3251];
     layer0_out[9506] <= ~(x[3866] | x[3867]);
     layer0_out[9507] <= x[8706] ^ x[8707];
     layer0_out[9508] <= ~(x[1599] & x[1601]);
     layer0_out[9509] <= ~(x[8922] & x[8923]);
     layer0_out[9510] <= x[81] & x[83];
     layer0_out[9511] <= ~x[8019];
     layer0_out[9512] <= x[7223];
     layer0_out[9513] <= ~x[927];
     layer0_out[9514] <= ~(x[2197] & x[2198]);
     layer0_out[9515] <= ~(x[164] & x[165]);
     layer0_out[9516] <= ~(x[4923] ^ x[4924]);
     layer0_out[9517] <= ~(x[1847] & x[1848]);
     layer0_out[9518] <= x[1137];
     layer0_out[9519] <= ~(x[7275] | x[7276]);
     layer0_out[9520] <= ~(x[2422] ^ x[2424]);
     layer0_out[9521] <= x[2668] ^ x[2669];
     layer0_out[9522] <= ~(x[3809] & x[3810]);
     layer0_out[9523] <= x[1112];
     layer0_out[9524] <= x[309] & ~x[308];
     layer0_out[9525] <= ~(x[6565] ^ x[6566]);
     layer0_out[9526] <= 1'b0;
     layer0_out[9527] <= x[6891] ^ x[6892];
     layer0_out[9528] <= ~(x[4498] | x[4499]);
     layer0_out[9529] <= ~x[1374];
     layer0_out[9530] <= ~(x[1043] & x[1045]);
     layer0_out[9531] <= ~(x[5307] & x[5308]);
     layer0_out[9532] <= x[8773] | x[8774];
     layer0_out[9533] <= 1'b1;
     layer0_out[9534] <= 1'b1;
     layer0_out[9535] <= x[5683] & x[5684];
     layer0_out[9536] <= ~(x[2110] & x[2112]);
     layer0_out[9537] <= ~x[2302] | x[2300];
     layer0_out[9538] <= x[6266] | x[6267];
     layer0_out[9539] <= ~x[916];
     layer0_out[9540] <= x[2602] & x[2604];
     layer0_out[9541] <= x[5777] ^ x[5778];
     layer0_out[9542] <= ~x[5823];
     layer0_out[9543] <= ~(x[2433] ^ x[2435]);
     layer0_out[9544] <= x[4535] ^ x[4536];
     layer0_out[9545] <= ~(x[1699] & x[1701]);
     layer0_out[9546] <= ~(x[1405] & x[1407]);
     layer0_out[9547] <= x[5697] & ~x[5696];
     layer0_out[9548] <= x[1602] & x[1604];
     layer0_out[9549] <= x[6707] & x[6708];
     layer0_out[9550] <= ~(x[7829] | x[7830]);
     layer0_out[9551] <= ~x[1113] | x[1112];
     layer0_out[9552] <= x[1933] ^ x[1935];
     layer0_out[9553] <= ~(x[131] & x[133]);
     layer0_out[9554] <= ~x[7600];
     layer0_out[9555] <= 1'b1;
     layer0_out[9556] <= x[4531];
     layer0_out[9557] <= ~(x[4573] & x[4574]);
     layer0_out[9558] <= x[3177] & x[3178];
     layer0_out[9559] <= x[5830] & x[5831];
     layer0_out[9560] <= ~(x[4570] & x[4571]);
     layer0_out[9561] <= ~(x[130] ^ x[131]);
     layer0_out[9562] <= ~x[5591];
     layer0_out[9563] <= ~x[2198];
     layer0_out[9564] <= ~x[1810];
     layer0_out[9565] <= x[7903];
     layer0_out[9566] <= x[5499];
     layer0_out[9567] <= x[3389] | x[3390];
     layer0_out[9568] <= x[8174] ^ x[8175];
     layer0_out[9569] <= ~(x[6965] ^ x[6966]);
     layer0_out[9570] <= x[2756] ^ x[2758];
     layer0_out[9571] <= x[7172] | x[7173];
     layer0_out[9572] <= ~x[8828];
     layer0_out[9573] <= x[4697] | x[4698];
     layer0_out[9574] <= ~(x[827] & x[829]);
     layer0_out[9575] <= x[93] & x[95];
     layer0_out[9576] <= x[8645];
     layer0_out[9577] <= ~(x[1803] & x[1805]);
     layer0_out[9578] <= ~(x[3058] & x[3059]);
     layer0_out[9579] <= ~(x[2453] & x[2454]);
     layer0_out[9580] <= 1'b0;
     layer0_out[9581] <= ~x[3121] | x[3120];
     layer0_out[9582] <= 1'b0;
     layer0_out[9583] <= ~(x[1613] & x[1615]);
     layer0_out[9584] <= x[8281] ^ x[8282];
     layer0_out[9585] <= ~x[5242];
     layer0_out[9586] <= x[507] ^ x[508];
     layer0_out[9587] <= x[7321] | x[7322];
     layer0_out[9588] <= x[915] & x[917];
     layer0_out[9589] <= ~x[1112];
     layer0_out[9590] <= ~(x[2484] & x[2486]);
     layer0_out[9591] <= ~(x[465] | x[466]);
     layer0_out[9592] <= x[2439] & x[2441];
     layer0_out[9593] <= x[957] & ~x[958];
     layer0_out[9594] <= ~(x[5680] | x[5681]);
     layer0_out[9595] <= x[2412] & x[2414];
     layer0_out[9596] <= ~x[1548];
     layer0_out[9597] <= ~(x[3176] & x[3177]);
     layer0_out[9598] <= ~(x[8872] | x[8873]);
     layer0_out[9599] <= ~x[8897];
     layer0_out[9600] <= x[734] ^ x[736];
     layer0_out[9601] <= ~(x[2318] | x[2319]);
     layer0_out[9602] <= ~(x[6183] | x[6184]);
     layer0_out[9603] <= x[1378] & x[1379];
     layer0_out[9604] <= x[7187] & ~x[7186];
     layer0_out[9605] <= x[5146] & x[5147];
     layer0_out[9606] <= ~x[9186];
     layer0_out[9607] <= ~x[2612];
     layer0_out[9608] <= ~(x[3649] & x[3650]);
     layer0_out[9609] <= x[8835] ^ x[8836];
     layer0_out[9610] <= x[8424] & x[8425];
     layer0_out[9611] <= x[3085] | x[3086];
     layer0_out[9612] <= x[5732] & x[5733];
     layer0_out[9613] <= x[5141];
     layer0_out[9614] <= x[2759] | x[2761];
     layer0_out[9615] <= ~(x[2466] ^ x[2468]);
     layer0_out[9616] <= ~(x[2745] ^ x[2746]);
     layer0_out[9617] <= x[9182] & x[9183];
     layer0_out[9618] <= x[2063];
     layer0_out[9619] <= x[772] | x[774];
     layer0_out[9620] <= x[1934] & x[1935];
     layer0_out[9621] <= x[7573];
     layer0_out[9622] <= ~(x[6876] ^ x[6877]);
     layer0_out[9623] <= ~(x[1130] ^ x[1131]);
     layer0_out[9624] <= ~(x[2654] ^ x[2656]);
     layer0_out[9625] <= ~x[7621] | x[7620];
     layer0_out[9626] <= ~(x[9202] & x[9203]);
     layer0_out[9627] <= x[3769] | x[3770];
     layer0_out[9628] <= ~(x[7280] | x[7281]);
     layer0_out[9629] <= x[1161];
     layer0_out[9630] <= ~(x[5395] & x[5396]);
     layer0_out[9631] <= ~(x[8363] ^ x[8364]);
     layer0_out[9632] <= ~x[8299];
     layer0_out[9633] <= ~x[1469] | x[1471];
     layer0_out[9634] <= ~(x[1865] & x[1867]);
     layer0_out[9635] <= ~(x[3301] ^ x[3302]);
     layer0_out[9636] <= ~(x[694] & x[695]);
     layer0_out[9637] <= x[2390];
     layer0_out[9638] <= ~(x[868] & x[870]);
     layer0_out[9639] <= ~(x[3091] | x[3092]);
     layer0_out[9640] <= x[4708] & x[4709];
     layer0_out[9641] <= ~(x[2586] & x[2587]);
     layer0_out[9642] <= x[3540] & x[3541];
     layer0_out[9643] <= ~(x[5676] | x[5677]);
     layer0_out[9644] <= 1'b0;
     layer0_out[9645] <= ~x[9150];
     layer0_out[9646] <= ~x[380];
     layer0_out[9647] <= ~x[1142];
     layer0_out[9648] <= x[2430] & ~x[2428];
     layer0_out[9649] <= x[3417] & x[3418];
     layer0_out[9650] <= ~x[680];
     layer0_out[9651] <= x[1706] & x[1708];
     layer0_out[9652] <= x[8345];
     layer0_out[9653] <= ~(x[2751] & x[2753]);
     layer0_out[9654] <= x[493];
     layer0_out[9655] <= ~(x[6881] & x[6882]);
     layer0_out[9656] <= ~(x[4403] & x[4404]);
     layer0_out[9657] <= ~x[3150];
     layer0_out[9658] <= 1'b1;
     layer0_out[9659] <= ~(x[7110] ^ x[7111]);
     layer0_out[9660] <= x[2315] ^ x[2317];
     layer0_out[9661] <= x[1707] | x[1709];
     layer0_out[9662] <= 1'b0;
     layer0_out[9663] <= x[7586] & x[7587];
     layer0_out[9664] <= x[1534] | x[1535];
     layer0_out[9665] <= ~(x[1170] & x[1172]);
     layer0_out[9666] <= ~x[4984];
     layer0_out[9667] <= ~x[3578];
     layer0_out[9668] <= x[8798] | x[8799];
     layer0_out[9669] <= ~x[4607];
     layer0_out[9670] <= x[8992] | x[8993];
     layer0_out[9671] <= ~x[3467];
     layer0_out[9672] <= ~(x[525] & x[526]);
     layer0_out[9673] <= x[1266] & x[1268];
     layer0_out[9674] <= x[4103] & x[4104];
     layer0_out[9675] <= ~(x[2178] & x[2180]);
     layer0_out[9676] <= ~(x[8738] ^ x[8739]);
     layer0_out[9677] <= ~(x[1901] & x[1903]);
     layer0_out[9678] <= x[2399];
     layer0_out[9679] <= x[668] & x[669];
     layer0_out[9680] <= x[3010];
     layer0_out[9681] <= x[1015] & x[1017];
     layer0_out[9682] <= x[7959] | x[7960];
     layer0_out[9683] <= ~(x[5788] ^ x[5789]);
     layer0_out[9684] <= x[6678] | x[6679];
     layer0_out[9685] <= ~(x[5654] & x[5655]);
     layer0_out[9686] <= x[1694];
     layer0_out[9687] <= x[6601];
     layer0_out[9688] <= ~(x[7439] | x[7440]);
     layer0_out[9689] <= ~(x[6990] & x[6991]);
     layer0_out[9690] <= ~(x[8475] | x[8476]);
     layer0_out[9691] <= ~(x[4846] | x[4847]);
     layer0_out[9692] <= ~(x[625] & x[627]);
     layer0_out[9693] <= 1'b0;
     layer0_out[9694] <= ~(x[7232] | x[7233]);
     layer0_out[9695] <= x[2247] & x[2248];
     layer0_out[9696] <= ~(x[7134] & x[7135]);
     layer0_out[9697] <= x[3775];
     layer0_out[9698] <= x[5577];
     layer0_out[9699] <= x[1612] & x[1613];
     layer0_out[9700] <= x[558] & x[559];
     layer0_out[9701] <= ~x[7582] | x[7583];
     layer0_out[9702] <= x[8613];
     layer0_out[9703] <= x[6595] & ~x[6596];
     layer0_out[9704] <= x[6882];
     layer0_out[9705] <= ~(x[7607] & x[7608]);
     layer0_out[9706] <= ~x[2176];
     layer0_out[9707] <= ~(x[2362] & x[2363]);
     layer0_out[9708] <= ~(x[8497] | x[8498]);
     layer0_out[9709] <= x[920] & x[921];
     layer0_out[9710] <= ~x[6033];
     layer0_out[9711] <= 1'b0;
     layer0_out[9712] <= x[2367] | x[2369];
     layer0_out[9713] <= x[2250] | x[2251];
     layer0_out[9714] <= x[2250] | x[2252];
     layer0_out[9715] <= ~x[1718];
     layer0_out[9716] <= x[570];
     layer0_out[9717] <= ~(x[7970] | x[7971]);
     layer0_out[9718] <= ~(x[1702] | x[1704]);
     layer0_out[9719] <= x[4215];
     layer0_out[9720] <= x[1163];
     layer0_out[9721] <= x[1689] & x[1691];
     layer0_out[9722] <= ~x[1356];
     layer0_out[9723] <= ~(x[332] & x[334]);
     layer0_out[9724] <= x[5570] & x[5571];
     layer0_out[9725] <= ~(x[1418] & x[1420]);
     layer0_out[9726] <= ~(x[6857] ^ x[6858]);
     layer0_out[9727] <= ~(x[3214] ^ x[3215]);
     layer0_out[9728] <= x[6993] | x[6994];
     layer0_out[9729] <= x[6211];
     layer0_out[9730] <= x[2290] & ~x[2291];
     layer0_out[9731] <= x[1904] & x[1905];
     layer0_out[9732] <= x[994] & x[995];
     layer0_out[9733] <= ~(x[5655] & x[5656]);
     layer0_out[9734] <= ~(x[1055] & x[1056]);
     layer0_out[9735] <= ~(x[3771] | x[3772]);
     layer0_out[9736] <= ~(x[4424] & x[4425]);
     layer0_out[9737] <= x[417];
     layer0_out[9738] <= x[4015] & x[4016];
     layer0_out[9739] <= ~(x[2579] & x[2580]);
     layer0_out[9740] <= x[8302] & x[8303];
     layer0_out[9741] <= ~(x[2095] & x[2097]);
     layer0_out[9742] <= ~(x[916] | x[917]);
     layer0_out[9743] <= x[6384] | x[6385];
     layer0_out[9744] <= ~(x[4349] | x[4350]);
     layer0_out[9745] <= ~(x[7296] | x[7297]);
     layer0_out[9746] <= x[5217] & x[5218];
     layer0_out[9747] <= ~(x[1711] & x[1713]);
     layer0_out[9748] <= x[1582] & x[1584];
     layer0_out[9749] <= ~x[7056];
     layer0_out[9750] <= ~(x[4463] & x[4464]);
     layer0_out[9751] <= ~x[1073];
     layer0_out[9752] <= 1'b0;
     layer0_out[9753] <= x[2135] & x[2137];
     layer0_out[9754] <= ~x[865];
     layer0_out[9755] <= ~x[1289];
     layer0_out[9756] <= x[4837] & x[4838];
     layer0_out[9757] <= 1'b1;
     layer0_out[9758] <= ~x[7695];
     layer0_out[9759] <= ~(x[1733] & x[1735]);
     layer0_out[9760] <= x[4609];
     layer0_out[9761] <= ~(x[343] & x[345]);
     layer0_out[9762] <= x[2591] & x[2593];
     layer0_out[9763] <= ~(x[311] | x[312]);
     layer0_out[9764] <= x[558] & x[560];
     layer0_out[9765] <= ~x[2491] | x[2493];
     layer0_out[9766] <= ~(x[2027] ^ x[2028]);
     layer0_out[9767] <= ~(x[1076] & x[1078]);
     layer0_out[9768] <= ~(x[330] | x[332]);
     layer0_out[9769] <= ~(x[9065] & x[9066]);
     layer0_out[9770] <= x[562] & x[563];
     layer0_out[9771] <= ~(x[769] ^ x[770]);
     layer0_out[9772] <= x[5794] & x[5795];
     layer0_out[9773] <= ~(x[2101] & x[2102]);
     layer0_out[9774] <= x[4568] | x[4569];
     layer0_out[9775] <= ~(x[311] & x[313]);
     layer0_out[9776] <= ~x[4941] | x[4942];
     layer0_out[9777] <= x[2504] & x[2506];
     layer0_out[9778] <= 1'b1;
     layer0_out[9779] <= x[7041] | x[7042];
     layer0_out[9780] <= x[5626] & x[5627];
     layer0_out[9781] <= x[251] | x[253];
     layer0_out[9782] <= ~x[7599];
     layer0_out[9783] <= x[2940] ^ x[2941];
     layer0_out[9784] <= x[6765] & x[6766];
     layer0_out[9785] <= 1'b1;
     layer0_out[9786] <= ~x[1985];
     layer0_out[9787] <= ~(x[8695] | x[8696]);
     layer0_out[9788] <= 1'b0;
     layer0_out[9789] <= x[8341];
     layer0_out[9790] <= ~x[2048];
     layer0_out[9791] <= x[3645] | x[3646];
     layer0_out[9792] <= ~(x[2667] | x[2668]);
     layer0_out[9793] <= 1'b0;
     layer0_out[9794] <= ~(x[669] | x[670]);
     layer0_out[9795] <= ~x[2133];
     layer0_out[9796] <= ~(x[4794] & x[4795]);
     layer0_out[9797] <= x[1812] | x[1813];
     layer0_out[9798] <= ~x[374];
     layer0_out[9799] <= x[1116] & ~x[1114];
     layer0_out[9800] <= x[2722] ^ x[2723];
     layer0_out[9801] <= x[1751] & x[1753];
     layer0_out[9802] <= ~x[5210];
     layer0_out[9803] <= x[167] | x[169];
     layer0_out[9804] <= ~x[6912] | x[6913];
     layer0_out[9805] <= x[2835] & x[2836];
     layer0_out[9806] <= x[8391] ^ x[8392];
     layer0_out[9807] <= ~x[6603];
     layer0_out[9808] <= ~(x[3793] | x[3794]);
     layer0_out[9809] <= x[648] | x[650];
     layer0_out[9810] <= ~(x[8319] | x[8320]);
     layer0_out[9811] <= ~(x[2771] ^ x[2772]);
     layer0_out[9812] <= ~(x[2675] & x[2677]);
     layer0_out[9813] <= x[6859];
     layer0_out[9814] <= ~(x[6894] | x[6895]);
     layer0_out[9815] <= ~(x[3892] | x[3893]);
     layer0_out[9816] <= ~(x[2388] & x[2389]);
     layer0_out[9817] <= x[5388];
     layer0_out[9818] <= x[7266] & ~x[7267];
     layer0_out[9819] <= ~x[7791];
     layer0_out[9820] <= ~(x[6041] & x[6042]);
     layer0_out[9821] <= 1'b1;
     layer0_out[9822] <= ~x[1777];
     layer0_out[9823] <= x[5394] ^ x[5395];
     layer0_out[9824] <= x[780] & x[782];
     layer0_out[9825] <= ~x[968];
     layer0_out[9826] <= x[1668] ^ x[1669];
     layer0_out[9827] <= x[6173] | x[6174];
     layer0_out[9828] <= ~x[1683] | x[1684];
     layer0_out[9829] <= x[5180] & x[5181];
     layer0_out[9830] <= 1'b0;
     layer0_out[9831] <= x[1586] & x[1587];
     layer0_out[9832] <= 1'b1;
     layer0_out[9833] <= ~x[1643];
     layer0_out[9834] <= ~(x[7001] | x[7002]);
     layer0_out[9835] <= ~(x[34] | x[35]);
     layer0_out[9836] <= ~(x[3357] | x[3358]);
     layer0_out[9837] <= x[2352] & ~x[2350];
     layer0_out[9838] <= ~x[8900];
     layer0_out[9839] <= x[2727] & x[2729];
     layer0_out[9840] <= x[299];
     layer0_out[9841] <= 1'b1;
     layer0_out[9842] <= x[5815] & ~x[5816];
     layer0_out[9843] <= ~x[8343];
     layer0_out[9844] <= x[1275] & x[1277];
     layer0_out[9845] <= x[5988] | x[5989];
     layer0_out[9846] <= ~(x[2814] | x[2815]);
     layer0_out[9847] <= ~x[8365];
     layer0_out[9848] <= x[138] ^ x[139];
     layer0_out[9849] <= ~(x[5684] | x[5685]);
     layer0_out[9850] <= ~x[1920];
     layer0_out[9851] <= ~(x[1074] ^ x[1076]);
     layer0_out[9852] <= ~(x[4047] | x[4048]);
     layer0_out[9853] <= x[40] | x[42];
     layer0_out[9854] <= ~(x[7210] & x[7211]);
     layer0_out[9855] <= ~(x[2712] & x[2714]);
     layer0_out[9856] <= ~(x[1122] ^ x[1124]);
     layer0_out[9857] <= x[890];
     layer0_out[9858] <= x[5656] ^ x[5657];
     layer0_out[9859] <= x[2156] & x[2157];
     layer0_out[9860] <= x[3609] | x[3610];
     layer0_out[9861] <= ~(x[1603] & x[1604]);
     layer0_out[9862] <= ~(x[6138] & x[6139]);
     layer0_out[9863] <= ~(x[6320] | x[6321]);
     layer0_out[9864] <= x[6100] & x[6101];
     layer0_out[9865] <= ~(x[2578] & x[2579]);
     layer0_out[9866] <= ~(x[55] & x[56]);
     layer0_out[9867] <= ~x[8600] | x[8601];
     layer0_out[9868] <= ~x[4127];
     layer0_out[9869] <= ~(x[8671] | x[8672]);
     layer0_out[9870] <= x[6038];
     layer0_out[9871] <= x[2172] | x[2174];
     layer0_out[9872] <= x[1062];
     layer0_out[9873] <= ~x[4101];
     layer0_out[9874] <= x[165] & x[167];
     layer0_out[9875] <= ~(x[4507] & x[4508]);
     layer0_out[9876] <= ~x[4720];
     layer0_out[9877] <= ~x[6840] | x[6839];
     layer0_out[9878] <= ~(x[783] & x[784]);
     layer0_out[9879] <= 1'b0;
     layer0_out[9880] <= x[5713];
     layer0_out[9881] <= ~x[1889] | x[1890];
     layer0_out[9882] <= ~x[3445] | x[3444];
     layer0_out[9883] <= ~x[2119];
     layer0_out[9884] <= ~(x[496] & x[497]);
     layer0_out[9885] <= x[3184] | x[3185];
     layer0_out[9886] <= ~x[7304];
     layer0_out[9887] <= x[4896] | x[4897];
     layer0_out[9888] <= x[4840];
     layer0_out[9889] <= ~(x[2974] & x[2975]);
     layer0_out[9890] <= ~(x[4049] ^ x[4050]);
     layer0_out[9891] <= x[2340] ^ x[2342];
     layer0_out[9892] <= x[3161] ^ x[3162];
     layer0_out[9893] <= 1'b1;
     layer0_out[9894] <= x[8765];
     layer0_out[9895] <= ~(x[5407] & x[5408]);
     layer0_out[9896] <= 1'b0;
     layer0_out[9897] <= x[1606] & x[1607];
     layer0_out[9898] <= x[8656] | x[8657];
     layer0_out[9899] <= ~(x[1143] | x[1145]);
     layer0_out[9900] <= ~(x[2495] ^ x[2496]);
     layer0_out[9901] <= x[65] & ~x[63];
     layer0_out[9902] <= x[2066] & x[2068];
     layer0_out[9903] <= ~(x[2463] & x[2465]);
     layer0_out[9904] <= x[8617] & ~x[8616];
     layer0_out[9905] <= ~(x[3267] | x[3268]);
     layer0_out[9906] <= x[45] & x[47];
     layer0_out[9907] <= x[3936] & ~x[3937];
     layer0_out[9908] <= ~x[7047];
     layer0_out[9909] <= 1'b1;
     layer0_out[9910] <= ~(x[1740] & x[1742]);
     layer0_out[9911] <= ~(x[2884] | x[2885]);
     layer0_out[9912] <= x[2032];
     layer0_out[9913] <= ~(x[260] ^ x[262]);
     layer0_out[9914] <= x[5694] & x[5695];
     layer0_out[9915] <= x[526] & ~x[524];
     layer0_out[9916] <= ~x[7413] | x[7414];
     layer0_out[9917] <= ~(x[1231] & x[1232]);
     layer0_out[9918] <= ~x[6907];
     layer0_out[9919] <= x[264];
     layer0_out[9920] <= x[488];
     layer0_out[9921] <= ~(x[5328] & x[5329]);
     layer0_out[9922] <= ~(x[1729] & x[1730]);
     layer0_out[9923] <= ~(x[3513] | x[3514]);
     layer0_out[9924] <= ~(x[2111] & x[2112]);
     layer0_out[9925] <= x[585] & x[586];
     layer0_out[9926] <= ~x[8826];
     layer0_out[9927] <= ~(x[8859] | x[8860]);
     layer0_out[9928] <= 1'b1;
     layer0_out[9929] <= ~(x[6207] | x[6208]);
     layer0_out[9930] <= ~(x[1371] & x[1373]);
     layer0_out[9931] <= x[966] & x[968];
     layer0_out[9932] <= x[2264];
     layer0_out[9933] <= ~(x[4097] & x[4098]);
     layer0_out[9934] <= ~(x[8275] & x[8276]);
     layer0_out[9935] <= x[950] & x[951];
     layer0_out[9936] <= ~x[8609];
     layer0_out[9937] <= ~x[519];
     layer0_out[9938] <= x[1783] & x[1784];
     layer0_out[9939] <= x[9170] & x[9171];
     layer0_out[9940] <= ~(x[5321] | x[5322]);
     layer0_out[9941] <= 1'b1;
     layer0_out[9942] <= ~(x[5269] & x[5270]);
     layer0_out[9943] <= ~(x[1799] & x[1801]);
     layer0_out[9944] <= ~(x[1739] & x[1741]);
     layer0_out[9945] <= ~(x[672] ^ x[674]);
     layer0_out[9946] <= x[7636] & x[7637];
     layer0_out[9947] <= x[4181] ^ x[4182];
     layer0_out[9948] <= ~(x[3125] | x[3126]);
     layer0_out[9949] <= 1'b1;
     layer0_out[9950] <= 1'b0;
     layer0_out[9951] <= 1'b1;
     layer0_out[9952] <= ~(x[7370] ^ x[7371]);
     layer0_out[9953] <= x[1834] & ~x[1832];
     layer0_out[9954] <= x[1955];
     layer0_out[9955] <= ~x[8300];
     layer0_out[9956] <= x[2595] & x[2597];
     layer0_out[9957] <= x[7363] | x[7364];
     layer0_out[9958] <= ~(x[5028] | x[5029]);
     layer0_out[9959] <= 1'b0;
     layer0_out[9960] <= ~(x[2665] ^ x[2667]);
     layer0_out[9961] <= x[1064] & x[1065];
     layer0_out[9962] <= ~(x[5421] & x[5422]);
     layer0_out[9963] <= x[7941] & ~x[7940];
     layer0_out[9964] <= ~(x[365] & x[367]);
     layer0_out[9965] <= ~(x[101] & x[103]);
     layer0_out[9966] <= ~(x[612] & x[614]);
     layer0_out[9967] <= x[3132] & x[3133];
     layer0_out[9968] <= ~(x[3024] & x[3025]);
     layer0_out[9969] <= x[900] & x[902];
     layer0_out[9970] <= x[1541] & x[1543];
     layer0_out[9971] <= ~(x[8444] ^ x[8445]);
     layer0_out[9972] <= x[4940] ^ x[4941];
     layer0_out[9973] <= x[2190] & x[2191];
     layer0_out[9974] <= x[2946] & x[2947];
     layer0_out[9975] <= x[1971] & x[1972];
     layer0_out[9976] <= ~(x[5254] & x[5255]);
     layer0_out[9977] <= x[6075] & x[6076];
     layer0_out[9978] <= 1'b0;
     layer0_out[9979] <= x[7499];
     layer0_out[9980] <= 1'b1;
     layer0_out[9981] <= ~(x[6233] | x[6234]);
     layer0_out[9982] <= ~(x[2622] | x[2624]);
     layer0_out[9983] <= ~(x[3881] | x[3882]);
     layer0_out[9984] <= x[1503] ^ x[1505];
     layer0_out[9985] <= x[1772] & x[1774];
     layer0_out[9986] <= ~x[909];
     layer0_out[9987] <= x[1198] & x[1199];
     layer0_out[9988] <= ~x[7802];
     layer0_out[9989] <= 1'b0;
     layer0_out[9990] <= x[2141] ^ x[2142];
     layer0_out[9991] <= ~x[6474] | x[6475];
     layer0_out[9992] <= x[6059] ^ x[6060];
     layer0_out[9993] <= ~(x[271] & x[272]);
     layer0_out[9994] <= ~x[6673];
     layer0_out[9995] <= x[1837] | x[1838];
     layer0_out[9996] <= x[375];
     layer0_out[9997] <= ~(x[598] & x[600]);
     layer0_out[9998] <= ~x[357];
     layer0_out[9999] <= x[2257] & x[2259];
     layer0_out[10000] <= ~(x[5905] & x[5906]);
     layer0_out[10001] <= ~(x[292] & x[294]);
     layer0_out[10002] <= x[7444] | x[7445];
     layer0_out[10003] <= 1'b0;
     layer0_out[10004] <= x[746] & x[748];
     layer0_out[10005] <= ~(x[708] & x[709]);
     layer0_out[10006] <= x[1197] & x[1198];
     layer0_out[10007] <= x[822] | x[824];
     layer0_out[10008] <= ~(x[7342] ^ x[7343]);
     layer0_out[10009] <= ~(x[8035] | x[8036]);
     layer0_out[10010] <= x[1309];
     layer0_out[10011] <= ~(x[5797] | x[5798]);
     layer0_out[10012] <= ~(x[5918] & x[5919]);
     layer0_out[10013] <= ~(x[5843] ^ x[5844]);
     layer0_out[10014] <= x[1655] & x[1656];
     layer0_out[10015] <= ~(x[3303] ^ x[3304]);
     layer0_out[10016] <= x[561] ^ x[563];
     layer0_out[10017] <= ~(x[5270] & x[5271]);
     layer0_out[10018] <= ~x[8858];
     layer0_out[10019] <= ~(x[6411] | x[6412]);
     layer0_out[10020] <= ~(x[2089] & x[2091]);
     layer0_out[10021] <= ~(x[364] & x[366]);
     layer0_out[10022] <= x[3673] & x[3674];
     layer0_out[10023] <= ~(x[8884] | x[8885]);
     layer0_out[10024] <= x[2777] & x[2778];
     layer0_out[10025] <= x[2982];
     layer0_out[10026] <= x[1624] & x[1625];
     layer0_out[10027] <= x[2396] | x[2397];
     layer0_out[10028] <= x[5398] & x[5399];
     layer0_out[10029] <= x[8741];
     layer0_out[10030] <= ~(x[2332] | x[2333]);
     layer0_out[10031] <= ~(x[3493] | x[3494]);
     layer0_out[10032] <= x[1185];
     layer0_out[10033] <= x[7547];
     layer0_out[10034] <= ~(x[5465] | x[5466]);
     layer0_out[10035] <= x[5010] | x[5011];
     layer0_out[10036] <= ~x[1171] | x[1169];
     layer0_out[10037] <= x[2064];
     layer0_out[10038] <= ~x[7524];
     layer0_out[10039] <= ~x[4542];
     layer0_out[10040] <= 1'b1;
     layer0_out[10041] <= x[1548];
     layer0_out[10042] <= ~x[8064];
     layer0_out[10043] <= x[2860] & x[2861];
     layer0_out[10044] <= ~x[609];
     layer0_out[10045] <= x[3566] | x[3567];
     layer0_out[10046] <= x[1681] | x[1683];
     layer0_out[10047] <= x[3311] & ~x[3310];
     layer0_out[10048] <= ~(x[402] & x[404]);
     layer0_out[10049] <= 1'b0;
     layer0_out[10050] <= x[95] | x[97];
     layer0_out[10051] <= ~(x[714] | x[715]);
     layer0_out[10052] <= ~(x[8135] ^ x[8136]);
     layer0_out[10053] <= 1'b0;
     layer0_out[10054] <= ~(x[4704] ^ x[4705]);
     layer0_out[10055] <= ~x[6551] | x[6552];
     layer0_out[10056] <= x[6403] | x[6404];
     layer0_out[10057] <= x[7090];
     layer0_out[10058] <= ~(x[2747] ^ x[2748]);
     layer0_out[10059] <= ~(x[1141] & x[1142]);
     layer0_out[10060] <= ~(x[777] & x[779]);
     layer0_out[10061] <= ~x[6910] | x[6911];
     layer0_out[10062] <= x[8759] | x[8760];
     layer0_out[10063] <= ~(x[7216] | x[7217]);
     layer0_out[10064] <= x[2803] & ~x[2802];
     layer0_out[10065] <= x[241] ^ x[243];
     layer0_out[10066] <= ~(x[7672] & x[7673]);
     layer0_out[10067] <= ~(x[895] & x[897]);
     layer0_out[10068] <= x[3736] & x[3737];
     layer0_out[10069] <= x[5549];
     layer0_out[10070] <= x[5488] & x[5489];
     layer0_out[10071] <= x[3276] ^ x[3277];
     layer0_out[10072] <= ~x[6598];
     layer0_out[10073] <= x[1192] ^ x[1193];
     layer0_out[10074] <= ~(x[1937] & x[1938]);
     layer0_out[10075] <= ~(x[3619] & x[3620]);
     layer0_out[10076] <= ~(x[6654] | x[6655]);
     layer0_out[10077] <= ~(x[8575] ^ x[8576]);
     layer0_out[10078] <= ~(x[7815] | x[7816]);
     layer0_out[10079] <= ~(x[608] ^ x[610]);
     layer0_out[10080] <= ~(x[927] & x[929]);
     layer0_out[10081] <= ~(x[397] & x[399]);
     layer0_out[10082] <= ~(x[6099] & x[6100]);
     layer0_out[10083] <= x[9194] & ~x[9195];
     layer0_out[10084] <= ~(x[7372] | x[7373]);
     layer0_out[10085] <= ~x[6328];
     layer0_out[10086] <= x[7291] & x[7292];
     layer0_out[10087] <= ~x[175] | x[177];
     layer0_out[10088] <= x[2469] ^ x[2470];
     layer0_out[10089] <= ~(x[6467] | x[6468]);
     layer0_out[10090] <= x[5882] & x[5883];
     layer0_out[10091] <= 1'b0;
     layer0_out[10092] <= ~x[6206] | x[6205];
     layer0_out[10093] <= ~x[5450];
     layer0_out[10094] <= x[3220] ^ x[3221];
     layer0_out[10095] <= 1'b0;
     layer0_out[10096] <= ~(x[5746] & x[5747]);
     layer0_out[10097] <= x[2453] & ~x[2455];
     layer0_out[10098] <= x[1402] & x[1404];
     layer0_out[10099] <= ~(x[4275] | x[4276]);
     layer0_out[10100] <= 1'b1;
     layer0_out[10101] <= x[5281] & x[5282];
     layer0_out[10102] <= ~(x[7012] ^ x[7013]);
     layer0_out[10103] <= ~(x[2687] ^ x[2688]);
     layer0_out[10104] <= ~(x[2418] | x[2419]);
     layer0_out[10105] <= ~(x[7005] | x[7006]);
     layer0_out[10106] <= ~x[7500];
     layer0_out[10107] <= ~(x[3397] | x[3398]);
     layer0_out[10108] <= ~(x[3602] | x[3603]);
     layer0_out[10109] <= x[7748] & ~x[7749];
     layer0_out[10110] <= ~x[5342];
     layer0_out[10111] <= ~(x[6605] | x[6606]);
     layer0_out[10112] <= x[7150] | x[7151];
     layer0_out[10113] <= ~(x[6297] | x[6298]);
     layer0_out[10114] <= x[7226];
     layer0_out[10115] <= ~x[8871];
     layer0_out[10116] <= ~(x[8227] | x[8228]);
     layer0_out[10117] <= ~(x[1232] & x[1233]);
     layer0_out[10118] <= x[1919] & x[1921];
     layer0_out[10119] <= x[6311] | x[6312];
     layer0_out[10120] <= x[8372];
     layer0_out[10121] <= x[6956] ^ x[6957];
     layer0_out[10122] <= x[6395];
     layer0_out[10123] <= x[4169];
     layer0_out[10124] <= x[1919];
     layer0_out[10125] <= x[358] | x[359];
     layer0_out[10126] <= ~x[8351];
     layer0_out[10127] <= x[3929] | x[3930];
     layer0_out[10128] <= ~x[137] | x[139];
     layer0_out[10129] <= x[2983] & x[2984];
     layer0_out[10130] <= ~(x[1152] & x[1153]);
     layer0_out[10131] <= x[1735] & x[1736];
     layer0_out[10132] <= x[1439] & x[1440];
     layer0_out[10133] <= ~(x[9171] & x[9172]);
     layer0_out[10134] <= 1'b0;
     layer0_out[10135] <= ~x[6801];
     layer0_out[10136] <= ~(x[442] ^ x[444]);
     layer0_out[10137] <= ~(x[6544] | x[6545]);
     layer0_out[10138] <= x[1637] ^ x[1639];
     layer0_out[10139] <= ~x[7151];
     layer0_out[10140] <= x[2354] & x[2355];
     layer0_out[10141] <= x[1333] & x[1334];
     layer0_out[10142] <= x[2551] & ~x[2550];
     layer0_out[10143] <= ~(x[817] | x[818]);
     layer0_out[10144] <= 1'b0;
     layer0_out[10145] <= ~(x[6639] | x[6640]);
     layer0_out[10146] <= x[5562] | x[5563];
     layer0_out[10147] <= x[461] & ~x[462];
     layer0_out[10148] <= x[5512] | x[5513];
     layer0_out[10149] <= x[2903] ^ x[2904];
     layer0_out[10150] <= x[6778] & ~x[6777];
     layer0_out[10151] <= ~x[3088];
     layer0_out[10152] <= x[3966] | x[3967];
     layer0_out[10153] <= x[2016] ^ x[2017];
     layer0_out[10154] <= ~(x[6583] | x[6584]);
     layer0_out[10155] <= x[682] & x[684];
     layer0_out[10156] <= ~(x[1027] & x[1029]);
     layer0_out[10157] <= ~(x[1508] ^ x[1510]);
     layer0_out[10158] <= x[4222] & x[4223];
     layer0_out[10159] <= x[1156] & x[1158];
     layer0_out[10160] <= x[3379] & ~x[3380];
     layer0_out[10161] <= x[8621] | x[8622];
     layer0_out[10162] <= ~(x[6046] & x[6047]);
     layer0_out[10163] <= ~(x[6184] ^ x[6185]);
     layer0_out[10164] <= x[2238];
     layer0_out[10165] <= x[1537] & x[1538];
     layer0_out[10166] <= ~(x[2146] | x[2148]);
     layer0_out[10167] <= ~x[2475];
     layer0_out[10168] <= x[934] | x[935];
     layer0_out[10169] <= x[8061] & x[8062];
     layer0_out[10170] <= ~x[1970];
     layer0_out[10171] <= ~(x[2768] ^ x[2770]);
     layer0_out[10172] <= ~(x[1498] ^ x[1500]);
     layer0_out[10173] <= x[8279] & ~x[8280];
     layer0_out[10174] <= x[6924] ^ x[6925];
     layer0_out[10175] <= ~(x[555] ^ x[556]);
     layer0_out[10176] <= x[5497] & x[5498];
     layer0_out[10177] <= ~(x[1709] ^ x[1710]);
     layer0_out[10178] <= ~x[45] | x[44];
     layer0_out[10179] <= 1'b0;
     layer0_out[10180] <= ~(x[1997] | x[1998]);
     layer0_out[10181] <= x[406] ^ x[407];
     layer0_out[10182] <= ~(x[6960] ^ x[6961]);
     layer0_out[10183] <= ~(x[2329] ^ x[2331]);
     layer0_out[10184] <= ~(x[5866] & x[5867]);
     layer0_out[10185] <= x[7875] & ~x[7874];
     layer0_out[10186] <= ~(x[463] & x[464]);
     layer0_out[10187] <= ~x[7333];
     layer0_out[10188] <= ~x[3114] | x[3113];
     layer0_out[10189] <= ~(x[6223] & x[6224]);
     layer0_out[10190] <= x[3549] | x[3550];
     layer0_out[10191] <= ~x[6782] | x[6781];
     layer0_out[10192] <= ~x[1883] | x[1882];
     layer0_out[10193] <= ~(x[3117] | x[3118]);
     layer0_out[10194] <= ~x[1417] | x[1416];
     layer0_out[10195] <= x[3873] ^ x[3874];
     layer0_out[10196] <= x[1592] & x[1594];
     layer0_out[10197] <= x[8994];
     layer0_out[10198] <= ~(x[3073] | x[3074]);
     layer0_out[10199] <= ~(x[2529] ^ x[2531]);
     layer0_out[10200] <= x[6578] & x[6579];
     layer0_out[10201] <= x[774] | x[776];
     layer0_out[10202] <= ~(x[6760] | x[6761]);
     layer0_out[10203] <= 1'b1;
     layer0_out[10204] <= ~x[1981] | x[1983];
     layer0_out[10205] <= ~x[3782];
     layer0_out[10206] <= ~(x[8655] & x[8656]);
     layer0_out[10207] <= ~x[2230] | x[2229];
     layer0_out[10208] <= ~(x[1276] ^ x[1278]);
     layer0_out[10209] <= x[625] ^ x[626];
     layer0_out[10210] <= ~x[1024];
     layer0_out[10211] <= ~(x[4585] ^ x[4586]);
     layer0_out[10212] <= x[2597] ^ x[2599];
     layer0_out[10213] <= ~(x[1740] & x[1741]);
     layer0_out[10214] <= ~x[2255] | x[2256];
     layer0_out[10215] <= ~x[4908];
     layer0_out[10216] <= 1'b0;
     layer0_out[10217] <= x[6798] & x[6799];
     layer0_out[10218] <= ~(x[992] | x[994]);
     layer0_out[10219] <= ~(x[8272] & x[8273]);
     layer0_out[10220] <= ~(x[247] | x[249]);
     layer0_out[10221] <= ~(x[8825] ^ x[8826]);
     layer0_out[10222] <= x[3251] & x[3252];
     layer0_out[10223] <= x[3867] | x[3868];
     layer0_out[10224] <= x[9084];
     layer0_out[10225] <= x[634] | x[636];
     layer0_out[10226] <= x[3100] ^ x[3101];
     layer0_out[10227] <= ~(x[5179] | x[5180]);
     layer0_out[10228] <= ~x[8594] | x[8595];
     layer0_out[10229] <= 1'b1;
     layer0_out[10230] <= ~(x[6657] ^ x[6658]);
     layer0_out[10231] <= x[4558] & x[4559];
     layer0_out[10232] <= x[3902];
     layer0_out[10233] <= x[1774] | x[1775];
     layer0_out[10234] <= x[2640] & x[2642];
     layer0_out[10235] <= ~(x[8321] & x[8322]);
     layer0_out[10236] <= x[4845] & ~x[4844];
     layer0_out[10237] <= ~(x[8161] | x[8162]);
     layer0_out[10238] <= x[1823] | x[1825];
     layer0_out[10239] <= ~x[2697] | x[2699];
     layer0_out[10240] <= 1'b1;
     layer0_out[10241] <= x[4230];
     layer0_out[10242] <= x[2402] & ~x[2400];
     layer0_out[10243] <= ~(x[5567] | x[5568]);
     layer0_out[10244] <= ~(x[2180] & x[2181]);
     layer0_out[10245] <= x[1502] ^ x[1503];
     layer0_out[10246] <= x[1561] ^ x[1562];
     layer0_out[10247] <= x[2535] ^ x[2536];
     layer0_out[10248] <= ~(x[5631] ^ x[5632]);
     layer0_out[10249] <= ~x[1715];
     layer0_out[10250] <= x[1575] ^ x[1576];
     layer0_out[10251] <= ~(x[5466] | x[5467]);
     layer0_out[10252] <= 1'b1;
     layer0_out[10253] <= x[462];
     layer0_out[10254] <= x[7696] & x[7697];
     layer0_out[10255] <= ~x[4233];
     layer0_out[10256] <= 1'b0;
     layer0_out[10257] <= x[8070] & ~x[8069];
     layer0_out[10258] <= ~(x[2780] ^ x[2781]);
     layer0_out[10259] <= ~(x[8990] & x[8991]);
     layer0_out[10260] <= x[2442] & x[2443];
     layer0_out[10261] <= ~(x[4058] | x[4059]);
     layer0_out[10262] <= x[2205] & x[2207];
     layer0_out[10263] <= x[61] & x[63];
     layer0_out[10264] <= x[3946] | x[3947];
     layer0_out[10265] <= x[2313] & ~x[2315];
     layer0_out[10266] <= ~(x[5040] & x[5041]);
     layer0_out[10267] <= ~(x[763] ^ x[764]);
     layer0_out[10268] <= ~x[6376];
     layer0_out[10269] <= ~x[3579];
     layer0_out[10270] <= ~(x[1240] & x[1242]);
     layer0_out[10271] <= ~(x[5310] & x[5311]);
     layer0_out[10272] <= ~x[2167];
     layer0_out[10273] <= x[8588] | x[8589];
     layer0_out[10274] <= ~(x[6556] & x[6557]);
     layer0_out[10275] <= 1'b1;
     layer0_out[10276] <= ~x[8239];
     layer0_out[10277] <= x[6663];
     layer0_out[10278] <= x[7725];
     layer0_out[10279] <= x[3304];
     layer0_out[10280] <= ~(x[1609] ^ x[1610]);
     layer0_out[10281] <= ~(x[4848] | x[4849]);
     layer0_out[10282] <= x[1877] & x[1879];
     layer0_out[10283] <= x[2575] | x[2576];
     layer0_out[10284] <= x[6515] | x[6516];
     layer0_out[10285] <= ~x[3223] | x[3224];
     layer0_out[10286] <= ~x[1855];
     layer0_out[10287] <= ~x[7777];
     layer0_out[10288] <= ~x[8071];
     layer0_out[10289] <= ~(x[3775] & x[3776]);
     layer0_out[10290] <= 1'b1;
     layer0_out[10291] <= ~(x[7369] & x[7370]);
     layer0_out[10292] <= x[3779] | x[3780];
     layer0_out[10293] <= ~(x[5101] | x[5102]);
     layer0_out[10294] <= x[1601] & x[1602];
     layer0_out[10295] <= ~(x[6949] & x[6950]);
     layer0_out[10296] <= x[2157] & x[2159];
     layer0_out[10297] <= x[3506] | x[3507];
     layer0_out[10298] <= ~(x[4713] | x[4714]);
     layer0_out[10299] <= 1'b0;
     layer0_out[10300] <= 1'b1;
     layer0_out[10301] <= ~(x[307] ^ x[309]);
     layer0_out[10302] <= x[7785] & ~x[7786];
     layer0_out[10303] <= x[1364] & x[1365];
     layer0_out[10304] <= ~(x[710] | x[712]);
     layer0_out[10305] <= ~(x[8599] & x[8600]);
     layer0_out[10306] <= x[8800] ^ x[8801];
     layer0_out[10307] <= ~x[3375];
     layer0_out[10308] <= x[2180];
     layer0_out[10309] <= x[2786] & x[2787];
     layer0_out[10310] <= ~x[1215];
     layer0_out[10311] <= ~(x[1040] | x[1041]);
     layer0_out[10312] <= ~(x[5392] & x[5393]);
     layer0_out[10313] <= ~(x[3285] & x[3286]);
     layer0_out[10314] <= x[4595] | x[4596];
     layer0_out[10315] <= 1'b0;
     layer0_out[10316] <= x[8368] & x[8369];
     layer0_out[10317] <= x[1245] & x[1246];
     layer0_out[10318] <= x[2987] ^ x[2988];
     layer0_out[10319] <= ~(x[1723] ^ x[1725]);
     layer0_out[10320] <= ~(x[6492] ^ x[6493]);
     layer0_out[10321] <= x[8206] | x[8207];
     layer0_out[10322] <= ~(x[3435] | x[3436]);
     layer0_out[10323] <= x[506] & x[508];
     layer0_out[10324] <= ~x[2280];
     layer0_out[10325] <= 1'b1;
     layer0_out[10326] <= x[4793] | x[4794];
     layer0_out[10327] <= ~(x[7019] | x[7020]);
     layer0_out[10328] <= ~(x[903] & x[905]);
     layer0_out[10329] <= 1'b1;
     layer0_out[10330] <= 1'b1;
     layer0_out[10331] <= ~(x[2047] ^ x[2049]);
     layer0_out[10332] <= x[2012] & x[2014];
     layer0_out[10333] <= x[7155] ^ x[7156];
     layer0_out[10334] <= 1'b0;
     layer0_out[10335] <= ~x[1807];
     layer0_out[10336] <= 1'b0;
     layer0_out[10337] <= x[8209];
     layer0_out[10338] <= x[2567] | x[2569];
     layer0_out[10339] <= x[1770];
     layer0_out[10340] <= 1'b1;
     layer0_out[10341] <= x[942] | x[944];
     layer0_out[10342] <= ~(x[5158] ^ x[5159]);
     layer0_out[10343] <= x[7824] & x[7825];
     layer0_out[10344] <= ~(x[8265] & x[8266]);
     layer0_out[10345] <= x[4931] & x[4932];
     layer0_out[10346] <= ~x[7317];
     layer0_out[10347] <= x[934];
     layer0_out[10348] <= 1'b1;
     layer0_out[10349] <= x[2116] & x[2118];
     layer0_out[10350] <= x[814] & x[816];
     layer0_out[10351] <= ~x[2846] | x[2847];
     layer0_out[10352] <= ~(x[4819] | x[4820]);
     layer0_out[10353] <= x[7206];
     layer0_out[10354] <= x[8900];
     layer0_out[10355] <= x[4554] & x[4555];
     layer0_out[10356] <= x[3049] & x[3050];
     layer0_out[10357] <= ~(x[3853] | x[3854]);
     layer0_out[10358] <= x[421];
     layer0_out[10359] <= x[4829] | x[4830];
     layer0_out[10360] <= ~x[1004];
     layer0_out[10361] <= x[9052] & x[9053];
     layer0_out[10362] <= 1'b1;
     layer0_out[10363] <= x[157] | x[159];
     layer0_out[10364] <= x[1778] & x[1780];
     layer0_out[10365] <= x[3558];
     layer0_out[10366] <= x[7218] ^ x[7219];
     layer0_out[10367] <= ~(x[1258] & x[1260]);
     layer0_out[10368] <= ~(x[1759] & x[1761]);
     layer0_out[10369] <= x[8886] ^ x[8887];
     layer0_out[10370] <= ~(x[2672] & x[2673]);
     layer0_out[10371] <= x[8376] & x[8377];
     layer0_out[10372] <= ~x[46] | x[48];
     layer0_out[10373] <= ~x[6270];
     layer0_out[10374] <= x[5373];
     layer0_out[10375] <= ~x[8152];
     layer0_out[10376] <= ~x[2401];
     layer0_out[10377] <= x[7617];
     layer0_out[10378] <= ~(x[1076] & x[1077]);
     layer0_out[10379] <= ~x[3891];
     layer0_out[10380] <= ~(x[3933] | x[3934]);
     layer0_out[10381] <= ~(x[8237] ^ x[8238]);
     layer0_out[10382] <= x[6704] | x[6705];
     layer0_out[10383] <= x[7937] & ~x[7936];
     layer0_out[10384] <= x[5303] & x[5304];
     layer0_out[10385] <= ~(x[7119] | x[7120]);
     layer0_out[10386] <= x[7803];
     layer0_out[10387] <= ~x[8544] | x[8545];
     layer0_out[10388] <= ~(x[2560] & x[2562]);
     layer0_out[10389] <= 1'b0;
     layer0_out[10390] <= x[2486] & x[2487];
     layer0_out[10391] <= x[1823];
     layer0_out[10392] <= ~x[4205];
     layer0_out[10393] <= x[6930] ^ x[6931];
     layer0_out[10394] <= x[1570] & x[1572];
     layer0_out[10395] <= ~x[6714];
     layer0_out[10396] <= x[8532] | x[8533];
     layer0_out[10397] <= x[3639] | x[3640];
     layer0_out[10398] <= x[1492];
     layer0_out[10399] <= ~x[2333];
     layer0_out[10400] <= x[7142] ^ x[7143];
     layer0_out[10401] <= ~(x[436] & x[437]);
     layer0_out[10402] <= x[1386];
     layer0_out[10403] <= ~(x[488] ^ x[489]);
     layer0_out[10404] <= 1'b1;
     layer0_out[10405] <= ~x[1469];
     layer0_out[10406] <= ~x[6116] | x[6117];
     layer0_out[10407] <= ~(x[5784] | x[5785]);
     layer0_out[10408] <= x[6675] | x[6676];
     layer0_out[10409] <= x[6933] & ~x[6934];
     layer0_out[10410] <= ~(x[4980] | x[4981]);
     layer0_out[10411] <= x[7643] & ~x[7644];
     layer0_out[10412] <= x[8778] | x[8779];
     layer0_out[10413] <= ~(x[2422] & x[2423]);
     layer0_out[10414] <= ~(x[2198] & x[2199]);
     layer0_out[10415] <= x[4769] ^ x[4770];
     layer0_out[10416] <= ~x[6027];
     layer0_out[10417] <= x[7469];
     layer0_out[10418] <= ~x[6418] | x[6417];
     layer0_out[10419] <= ~x[4943];
     layer0_out[10420] <= ~(x[1662] & x[1664]);
     layer0_out[10421] <= ~x[1213] | x[1214];
     layer0_out[10422] <= ~(x[1018] & x[1020]);
     layer0_out[10423] <= x[1077] ^ x[1078];
     layer0_out[10424] <= ~(x[712] ^ x[713]);
     layer0_out[10425] <= ~(x[2592] & x[2593]);
     layer0_out[10426] <= ~x[37];
     layer0_out[10427] <= x[6001];
     layer0_out[10428] <= x[1149];
     layer0_out[10429] <= ~(x[2774] ^ x[2776]);
     layer0_out[10430] <= x[8806] | x[8807];
     layer0_out[10431] <= x[8030];
     layer0_out[10432] <= ~(x[2116] & x[2117]);
     layer0_out[10433] <= ~x[4981];
     layer0_out[10434] <= ~x[9167];
     layer0_out[10435] <= ~x[7506] | x[7507];
     layer0_out[10436] <= 1'b0;
     layer0_out[10437] <= ~x[309];
     layer0_out[10438] <= 1'b1;
     layer0_out[10439] <= ~(x[1475] & x[1477]);
     layer0_out[10440] <= ~x[1069] | x[1067];
     layer0_out[10441] <= ~x[898];
     layer0_out[10442] <= x[6668] | x[6669];
     layer0_out[10443] <= x[3695] & x[3696];
     layer0_out[10444] <= ~(x[4836] ^ x[4837]);
     layer0_out[10445] <= ~x[3631];
     layer0_out[10446] <= ~(x[1402] & x[1403]);
     layer0_out[10447] <= ~(x[5143] | x[5144]);
     layer0_out[10448] <= ~(x[402] ^ x[403]);
     layer0_out[10449] <= ~(x[1721] & x[1722]);
     layer0_out[10450] <= ~(x[5357] & x[5358]);
     layer0_out[10451] <= ~(x[155] & x[157]);
     layer0_out[10452] <= x[8077] & ~x[8078];
     layer0_out[10453] <= ~(x[2181] & x[2182]);
     layer0_out[10454] <= x[479] ^ x[480];
     layer0_out[10455] <= x[1274] & x[1275];
     layer0_out[10456] <= x[4343] | x[4344];
     layer0_out[10457] <= ~(x[2285] & x[2286]);
     layer0_out[10458] <= 1'b1;
     layer0_out[10459] <= ~(x[1722] & x[1723]);
     layer0_out[10460] <= ~(x[9105] ^ x[9106]);
     layer0_out[10461] <= ~(x[995] ^ x[997]);
     layer0_out[10462] <= ~(x[2796] & x[2797]);
     layer0_out[10463] <= x[6866];
     layer0_out[10464] <= ~x[6015];
     layer0_out[10465] <= x[7204];
     layer0_out[10466] <= ~(x[3572] & x[3573]);
     layer0_out[10467] <= ~(x[6914] & x[6915]);
     layer0_out[10468] <= ~(x[8870] | x[8871]);
     layer0_out[10469] <= ~x[6005];
     layer0_out[10470] <= ~(x[2500] | x[2502]);
     layer0_out[10471] <= x[8418];
     layer0_out[10472] <= ~x[2117];
     layer0_out[10473] <= ~(x[554] ^ x[555]);
     layer0_out[10474] <= ~x[2120];
     layer0_out[10475] <= ~(x[205] & x[206]);
     layer0_out[10476] <= ~(x[7437] & x[7438]);
     layer0_out[10477] <= ~(x[4672] & x[4673]);
     layer0_out[10478] <= 1'b1;
     layer0_out[10479] <= x[6769] & x[6770];
     layer0_out[10480] <= 1'b1;
     layer0_out[10481] <= x[2955] & ~x[2956];
     layer0_out[10482] <= ~(x[5781] & x[5782]);
     layer0_out[10483] <= ~x[1507] | x[1508];
     layer0_out[10484] <= x[1484] & x[1486];
     layer0_out[10485] <= 1'b0;
     layer0_out[10486] <= ~(x[1433] | x[1435]);
     layer0_out[10487] <= ~x[8447];
     layer0_out[10488] <= ~(x[8693] | x[8694]);
     layer0_out[10489] <= x[4496] | x[4497];
     layer0_out[10490] <= ~(x[7034] | x[7035]);
     layer0_out[10491] <= x[1178];
     layer0_out[10492] <= x[9050] & ~x[9051];
     layer0_out[10493] <= x[1390] & x[1391];
     layer0_out[10494] <= 1'b0;
     layer0_out[10495] <= x[6434];
     layer0_out[10496] <= ~(x[2225] | x[2227]);
     layer0_out[10497] <= x[3346] | x[3347];
     layer0_out[10498] <= x[6141] | x[6142];
     layer0_out[10499] <= x[1399] & x[1400];
     layer0_out[10500] <= x[7508];
     layer0_out[10501] <= x[2049] & x[2050];
     layer0_out[10502] <= x[1467] ^ x[1468];
     layer0_out[10503] <= 1'b1;
     layer0_out[10504] <= x[1381] | x[1383];
     layer0_out[10505] <= x[7485] | x[7486];
     layer0_out[10506] <= 1'b1;
     layer0_out[10507] <= x[7841] & x[7842];
     layer0_out[10508] <= 1'b0;
     layer0_out[10509] <= 1'b0;
     layer0_out[10510] <= ~x[824];
     layer0_out[10511] <= x[968] & ~x[969];
     layer0_out[10512] <= x[1439];
     layer0_out[10513] <= 1'b1;
     layer0_out[10514] <= x[7642] | x[7643];
     layer0_out[10515] <= ~(x[1020] & x[1022]);
     layer0_out[10516] <= x[1682] & x[1684];
     layer0_out[10517] <= x[8084] & ~x[8083];
     layer0_out[10518] <= x[5483];
     layer0_out[10519] <= ~(x[441] ^ x[443]);
     layer0_out[10520] <= x[1578] & x[1579];
     layer0_out[10521] <= 1'b1;
     layer0_out[10522] <= ~(x[1568] & x[1569]);
     layer0_out[10523] <= x[113] & x[114];
     layer0_out[10524] <= x[4479] ^ x[4480];
     layer0_out[10525] <= ~x[2449];
     layer0_out[10526] <= 1'b0;
     layer0_out[10527] <= x[5296] & x[5297];
     layer0_out[10528] <= ~(x[5706] & x[5707]);
     layer0_out[10529] <= x[3637] ^ x[3638];
     layer0_out[10530] <= x[7844] | x[7845];
     layer0_out[10531] <= ~(x[4863] ^ x[4864]);
     layer0_out[10532] <= x[4696] & x[4697];
     layer0_out[10533] <= x[2271] | x[2273];
     layer0_out[10534] <= x[2539] & x[2540];
     layer0_out[10535] <= x[1543] ^ x[1544];
     layer0_out[10536] <= ~x[606];
     layer0_out[10537] <= x[3962] & ~x[3963];
     layer0_out[10538] <= ~x[6148];
     layer0_out[10539] <= x[169] ^ x[171];
     layer0_out[10540] <= 1'b0;
     layer0_out[10541] <= ~x[8121];
     layer0_out[10542] <= ~(x[1826] ^ x[1828]);
     layer0_out[10543] <= x[1854] ^ x[1856];
     layer0_out[10544] <= x[3965];
     layer0_out[10545] <= ~(x[2539] & x[2541]);
     layer0_out[10546] <= ~(x[1269] | x[1270]);
     layer0_out[10547] <= ~(x[8291] | x[8292]);
     layer0_out[10548] <= 1'b1;
     layer0_out[10549] <= ~(x[6827] | x[6828]);
     layer0_out[10550] <= 1'b0;
     layer0_out[10551] <= ~(x[7163] | x[7164]);
     layer0_out[10552] <= ~x[7471] | x[7470];
     layer0_out[10553] <= x[5736] ^ x[5737];
     layer0_out[10554] <= x[3127] | x[3128];
     layer0_out[10555] <= ~(x[8420] & x[8421]);
     layer0_out[10556] <= x[3452] | x[3453];
     layer0_out[10557] <= x[589];
     layer0_out[10558] <= ~x[6815];
     layer0_out[10559] <= x[8175];
     layer0_out[10560] <= x[3545] ^ x[3546];
     layer0_out[10561] <= x[4746] | x[4747];
     layer0_out[10562] <= x[4484] & x[4485];
     layer0_out[10563] <= ~x[1334];
     layer0_out[10564] <= x[7263] | x[7264];
     layer0_out[10565] <= ~x[2649] | x[2650];
     layer0_out[10566] <= ~(x[296] & x[297]);
     layer0_out[10567] <= x[2934] ^ x[2935];
     layer0_out[10568] <= x[2055] & x[2056];
     layer0_out[10569] <= x[6569] & ~x[6568];
     layer0_out[10570] <= ~(x[8732] | x[8733]);
     layer0_out[10571] <= x[5138] & x[5139];
     layer0_out[10572] <= x[2863] & x[2864];
     layer0_out[10573] <= x[1082];
     layer0_out[10574] <= ~(x[4088] & x[4089]);
     layer0_out[10575] <= x[2436];
     layer0_out[10576] <= ~(x[6425] | x[6426]);
     layer0_out[10577] <= x[7178];
     layer0_out[10578] <= x[4874];
     layer0_out[10579] <= x[8640];
     layer0_out[10580] <= ~(x[1212] & x[1213]);
     layer0_out[10581] <= ~(x[4543] & x[4544]);
     layer0_out[10582] <= x[3612] & x[3613];
     layer0_out[10583] <= x[3999] & x[4000];
     layer0_out[10584] <= ~(x[1491] ^ x[1493]);
     layer0_out[10585] <= ~x[9203];
     layer0_out[10586] <= x[2645] ^ x[2646];
     layer0_out[10587] <= x[4949] ^ x[4950];
     layer0_out[10588] <= ~(x[1350] ^ x[1351]);
     layer0_out[10589] <= ~(x[4590] & x[4591]);
     layer0_out[10590] <= ~(x[3239] | x[3240]);
     layer0_out[10591] <= x[5400] | x[5401];
     layer0_out[10592] <= ~(x[1000] & x[1001]);
     layer0_out[10593] <= ~x[4122];
     layer0_out[10594] <= x[1830] & x[1831];
     layer0_out[10595] <= 1'b1;
     layer0_out[10596] <= x[502] & x[504];
     layer0_out[10597] <= ~x[6968];
     layer0_out[10598] <= x[1817] & x[1818];
     layer0_out[10599] <= ~(x[1908] ^ x[1910]);
     layer0_out[10600] <= x[1016] ^ x[1018];
     layer0_out[10601] <= ~(x[4527] | x[4528]);
     layer0_out[10602] <= x[1316] & x[1317];
     layer0_out[10603] <= x[927] ^ x[928];
     layer0_out[10604] <= ~x[1252];
     layer0_out[10605] <= ~(x[3984] | x[3985]);
     layer0_out[10606] <= x[234] ^ x[235];
     layer0_out[10607] <= x[8487] | x[8488];
     layer0_out[10608] <= ~(x[754] ^ x[756]);
     layer0_out[10609] <= ~(x[2690] ^ x[2691]);
     layer0_out[10610] <= ~(x[1956] ^ x[1957]);
     layer0_out[10611] <= ~(x[1870] & x[1872]);
     layer0_out[10612] <= x[2888] & x[2889];
     layer0_out[10613] <= x[4032];
     layer0_out[10614] <= ~(x[7174] & x[7175]);
     layer0_out[10615] <= ~(x[1349] | x[1350]);
     layer0_out[10616] <= ~x[8043];
     layer0_out[10617] <= ~(x[3258] & x[3259]);
     layer0_out[10618] <= ~x[7717] | x[7716];
     layer0_out[10619] <= ~(x[2208] & x[2209]);
     layer0_out[10620] <= ~(x[7053] | x[7054]);
     layer0_out[10621] <= x[688];
     layer0_out[10622] <= x[8515] & x[8516];
     layer0_out[10623] <= x[1774] & x[1776];
     layer0_out[10624] <= ~x[174] | x[173];
     layer0_out[10625] <= x[6887] | x[6888];
     layer0_out[10626] <= ~(x[2310] & x[2311]);
     layer0_out[10627] <= x[223] & x[225];
     layer0_out[10628] <= ~(x[8592] | x[8593]);
     layer0_out[10629] <= ~(x[251] ^ x[252]);
     layer0_out[10630] <= ~x[7976];
     layer0_out[10631] <= ~x[803];
     layer0_out[10632] <= x[449] & x[451];
     layer0_out[10633] <= ~x[893];
     layer0_out[10634] <= ~x[7263];
     layer0_out[10635] <= ~(x[8702] ^ x[8703]);
     layer0_out[10636] <= ~(x[5137] & x[5138]);
     layer0_out[10637] <= ~x[8096] | x[8095];
     layer0_out[10638] <= ~(x[1334] | x[1336]);
     layer0_out[10639] <= x[1820] & x[1822];
     layer0_out[10640] <= ~x[71];
     layer0_out[10641] <= ~(x[8358] & x[8359]);
     layer0_out[10642] <= ~x[2007];
     layer0_out[10643] <= x[6852] ^ x[6853];
     layer0_out[10644] <= x[7461] ^ x[7462];
     layer0_out[10645] <= x[1692] ^ x[1693];
     layer0_out[10646] <= x[452] ^ x[454];
     layer0_out[10647] <= x[9059] | x[9060];
     layer0_out[10648] <= x[29] & x[31];
     layer0_out[10649] <= x[7896] | x[7897];
     layer0_out[10650] <= ~(x[8055] | x[8056]);
     layer0_out[10651] <= ~(x[5192] & x[5193]);
     layer0_out[10652] <= ~(x[645] & x[646]);
     layer0_out[10653] <= ~(x[6434] | x[6435]);
     layer0_out[10654] <= x[1033] & x[1035];
     layer0_out[10655] <= ~(x[6357] | x[6358]);
     layer0_out[10656] <= x[65] & x[67];
     layer0_out[10657] <= x[3155] | x[3156];
     layer0_out[10658] <= ~x[5669];
     layer0_out[10659] <= ~x[2285];
     layer0_out[10660] <= ~x[347];
     layer0_out[10661] <= ~(x[8863] ^ x[8864]);
     layer0_out[10662] <= x[1824] | x[1825];
     layer0_out[10663] <= x[1283] ^ x[1284];
     layer0_out[10664] <= ~x[457];
     layer0_out[10665] <= x[556] | x[557];
     layer0_out[10666] <= x[4487] | x[4488];
     layer0_out[10667] <= x[4860] | x[4861];
     layer0_out[10668] <= ~(x[1722] ^ x[1724]);
     layer0_out[10669] <= ~(x[3894] | x[3895]);
     layer0_out[10670] <= ~(x[911] | x[913]);
     layer0_out[10671] <= x[134];
     layer0_out[10672] <= x[2374] & x[2376];
     layer0_out[10673] <= x[3705] & ~x[3706];
     layer0_out[10674] <= ~(x[875] & x[876]);
     layer0_out[10675] <= ~(x[3959] | x[3960]);
     layer0_out[10676] <= x[4246] | x[4247];
     layer0_out[10677] <= ~x[3982];
     layer0_out[10678] <= ~x[2193] | x[2194];
     layer0_out[10679] <= x[8606] | x[8607];
     layer0_out[10680] <= ~(x[2159] ^ x[2160]);
     layer0_out[10681] <= ~(x[6015] | x[6016]);
     layer0_out[10682] <= x[8158] | x[8159];
     layer0_out[10683] <= x[8421] | x[8422];
     layer0_out[10684] <= x[792];
     layer0_out[10685] <= ~x[509];
     layer0_out[10686] <= ~(x[494] | x[496]);
     layer0_out[10687] <= x[2631] & x[2633];
     layer0_out[10688] <= x[6495];
     layer0_out[10689] <= x[3599];
     layer0_out[10690] <= 1'b0;
     layer0_out[10691] <= x[223] ^ x[224];
     layer0_out[10692] <= ~x[4899];
     layer0_out[10693] <= x[1306] ^ x[1308];
     layer0_out[10694] <= ~(x[435] ^ x[437]);
     layer0_out[10695] <= ~(x[3256] ^ x[3257]);
     layer0_out[10696] <= 1'b1;
     layer0_out[10697] <= x[5207] & x[5208];
     layer0_out[10698] <= x[8185] ^ x[8186];
     layer0_out[10699] <= ~(x[999] & x[1001]);
     layer0_out[10700] <= ~(x[584] ^ x[586]);
     layer0_out[10701] <= ~(x[219] & x[220]);
     layer0_out[10702] <= x[8524] & ~x[8523];
     layer0_out[10703] <= x[1020] & x[1021];
     layer0_out[10704] <= ~(x[8129] & x[8130]);
     layer0_out[10705] <= x[4385] & x[4386];
     layer0_out[10706] <= x[1813];
     layer0_out[10707] <= x[2419] & x[2420];
     layer0_out[10708] <= x[2107] & x[2109];
     layer0_out[10709] <= x[4307];
     layer0_out[10710] <= ~(x[3068] & x[3069]);
     layer0_out[10711] <= ~x[2980];
     layer0_out[10712] <= ~x[4147] | x[4148];
     layer0_out[10713] <= ~x[166];
     layer0_out[10714] <= ~(x[5115] ^ x[5116]);
     layer0_out[10715] <= ~(x[658] & x[660]);
     layer0_out[10716] <= ~(x[9197] & x[9198]);
     layer0_out[10717] <= x[477];
     layer0_out[10718] <= ~(x[4425] & x[4426]);
     layer0_out[10719] <= x[2461] & x[2463];
     layer0_out[10720] <= x[1260] ^ x[1262];
     layer0_out[10721] <= x[1170] ^ x[1171];
     layer0_out[10722] <= ~(x[6773] | x[6774]);
     layer0_out[10723] <= ~(x[6089] & x[6090]);
     layer0_out[10724] <= x[661] ^ x[662];
     layer0_out[10725] <= x[2189] & x[2190];
     layer0_out[10726] <= x[941] | x[943];
     layer0_out[10727] <= x[5184] & x[5185];
     layer0_out[10728] <= x[8286] | x[8287];
     layer0_out[10729] <= ~(x[1200] | x[1201]);
     layer0_out[10730] <= x[7888];
     layer0_out[10731] <= x[8854];
     layer0_out[10732] <= x[3039] & x[3040];
     layer0_out[10733] <= x[2409] ^ x[2411];
     layer0_out[10734] <= x[7630] ^ x[7631];
     layer0_out[10735] <= ~(x[6428] ^ x[6429]);
     layer0_out[10736] <= x[4575] & x[4576];
     layer0_out[10737] <= x[8463] | x[8464];
     layer0_out[10738] <= 1'b0;
     layer0_out[10739] <= x[8426] | x[8427];
     layer0_out[10740] <= ~(x[914] | x[915]);
     layer0_out[10741] <= x[2435] & x[2437];
     layer0_out[10742] <= x[1130] & ~x[1128];
     layer0_out[10743] <= ~x[274];
     layer0_out[10744] <= ~x[1240] | x[1241];
     layer0_out[10745] <= ~x[481] | x[483];
     layer0_out[10746] <= x[6611] | x[6612];
     layer0_out[10747] <= x[666] & x[667];
     layer0_out[10748] <= ~(x[9048] | x[9049]);
     layer0_out[10749] <= 1'b0;
     layer0_out[10750] <= ~x[7729];
     layer0_out[10751] <= x[6179];
     layer0_out[10752] <= 1'b1;
     layer0_out[10753] <= 1'b1;
     layer0_out[10754] <= ~(x[5492] | x[5493]);
     layer0_out[10755] <= x[6165] | x[6166];
     layer0_out[10756] <= 1'b1;
     layer0_out[10757] <= x[3048];
     layer0_out[10758] <= 1'b1;
     layer0_out[10759] <= x[6698] & x[6699];
     layer0_out[10760] <= ~(x[5104] & x[5105]);
     layer0_out[10761] <= x[6169] | x[6170];
     layer0_out[10762] <= x[7719];
     layer0_out[10763] <= x[157] & ~x[156];
     layer0_out[10764] <= x[831];
     layer0_out[10765] <= x[2160] ^ x[2162];
     layer0_out[10766] <= ~(x[7726] & x[7727]);
     layer0_out[10767] <= ~(x[8585] | x[8586]);
     layer0_out[10768] <= 1'b0;
     layer0_out[10769] <= ~x[5819];
     layer0_out[10770] <= x[3980] ^ x[3981];
     layer0_out[10771] <= x[6812] & x[6813];
     layer0_out[10772] <= x[7121] & x[7122];
     layer0_out[10773] <= x[6147];
     layer0_out[10774] <= x[2839] & x[2840];
     layer0_out[10775] <= ~(x[2613] & x[2615]);
     layer0_out[10776] <= x[1218] & x[1219];
     layer0_out[10777] <= 1'b1;
     layer0_out[10778] <= x[1939] | x[1940];
     layer0_out[10779] <= ~(x[623] & x[624]);
     layer0_out[10780] <= x[2578];
     layer0_out[10781] <= x[8138] & x[8139];
     layer0_out[10782] <= x[7199] | x[7200];
     layer0_out[10783] <= ~x[7040];
     layer0_out[10784] <= x[2249];
     layer0_out[10785] <= x[1008] & x[1010];
     layer0_out[10786] <= 1'b1;
     layer0_out[10787] <= ~x[2194];
     layer0_out[10788] <= x[859] | x[861];
     layer0_out[10789] <= ~x[3211];
     layer0_out[10790] <= ~(x[4141] & x[4142]);
     layer0_out[10791] <= ~(x[4235] & x[4236]);
     layer0_out[10792] <= x[2631] | x[2632];
     layer0_out[10793] <= x[6945] ^ x[6946];
     layer0_out[10794] <= x[6482] | x[6483];
     layer0_out[10795] <= ~(x[7701] | x[7702]);
     layer0_out[10796] <= ~(x[7509] & x[7510]);
     layer0_out[10797] <= x[2671] | x[2673];
     layer0_out[10798] <= ~(x[4600] ^ x[4601]);
     layer0_out[10799] <= ~x[1912];
     layer0_out[10800] <= x[2004] & x[2006];
     layer0_out[10801] <= x[1234];
     layer0_out[10802] <= ~(x[619] ^ x[620]);
     layer0_out[10803] <= x[4712] & x[4713];
     layer0_out[10804] <= x[639] & x[641];
     layer0_out[10805] <= ~(x[8243] | x[8244]);
     layer0_out[10806] <= x[5940] & ~x[5941];
     layer0_out[10807] <= ~(x[5662] ^ x[5663]);
     layer0_out[10808] <= x[1963] | x[1965];
     layer0_out[10809] <= ~x[8127];
     layer0_out[10810] <= ~x[3879];
     layer0_out[10811] <= ~x[5553];
     layer0_out[10812] <= ~(x[2256] | x[2257]);
     layer0_out[10813] <= x[8145];
     layer0_out[10814] <= x[186] & ~x[185];
     layer0_out[10815] <= ~x[5348];
     layer0_out[10816] <= x[8514];
     layer0_out[10817] <= ~x[7074];
     layer0_out[10818] <= x[2790];
     layer0_out[10819] <= x[8461] & ~x[8460];
     layer0_out[10820] <= ~(x[1472] & x[1473]);
     layer0_out[10821] <= ~(x[1092] & x[1094]);
     layer0_out[10822] <= x[7306];
     layer0_out[10823] <= ~(x[1649] ^ x[1651]);
     layer0_out[10824] <= x[7046] | x[7047];
     layer0_out[10825] <= ~x[2337];
     layer0_out[10826] <= x[784] & x[786];
     layer0_out[10827] <= x[1784] & x[1786];
     layer0_out[10828] <= 1'b1;
     layer0_out[10829] <= x[6462];
     layer0_out[10830] <= ~(x[3318] | x[3319]);
     layer0_out[10831] <= ~(x[1831] & x[1833]);
     layer0_out[10832] <= ~(x[1126] & x[1128]);
     layer0_out[10833] <= ~x[3263];
     layer0_out[10834] <= ~(x[4799] & x[4800]);
     layer0_out[10835] <= ~x[7510];
     layer0_out[10836] <= ~(x[7445] & x[7446]);
     layer0_out[10837] <= ~(x[2614] ^ x[2616]);
     layer0_out[10838] <= x[4025] | x[4026];
     layer0_out[10839] <= x[2305];
     layer0_out[10840] <= ~(x[375] ^ x[377]);
     layer0_out[10841] <= x[6938] | x[6939];
     layer0_out[10842] <= x[7808];
     layer0_out[10843] <= x[724] | x[725];
     layer0_out[10844] <= ~(x[895] | x[896]);
     layer0_out[10845] <= 1'b1;
     layer0_out[10846] <= ~x[2894];
     layer0_out[10847] <= x[3554] & ~x[3555];
     layer0_out[10848] <= x[850] & x[852];
     layer0_out[10849] <= ~(x[6477] | x[6478]);
     layer0_out[10850] <= ~(x[8699] & x[8700]);
     layer0_out[10851] <= x[2545];
     layer0_out[10852] <= 1'b1;
     layer0_out[10853] <= ~(x[647] | x[649]);
     layer0_out[10854] <= ~x[3130];
     layer0_out[10855] <= ~x[2375];
     layer0_out[10856] <= ~x[4105];
     layer0_out[10857] <= x[6560] & x[6561];
     layer0_out[10858] <= x[1199] ^ x[1201];
     layer0_out[10859] <= x[6932] & x[6933];
     layer0_out[10860] <= x[97];
     layer0_out[10861] <= x[2206];
     layer0_out[10862] <= ~(x[3047] & x[3048]);
     layer0_out[10863] <= x[1095] | x[1097];
     layer0_out[10864] <= ~(x[8498] | x[8499]);
     layer0_out[10865] <= ~(x[1664] ^ x[1665]);
     layer0_out[10866] <= ~x[1052];
     layer0_out[10867] <= ~(x[2853] & x[2854]);
     layer0_out[10868] <= x[2652];
     layer0_out[10869] <= x[59] & ~x[60];
     layer0_out[10870] <= x[7902];
     layer0_out[10871] <= ~(x[1218] & x[1220]);
     layer0_out[10872] <= ~(x[1263] & x[1264]);
     layer0_out[10873] <= x[2274] | x[2276];
     layer0_out[10874] <= x[421] | x[422];
     layer0_out[10875] <= ~(x[6505] | x[6506]);
     layer0_out[10876] <= ~(x[7589] ^ x[7590]);
     layer0_out[10877] <= 1'b1;
     layer0_out[10878] <= x[4111] ^ x[4112];
     layer0_out[10879] <= x[8891] ^ x[8892];
     layer0_out[10880] <= ~(x[6127] & x[6128]);
     layer0_out[10881] <= ~(x[7953] | x[7954]);
     layer0_out[10882] <= ~(x[8919] | x[8920]);
     layer0_out[10883] <= x[88] ^ x[90];
     layer0_out[10884] <= x[1082] & ~x[1081];
     layer0_out[10885] <= ~(x[286] & x[287]);
     layer0_out[10886] <= ~(x[1598] & x[1600]);
     layer0_out[10887] <= x[656] & ~x[655];
     layer0_out[10888] <= x[1055] & x[1057];
     layer0_out[10889] <= ~x[317];
     layer0_out[10890] <= x[3084] & x[3085];
     layer0_out[10891] <= x[4335] | x[4336];
     layer0_out[10892] <= ~x[3658];
     layer0_out[10893] <= x[6283] | x[6284];
     layer0_out[10894] <= x[1899] & x[1900];
     layer0_out[10895] <= 1'b0;
     layer0_out[10896] <= x[7235];
     layer0_out[10897] <= ~(x[8524] | x[8525]);
     layer0_out[10898] <= ~(x[8020] | x[8021]);
     layer0_out[10899] <= ~(x[8933] & x[8934]);
     layer0_out[10900] <= ~(x[4607] & x[4608]);
     layer0_out[10901] <= x[965] ^ x[967];
     layer0_out[10902] <= ~(x[2356] & x[2357]);
     layer0_out[10903] <= ~(x[1093] & x[1094]);
     layer0_out[10904] <= x[3230] & x[3231];
     layer0_out[10905] <= x[1753] & x[1755];
     layer0_out[10906] <= ~(x[192] ^ x[194]);
     layer0_out[10907] <= ~(x[7351] ^ x[7352]);
     layer0_out[10908] <= ~(x[5412] ^ x[5413]);
     layer0_out[10909] <= ~(x[7114] ^ x[7115]);
     layer0_out[10910] <= ~(x[2551] & x[2552]);
     layer0_out[10911] <= x[595] ^ x[597];
     layer0_out[10912] <= ~(x[2244] & x[2246]);
     layer0_out[10913] <= ~(x[2773] & x[2775]);
     layer0_out[10914] <= x[2149] | x[2151];
     layer0_out[10915] <= x[4536] & x[4537];
     layer0_out[10916] <= x[5484] & ~x[5483];
     layer0_out[10917] <= x[5322] & x[5323];
     layer0_out[10918] <= ~x[4054];
     layer0_out[10919] <= ~(x[3826] | x[3827]);
     layer0_out[10920] <= ~(x[8195] & x[8196]);
     layer0_out[10921] <= ~(x[773] & x[775]);
     layer0_out[10922] <= ~(x[392] ^ x[394]);
     layer0_out[10923] <= ~(x[5340] & x[5341]);
     layer0_out[10924] <= x[2000] | x[2002];
     layer0_out[10925] <= ~(x[1660] & x[1661]);
     layer0_out[10926] <= x[6163] | x[6164];
     layer0_out[10927] <= ~(x[1349] & x[1351]);
     layer0_out[10928] <= ~(x[2253] & x[2255]);
     layer0_out[10929] <= ~(x[503] | x[505]);
     layer0_out[10930] <= ~(x[2431] & x[2433]);
     layer0_out[10931] <= x[2257];
     layer0_out[10932] <= ~(x[8461] ^ x[8462]);
     layer0_out[10933] <= x[2594] & x[2595];
     layer0_out[10934] <= ~(x[5098] & x[5099]);
     layer0_out[10935] <= x[2284] & x[2285];
     layer0_out[10936] <= 1'b1;
     layer0_out[10937] <= ~(x[984] | x[985]);
     layer0_out[10938] <= ~x[2512];
     layer0_out[10939] <= 1'b0;
     layer0_out[10940] <= x[1526];
     layer0_out[10941] <= x[2174] & x[2176];
     layer0_out[10942] <= ~(x[2789] ^ x[2790]);
     layer0_out[10943] <= x[6860];
     layer0_out[10944] <= x[6369] | x[6370];
     layer0_out[10945] <= ~x[3421];
     layer0_out[10946] <= ~x[7066] | x[7067];
     layer0_out[10947] <= ~x[5860];
     layer0_out[10948] <= x[2222] & x[2224];
     layer0_out[10949] <= x[4892];
     layer0_out[10950] <= ~x[6164];
     layer0_out[10951] <= ~(x[43] ^ x[44]);
     layer0_out[10952] <= 1'b0;
     layer0_out[10953] <= x[8471] & x[8472];
     layer0_out[10954] <= ~(x[4129] ^ x[4130]);
     layer0_out[10955] <= x[3904] | x[3905];
     layer0_out[10956] <= x[8793] ^ x[8794];
     layer0_out[10957] <= 1'b1;
     layer0_out[10958] <= ~(x[1543] | x[1545]);
     layer0_out[10959] <= x[5019] & ~x[5018];
     layer0_out[10960] <= ~x[419];
     layer0_out[10961] <= ~(x[9010] ^ x[9011]);
     layer0_out[10962] <= x[4951] ^ x[4952];
     layer0_out[10963] <= x[2680] ^ x[2681];
     layer0_out[10964] <= x[7320] | x[7321];
     layer0_out[10965] <= ~(x[8827] | x[8828]);
     layer0_out[10966] <= ~x[6973];
     layer0_out[10967] <= x[3237] ^ x[3238];
     layer0_out[10968] <= ~x[1619] | x[1620];
     layer0_out[10969] <= x[6662];
     layer0_out[10970] <= x[2462];
     layer0_out[10971] <= ~x[5951];
     layer0_out[10972] <= x[5146];
     layer0_out[10973] <= x[2762] ^ x[2763];
     layer0_out[10974] <= x[7686] | x[7687];
     layer0_out[10975] <= ~(x[321] ^ x[322]);
     layer0_out[10976] <= ~(x[3570] ^ x[3571]);
     layer0_out[10977] <= x[8193] | x[8194];
     layer0_out[10978] <= x[1461] & x[1463];
     layer0_out[10979] <= ~(x[446] & x[447]);
     layer0_out[10980] <= ~x[2732] | x[2730];
     layer0_out[10981] <= x[2765] ^ x[2766];
     layer0_out[10982] <= x[8256] | x[8257];
     layer0_out[10983] <= ~(x[9165] & x[9166]);
     layer0_out[10984] <= ~(x[5448] & x[5449]);
     layer0_out[10985] <= x[4] & x[5];
     layer0_out[10986] <= ~(x[7233] | x[7234]);
     layer0_out[10987] <= x[271] & x[273];
     layer0_out[10988] <= x[2559] ^ x[2560];
     layer0_out[10989] <= 1'b1;
     layer0_out[10990] <= ~(x[701] | x[702]);
     layer0_out[10991] <= x[1517] & x[1518];
     layer0_out[10992] <= x[2735] & x[2736];
     layer0_out[10993] <= x[2190] ^ x[2192];
     layer0_out[10994] <= x[8068];
     layer0_out[10995] <= x[4008] & ~x[4007];
     layer0_out[10996] <= ~(x[5912] & x[5913]);
     layer0_out[10997] <= ~x[1083] | x[1085];
     layer0_out[10998] <= x[2583] & x[2584];
     layer0_out[10999] <= x[7278] & x[7279];
     layer0_out[11000] <= x[997] & x[999];
     layer0_out[11001] <= ~(x[4845] | x[4846]);
     layer0_out[11002] <= ~x[678] | x[679];
     layer0_out[11003] <= ~(x[3341] | x[3342]);
     layer0_out[11004] <= ~x[1941];
     layer0_out[11005] <= x[1616] ^ x[1618];
     layer0_out[11006] <= x[4059] ^ x[4060];
     layer0_out[11007] <= ~x[5648];
     layer0_out[11008] <= x[6639];
     layer0_out[11009] <= ~(x[10] & x[12]);
     layer0_out[11010] <= ~(x[2937] & x[2938]);
     layer0_out[11011] <= ~(x[1310] & x[1311]);
     layer0_out[11012] <= ~(x[3075] & x[3076]);
     layer0_out[11013] <= x[2698] & x[2700];
     layer0_out[11014] <= x[602] ^ x[604];
     layer0_out[11015] <= ~x[8350];
     layer0_out[11016] <= x[4751] & ~x[4752];
     layer0_out[11017] <= ~(x[1430] ^ x[1432]);
     layer0_out[11018] <= 1'b1;
     layer0_out[11019] <= x[2248] & x[2249];
     layer0_out[11020] <= ~(x[5133] & x[5134]);
     layer0_out[11021] <= ~(x[1105] & x[1107]);
     layer0_out[11022] <= ~(x[4327] & x[4328]);
     layer0_out[11023] <= ~(x[6862] | x[6863]);
     layer0_out[11024] <= x[4766] ^ x[4767];
     layer0_out[11025] <= x[4766];
     layer0_out[11026] <= ~(x[4163] ^ x[4164]);
     layer0_out[11027] <= 1'b0;
     layer0_out[11028] <= x[2077];
     layer0_out[11029] <= x[7104];
     layer0_out[11030] <= 1'b1;
     layer0_out[11031] <= x[618] & x[619];
     layer0_out[11032] <= x[2971] | x[2972];
     layer0_out[11033] <= ~x[2354];
     layer0_out[11034] <= ~(x[111] ^ x[112]);
     layer0_out[11035] <= ~(x[1817] & x[1819]);
     layer0_out[11036] <= ~x[1990];
     layer0_out[11037] <= ~(x[7782] | x[7783]);
     layer0_out[11038] <= ~(x[7185] | x[7186]);
     layer0_out[11039] <= ~(x[8314] | x[8315]);
     layer0_out[11040] <= ~(x[2504] ^ x[2505]);
     layer0_out[11041] <= ~(x[1447] & x[1449]);
     layer0_out[11042] <= x[3399] | x[3400];
     layer0_out[11043] <= x[8022] ^ x[8023];
     layer0_out[11044] <= ~x[1775];
     layer0_out[11045] <= ~(x[482] | x[483]);
     layer0_out[11046] <= 1'b0;
     layer0_out[11047] <= 1'b1;
     layer0_out[11048] <= ~x[5461];
     layer0_out[11049] <= ~(x[294] | x[295]);
     layer0_out[11050] <= x[5926];
     layer0_out[11051] <= x[267] & ~x[266];
     layer0_out[11052] <= x[4295] ^ x[4296];
     layer0_out[11053] <= ~x[8411];
     layer0_out[11054] <= ~x[3029] | x[3028];
     layer0_out[11055] <= ~(x[3050] & x[3051]);
     layer0_out[11056] <= x[3365] | x[3366];
     layer0_out[11057] <= ~(x[5485] & x[5486]);
     layer0_out[11058] <= 1'b0;
     layer0_out[11059] <= ~x[1441];
     layer0_out[11060] <= x[758] & x[759];
     layer0_out[11061] <= x[6162];
     layer0_out[11062] <= ~(x[1701] & x[1702]);
     layer0_out[11063] <= x[9166] | x[9167];
     layer0_out[11064] <= x[4671] | x[4672];
     layer0_out[11065] <= x[5266] ^ x[5267];
     layer0_out[11066] <= x[1321] | x[1322];
     layer0_out[11067] <= x[7862] ^ x[7863];
     layer0_out[11068] <= 1'b1;
     layer0_out[11069] <= x[7888] | x[7889];
     layer0_out[11070] <= ~(x[708] ^ x[710]);
     layer0_out[11071] <= x[117] | x[118];
     layer0_out[11072] <= ~(x[2560] & x[2561]);
     layer0_out[11073] <= x[4236] & ~x[4237];
     layer0_out[11074] <= x[8261] | x[8262];
     layer0_out[11075] <= ~x[7744];
     layer0_out[11076] <= x[2632];
     layer0_out[11077] <= x[6535] | x[6536];
     layer0_out[11078] <= ~x[1580];
     layer0_out[11079] <= ~(x[805] & x[807]);
     layer0_out[11080] <= ~(x[2103] | x[2105]);
     layer0_out[11081] <= 1'b1;
     layer0_out[11082] <= x[5709];
     layer0_out[11083] <= 1'b0;
     layer0_out[11084] <= ~(x[3889] | x[3890]);
     layer0_out[11085] <= 1'b0;
     layer0_out[11086] <= x[468] & x[469];
     layer0_out[11087] <= 1'b1;
     layer0_out[11088] <= ~(x[1807] & x[1809]);
     layer0_out[11089] <= x[6118] & x[6119];
     layer0_out[11090] <= ~x[3021];
     layer0_out[11091] <= x[3969] & x[3970];
     layer0_out[11092] <= x[4986];
     layer0_out[11093] <= ~(x[2166] | x[2167]);
     layer0_out[11094] <= x[3097] | x[3098];
     layer0_out[11095] <= x[2736] | x[2737];
     layer0_out[11096] <= x[195] & x[196];
     layer0_out[11097] <= x[3098];
     layer0_out[11098] <= 1'b0;
     layer0_out[11099] <= x[1060] & ~x[1058];
     layer0_out[11100] <= 1'b0;
     layer0_out[11101] <= ~(x[7549] & x[7550]);
     layer0_out[11102] <= ~(x[2969] ^ x[2970]);
     layer0_out[11103] <= x[4342] | x[4343];
     layer0_out[11104] <= ~(x[2287] | x[2288]);
     layer0_out[11105] <= ~(x[2822] | x[2823]);
     layer0_out[11106] <= x[7556] & ~x[7555];
     layer0_out[11107] <= x[1838] | x[1839];
     layer0_out[11108] <= x[6514] | x[6515];
     layer0_out[11109] <= ~(x[6673] & x[6674]);
     layer0_out[11110] <= 1'b0;
     layer0_out[11111] <= ~(x[5504] ^ x[5505]);
     layer0_out[11112] <= x[7853] & x[7854];
     layer0_out[11113] <= ~(x[6186] | x[6187]);
     layer0_out[11114] <= ~(x[2961] ^ x[2962]);
     layer0_out[11115] <= x[2625] & x[2626];
     layer0_out[11116] <= x[1850] & x[1852];
     layer0_out[11117] <= ~(x[5922] & x[5923]);
     layer0_out[11118] <= ~(x[2890] & x[2891]);
     layer0_out[11119] <= 1'b1;
     layer0_out[11120] <= ~(x[5366] & x[5367]);
     layer0_out[11121] <= ~(x[1277] | x[1278]);
     layer0_out[11122] <= x[7307] | x[7308];
     layer0_out[11123] <= x[2079] & x[2080];
     layer0_out[11124] <= x[1158] & x[1160];
     layer0_out[11125] <= x[1518] ^ x[1519];
     layer0_out[11126] <= x[6071] & x[6072];
     layer0_out[11127] <= ~(x[4715] ^ x[4716]);
     layer0_out[11128] <= x[8704];
     layer0_out[11129] <= x[328] & x[329];
     layer0_out[11130] <= x[2135] | x[2136];
     layer0_out[11131] <= ~(x[3046] & x[3047]);
     layer0_out[11132] <= x[2662] & x[2664];
     layer0_out[11133] <= ~(x[602] & x[603]);
     layer0_out[11134] <= ~(x[1507] & x[1509]);
     layer0_out[11135] <= ~x[1608] | x[1609];
     layer0_out[11136] <= ~x[7986] | x[7987];
     layer0_out[11137] <= x[8106];
     layer0_out[11138] <= ~(x[7243] | x[7244]);
     layer0_out[11139] <= x[8987] & x[8988];
     layer0_out[11140] <= ~x[2763];
     layer0_out[11141] <= x[1864] & x[1865];
     layer0_out[11142] <= ~(x[4938] | x[4939]);
     layer0_out[11143] <= x[2075] & x[2077];
     layer0_out[11144] <= 1'b1;
     layer0_out[11145] <= ~(x[3064] & x[3065]);
     layer0_out[11146] <= x[7957];
     layer0_out[11147] <= ~(x[5178] & x[5179]);
     layer0_out[11148] <= ~(x[2270] | x[2272]);
     layer0_out[11149] <= ~(x[3829] | x[3830]);
     layer0_out[11150] <= ~(x[8001] | x[8002]);
     layer0_out[11151] <= x[1224] & x[1225];
     layer0_out[11152] <= ~(x[1026] & x[1027]);
     layer0_out[11153] <= ~(x[4526] | x[4527]);
     layer0_out[11154] <= ~(x[8537] | x[8538]);
     layer0_out[11155] <= ~x[2643];
     layer0_out[11156] <= x[5608] & x[5609];
     layer0_out[11157] <= ~(x[8483] ^ x[8484]);
     layer0_out[11158] <= x[1625] | x[1626];
     layer0_out[11159] <= x[476];
     layer0_out[11160] <= x[8712] | x[8713];
     layer0_out[11161] <= x[1084] | x[1085];
     layer0_out[11162] <= ~(x[2336] | x[2337]);
     layer0_out[11163] <= x[5471] & x[5472];
     layer0_out[11164] <= x[6047] | x[6048];
     layer0_out[11165] <= ~(x[2738] & x[2739]);
     layer0_out[11166] <= ~(x[5901] & x[5902]);
     layer0_out[11167] <= ~(x[584] ^ x[585]);
     layer0_out[11168] <= x[227] & ~x[229];
     layer0_out[11169] <= ~(x[2364] | x[2365]);
     layer0_out[11170] <= ~(x[2759] ^ x[2760]);
     layer0_out[11171] <= x[5991];
     layer0_out[11172] <= x[7440] | x[7441];
     layer0_out[11173] <= x[4811];
     layer0_out[11174] <= ~x[1082];
     layer0_out[11175] <= ~(x[1335] & x[1336]);
     layer0_out[11176] <= ~(x[2214] & x[2215]);
     layer0_out[11177] <= ~x[7666];
     layer0_out[11178] <= ~x[3456];
     layer0_out[11179] <= x[384] & x[385];
     layer0_out[11180] <= x[3912] | x[3913];
     layer0_out[11181] <= x[6948] ^ x[6949];
     layer0_out[11182] <= x[9101] & x[9102];
     layer0_out[11183] <= ~(x[1246] & x[1247]);
     layer0_out[11184] <= ~(x[2708] ^ x[2710]);
     layer0_out[11185] <= ~(x[2377] & x[2378]);
     layer0_out[11186] <= ~(x[3186] & x[3187]);
     layer0_out[11187] <= ~(x[6988] ^ x[6989]);
     layer0_out[11188] <= 1'b0;
     layer0_out[11189] <= ~x[5460];
     layer0_out[11190] <= 1'b0;
     layer0_out[11191] <= x[2311] & x[2312];
     layer0_out[11192] <= x[6082] ^ x[6083];
     layer0_out[11193] <= x[2318] & x[2320];
     layer0_out[11194] <= ~(x[6754] & x[6755]);
     layer0_out[11195] <= ~(x[197] | x[199]);
     layer0_out[11196] <= x[7932];
     layer0_out[11197] <= x[9193];
     layer0_out[11198] <= x[3297] | x[3298];
     layer0_out[11199] <= ~(x[6192] | x[6193]);
     layer0_out[11200] <= x[1411] & ~x[1412];
     layer0_out[11201] <= x[3357];
     layer0_out[11202] <= ~x[330] | x[328];
     layer0_out[11203] <= x[7585] & x[7586];
     layer0_out[11204] <= ~(x[2859] & x[2860]);
     layer0_out[11205] <= ~x[28] | x[27];
     layer0_out[11206] <= ~(x[1351] & x[1353]);
     layer0_out[11207] <= ~(x[4228] ^ x[4229]);
     layer0_out[11208] <= ~(x[1697] ^ x[1698]);
     layer0_out[11209] <= ~(x[5247] & x[5248]);
     layer0_out[11210] <= x[8112];
     layer0_out[11211] <= ~(x[7669] | x[7670]);
     layer0_out[11212] <= ~(x[1693] ^ x[1695]);
     layer0_out[11213] <= ~(x[876] & x[878]);
     layer0_out[11214] <= x[6705];
     layer0_out[11215] <= x[8569];
     layer0_out[11216] <= x[5132] & x[5133];
     layer0_out[11217] <= x[878] & x[880];
     layer0_out[11218] <= x[355];
     layer0_out[11219] <= x[3332] | x[3333];
     layer0_out[11220] <= x[1494] | x[1495];
     layer0_out[11221] <= ~(x[1510] | x[1512]);
     layer0_out[11222] <= x[4304] ^ x[4305];
     layer0_out[11223] <= x[2454] & x[2456];
     layer0_out[11224] <= ~x[7385];
     layer0_out[11225] <= x[79] | x[80];
     layer0_out[11226] <= ~(x[9037] | x[9038]);
     layer0_out[11227] <= ~x[1904];
     layer0_out[11228] <= x[1057] | x[1058];
     layer0_out[11229] <= ~(x[8332] | x[8333]);
     layer0_out[11230] <= 1'b1;
     layer0_out[11231] <= x[4068];
     layer0_out[11232] <= x[4514] & ~x[4513];
     layer0_out[11233] <= ~(x[851] & x[853]);
     layer0_out[11234] <= ~x[436];
     layer0_out[11235] <= 1'b0;
     layer0_out[11236] <= x[6471] ^ x[6472];
     layer0_out[11237] <= x[2150] & x[2152];
     layer0_out[11238] <= x[2927] & x[2928];
     layer0_out[11239] <= ~(x[4196] & x[4197]);
     layer0_out[11240] <= ~x[3426] | x[3427];
     layer0_out[11241] <= x[9072] | x[9073];
     layer0_out[11242] <= x[6210] | x[6211];
     layer0_out[11243] <= ~(x[5230] ^ x[5231]);
     layer0_out[11244] <= x[7655];
     layer0_out[11245] <= ~(x[2688] & x[2690]);
     layer0_out[11246] <= x[2514] & x[2516];
     layer0_out[11247] <= x[2645] ^ x[2647];
     layer0_out[11248] <= x[7825] | x[7826];
     layer0_out[11249] <= ~(x[1564] & x[1565]);
     layer0_out[11250] <= x[947] | x[949];
     layer0_out[11251] <= x[4501] | x[4502];
     layer0_out[11252] <= ~(x[8015] | x[8016]);
     layer0_out[11253] <= x[177];
     layer0_out[11254] <= ~(x[1717] & x[1719]);
     layer0_out[11255] <= x[3298] ^ x[3299];
     layer0_out[11256] <= x[8467] & x[8468];
     layer0_out[11257] <= x[1870];
     layer0_out[11258] <= ~x[7974];
     layer0_out[11259] <= ~(x[4174] & x[4175]);
     layer0_out[11260] <= ~x[5122];
     layer0_out[11261] <= ~x[7662];
     layer0_out[11262] <= x[1865] & x[1866];
     layer0_out[11263] <= ~x[2896] | x[2897];
     layer0_out[11264] <= x[9164] | x[9165];
     layer0_out[11265] <= 1'b1;
     layer0_out[11266] <= x[3445] | x[3446];
     layer0_out[11267] <= x[2385] & x[2386];
     layer0_out[11268] <= x[3842] | x[3843];
     layer0_out[11269] <= ~(x[5924] ^ x[5925]);
     layer0_out[11270] <= ~x[2315] | x[2316];
     layer0_out[11271] <= ~(x[2139] & x[2140]);
     layer0_out[11272] <= x[1007] | x[1008];
     layer0_out[11273] <= x[5506] & x[5507];
     layer0_out[11274] <= ~(x[1398] & x[1400]);
     layer0_out[11275] <= x[8176] | x[8177];
     layer0_out[11276] <= ~(x[1336] & x[1337]);
     layer0_out[11277] <= ~x[6602];
     layer0_out[11278] <= x[4176] & x[4177];
     layer0_out[11279] <= ~(x[403] ^ x[405]);
     layer0_out[11280] <= ~x[80];
     layer0_out[11281] <= ~x[2816];
     layer0_out[11282] <= x[5726];
     layer0_out[11283] <= x[753] ^ x[755];
     layer0_out[11284] <= x[7779] & ~x[7778];
     layer0_out[11285] <= ~(x[3898] & x[3899]);
     layer0_out[11286] <= ~x[2346] | x[2344];
     layer0_out[11287] <= ~x[6318] | x[6319];
     layer0_out[11288] <= x[1172] ^ x[1174];
     layer0_out[11289] <= x[3371] | x[3372];
     layer0_out[11290] <= ~(x[3708] ^ x[3709]);
     layer0_out[11291] <= ~x[4136] | x[4137];
     layer0_out[11292] <= ~(x[1643] ^ x[1644]);
     layer0_out[11293] <= ~x[190] | x[189];
     layer0_out[11294] <= ~(x[9120] ^ x[9121]);
     layer0_out[11295] <= ~(x[7593] | x[7594]);
     layer0_out[11296] <= x[5832];
     layer0_out[11297] <= x[925] & x[926];
     layer0_out[11298] <= x[7424] ^ x[7425];
     layer0_out[11299] <= x[1505] & ~x[1506];
     layer0_out[11300] <= 1'b0;
     layer0_out[11301] <= ~x[7759];
     layer0_out[11302] <= 1'b0;
     layer0_out[11303] <= 1'b1;
     layer0_out[11304] <= ~x[6643];
     layer0_out[11305] <= ~x[6422];
     layer0_out[11306] <= x[333] & x[335];
     layer0_out[11307] <= 1'b0;
     layer0_out[11308] <= ~(x[2209] & x[2210]);
     layer0_out[11309] <= ~(x[365] & x[366]);
     layer0_out[11310] <= ~x[2480];
     layer0_out[11311] <= ~x[3789];
     layer0_out[11312] <= ~x[1547];
     layer0_out[11313] <= 1'b1;
     layer0_out[11314] <= x[5073] ^ x[5074];
     layer0_out[11315] <= ~(x[2598] & x[2600]);
     layer0_out[11316] <= ~(x[649] ^ x[650]);
     layer0_out[11317] <= x[1162] & ~x[1160];
     layer0_out[11318] <= ~x[368] | x[370];
     layer0_out[11319] <= x[2788] & x[2789];
     layer0_out[11320] <= x[4990] ^ x[4991];
     layer0_out[11321] <= x[1759] & x[1760];
     layer0_out[11322] <= ~(x[2073] & x[2074]);
     layer0_out[11323] <= x[1047] ^ x[1048];
     layer0_out[11324] <= ~(x[2140] & x[2141]);
     layer0_out[11325] <= 1'b1;
     layer0_out[11326] <= x[6570] | x[6571];
     layer0_out[11327] <= ~(x[3398] ^ x[3399]);
     layer0_out[11328] <= ~x[27] | x[29];
     layer0_out[11329] <= x[1963] | x[1964];
     layer0_out[11330] <= x[540] | x[541];
     layer0_out[11331] <= 1'b1;
     layer0_out[11332] <= 1'b1;
     layer0_out[11333] <= x[768] | x[769];
     layer0_out[11334] <= ~(x[2246] & x[2248]);
     layer0_out[11335] <= ~x[2629] | x[2630];
     layer0_out[11336] <= 1'b0;
     layer0_out[11337] <= 1'b0;
     layer0_out[11338] <= ~(x[1206] ^ x[1207]);
     layer0_out[11339] <= ~(x[350] | x[352]);
     layer0_out[11340] <= x[2767] ^ x[2769];
     layer0_out[11341] <= x[3158] ^ x[3159];
     layer0_out[11342] <= ~x[2352];
     layer0_out[11343] <= x[4157];
     layer0_out[11344] <= 1'b1;
     layer0_out[11345] <= x[2930] & x[2931];
     layer0_out[11346] <= ~(x[1700] & x[1702]);
     layer0_out[11347] <= x[6656] & x[6657];
     layer0_out[11348] <= ~(x[7389] | x[7390]);
     layer0_out[11349] <= x[6609] | x[6610];
     layer0_out[11350] <= ~x[9090];
     layer0_out[11351] <= x[4992] ^ x[4993];
     layer0_out[11352] <= x[2024] & x[2025];
     layer0_out[11353] <= ~(x[6190] ^ x[6191]);
     layer0_out[11354] <= ~(x[1628] & x[1630]);
     layer0_out[11355] <= ~(x[2176] & x[2177]);
     layer0_out[11356] <= x[3441] | x[3442];
     layer0_out[11357] <= x[3165] ^ x[3166];
     layer0_out[11358] <= ~(x[4038] | x[4039]);
     layer0_out[11359] <= x[3680] & x[3681];
     layer0_out[11360] <= ~(x[5410] & x[5411]);
     layer0_out[11361] <= ~(x[1571] ^ x[1572]);
     layer0_out[11362] <= ~(x[23] | x[24]);
     layer0_out[11363] <= x[229] ^ x[230];
     layer0_out[11364] <= x[5771] | x[5772];
     layer0_out[11365] <= ~x[2731] | x[2732];
     layer0_out[11366] <= ~x[1072];
     layer0_out[11367] <= x[6315] | x[6316];
     layer0_out[11368] <= ~x[2875];
     layer0_out[11369] <= ~(x[1861] ^ x[1863]);
     layer0_out[11370] <= x[1520] & x[1521];
     layer0_out[11371] <= ~(x[4368] ^ x[4369]);
     layer0_out[11372] <= x[1334] & x[1335];
     layer0_out[11373] <= ~x[8662];
     layer0_out[11374] <= 1'b0;
     layer0_out[11375] <= x[2957] | x[2958];
     layer0_out[11376] <= ~x[1911];
     layer0_out[11377] <= ~x[996];
     layer0_out[11378] <= x[3416] | x[3417];
     layer0_out[11379] <= ~(x[3578] ^ x[3579]);
     layer0_out[11380] <= ~(x[2168] & x[2170]);
     layer0_out[11381] <= ~x[3133];
     layer0_out[11382] <= x[7426] | x[7427];
     layer0_out[11383] <= ~x[1435] | x[1434];
     layer0_out[11384] <= x[5167] | x[5168];
     layer0_out[11385] <= x[1859] & x[1861];
     layer0_out[11386] <= ~x[9200];
     layer0_out[11387] <= ~(x[6359] ^ x[6360]);
     layer0_out[11388] <= x[4684] | x[4685];
     layer0_out[11389] <= x[4610] & x[4611];
     layer0_out[11390] <= 1'b0;
     layer0_out[11391] <= x[5150] & x[5151];
     layer0_out[11392] <= x[3095];
     layer0_out[11393] <= ~(x[5346] | x[5347]);
     layer0_out[11394] <= ~x[2455] | x[2457];
     layer0_out[11395] <= ~(x[2126] & x[2128]);
     layer0_out[11396] <= x[2288] & x[2289];
     layer0_out[11397] <= x[4457] ^ x[4458];
     layer0_out[11398] <= ~x[3075];
     layer0_out[11399] <= ~(x[1458] & x[1460]);
     layer0_out[11400] <= x[2652] & ~x[2650];
     layer0_out[11401] <= ~(x[2182] & x[2184]);
     layer0_out[11402] <= x[5481] & ~x[5482];
     layer0_out[11403] <= ~(x[2262] & x[2263]);
     layer0_out[11404] <= ~x[2401];
     layer0_out[11405] <= ~(x[1276] & x[1277]);
     layer0_out[11406] <= ~(x[104] | x[105]);
     layer0_out[11407] <= ~x[7260];
     layer0_out[11408] <= ~(x[7969] & x[7970]);
     layer0_out[11409] <= ~(x[668] | x[670]);
     layer0_out[11410] <= x[7811];
     layer0_out[11411] <= ~(x[2415] & x[2417]);
     layer0_out[11412] <= ~(x[7377] | x[7378]);
     layer0_out[11413] <= x[1589] | x[1591];
     layer0_out[11414] <= ~(x[5858] ^ x[5859]);
     layer0_out[11415] <= ~(x[1743] & x[1745]);
     layer0_out[11416] <= x[857];
     layer0_out[11417] <= x[1223];
     layer0_out[11418] <= x[1108] | x[1110];
     layer0_out[11419] <= x[1839] & x[1841];
     layer0_out[11420] <= ~(x[292] & x[293]);
     layer0_out[11421] <= x[146] & x[147];
     layer0_out[11422] <= ~(x[4714] ^ x[4715]);
     layer0_out[11423] <= ~x[1576];
     layer0_out[11424] <= x[6205] & ~x[6204];
     layer0_out[11425] <= ~(x[2547] & x[2548]);
     layer0_out[11426] <= x[3950] & ~x[3949];
     layer0_out[11427] <= x[2339] & ~x[2337];
     layer0_out[11428] <= ~(x[1454] & x[1456]);
     layer0_out[11429] <= ~(x[1376] & x[1377]);
     layer0_out[11430] <= x[2670] & x[2671];
     layer0_out[11431] <= ~(x[5276] & x[5277]);
     layer0_out[11432] <= x[8761] | x[8762];
     layer0_out[11433] <= ~(x[6735] | x[6736]);
     layer0_out[11434] <= x[6488];
     layer0_out[11435] <= ~x[2046] | x[2048];
     layer0_out[11436] <= x[5889] & x[5890];
     layer0_out[11437] <= 1'b0;
     layer0_out[11438] <= x[3907];
     layer0_out[11439] <= ~(x[289] & x[290]);
     layer0_out[11440] <= x[5774] & ~x[5773];
     layer0_out[11441] <= ~(x[4858] & x[4859]);
     layer0_out[11442] <= x[6920] | x[6921];
     layer0_out[11443] <= x[1297] & x[1299];
     layer0_out[11444] <= ~x[7657];
     layer0_out[11445] <= x[3662];
     layer0_out[11446] <= ~(x[2435] & x[2436]);
     layer0_out[11447] <= ~x[2222];
     layer0_out[11448] <= ~(x[487] ^ x[489]);
     layer0_out[11449] <= ~(x[6917] & x[6918]);
     layer0_out[11450] <= ~x[8466];
     layer0_out[11451] <= x[7391] | x[7392];
     layer0_out[11452] <= ~x[8145] | x[8146];
     layer0_out[11453] <= ~(x[5954] | x[5955]);
     layer0_out[11454] <= x[7362] & ~x[7361];
     layer0_out[11455] <= x[1326] & x[1328];
     layer0_out[11456] <= x[1026] & x[1028];
     layer0_out[11457] <= ~x[1541] | x[1542];
     layer0_out[11458] <= x[3987] | x[3988];
     layer0_out[11459] <= ~x[3489] | x[3490];
     layer0_out[11460] <= x[4907];
     layer0_out[11461] <= ~x[4195];
     layer0_out[11462] <= x[4208];
     layer0_out[11463] <= ~(x[1800] & x[1802]);
     layer0_out[11464] <= x[1639] & x[1640];
     layer0_out[11465] <= ~x[74];
     layer0_out[11466] <= ~(x[2773] | x[2774]);
     layer0_out[11467] <= x[3396] ^ x[3397];
     layer0_out[11468] <= x[4337] & x[4338];
     layer0_out[11469] <= ~(x[192] & x[193]);
     layer0_out[11470] <= 1'b0;
     layer0_out[11471] <= x[5418] & x[5419];
     layer0_out[11472] <= ~(x[5865] & x[5866]);
     layer0_out[11473] <= ~(x[7365] & x[7366]);
     layer0_out[11474] <= x[9098] ^ x[9099];
     layer0_out[11475] <= ~(x[3330] | x[3331]);
     layer0_out[11476] <= ~(x[2686] ^ x[2687]);
     layer0_out[11477] <= x[3243] & ~x[3244];
     layer0_out[11478] <= x[145];
     layer0_out[11479] <= ~x[2131];
     layer0_out[11480] <= x[6229] & ~x[6228];
     layer0_out[11481] <= 1'b1;
     layer0_out[11482] <= ~x[8491];
     layer0_out[11483] <= ~(x[492] ^ x[494]);
     layer0_out[11484] <= x[1556] & x[1557];
     layer0_out[11485] <= ~(x[6512] ^ x[6513]);
     layer0_out[11486] <= ~(x[5308] & x[5309]);
     layer0_out[11487] <= 1'b0;
     layer0_out[11488] <= ~x[3734];
     layer0_out[11489] <= ~(x[2438] & x[2439]);
     layer0_out[11490] <= x[221] ^ x[222];
     layer0_out[11491] <= x[9017] & ~x[9016];
     layer0_out[11492] <= x[6630];
     layer0_out[11493] <= x[1676] ^ x[1678];
     layer0_out[11494] <= x[3985] | x[3986];
     layer0_out[11495] <= ~(x[1600] | x[1602]);
     layer0_out[11496] <= x[7663] & x[7664];
     layer0_out[11497] <= ~(x[8554] | x[8555]);
     layer0_out[11498] <= 1'b1;
     layer0_out[11499] <= ~x[1516];
     layer0_out[11500] <= ~(x[2573] | x[2574]);
     layer0_out[11501] <= x[4961] & ~x[4960];
     layer0_out[11502] <= ~x[1096] | x[1098];
     layer0_out[11503] <= ~(x[7011] ^ x[7012]);
     layer0_out[11504] <= x[1] ^ x[2];
     layer0_out[11505] <= x[6830];
     layer0_out[11506] <= ~x[5610];
     layer0_out[11507] <= x[7390] ^ x[7391];
     layer0_out[11508] <= ~(x[1535] & x[1537]);
     layer0_out[11509] <= x[1275];
     layer0_out[11510] <= x[1803] & x[1804];
     layer0_out[11511] <= ~(x[2108] & x[2110]);
     layer0_out[11512] <= ~(x[2441] | x[2443]);
     layer0_out[11513] <= x[8711] | x[8712];
     layer0_out[11514] <= x[7293] ^ x[7294];
     layer0_out[11515] <= x[2118] & x[2119];
     layer0_out[11516] <= x[545] ^ x[547];
     layer0_out[11517] <= x[1099] & x[1100];
     layer0_out[11518] <= ~(x[4180] ^ x[4181]);
     layer0_out[11519] <= ~(x[1565] & x[1567]);
     layer0_out[11520] <= x[7334] ^ x[7335];
     layer0_out[11521] <= ~(x[1154] ^ x[1156]);
     layer0_out[11522] <= ~(x[499] ^ x[501]);
     layer0_out[11523] <= ~(x[5468] & x[5469]);
     layer0_out[11524] <= x[1240];
     layer0_out[11525] <= ~(x[1862] & x[1864]);
     layer0_out[11526] <= x[2598];
     layer0_out[11527] <= 1'b0;
     layer0_out[11528] <= ~x[1541] | x[1539];
     layer0_out[11529] <= x[238] & x[239];
     layer0_out[11530] <= 1'b0;
     layer0_out[11531] <= x[8379] & x[8380];
     layer0_out[11532] <= x[4093] ^ x[4094];
     layer0_out[11533] <= x[7878] | x[7879];
     layer0_out[11534] <= x[2009] | x[2011];
     layer0_out[11535] <= x[8667] | x[8668];
     layer0_out[11536] <= x[5320] & x[5321];
     layer0_out[11537] <= ~x[3334] | x[3335];
     layer0_out[11538] <= x[485] & x[487];
     layer0_out[11539] <= ~(x[8396] & x[8397]);
     layer0_out[11540] <= x[5872] & x[5873];
     layer0_out[11541] <= ~(x[6423] | x[6424]);
     layer0_out[11542] <= x[472];
     layer0_out[11543] <= x[3561];
     layer0_out[11544] <= x[5437] & ~x[5436];
     layer0_out[11545] <= x[6106] | x[6107];
     layer0_out[11546] <= x[1343] & x[1344];
     layer0_out[11547] <= x[4688] & x[4689];
     layer0_out[11548] <= x[923] ^ x[924];
     layer0_out[11549] <= x[2206] & x[2208];
     layer0_out[11550] <= ~(x[7284] ^ x[7285]);
     layer0_out[11551] <= x[4868];
     layer0_out[11552] <= ~(x[177] & x[179]);
     layer0_out[11553] <= ~(x[7533] & x[7534]);
     layer0_out[11554] <= x[2233] & ~x[2235];
     layer0_out[11555] <= ~(x[5080] | x[5081]);
     layer0_out[11556] <= ~x[1588] | x[1587];
     layer0_out[11557] <= ~(x[3069] ^ x[3070]);
     layer0_out[11558] <= x[1916] & x[1917];
     layer0_out[11559] <= x[8004] & ~x[8005];
     layer0_out[11560] <= ~(x[5033] | x[5034]);
     layer0_out[11561] <= 1'b1;
     layer0_out[11562] <= x[2791] ^ x[2792];
     layer0_out[11563] <= ~x[6269];
     layer0_out[11564] <= x[3162] | x[3163];
     layer0_out[11565] <= ~x[6999];
     layer0_out[11566] <= x[5895] | x[5896];
     layer0_out[11567] <= ~(x[1595] & x[1596]);
     layer0_out[11568] <= x[8741];
     layer0_out[11569] <= ~(x[7692] & x[7693]);
     layer0_out[11570] <= x[1470] & x[1471];
     layer0_out[11571] <= ~(x[1533] & x[1535]);
     layer0_out[11572] <= x[6951] & x[6952];
     layer0_out[11573] <= x[3686] ^ x[3687];
     layer0_out[11574] <= ~(x[2905] & x[2906]);
     layer0_out[11575] <= x[5938] & x[5939];
     layer0_out[11576] <= x[5017] | x[5018];
     layer0_out[11577] <= 1'b0;
     layer0_out[11578] <= x[8086] ^ x[8087];
     layer0_out[11579] <= ~(x[1290] ^ x[1292]);
     layer0_out[11580] <= x[5120];
     layer0_out[11581] <= 1'b1;
     layer0_out[11582] <= x[369] & x[371];
     layer0_out[11583] <= ~(x[7608] & x[7609]);
     layer0_out[11584] <= ~(x[1792] & x[1794]);
     layer0_out[11585] <= ~(x[8593] | x[8594]);
     layer0_out[11586] <= ~x[8032];
     layer0_out[11587] <= ~x[8864];
     layer0_out[11588] <= ~(x[8259] | x[8260]);
     layer0_out[11589] <= ~x[8323];
     layer0_out[11590] <= ~(x[7623] & x[7624]);
     layer0_out[11591] <= ~(x[7331] | x[7332]);
     layer0_out[11592] <= x[1788];
     layer0_out[11593] <= x[3412];
     layer0_out[11594] <= x[567] ^ x[569];
     layer0_out[11595] <= x[6356];
     layer0_out[11596] <= ~(x[7863] | x[7864]);
     layer0_out[11597] <= x[2603] & x[2604];
     layer0_out[11598] <= x[1594] & x[1595];
     layer0_out[11599] <= ~(x[12] ^ x[14]);
     layer0_out[11600] <= ~(x[2858] & x[2859]);
     layer0_out[11601] <= x[1736] & x[1737];
     layer0_out[11602] <= x[3409] | x[3410];
     layer0_out[11603] <= ~(x[6146] | x[6147]);
     layer0_out[11604] <= x[1233] & x[1234];
     layer0_out[11605] <= ~x[15];
     layer0_out[11606] <= x[7568] | x[7569];
     layer0_out[11607] <= ~(x[9206] | x[9207]);
     layer0_out[11608] <= x[5350];
     layer0_out[11609] <= x[405] ^ x[407];
     layer0_out[11610] <= ~(x[4122] & x[4123]);
     layer0_out[11611] <= ~x[7733];
     layer0_out[11612] <= ~x[6530];
     layer0_out[11613] <= x[379] & x[380];
     layer0_out[11614] <= ~x[867];
     layer0_out[11615] <= x[164];
     layer0_out[11616] <= x[7914] | x[7915];
     layer0_out[11617] <= ~(x[8034] | x[8035]);
     layer0_out[11618] <= x[1782] & x[1784];
     layer0_out[11619] <= ~(x[1801] ^ x[1803]);
     layer0_out[11620] <= x[6909] | x[6910];
     layer0_out[11621] <= x[2532] ^ x[2533];
     layer0_out[11622] <= ~(x[5780] | x[5781]);
     layer0_out[11623] <= x[6676] | x[6677];
     layer0_out[11624] <= x[2653] | x[2655];
     layer0_out[11625] <= x[975] & x[977];
     layer0_out[11626] <= x[7092] | x[7093];
     layer0_out[11627] <= x[2360] & ~x[2359];
     layer0_out[11628] <= ~x[525];
     layer0_out[11629] <= x[1499] & x[1501];
     layer0_out[11630] <= ~(x[8581] | x[8582]);
     layer0_out[11631] <= x[594] & ~x[596];
     layer0_out[11632] <= x[2772] & ~x[2770];
     layer0_out[11633] <= x[3023] | x[3024];
     layer0_out[11634] <= x[1348] ^ x[1350];
     layer0_out[11635] <= ~(x[5300] | x[5301]);
     layer0_out[11636] <= ~x[6581];
     layer0_out[11637] <= 1'b0;
     layer0_out[11638] <= x[4528] & x[4529];
     layer0_out[11639] <= 1'b0;
     layer0_out[11640] <= ~x[8716];
     layer0_out[11641] <= ~(x[6198] | x[6199]);
     layer0_out[11642] <= 1'b1;
     layer0_out[11643] <= ~(x[359] | x[360]);
     layer0_out[11644] <= ~(x[8472] | x[8473]);
     layer0_out[11645] <= x[2785] & ~x[2786];
     layer0_out[11646] <= x[900] | x[901];
     layer0_out[11647] <= x[4399] | x[4400];
     layer0_out[11648] <= x[3917] & ~x[3918];
     layer0_out[11649] <= x[5535];
     layer0_out[11650] <= ~x[6174];
     layer0_out[11651] <= x[4808] | x[4809];
     layer0_out[11652] <= ~(x[854] & x[856]);
     layer0_out[11653] <= 1'b0;
     layer0_out[11654] <= ~x[2318];
     layer0_out[11655] <= x[8482] & x[8483];
     layer0_out[11656] <= ~x[7422] | x[7423];
     layer0_out[11657] <= x[1582];
     layer0_out[11658] <= x[3151] | x[3152];
     layer0_out[11659] <= x[4022] ^ x[4023];
     layer0_out[11660] <= ~(x[699] | x[700]);
     layer0_out[11661] <= 1'b0;
     layer0_out[11662] <= x[1561] & ~x[1559];
     layer0_out[11663] <= ~(x[3110] & x[3111]);
     layer0_out[11664] <= x[3344];
     layer0_out[11665] <= 1'b1;
     layer0_out[11666] <= ~(x[4218] ^ x[4219]);
     layer0_out[11667] <= x[6763] & ~x[6762];
     layer0_out[11668] <= ~(x[4930] | x[4931]);
     layer0_out[11669] <= x[2711];
     layer0_out[11670] <= ~x[145] | x[144];
     layer0_out[11671] <= x[6034] & x[6035];
     layer0_out[11672] <= x[2312] | x[2313];
     layer0_out[11673] <= x[1199] & x[1200];
     layer0_out[11674] <= ~(x[9134] | x[9135]);
     layer0_out[11675] <= x[1140] & x[1142];
     layer0_out[11676] <= x[1466] | x[1468];
     layer0_out[11677] <= x[224] & ~x[222];
     layer0_out[11678] <= 1'b0;
     layer0_out[11679] <= ~(x[211] & x[212]);
     layer0_out[11680] <= ~x[5374];
     layer0_out[11681] <= x[845] | x[846];
     layer0_out[11682] <= x[852] ^ x[853];
     layer0_out[11683] <= ~(x[55] ^ x[57]);
     layer0_out[11684] <= x[3092] & x[3093];
     layer0_out[11685] <= x[2443];
     layer0_out[11686] <= x[2850] & x[2851];
     layer0_out[11687] <= x[1410];
     layer0_out[11688] <= ~(x[2387] & x[2388]);
     layer0_out[11689] <= x[1047];
     layer0_out[11690] <= ~x[1409] | x[1408];
     layer0_out[11691] <= ~x[8746] | x[8747];
     layer0_out[11692] <= 1'b1;
     layer0_out[11693] <= x[9070] | x[9071];
     layer0_out[11694] <= ~(x[4336] & x[4337]);
     layer0_out[11695] <= ~(x[1423] & x[1424]);
     layer0_out[11696] <= ~(x[999] ^ x[1000]);
     layer0_out[11697] <= x[2454] & x[2455];
     layer0_out[11698] <= x[2556] | x[2558];
     layer0_out[11699] <= ~x[1307] | x[1308];
     layer0_out[11700] <= x[3596] | x[3597];
     layer0_out[11701] <= x[5274] | x[5275];
     layer0_out[11702] <= x[2582] ^ x[2583];
     layer0_out[11703] <= ~(x[5751] & x[5752]);
     layer0_out[11704] <= x[1278];
     layer0_out[11705] <= x[1372] & ~x[1370];
     layer0_out[11706] <= ~x[3102];
     layer0_out[11707] <= ~(x[2372] & x[2374]);
     layer0_out[11708] <= x[9145] ^ x[9146];
     layer0_out[11709] <= x[1707] | x[1708];
     layer0_out[11710] <= 1'b0;
     layer0_out[11711] <= x[2638] & x[2639];
     layer0_out[11712] <= x[7270] ^ x[7271];
     layer0_out[11713] <= ~(x[2493] ^ x[2495]);
     layer0_out[11714] <= x[7393];
     layer0_out[11715] <= ~(x[195] | x[197]);
     layer0_out[11716] <= ~(x[5343] & x[5344]);
     layer0_out[11717] <= ~x[2726] | x[2724];
     layer0_out[11718] <= ~(x[4313] ^ x[4314]);
     layer0_out[11719] <= x[9210] | x[9211];
     layer0_out[11720] <= ~(x[3403] & x[3404]);
     layer0_out[11721] <= x[1328];
     layer0_out[11722] <= x[2097] & ~x[2096];
     layer0_out[11723] <= ~(x[2331] & x[2332]);
     layer0_out[11724] <= x[4975];
     layer0_out[11725] <= ~(x[556] & x[558]);
     layer0_out[11726] <= x[204];
     layer0_out[11727] <= ~x[7518] | x[7519];
     layer0_out[11728] <= x[2488] & x[2489];
     layer0_out[11729] <= 1'b1;
     layer0_out[11730] <= x[8662];
     layer0_out[11731] <= ~x[1492];
     layer0_out[11732] <= ~(x[8428] ^ x[8429]);
     layer0_out[11733] <= ~(x[284] ^ x[285]);
     layer0_out[11734] <= ~(x[2844] & x[2845]);
     layer0_out[11735] <= ~(x[5015] ^ x[5016]);
     layer0_out[11736] <= x[984] & x[986];
     layer0_out[11737] <= x[2220] | x[2222];
     layer0_out[11738] <= x[1899] & x[1901];
     layer0_out[11739] <= ~x[464];
     layer0_out[11740] <= ~x[119];
     layer0_out[11741] <= x[5237] & x[5238];
     layer0_out[11742] <= ~(x[5903] & x[5904]);
     layer0_out[11743] <= x[8091] | x[8092];
     layer0_out[11744] <= x[50];
     layer0_out[11745] <= ~(x[1701] ^ x[1703]);
     layer0_out[11746] <= ~x[1404] | x[1405];
     layer0_out[11747] <= x[380] & ~x[378];
     layer0_out[11748] <= ~(x[1834] & x[1836]);
     layer0_out[11749] <= ~x[3675];
     layer0_out[11750] <= x[3928];
     layer0_out[11751] <= ~(x[2592] & x[2594]);
     layer0_out[11752] <= ~(x[3201] | x[3202]);
     layer0_out[11753] <= ~(x[5943] ^ x[5944]);
     layer0_out[11754] <= x[1766] & x[1768];
     layer0_out[11755] <= ~x[3423];
     layer0_out[11756] <= ~x[546];
     layer0_out[11757] <= ~(x[1516] & x[1518]);
     layer0_out[11758] <= x[1152];
     layer0_out[11759] <= ~(x[3043] ^ x[3044]);
     layer0_out[11760] <= ~(x[7856] | x[7857]);
     layer0_out[11761] <= ~x[349] | x[350];
     layer0_out[11762] <= ~(x[2476] ^ x[2478]);
     layer0_out[11763] <= x[616] | x[617];
     layer0_out[11764] <= ~x[5053];
     layer0_out[11765] <= ~(x[7060] | x[7061]);
     layer0_out[11766] <= x[2058] & x[2060];
     layer0_out[11767] <= x[2634] ^ x[2636];
     layer0_out[11768] <= x[4894] | x[4895];
     layer0_out[11769] <= 1'b0;
     layer0_out[11770] <= ~(x[8653] | x[8654]);
     layer0_out[11771] <= ~(x[1855] ^ x[1857]);
     layer0_out[11772] <= x[5667] ^ x[5668];
     layer0_out[11773] <= 1'b1;
     layer0_out[11774] <= ~(x[1565] | x[1566]);
     layer0_out[11775] <= ~(x[3170] & x[3171]);
     layer0_out[11776] <= ~(x[6345] | x[6346]);
     layer0_out[11777] <= 1'b1;
     layer0_out[11778] <= ~(x[87] ^ x[89]);
     layer0_out[11779] <= x[1538];
     layer0_out[11780] <= x[7634] ^ x[7635];
     layer0_out[11781] <= ~(x[3054] & x[3055]);
     layer0_out[11782] <= ~(x[57] ^ x[59]);
     layer0_out[11783] <= x[1857] & ~x[1859];
     layer0_out[11784] <= ~(x[4743] ^ x[4744]);
     layer0_out[11785] <= x[5100] & ~x[5099];
     layer0_out[11786] <= x[963] | x[964];
     layer0_out[11787] <= ~(x[2302] | x[2303]);
     layer0_out[11788] <= x[7645];
     layer0_out[11789] <= x[1413] & x[1415];
     layer0_out[11790] <= ~(x[7792] & x[7793]);
     layer0_out[11791] <= ~(x[1260] & x[1261]);
     layer0_out[11792] <= ~(x[3486] ^ x[3487]);
     layer0_out[11793] <= x[7641] ^ x[7642];
     layer0_out[11794] <= x[7107] & x[7108];
     layer0_out[11795] <= ~(x[4229] & x[4230]);
     layer0_out[11796] <= ~(x[262] ^ x[264]);
     layer0_out[11797] <= x[2021] & x[2023];
     layer0_out[11798] <= x[2563] ^ x[2565];
     layer0_out[11799] <= ~(x[4381] ^ x[4382]);
     layer0_out[11800] <= ~x[324] | x[323];
     layer0_out[11801] <= x[3406] | x[3407];
     layer0_out[11802] <= ~(x[6610] ^ x[6611]);
     layer0_out[11803] <= ~x[865];
     layer0_out[11804] <= ~x[2693];
     layer0_out[11805] <= x[2776] & x[2777];
     layer0_out[11806] <= x[3733] | x[3734];
     layer0_out[11807] <= x[1766] | x[1767];
     layer0_out[11808] <= x[1818] & ~x[1816];
     layer0_out[11809] <= ~x[2976];
     layer0_out[11810] <= ~x[8539] | x[8538];
     layer0_out[11811] <= x[2276] & ~x[2278];
     layer0_out[11812] <= x[5303];
     layer0_out[11813] <= x[8405] & ~x[8406];
     layer0_out[11814] <= x[2561] ^ x[2563];
     layer0_out[11815] <= x[8638] ^ x[8639];
     layer0_out[11816] <= x[983] | x[985];
     layer0_out[11817] <= x[1515];
     layer0_out[11818] <= ~x[7623];
     layer0_out[11819] <= ~x[3208];
     layer0_out[11820] <= ~x[1296] | x[1297];
     layer0_out[11821] <= ~x[68];
     layer0_out[11822] <= ~(x[1396] & x[1397]);
     layer0_out[11823] <= x[6333] & ~x[6332];
     layer0_out[11824] <= x[1065] & x[1067];
     layer0_out[11825] <= ~(x[2316] & x[2317]);
     layer0_out[11826] <= ~(x[2264] | x[2266]);
     layer0_out[11827] <= 1'b1;
     layer0_out[11828] <= x[4331];
     layer0_out[11829] <= x[1002] | x[1003];
     layer0_out[11830] <= ~(x[3641] & x[3642]);
     layer0_out[11831] <= x[2641] ^ x[2643];
     layer0_out[11832] <= ~(x[5904] & x[5905]);
     layer0_out[11833] <= ~(x[5975] & x[5976]);
     layer0_out[11834] <= ~x[4639] | x[4640];
     layer0_out[11835] <= ~(x[8297] & x[8298]);
     layer0_out[11836] <= ~x[7228] | x[7229];
     layer0_out[11837] <= x[7998] | x[7999];
     layer0_out[11838] <= ~x[6661];
     layer0_out[11839] <= ~(x[5561] & x[5562]);
     layer0_out[11840] <= ~x[8570] | x[8571];
     layer0_out[11841] <= x[8346] ^ x[8347];
     layer0_out[11842] <= x[6454] & x[6455];
     layer0_out[11843] <= ~x[692];
     layer0_out[11844] <= ~(x[856] & x[858]);
     layer0_out[11845] <= x[2053] & x[2055];
     layer0_out[11846] <= 1'b0;
     layer0_out[11847] <= ~x[5249];
     layer0_out[11848] <= x[6519] | x[6520];
     layer0_out[11849] <= 1'b1;
     layer0_out[11850] <= x[3824] | x[3825];
     layer0_out[11851] <= x[2583];
     layer0_out[11852] <= ~x[3246];
     layer0_out[11853] <= x[7354];
     layer0_out[11854] <= ~x[3191];
     layer0_out[11855] <= x[4646] & x[4647];
     layer0_out[11856] <= x[726] ^ x[727];
     layer0_out[11857] <= x[1257];
     layer0_out[11858] <= ~(x[3772] & x[3773]);
     layer0_out[11859] <= x[5531] | x[5532];
     layer0_out[11860] <= 1'b1;
     layer0_out[11861] <= x[8408] & x[8409];
     layer0_out[11862] <= x[543] ^ x[545];
     layer0_out[11863] <= ~x[1216];
     layer0_out[11864] <= ~x[587];
     layer0_out[11865] <= x[2000] & ~x[2001];
     layer0_out[11866] <= x[6413] ^ x[6414];
     layer0_out[11867] <= ~(x[2128] & x[2130]);
     layer0_out[11868] <= x[148] | x[149];
     layer0_out[11869] <= x[985];
     layer0_out[11870] <= x[5763] & x[5764];
     layer0_out[11871] <= x[8634] & ~x[8633];
     layer0_out[11872] <= ~x[4193];
     layer0_out[11873] <= x[275] & x[277];
     layer0_out[11874] <= ~(x[3103] & x[3104]);
     layer0_out[11875] <= ~(x[3848] | x[3849]);
     layer0_out[11876] <= ~(x[7127] | x[7128]);
     layer0_out[11877] <= ~x[1738];
     layer0_out[11878] <= ~(x[2606] & x[2608]);
     layer0_out[11879] <= ~(x[329] ^ x[330]);
     layer0_out[11880] <= x[2005] | x[2006];
     layer0_out[11881] <= ~(x[6637] & x[6638]);
     layer0_out[11882] <= 1'b1;
     layer0_out[11883] <= x[2289] ^ x[2291];
     layer0_out[11884] <= ~(x[785] ^ x[786]);
     layer0_out[11885] <= ~(x[7804] & x[7805]);
     layer0_out[11886] <= ~(x[921] ^ x[923]);
     layer0_out[11887] <= x[2069] | x[2071];
     layer0_out[11888] <= x[348] ^ x[349];
     layer0_out[11889] <= ~(x[893] | x[895]);
     layer0_out[11890] <= ~x[2310];
     layer0_out[11891] <= ~(x[1644] & x[1645]);
     layer0_out[11892] <= ~(x[1845] & x[1847]);
     layer0_out[11893] <= x[7605] | x[7606];
     layer0_out[11894] <= x[7983] | x[7984];
     layer0_out[11895] <= x[8007] | x[8008];
     layer0_out[11896] <= x[6690];
     layer0_out[11897] <= x[8649] | x[8650];
     layer0_out[11898] <= x[5325] & x[5326];
     layer0_out[11899] <= ~x[3808];
     layer0_out[11900] <= ~(x[2769] & x[2770]);
     layer0_out[11901] <= x[702] ^ x[703];
     layer0_out[11902] <= ~(x[2517] & x[2519]);
     layer0_out[11903] <= x[5005];
     layer0_out[11904] <= ~(x[2713] & x[2714]);
     layer0_out[11905] <= 1'b0;
     layer0_out[11906] <= ~x[5856];
     layer0_out[11907] <= x[688] & x[690];
     layer0_out[11908] <= ~x[4494];
     layer0_out[11909] <= ~(x[3061] ^ x[3062]);
     layer0_out[11910] <= ~(x[5408] & x[5409]);
     layer0_out[11911] <= ~x[948] | x[950];
     layer0_out[11912] <= ~x[7331];
     layer0_out[11913] <= ~(x[4297] & x[4298]);
     layer0_out[11914] <= x[3714] & x[3715];
     layer0_out[11915] <= x[1464];
     layer0_out[11916] <= ~(x[5212] & x[5213]);
     layer0_out[11917] <= ~x[1221];
     layer0_out[11918] <= ~(x[8305] & x[8306]);
     layer0_out[11919] <= x[4426] & x[4427];
     layer0_out[11920] <= x[7845] ^ x[7846];
     layer0_out[11921] <= ~x[6617] | x[6618];
     layer0_out[11922] <= x[7132] ^ x[7133];
     layer0_out[11923] <= x[449] & x[450];
     layer0_out[11924] <= x[5951] ^ x[5952];
     layer0_out[11925] <= x[2120] & x[2122];
     layer0_out[11926] <= ~(x[3226] | x[3227]);
     layer0_out[11927] <= ~x[2485] | x[2487];
     layer0_out[11928] <= x[1147];
     layer0_out[11929] <= x[947];
     layer0_out[11930] <= x[1685] & x[1687];
     layer0_out[11931] <= x[5816] & x[5817];
     layer0_out[11932] <= ~x[2886];
     layer0_out[11933] <= x[3640] | x[3641];
     layer0_out[11934] <= ~x[4765];
     layer0_out[11935] <= ~x[4683];
     layer0_out[11936] <= ~x[6691] | x[6692];
     layer0_out[11937] <= x[7478] | x[7479];
     layer0_out[11938] <= x[6808] & x[6809];
     layer0_out[11939] <= x[544] | x[545];
     layer0_out[11940] <= ~x[2059];
     layer0_out[11941] <= ~(x[612] & x[613]);
     layer0_out[11942] <= ~(x[7164] | x[7165]);
     layer0_out[11943] <= x[582] ^ x[583];
     layer0_out[11944] <= x[6201] | x[6202];
     layer0_out[11945] <= ~(x[3015] & x[3016]);
     layer0_out[11946] <= ~(x[566] & x[567]);
     layer0_out[11947] <= x[1266] & x[1267];
     layer0_out[11948] <= 1'b0;
     layer0_out[11949] <= ~x[6731] | x[6732];
     layer0_out[11950] <= x[1458] & x[1459];
     layer0_out[11951] <= 1'b0;
     layer0_out[11952] <= ~(x[1614] & x[1616]);
     layer0_out[11953] <= x[2556] & x[2557];
     layer0_out[11954] <= ~x[4132];
     layer0_out[11955] <= x[5553] & x[5554];
     layer0_out[11956] <= ~(x[5330] & x[5331]);
     layer0_out[11957] <= ~x[7652];
     layer0_out[11958] <= x[2054] & x[2056];
     layer0_out[11959] <= ~(x[1155] & x[1156]);
     layer0_out[11960] <= ~(x[2715] ^ x[2717]);
     layer0_out[11961] <= ~(x[2537] ^ x[2538]);
     layer0_out[11962] <= ~(x[3526] & x[3527]);
     layer0_out[11963] <= ~x[8792];
     layer0_out[11964] <= ~(x[5842] & x[5843]);
     layer0_out[11965] <= ~(x[9125] | x[9126]);
     layer0_out[11966] <= 1'b0;
     layer0_out[11967] <= ~(x[4239] & x[4240]);
     layer0_out[11968] <= x[5750] ^ x[5751];
     layer0_out[11969] <= x[4398];
     layer0_out[11970] <= x[6134];
     layer0_out[11971] <= x[332];
     layer0_out[11972] <= x[1061] & x[1063];
     layer0_out[11973] <= x[1202] & x[1203];
     layer0_out[11974] <= ~x[6203];
     layer0_out[11975] <= x[3827] & x[3828];
     layer0_out[11976] <= ~x[8441];
     layer0_out[11977] <= ~(x[4495] & x[4496]);
     layer0_out[11978] <= x[1987] & ~x[1988];
     layer0_out[11979] <= x[2812] | x[2813];
     layer0_out[11980] <= x[1959] & x[1961];
     layer0_out[11981] <= ~(x[6222] & x[6223]);
     layer0_out[11982] <= ~(x[522] | x[523]);
     layer0_out[11983] <= ~x[6048];
     layer0_out[11984] <= x[409];
     layer0_out[11985] <= ~x[5544];
     layer0_out[11986] <= ~(x[1302] ^ x[1304]);
     layer0_out[11987] <= ~x[2439] | x[2437];
     layer0_out[11988] <= ~x[9130];
     layer0_out[11989] <= x[9116] ^ x[9117];
     layer0_out[11990] <= ~x[8715];
     layer0_out[11991] <= ~(x[7481] | x[7482]);
     layer0_out[11992] <= ~(x[2105] | x[2107]);
     layer0_out[11993] <= x[5160];
     layer0_out[11994] <= 1'b0;
     layer0_out[11995] <= x[3896] | x[3897];
     layer0_out[11996] <= x[1912];
     layer0_out[11997] <= x[3083] & x[3084];
     layer0_out[11998] <= ~x[563];
     layer0_out[11999] <= 1'b0;
     layer1_out[0] <= ~layer0_out[7185];
     layer1_out[1] <= 1'b0;
     layer1_out[2] <= ~layer0_out[9645];
     layer1_out[3] <= ~layer0_out[6018];
     layer1_out[4] <= ~(layer0_out[3173] | layer0_out[3174]);
     layer1_out[5] <= layer0_out[3540];
     layer1_out[6] <= ~layer0_out[5348] | layer0_out[5347];
     layer1_out[7] <= ~layer0_out[145] | layer0_out[144];
     layer1_out[8] <= ~layer0_out[5864] | layer0_out[5863];
     layer1_out[9] <= layer0_out[1581] & layer0_out[1582];
     layer1_out[10] <= ~layer0_out[3197] | layer0_out[3196];
     layer1_out[11] <= ~layer0_out[4462] | layer0_out[4463];
     layer1_out[12] <= layer0_out[10492] ^ layer0_out[10493];
     layer1_out[13] <= ~(layer0_out[7072] & layer0_out[7073]);
     layer1_out[14] <= 1'b0;
     layer1_out[15] <= ~layer0_out[320];
     layer1_out[16] <= layer0_out[6506] | layer0_out[6507];
     layer1_out[17] <= layer0_out[10377] | layer0_out[10378];
     layer1_out[18] <= ~(layer0_out[10358] ^ layer0_out[10359]);
     layer1_out[19] <= ~layer0_out[1232] | layer0_out[1231];
     layer1_out[20] <= layer0_out[2994];
     layer1_out[21] <= ~layer0_out[11850];
     layer1_out[22] <= ~layer0_out[6676];
     layer1_out[23] <= ~layer0_out[10827];
     layer1_out[24] <= ~layer0_out[4256];
     layer1_out[25] <= ~layer0_out[8919] | layer0_out[8918];
     layer1_out[26] <= layer0_out[4688] | layer0_out[4689];
     layer1_out[27] <= ~layer0_out[1927] | layer0_out[1926];
     layer1_out[28] <= ~layer0_out[5106] | layer0_out[5105];
     layer1_out[29] <= 1'b0;
     layer1_out[30] <= layer0_out[928] & ~layer0_out[927];
     layer1_out[31] <= ~(layer0_out[4574] | layer0_out[4575]);
     layer1_out[32] <= layer0_out[7240] | layer0_out[7241];
     layer1_out[33] <= layer0_out[3659] & ~layer0_out[3660];
     layer1_out[34] <= ~layer0_out[9359] | layer0_out[9360];
     layer1_out[35] <= ~(layer0_out[1956] ^ layer0_out[1957]);
     layer1_out[36] <= layer0_out[720];
     layer1_out[37] <= ~layer0_out[5625];
     layer1_out[38] <= ~layer0_out[1084];
     layer1_out[39] <= layer0_out[11547];
     layer1_out[40] <= ~layer0_out[1459] | layer0_out[1458];
     layer1_out[41] <= layer0_out[5738] & layer0_out[5739];
     layer1_out[42] <= layer0_out[1127];
     layer1_out[43] <= layer0_out[5888];
     layer1_out[44] <= ~layer0_out[4384] | layer0_out[4385];
     layer1_out[45] <= ~(layer0_out[9176] | layer0_out[9177]);
     layer1_out[46] <= layer0_out[2552] | layer0_out[2553];
     layer1_out[47] <= ~layer0_out[2219];
     layer1_out[48] <= ~layer0_out[6371];
     layer1_out[49] <= ~layer0_out[583] | layer0_out[582];
     layer1_out[50] <= ~layer0_out[2249] | layer0_out[2250];
     layer1_out[51] <= layer0_out[7360];
     layer1_out[52] <= ~(layer0_out[6813] ^ layer0_out[6814]);
     layer1_out[53] <= ~layer0_out[1532];
     layer1_out[54] <= ~layer0_out[1860] | layer0_out[1861];
     layer1_out[55] <= layer0_out[8013];
     layer1_out[56] <= ~(layer0_out[1391] & layer0_out[1392]);
     layer1_out[57] <= ~(layer0_out[7909] | layer0_out[7910]);
     layer1_out[58] <= layer0_out[10445];
     layer1_out[59] <= ~layer0_out[10259];
     layer1_out[60] <= layer0_out[3877];
     layer1_out[61] <= ~(layer0_out[11866] & layer0_out[11867]);
     layer1_out[62] <= ~layer0_out[3081];
     layer1_out[63] <= ~layer0_out[10461] | layer0_out[10460];
     layer1_out[64] <= layer0_out[10200] | layer0_out[10201];
     layer1_out[65] <= layer0_out[6137] & ~layer0_out[6136];
     layer1_out[66] <= ~layer0_out[6318] | layer0_out[6319];
     layer1_out[67] <= ~layer0_out[11641];
     layer1_out[68] <= layer0_out[8805] | layer0_out[8806];
     layer1_out[69] <= ~layer0_out[5985];
     layer1_out[70] <= layer0_out[9753];
     layer1_out[71] <= ~(layer0_out[4424] & layer0_out[4425]);
     layer1_out[72] <= ~layer0_out[8715] | layer0_out[8714];
     layer1_out[73] <= ~layer0_out[10883] | layer0_out[10882];
     layer1_out[74] <= ~layer0_out[3035];
     layer1_out[75] <= layer0_out[2721] & layer0_out[2722];
     layer1_out[76] <= layer0_out[2234] & ~layer0_out[2235];
     layer1_out[77] <= layer0_out[11178] | layer0_out[11179];
     layer1_out[78] <= layer0_out[10273];
     layer1_out[79] <= layer0_out[1068];
     layer1_out[80] <= layer0_out[8560];
     layer1_out[81] <= ~(layer0_out[5743] & layer0_out[5744]);
     layer1_out[82] <= ~layer0_out[11959] | layer0_out[11960];
     layer1_out[83] <= layer0_out[3146] & ~layer0_out[3145];
     layer1_out[84] <= layer0_out[6957] ^ layer0_out[6958];
     layer1_out[85] <= ~(layer0_out[1645] ^ layer0_out[1646]);
     layer1_out[86] <= ~layer0_out[11476] | layer0_out[11477];
     layer1_out[87] <= layer0_out[525] ^ layer0_out[526];
     layer1_out[88] <= layer0_out[8491] | layer0_out[8492];
     layer1_out[89] <= layer0_out[4363] | layer0_out[4364];
     layer1_out[90] <= layer0_out[2980] & ~layer0_out[2979];
     layer1_out[91] <= ~(layer0_out[9340] | layer0_out[9341]);
     layer1_out[92] <= ~(layer0_out[3883] | layer0_out[3884]);
     layer1_out[93] <= layer0_out[7805] | layer0_out[7806];
     layer1_out[94] <= ~layer0_out[3029];
     layer1_out[95] <= layer0_out[4664] & ~layer0_out[4665];
     layer1_out[96] <= ~(layer0_out[44] & layer0_out[45]);
     layer1_out[97] <= ~layer0_out[6949];
     layer1_out[98] <= layer0_out[3182] ^ layer0_out[3183];
     layer1_out[99] <= ~(layer0_out[7903] & layer0_out[7904]);
     layer1_out[100] <= layer0_out[4218];
     layer1_out[101] <= ~(layer0_out[8854] | layer0_out[8855]);
     layer1_out[102] <= ~layer0_out[7760];
     layer1_out[103] <= layer0_out[5635] | layer0_out[5636];
     layer1_out[104] <= layer0_out[2924];
     layer1_out[105] <= layer0_out[7230];
     layer1_out[106] <= layer0_out[3933] & ~layer0_out[3932];
     layer1_out[107] <= layer0_out[8312] ^ layer0_out[8313];
     layer1_out[108] <= layer0_out[5846] ^ layer0_out[5847];
     layer1_out[109] <= layer0_out[10479] & layer0_out[10480];
     layer1_out[110] <= layer0_out[1358] & layer0_out[1359];
     layer1_out[111] <= ~(layer0_out[1354] & layer0_out[1355]);
     layer1_out[112] <= layer0_out[212] & ~layer0_out[213];
     layer1_out[113] <= layer0_out[954] & ~layer0_out[955];
     layer1_out[114] <= 1'b1;
     layer1_out[115] <= ~layer0_out[8428];
     layer1_out[116] <= ~layer0_out[7914];
     layer1_out[117] <= layer0_out[1089] & ~layer0_out[1090];
     layer1_out[118] <= ~(layer0_out[8586] | layer0_out[8587]);
     layer1_out[119] <= 1'b1;
     layer1_out[120] <= layer0_out[1000] & ~layer0_out[999];
     layer1_out[121] <= 1'b0;
     layer1_out[122] <= layer0_out[5264] & ~layer0_out[5263];
     layer1_out[123] <= layer0_out[9455];
     layer1_out[124] <= ~layer0_out[6153];
     layer1_out[125] <= layer0_out[11956];
     layer1_out[126] <= layer0_out[4192];
     layer1_out[127] <= layer0_out[4757];
     layer1_out[128] <= 1'b1;
     layer1_out[129] <= ~layer0_out[1876] | layer0_out[1877];
     layer1_out[130] <= layer0_out[10250] & ~layer0_out[10251];
     layer1_out[131] <= ~layer0_out[9712] | layer0_out[9711];
     layer1_out[132] <= 1'b0;
     layer1_out[133] <= ~layer0_out[1793];
     layer1_out[134] <= layer0_out[1892] & ~layer0_out[1893];
     layer1_out[135] <= ~layer0_out[11847] | layer0_out[11848];
     layer1_out[136] <= 1'b0;
     layer1_out[137] <= layer0_out[1884] | layer0_out[1885];
     layer1_out[138] <= ~layer0_out[3287] | layer0_out[3286];
     layer1_out[139] <= layer0_out[10162] & layer0_out[10163];
     layer1_out[140] <= ~layer0_out[7337] | layer0_out[7336];
     layer1_out[141] <= ~(layer0_out[5633] | layer0_out[5634]);
     layer1_out[142] <= ~layer0_out[9351] | layer0_out[9350];
     layer1_out[143] <= layer0_out[8679] | layer0_out[8680];
     layer1_out[144] <= layer0_out[38];
     layer1_out[145] <= ~(layer0_out[1133] | layer0_out[1134]);
     layer1_out[146] <= layer0_out[7074] ^ layer0_out[7075];
     layer1_out[147] <= ~layer0_out[70] | layer0_out[71];
     layer1_out[148] <= layer0_out[4715] ^ layer0_out[4716];
     layer1_out[149] <= layer0_out[6617];
     layer1_out[150] <= ~layer0_out[9304];
     layer1_out[151] <= layer0_out[9193] & ~layer0_out[9194];
     layer1_out[152] <= layer0_out[8221];
     layer1_out[153] <= layer0_out[5341];
     layer1_out[154] <= 1'b1;
     layer1_out[155] <= ~layer0_out[8390] | layer0_out[8391];
     layer1_out[156] <= layer0_out[1857];
     layer1_out[157] <= ~layer0_out[2741];
     layer1_out[158] <= ~layer0_out[9508];
     layer1_out[159] <= layer0_out[10216] & ~layer0_out[10215];
     layer1_out[160] <= 1'b1;
     layer1_out[161] <= ~(layer0_out[7970] | layer0_out[7971]);
     layer1_out[162] <= ~layer0_out[10235];
     layer1_out[163] <= layer0_out[8524] & ~layer0_out[8525];
     layer1_out[164] <= layer0_out[1755];
     layer1_out[165] <= layer0_out[7187] & ~layer0_out[7188];
     layer1_out[166] <= layer0_out[8596] & ~layer0_out[8595];
     layer1_out[167] <= layer0_out[1100] & ~layer0_out[1099];
     layer1_out[168] <= ~layer0_out[6790];
     layer1_out[169] <= ~layer0_out[3479];
     layer1_out[170] <= layer0_out[8418];
     layer1_out[171] <= ~(layer0_out[11258] & layer0_out[11259]);
     layer1_out[172] <= ~layer0_out[8940];
     layer1_out[173] <= ~layer0_out[2987] | layer0_out[2986];
     layer1_out[174] <= layer0_out[6845] | layer0_out[6846];
     layer1_out[175] <= 1'b1;
     layer1_out[176] <= ~layer0_out[11202];
     layer1_out[177] <= layer0_out[11699] & ~layer0_out[11700];
     layer1_out[178] <= layer0_out[11703];
     layer1_out[179] <= 1'b1;
     layer1_out[180] <= ~(layer0_out[11153] ^ layer0_out[11154]);
     layer1_out[181] <= ~layer0_out[86] | layer0_out[85];
     layer1_out[182] <= ~layer0_out[9520] | layer0_out[9521];
     layer1_out[183] <= layer0_out[8464] | layer0_out[8465];
     layer1_out[184] <= layer0_out[1710];
     layer1_out[185] <= ~(layer0_out[1143] ^ layer0_out[1144]);
     layer1_out[186] <= layer0_out[4869];
     layer1_out[187] <= layer0_out[6363] & ~layer0_out[6362];
     layer1_out[188] <= ~layer0_out[10044];
     layer1_out[189] <= 1'b0;
     layer1_out[190] <= ~layer0_out[1607] | layer0_out[1608];
     layer1_out[191] <= ~layer0_out[7071] | layer0_out[7070];
     layer1_out[192] <= ~(layer0_out[60] ^ layer0_out[61]);
     layer1_out[193] <= 1'b1;
     layer1_out[194] <= ~(layer0_out[5207] ^ layer0_out[5208]);
     layer1_out[195] <= layer0_out[9665] | layer0_out[9666];
     layer1_out[196] <= ~layer0_out[2405];
     layer1_out[197] <= layer0_out[4461] | layer0_out[4462];
     layer1_out[198] <= layer0_out[3191] & layer0_out[3192];
     layer1_out[199] <= ~layer0_out[2462] | layer0_out[2463];
     layer1_out[200] <= ~layer0_out[9810];
     layer1_out[201] <= ~(layer0_out[3463] | layer0_out[3464]);
     layer1_out[202] <= layer0_out[6372];
     layer1_out[203] <= ~(layer0_out[5974] & layer0_out[5975]);
     layer1_out[204] <= ~layer0_out[9779];
     layer1_out[205] <= ~(layer0_out[10807] & layer0_out[10808]);
     layer1_out[206] <= ~layer0_out[2304];
     layer1_out[207] <= layer0_out[8086];
     layer1_out[208] <= ~(layer0_out[8326] | layer0_out[8327]);
     layer1_out[209] <= layer0_out[617];
     layer1_out[210] <= layer0_out[3653] & ~layer0_out[3652];
     layer1_out[211] <= ~layer0_out[5508];
     layer1_out[212] <= layer0_out[11089] ^ layer0_out[11090];
     layer1_out[213] <= layer0_out[3808];
     layer1_out[214] <= layer0_out[9020] & ~layer0_out[9019];
     layer1_out[215] <= layer0_out[2283];
     layer1_out[216] <= layer0_out[10009] & layer0_out[10010];
     layer1_out[217] <= ~(layer0_out[1533] & layer0_out[1534]);
     layer1_out[218] <= 1'b0;
     layer1_out[219] <= ~layer0_out[10826];
     layer1_out[220] <= ~layer0_out[8037];
     layer1_out[221] <= layer0_out[6163] ^ layer0_out[6164];
     layer1_out[222] <= ~(layer0_out[1971] | layer0_out[1972]);
     layer1_out[223] <= ~(layer0_out[11490] | layer0_out[11491]);
     layer1_out[224] <= layer0_out[11998];
     layer1_out[225] <= layer0_out[5628];
     layer1_out[226] <= ~layer0_out[7316];
     layer1_out[227] <= ~layer0_out[10611];
     layer1_out[228] <= ~layer0_out[11628] | layer0_out[11627];
     layer1_out[229] <= layer0_out[10621] & ~layer0_out[10622];
     layer1_out[230] <= ~layer0_out[1664] | layer0_out[1663];
     layer1_out[231] <= ~layer0_out[9173];
     layer1_out[232] <= layer0_out[6607] & layer0_out[6608];
     layer1_out[233] <= layer0_out[11984];
     layer1_out[234] <= ~(layer0_out[1334] | layer0_out[1335]);
     layer1_out[235] <= ~(layer0_out[4982] ^ layer0_out[4983]);
     layer1_out[236] <= layer0_out[8305];
     layer1_out[237] <= ~layer0_out[3627] | layer0_out[3626];
     layer1_out[238] <= ~layer0_out[2278];
     layer1_out[239] <= layer0_out[6116] | layer0_out[6117];
     layer1_out[240] <= layer0_out[3513] | layer0_out[3514];
     layer1_out[241] <= ~layer0_out[2838];
     layer1_out[242] <= layer0_out[3311];
     layer1_out[243] <= ~layer0_out[11597];
     layer1_out[244] <= layer0_out[9084] | layer0_out[9085];
     layer1_out[245] <= layer0_out[4051];
     layer1_out[246] <= ~layer0_out[10023] | layer0_out[10022];
     layer1_out[247] <= ~layer0_out[2778];
     layer1_out[248] <= ~layer0_out[10092] | layer0_out[10093];
     layer1_out[249] <= ~(layer0_out[11288] | layer0_out[11289]);
     layer1_out[250] <= layer0_out[10537] ^ layer0_out[10538];
     layer1_out[251] <= layer0_out[4852] & layer0_out[4853];
     layer1_out[252] <= layer0_out[8536] & ~layer0_out[8537];
     layer1_out[253] <= layer0_out[7395] & ~layer0_out[7394];
     layer1_out[254] <= ~(layer0_out[10796] | layer0_out[10797]);
     layer1_out[255] <= ~(layer0_out[9086] ^ layer0_out[9087]);
     layer1_out[256] <= ~layer0_out[8109] | layer0_out[8110];
     layer1_out[257] <= layer0_out[9145] & ~layer0_out[9146];
     layer1_out[258] <= layer0_out[2859] | layer0_out[2860];
     layer1_out[259] <= ~layer0_out[3326];
     layer1_out[260] <= ~layer0_out[11726];
     layer1_out[261] <= layer0_out[406];
     layer1_out[262] <= layer0_out[8568] & ~layer0_out[8569];
     layer1_out[263] <= ~(layer0_out[2601] | layer0_out[2602]);
     layer1_out[264] <= ~(layer0_out[132] ^ layer0_out[133]);
     layer1_out[265] <= ~(layer0_out[1401] | layer0_out[1402]);
     layer1_out[266] <= ~layer0_out[2478];
     layer1_out[267] <= layer0_out[11615];
     layer1_out[268] <= 1'b0;
     layer1_out[269] <= ~layer0_out[10418];
     layer1_out[270] <= ~layer0_out[112];
     layer1_out[271] <= ~layer0_out[9058];
     layer1_out[272] <= layer0_out[10865] & ~layer0_out[10864];
     layer1_out[273] <= ~layer0_out[9915];
     layer1_out[274] <= layer0_out[8417];
     layer1_out[275] <= layer0_out[8565] & layer0_out[8566];
     layer1_out[276] <= ~layer0_out[11177] | layer0_out[11178];
     layer1_out[277] <= ~(layer0_out[2692] ^ layer0_out[2693]);
     layer1_out[278] <= layer0_out[7966] & ~layer0_out[7967];
     layer1_out[279] <= layer0_out[11015] | layer0_out[11016];
     layer1_out[280] <= layer0_out[11616] & ~layer0_out[11617];
     layer1_out[281] <= layer0_out[6671];
     layer1_out[282] <= ~layer0_out[10524] | layer0_out[10525];
     layer1_out[283] <= ~(layer0_out[5966] | layer0_out[5967]);
     layer1_out[284] <= layer0_out[8057] & layer0_out[8058];
     layer1_out[285] <= ~layer0_out[10322] | layer0_out[10321];
     layer1_out[286] <= layer0_out[2312] & layer0_out[2313];
     layer1_out[287] <= ~layer0_out[11359];
     layer1_out[288] <= layer0_out[10926];
     layer1_out[289] <= layer0_out[11845];
     layer1_out[290] <= layer0_out[1289] & layer0_out[1290];
     layer1_out[291] <= layer0_out[9396] & layer0_out[9397];
     layer1_out[292] <= layer0_out[795] ^ layer0_out[796];
     layer1_out[293] <= ~layer0_out[8161];
     layer1_out[294] <= ~layer0_out[4386];
     layer1_out[295] <= 1'b0;
     layer1_out[296] <= ~(layer0_out[10863] & layer0_out[10864]);
     layer1_out[297] <= ~layer0_out[10599];
     layer1_out[298] <= ~layer0_out[7347];
     layer1_out[299] <= ~(layer0_out[526] & layer0_out[527]);
     layer1_out[300] <= ~(layer0_out[10858] | layer0_out[10859]);
     layer1_out[301] <= ~(layer0_out[10560] | layer0_out[10561]);
     layer1_out[302] <= layer0_out[7956] | layer0_out[7957];
     layer1_out[303] <= layer0_out[10413] ^ layer0_out[10414];
     layer1_out[304] <= layer0_out[8406] & layer0_out[8407];
     layer1_out[305] <= layer0_out[7552] & ~layer0_out[7551];
     layer1_out[306] <= ~layer0_out[2572] | layer0_out[2573];
     layer1_out[307] <= layer0_out[10159] | layer0_out[10160];
     layer1_out[308] <= layer0_out[1094] & ~layer0_out[1093];
     layer1_out[309] <= ~layer0_out[2404] | layer0_out[2405];
     layer1_out[310] <= ~(layer0_out[7076] & layer0_out[7077]);
     layer1_out[311] <= ~layer0_out[6584] | layer0_out[6583];
     layer1_out[312] <= 1'b0;
     layer1_out[313] <= layer0_out[8447] ^ layer0_out[8448];
     layer1_out[314] <= ~layer0_out[10190] | layer0_out[10191];
     layer1_out[315] <= ~layer0_out[11012];
     layer1_out[316] <= ~(layer0_out[8203] & layer0_out[8204]);
     layer1_out[317] <= ~layer0_out[7635] | layer0_out[7634];
     layer1_out[318] <= layer0_out[6375] & ~layer0_out[6374];
     layer1_out[319] <= ~layer0_out[102] | layer0_out[101];
     layer1_out[320] <= ~layer0_out[10967];
     layer1_out[321] <= layer0_out[11140] ^ layer0_out[11141];
     layer1_out[322] <= 1'b1;
     layer1_out[323] <= layer0_out[1927] | layer0_out[1928];
     layer1_out[324] <= layer0_out[6337];
     layer1_out[325] <= layer0_out[9613] & ~layer0_out[9612];
     layer1_out[326] <= ~(layer0_out[5311] & layer0_out[5312]);
     layer1_out[327] <= ~layer0_out[11902];
     layer1_out[328] <= layer0_out[7734] & layer0_out[7735];
     layer1_out[329] <= layer0_out[8649] & ~layer0_out[8650];
     layer1_out[330] <= ~layer0_out[11284] | layer0_out[11283];
     layer1_out[331] <= ~layer0_out[4515] | layer0_out[4514];
     layer1_out[332] <= layer0_out[204];
     layer1_out[333] <= ~layer0_out[6159];
     layer1_out[334] <= ~layer0_out[1478];
     layer1_out[335] <= ~layer0_out[4418] | layer0_out[4417];
     layer1_out[336] <= layer0_out[10778] ^ layer0_out[10779];
     layer1_out[337] <= layer0_out[11221] & ~layer0_out[11220];
     layer1_out[338] <= layer0_out[2105] & ~layer0_out[2106];
     layer1_out[339] <= layer0_out[1563] | layer0_out[1564];
     layer1_out[340] <= layer0_out[10431] | layer0_out[10432];
     layer1_out[341] <= layer0_out[8792] ^ layer0_out[8793];
     layer1_out[342] <= layer0_out[1107] & ~layer0_out[1108];
     layer1_out[343] <= layer0_out[3510] & ~layer0_out[3509];
     layer1_out[344] <= ~layer0_out[4759];
     layer1_out[345] <= layer0_out[4861] | layer0_out[4862];
     layer1_out[346] <= layer0_out[7355];
     layer1_out[347] <= ~(layer0_out[10266] & layer0_out[10267]);
     layer1_out[348] <= ~(layer0_out[1268] | layer0_out[1269]);
     layer1_out[349] <= ~(layer0_out[5994] | layer0_out[5995]);
     layer1_out[350] <= layer0_out[11455];
     layer1_out[351] <= layer0_out[8219] ^ layer0_out[8220];
     layer1_out[352] <= layer0_out[4818] ^ layer0_out[4819];
     layer1_out[353] <= ~layer0_out[6355] | layer0_out[6356];
     layer1_out[354] <= layer0_out[6451] & layer0_out[6452];
     layer1_out[355] <= layer0_out[6897];
     layer1_out[356] <= layer0_out[7472];
     layer1_out[357] <= layer0_out[7317];
     layer1_out[358] <= 1'b0;
     layer1_out[359] <= ~layer0_out[566] | layer0_out[567];
     layer1_out[360] <= layer0_out[5313] & ~layer0_out[5314];
     layer1_out[361] <= layer0_out[123] ^ layer0_out[124];
     layer1_out[362] <= ~(layer0_out[2458] & layer0_out[2459]);
     layer1_out[363] <= layer0_out[1905] & ~layer0_out[1906];
     layer1_out[364] <= ~layer0_out[11817] | layer0_out[11818];
     layer1_out[365] <= layer0_out[8674];
     layer1_out[366] <= layer0_out[11623];
     layer1_out[367] <= layer0_out[8631];
     layer1_out[368] <= 1'b0;
     layer1_out[369] <= ~(layer0_out[7664] | layer0_out[7665]);
     layer1_out[370] <= 1'b0;
     layer1_out[371] <= 1'b1;
     layer1_out[372] <= layer0_out[3579];
     layer1_out[373] <= ~layer0_out[8531];
     layer1_out[374] <= ~layer0_out[10065] | layer0_out[10064];
     layer1_out[375] <= layer0_out[5566];
     layer1_out[376] <= ~(layer0_out[5734] | layer0_out[5735]);
     layer1_out[377] <= ~(layer0_out[3293] | layer0_out[3294]);
     layer1_out[378] <= ~layer0_out[4526] | layer0_out[4527];
     layer1_out[379] <= layer0_out[3519];
     layer1_out[380] <= layer0_out[5271] & layer0_out[5272];
     layer1_out[381] <= layer0_out[4103];
     layer1_out[382] <= 1'b1;
     layer1_out[383] <= layer0_out[2310] & ~layer0_out[2311];
     layer1_out[384] <= ~(layer0_out[8950] & layer0_out[8951]);
     layer1_out[385] <= layer0_out[4681] ^ layer0_out[4682];
     layer1_out[386] <= ~layer0_out[2682] | layer0_out[2681];
     layer1_out[387] <= ~(layer0_out[8342] | layer0_out[8343]);
     layer1_out[388] <= layer0_out[1721] & ~layer0_out[1722];
     layer1_out[389] <= layer0_out[3957] & ~layer0_out[3958];
     layer1_out[390] <= 1'b1;
     layer1_out[391] <= ~layer0_out[3404];
     layer1_out[392] <= ~(layer0_out[2748] | layer0_out[2749]);
     layer1_out[393] <= ~layer0_out[1903];
     layer1_out[394] <= ~layer0_out[5016];
     layer1_out[395] <= ~layer0_out[7183] | layer0_out[7184];
     layer1_out[396] <= layer0_out[1618] & layer0_out[1619];
     layer1_out[397] <= ~layer0_out[11306];
     layer1_out[398] <= ~(layer0_out[11147] | layer0_out[11148]);
     layer1_out[399] <= ~(layer0_out[9006] & layer0_out[9007]);
     layer1_out[400] <= layer0_out[685];
     layer1_out[401] <= ~layer0_out[10150];
     layer1_out[402] <= ~(layer0_out[11946] ^ layer0_out[11947]);
     layer1_out[403] <= ~(layer0_out[278] | layer0_out[279]);
     layer1_out[404] <= ~(layer0_out[213] ^ layer0_out[214]);
     layer1_out[405] <= ~layer0_out[10667] | layer0_out[10666];
     layer1_out[406] <= layer0_out[9717];
     layer1_out[407] <= ~layer0_out[1222] | layer0_out[1221];
     layer1_out[408] <= layer0_out[9037];
     layer1_out[409] <= ~layer0_out[4625];
     layer1_out[410] <= ~(layer0_out[261] | layer0_out[262]);
     layer1_out[411] <= ~layer0_out[8393];
     layer1_out[412] <= layer0_out[10264];
     layer1_out[413] <= layer0_out[2351] & ~layer0_out[2352];
     layer1_out[414] <= ~layer0_out[11381] | layer0_out[11382];
     layer1_out[415] <= layer0_out[5748] & layer0_out[5749];
     layer1_out[416] <= layer0_out[9802];
     layer1_out[417] <= 1'b1;
     layer1_out[418] <= layer0_out[3274];
     layer1_out[419] <= layer0_out[11737] & layer0_out[11738];
     layer1_out[420] <= ~layer0_out[3477];
     layer1_out[421] <= ~layer0_out[1158];
     layer1_out[422] <= ~layer0_out[8709];
     layer1_out[423] <= ~layer0_out[3247] | layer0_out[3246];
     layer1_out[424] <= layer0_out[4396];
     layer1_out[425] <= ~layer0_out[1718];
     layer1_out[426] <= ~layer0_out[11706];
     layer1_out[427] <= layer0_out[9175] & ~layer0_out[9176];
     layer1_out[428] <= layer0_out[11584];
     layer1_out[429] <= layer0_out[5740];
     layer1_out[430] <= 1'b0;
     layer1_out[431] <= layer0_out[974] & ~layer0_out[975];
     layer1_out[432] <= ~layer0_out[5214];
     layer1_out[433] <= layer0_out[2670];
     layer1_out[434] <= ~layer0_out[4554] | layer0_out[4555];
     layer1_out[435] <= 1'b1;
     layer1_out[436] <= ~(layer0_out[353] ^ layer0_out[354]);
     layer1_out[437] <= layer0_out[11807];
     layer1_out[438] <= ~layer0_out[5685];
     layer1_out[439] <= layer0_out[867] | layer0_out[868];
     layer1_out[440] <= layer0_out[265] ^ layer0_out[266];
     layer1_out[441] <= layer0_out[104] & ~layer0_out[103];
     layer1_out[442] <= ~(layer0_out[11310] ^ layer0_out[11311]);
     layer1_out[443] <= layer0_out[10555];
     layer1_out[444] <= layer0_out[9082];
     layer1_out[445] <= layer0_out[6563] | layer0_out[6564];
     layer1_out[446] <= layer0_out[4997];
     layer1_out[447] <= ~layer0_out[10351] | layer0_out[10350];
     layer1_out[448] <= layer0_out[11550] & layer0_out[11551];
     layer1_out[449] <= ~layer0_out[1245] | layer0_out[1246];
     layer1_out[450] <= layer0_out[7653] | layer0_out[7654];
     layer1_out[451] <= ~layer0_out[6267] | layer0_out[6268];
     layer1_out[452] <= 1'b0;
     layer1_out[453] <= ~layer0_out[2269];
     layer1_out[454] <= layer0_out[632] & ~layer0_out[631];
     layer1_out[455] <= layer0_out[11127] & ~layer0_out[11128];
     layer1_out[456] <= ~(layer0_out[7134] | layer0_out[7135]);
     layer1_out[457] <= layer0_out[6384];
     layer1_out[458] <= layer0_out[3520];
     layer1_out[459] <= ~(layer0_out[2892] | layer0_out[2893]);
     layer1_out[460] <= layer0_out[8382];
     layer1_out[461] <= ~layer0_out[2057];
     layer1_out[462] <= layer0_out[5754];
     layer1_out[463] <= layer0_out[11659] & ~layer0_out[11660];
     layer1_out[464] <= layer0_out[6434];
     layer1_out[465] <= ~layer0_out[6347] | layer0_out[6346];
     layer1_out[466] <= layer0_out[9756];
     layer1_out[467] <= ~layer0_out[7103];
     layer1_out[468] <= layer0_out[11512] ^ layer0_out[11513];
     layer1_out[469] <= layer0_out[1175] & ~layer0_out[1174];
     layer1_out[470] <= ~layer0_out[8351];
     layer1_out[471] <= layer0_out[3736];
     layer1_out[472] <= ~(layer0_out[9470] & layer0_out[9471]);
     layer1_out[473] <= layer0_out[6670] & layer0_out[6671];
     layer1_out[474] <= layer0_out[10364];
     layer1_out[475] <= ~(layer0_out[3354] ^ layer0_out[3355]);
     layer1_out[476] <= layer0_out[9399] & ~layer0_out[9400];
     layer1_out[477] <= ~(layer0_out[55] ^ layer0_out[56]);
     layer1_out[478] <= layer0_out[9326] & ~layer0_out[9325];
     layer1_out[479] <= ~(layer0_out[11820] ^ layer0_out[11821]);
     layer1_out[480] <= ~layer0_out[193] | layer0_out[194];
     layer1_out[481] <= ~layer0_out[3525] | layer0_out[3526];
     layer1_out[482] <= ~(layer0_out[9367] & layer0_out[9368]);
     layer1_out[483] <= ~(layer0_out[6792] ^ layer0_out[6793]);
     layer1_out[484] <= layer0_out[10611];
     layer1_out[485] <= layer0_out[10046];
     layer1_out[486] <= ~(layer0_out[11742] | layer0_out[11743]);
     layer1_out[487] <= ~(layer0_out[9467] & layer0_out[9468]);
     layer1_out[488] <= layer0_out[8345] ^ layer0_out[8346];
     layer1_out[489] <= layer0_out[5977];
     layer1_out[490] <= ~layer0_out[899] | layer0_out[898];
     layer1_out[491] <= ~layer0_out[6131] | layer0_out[6132];
     layer1_out[492] <= layer0_out[9974];
     layer1_out[493] <= ~layer0_out[11507] | layer0_out[11508];
     layer1_out[494] <= layer0_out[1886];
     layer1_out[495] <= ~layer0_out[3727];
     layer1_out[496] <= ~layer0_out[2679];
     layer1_out[497] <= layer0_out[3545] & ~layer0_out[3546];
     layer1_out[498] <= layer0_out[3095] & layer0_out[3096];
     layer1_out[499] <= layer0_out[7373];
     layer1_out[500] <= ~(layer0_out[4849] | layer0_out[4850]);
     layer1_out[501] <= ~layer0_out[8597];
     layer1_out[502] <= layer0_out[10143] & ~layer0_out[10144];
     layer1_out[503] <= layer0_out[6230] ^ layer0_out[6231];
     layer1_out[504] <= ~layer0_out[3996];
     layer1_out[505] <= ~layer0_out[9022];
     layer1_out[506] <= layer0_out[9871] ^ layer0_out[9872];
     layer1_out[507] <= layer0_out[3119] | layer0_out[3120];
     layer1_out[508] <= ~layer0_out[4039] | layer0_out[4038];
     layer1_out[509] <= layer0_out[7132];
     layer1_out[510] <= layer0_out[5447] & layer0_out[5448];
     layer1_out[511] <= layer0_out[1909];
     layer1_out[512] <= layer0_out[543] | layer0_out[544];
     layer1_out[513] <= layer0_out[2482] | layer0_out[2483];
     layer1_out[514] <= ~layer0_out[3601];
     layer1_out[515] <= ~layer0_out[2519] | layer0_out[2520];
     layer1_out[516] <= ~layer0_out[80] | layer0_out[81];
     layer1_out[517] <= ~(layer0_out[2324] | layer0_out[2325]);
     layer1_out[518] <= ~(layer0_out[346] & layer0_out[347]);
     layer1_out[519] <= layer0_out[11887];
     layer1_out[520] <= layer0_out[770] & ~layer0_out[769];
     layer1_out[521] <= ~layer0_out[10805];
     layer1_out[522] <= ~(layer0_out[8377] | layer0_out[8378]);
     layer1_out[523] <= layer0_out[2017] & ~layer0_out[2016];
     layer1_out[524] <= ~layer0_out[5260] | layer0_out[5261];
     layer1_out[525] <= ~layer0_out[3640];
     layer1_out[526] <= layer0_out[6726] | layer0_out[6727];
     layer1_out[527] <= layer0_out[8814];
     layer1_out[528] <= layer0_out[8559];
     layer1_out[529] <= layer0_out[9363];
     layer1_out[530] <= layer0_out[10158] & layer0_out[10159];
     layer1_out[531] <= ~layer0_out[4878] | layer0_out[4879];
     layer1_out[532] <= layer0_out[9490] & layer0_out[9491];
     layer1_out[533] <= layer0_out[8590];
     layer1_out[534] <= layer0_out[4779];
     layer1_out[535] <= ~layer0_out[10908] | layer0_out[10907];
     layer1_out[536] <= layer0_out[6008];
     layer1_out[537] <= layer0_out[5176];
     layer1_out[538] <= ~layer0_out[6130];
     layer1_out[539] <= ~layer0_out[2017] | layer0_out[2018];
     layer1_out[540] <= 1'b0;
     layer1_out[541] <= ~layer0_out[6294];
     layer1_out[542] <= ~layer0_out[7031];
     layer1_out[543] <= layer0_out[5201] & ~layer0_out[5202];
     layer1_out[544] <= ~layer0_out[10820];
     layer1_out[545] <= 1'b1;
     layer1_out[546] <= layer0_out[11443] & ~layer0_out[11442];
     layer1_out[547] <= layer0_out[8212];
     layer1_out[548] <= ~layer0_out[8033] | layer0_out[8034];
     layer1_out[549] <= layer0_out[5737] & layer0_out[5738];
     layer1_out[550] <= layer0_out[4860] | layer0_out[4861];
     layer1_out[551] <= ~layer0_out[6862] | layer0_out[6861];
     layer1_out[552] <= ~layer0_out[7223];
     layer1_out[553] <= layer0_out[2565];
     layer1_out[554] <= ~(layer0_out[2636] | layer0_out[2637]);
     layer1_out[555] <= layer0_out[344];
     layer1_out[556] <= layer0_out[5902] & ~layer0_out[5901];
     layer1_out[557] <= layer0_out[8867];
     layer1_out[558] <= ~layer0_out[2668];
     layer1_out[559] <= 1'b0;
     layer1_out[560] <= ~(layer0_out[6516] ^ layer0_out[6517]);
     layer1_out[561] <= ~layer0_out[5125] | layer0_out[5126];
     layer1_out[562] <= 1'b1;
     layer1_out[563] <= layer0_out[9010];
     layer1_out[564] <= layer0_out[712];
     layer1_out[565] <= layer0_out[5333];
     layer1_out[566] <= ~layer0_out[5100];
     layer1_out[567] <= ~(layer0_out[2888] | layer0_out[2889]);
     layer1_out[568] <= layer0_out[9998] | layer0_out[9999];
     layer1_out[569] <= ~(layer0_out[1321] & layer0_out[1322]);
     layer1_out[570] <= ~(layer0_out[1153] ^ layer0_out[1154]);
     layer1_out[571] <= layer0_out[4937] | layer0_out[4938];
     layer1_out[572] <= layer0_out[5809] & layer0_out[5810];
     layer1_out[573] <= layer0_out[4717];
     layer1_out[574] <= ~layer0_out[1044] | layer0_out[1045];
     layer1_out[575] <= layer0_out[11573] | layer0_out[11574];
     layer1_out[576] <= layer0_out[1874];
     layer1_out[577] <= ~(layer0_out[2684] & layer0_out[2685]);
     layer1_out[578] <= layer0_out[8179] & layer0_out[8180];
     layer1_out[579] <= ~layer0_out[7186];
     layer1_out[580] <= ~layer0_out[1480] | layer0_out[1479];
     layer1_out[581] <= ~layer0_out[7008] | layer0_out[7007];
     layer1_out[582] <= layer0_out[7724];
     layer1_out[583] <= ~layer0_out[10167];
     layer1_out[584] <= ~(layer0_out[7311] ^ layer0_out[7312]);
     layer1_out[585] <= ~layer0_out[9178];
     layer1_out[586] <= layer0_out[9040] & ~layer0_out[9041];
     layer1_out[587] <= layer0_out[11520];
     layer1_out[588] <= ~layer0_out[3227] | layer0_out[3226];
     layer1_out[589] <= layer0_out[10394] & ~layer0_out[10393];
     layer1_out[590] <= layer0_out[6329] & ~layer0_out[6330];
     layer1_out[591] <= ~(layer0_out[1665] & layer0_out[1666]);
     layer1_out[592] <= layer0_out[9622] ^ layer0_out[9623];
     layer1_out[593] <= ~layer0_out[4216] | layer0_out[4217];
     layer1_out[594] <= ~layer0_out[5233];
     layer1_out[595] <= ~layer0_out[1970] | layer0_out[1971];
     layer1_out[596] <= ~(layer0_out[8177] | layer0_out[8178]);
     layer1_out[597] <= ~(layer0_out[915] ^ layer0_out[916]);
     layer1_out[598] <= ~(layer0_out[7657] | layer0_out[7658]);
     layer1_out[599] <= layer0_out[6797] & layer0_out[6798];
     layer1_out[600] <= layer0_out[1391];
     layer1_out[601] <= ~(layer0_out[6406] | layer0_out[6407]);
     layer1_out[602] <= ~layer0_out[3937];
     layer1_out[603] <= ~(layer0_out[8001] & layer0_out[8002]);
     layer1_out[604] <= layer0_out[1418] | layer0_out[1419];
     layer1_out[605] <= layer0_out[5674] | layer0_out[5675];
     layer1_out[606] <= ~layer0_out[6747] | layer0_out[6746];
     layer1_out[607] <= ~layer0_out[7927];
     layer1_out[608] <= layer0_out[4014];
     layer1_out[609] <= ~layer0_out[9924];
     layer1_out[610] <= layer0_out[6877];
     layer1_out[611] <= layer0_out[5091];
     layer1_out[612] <= ~(layer0_out[8149] | layer0_out[8150]);
     layer1_out[613] <= 1'b0;
     layer1_out[614] <= layer0_out[5240];
     layer1_out[615] <= ~(layer0_out[6749] | layer0_out[6750]);
     layer1_out[616] <= layer0_out[2795] | layer0_out[2796];
     layer1_out[617] <= layer0_out[6170] | layer0_out[6171];
     layer1_out[618] <= layer0_out[9996] ^ layer0_out[9997];
     layer1_out[619] <= 1'b0;
     layer1_out[620] <= ~layer0_out[11385];
     layer1_out[621] <= layer0_out[3886] & layer0_out[3887];
     layer1_out[622] <= layer0_out[7586];
     layer1_out[623] <= layer0_out[11936];
     layer1_out[624] <= ~layer0_out[2012];
     layer1_out[625] <= layer0_out[10742] & ~layer0_out[10741];
     layer1_out[626] <= layer0_out[3673];
     layer1_out[627] <= layer0_out[11788] & layer0_out[11789];
     layer1_out[628] <= ~(layer0_out[4622] ^ layer0_out[4623]);
     layer1_out[629] <= ~layer0_out[8969] | layer0_out[8970];
     layer1_out[630] <= layer0_out[5301] | layer0_out[5302];
     layer1_out[631] <= layer0_out[2619];
     layer1_out[632] <= ~layer0_out[7740] | layer0_out[7739];
     layer1_out[633] <= ~(layer0_out[1236] & layer0_out[1237]);
     layer1_out[634] <= ~layer0_out[616];
     layer1_out[635] <= layer0_out[9051];
     layer1_out[636] <= ~(layer0_out[6989] ^ layer0_out[6990]);
     layer1_out[637] <= ~layer0_out[8863] | layer0_out[8864];
     layer1_out[638] <= layer0_out[2058];
     layer1_out[639] <= layer0_out[1210] & ~layer0_out[1211];
     layer1_out[640] <= ~layer0_out[7402];
     layer1_out[641] <= ~layer0_out[7522] | layer0_out[7523];
     layer1_out[642] <= 1'b0;
     layer1_out[643] <= ~(layer0_out[7639] & layer0_out[7640]);
     layer1_out[644] <= layer0_out[5074] & ~layer0_out[5073];
     layer1_out[645] <= ~layer0_out[267];
     layer1_out[646] <= layer0_out[3301];
     layer1_out[647] <= ~layer0_out[4306] | layer0_out[4307];
     layer1_out[648] <= layer0_out[5053] & ~layer0_out[5054];
     layer1_out[649] <= layer0_out[2869];
     layer1_out[650] <= layer0_out[10818];
     layer1_out[651] <= layer0_out[7214] & layer0_out[7215];
     layer1_out[652] <= layer0_out[7155];
     layer1_out[653] <= layer0_out[3482] & ~layer0_out[3483];
     layer1_out[654] <= ~(layer0_out[8196] | layer0_out[8197]);
     layer1_out[655] <= layer0_out[42] & ~layer0_out[43];
     layer1_out[656] <= ~(layer0_out[845] | layer0_out[846]);
     layer1_out[657] <= layer0_out[11389];
     layer1_out[658] <= layer0_out[8257] & ~layer0_out[8258];
     layer1_out[659] <= layer0_out[1366] & ~layer0_out[1367];
     layer1_out[660] <= ~(layer0_out[2230] | layer0_out[2231]);
     layer1_out[661] <= layer0_out[7615] & ~layer0_out[7614];
     layer1_out[662] <= layer0_out[9448] & ~layer0_out[9449];
     layer1_out[663] <= layer0_out[969];
     layer1_out[664] <= ~layer0_out[7827] | layer0_out[7828];
     layer1_out[665] <= ~layer0_out[2675];
     layer1_out[666] <= ~layer0_out[5389] | layer0_out[5390];
     layer1_out[667] <= ~(layer0_out[949] | layer0_out[950]);
     layer1_out[668] <= ~(layer0_out[3373] | layer0_out[3374]);
     layer1_out[669] <= layer0_out[3396];
     layer1_out[670] <= layer0_out[6646];
     layer1_out[671] <= ~(layer0_out[3727] & layer0_out[3728]);
     layer1_out[672] <= ~layer0_out[8571];
     layer1_out[673] <= ~layer0_out[3444] | layer0_out[3445];
     layer1_out[674] <= layer0_out[11431] & ~layer0_out[11430];
     layer1_out[675] <= layer0_out[11435];
     layer1_out[676] <= layer0_out[9422] ^ layer0_out[9423];
     layer1_out[677] <= layer0_out[4067];
     layer1_out[678] <= layer0_out[9796] & ~layer0_out[9795];
     layer1_out[679] <= 1'b1;
     layer1_out[680] <= layer0_out[10637] & ~layer0_out[10636];
     layer1_out[681] <= ~(layer0_out[6698] | layer0_out[6699]);
     layer1_out[682] <= ~layer0_out[7851];
     layer1_out[683] <= layer0_out[4568];
     layer1_out[684] <= ~(layer0_out[10949] | layer0_out[10950]);
     layer1_out[685] <= ~layer0_out[11112] | layer0_out[11113];
     layer1_out[686] <= layer0_out[7673] ^ layer0_out[7674];
     layer1_out[687] <= ~layer0_out[1888];
     layer1_out[688] <= layer0_out[10408] & ~layer0_out[10409];
     layer1_out[689] <= ~(layer0_out[10678] & layer0_out[10679]);
     layer1_out[690] <= layer0_out[8094];
     layer1_out[691] <= ~(layer0_out[2882] & layer0_out[2883]);
     layer1_out[692] <= layer0_out[848] & ~layer0_out[847];
     layer1_out[693] <= ~layer0_out[11905];
     layer1_out[694] <= ~layer0_out[5959];
     layer1_out[695] <= layer0_out[491] & layer0_out[492];
     layer1_out[696] <= ~(layer0_out[1441] | layer0_out[1442]);
     layer1_out[697] <= ~layer0_out[7317];
     layer1_out[698] <= ~(layer0_out[3615] ^ layer0_out[3616]);
     layer1_out[699] <= layer0_out[9952];
     layer1_out[700] <= ~(layer0_out[5185] ^ layer0_out[5186]);
     layer1_out[701] <= layer0_out[3014];
     layer1_out[702] <= ~(layer0_out[11257] ^ layer0_out[11258]);
     layer1_out[703] <= ~(layer0_out[6943] ^ layer0_out[6944]);
     layer1_out[704] <= layer0_out[3636] & ~layer0_out[3637];
     layer1_out[705] <= ~layer0_out[9337] | layer0_out[9336];
     layer1_out[706] <= ~layer0_out[1015] | layer0_out[1016];
     layer1_out[707] <= ~layer0_out[6460] | layer0_out[6459];
     layer1_out[708] <= layer0_out[8221];
     layer1_out[709] <= layer0_out[2891] ^ layer0_out[2892];
     layer1_out[710] <= layer0_out[1423] & ~layer0_out[1424];
     layer1_out[711] <= layer0_out[6930] & ~layer0_out[6931];
     layer1_out[712] <= 1'b1;
     layer1_out[713] <= ~(layer0_out[2027] ^ layer0_out[2028]);
     layer1_out[714] <= layer0_out[9885] ^ layer0_out[9886];
     layer1_out[715] <= ~layer0_out[914];
     layer1_out[716] <= layer0_out[9918];
     layer1_out[717] <= ~layer0_out[11513];
     layer1_out[718] <= ~(layer0_out[2318] ^ layer0_out[2319]);
     layer1_out[719] <= layer0_out[6811] ^ layer0_out[6812];
     layer1_out[720] <= 1'b1;
     layer1_out[721] <= ~(layer0_out[8136] | layer0_out[8137]);
     layer1_out[722] <= layer0_out[6206] & ~layer0_out[6207];
     layer1_out[723] <= ~layer0_out[3202] | layer0_out[3203];
     layer1_out[724] <= ~(layer0_out[9922] | layer0_out[9923]);
     layer1_out[725] <= ~(layer0_out[5307] & layer0_out[5308]);
     layer1_out[726] <= ~layer0_out[10843] | layer0_out[10844];
     layer1_out[727] <= layer0_out[4371];
     layer1_out[728] <= ~(layer0_out[2836] ^ layer0_out[2837]);
     layer1_out[729] <= 1'b1;
     layer1_out[730] <= layer0_out[2238] & ~layer0_out[2237];
     layer1_out[731] <= layer0_out[6250] & layer0_out[6251];
     layer1_out[732] <= 1'b1;
     layer1_out[733] <= layer0_out[1007] ^ layer0_out[1008];
     layer1_out[734] <= layer0_out[6794] & ~layer0_out[6793];
     layer1_out[735] <= layer0_out[9921];
     layer1_out[736] <= layer0_out[1110];
     layer1_out[737] <= ~layer0_out[3849] | layer0_out[3848];
     layer1_out[738] <= layer0_out[10590];
     layer1_out[739] <= ~layer0_out[1668] | layer0_out[1669];
     layer1_out[740] <= 1'b1;
     layer1_out[741] <= ~(layer0_out[7687] ^ layer0_out[7688]);
     layer1_out[742] <= ~(layer0_out[4811] & layer0_out[4812]);
     layer1_out[743] <= layer0_out[893] & ~layer0_out[892];
     layer1_out[744] <= layer0_out[1805];
     layer1_out[745] <= layer0_out[10442] & ~layer0_out[10443];
     layer1_out[746] <= layer0_out[3341] | layer0_out[3342];
     layer1_out[747] <= ~layer0_out[1465];
     layer1_out[748] <= ~(layer0_out[9122] & layer0_out[9123]);
     layer1_out[749] <= ~(layer0_out[10246] | layer0_out[10247]);
     layer1_out[750] <= layer0_out[11960] & layer0_out[11961];
     layer1_out[751] <= layer0_out[7204];
     layer1_out[752] <= ~(layer0_out[11668] & layer0_out[11669]);
     layer1_out[753] <= ~(layer0_out[8545] | layer0_out[8546]);
     layer1_out[754] <= ~layer0_out[5765] | layer0_out[5766];
     layer1_out[755] <= layer0_out[11492];
     layer1_out[756] <= ~layer0_out[3986];
     layer1_out[757] <= ~(layer0_out[11778] | layer0_out[11779]);
     layer1_out[758] <= layer0_out[10822];
     layer1_out[759] <= ~(layer0_out[1325] & layer0_out[1326]);
     layer1_out[760] <= layer0_out[6179] | layer0_out[6180];
     layer1_out[761] <= layer0_out[3747];
     layer1_out[762] <= ~layer0_out[4964] | layer0_out[4965];
     layer1_out[763] <= ~(layer0_out[4081] | layer0_out[4082]);
     layer1_out[764] <= layer0_out[10263] ^ layer0_out[10264];
     layer1_out[765] <= layer0_out[1535] & ~layer0_out[1534];
     layer1_out[766] <= layer0_out[1031] | layer0_out[1032];
     layer1_out[767] <= ~(layer0_out[9720] & layer0_out[9721]);
     layer1_out[768] <= ~(layer0_out[5490] | layer0_out[5491]);
     layer1_out[769] <= layer0_out[1200] & ~layer0_out[1201];
     layer1_out[770] <= ~layer0_out[5434];
     layer1_out[771] <= ~layer0_out[3329];
     layer1_out[772] <= layer0_out[3214] & ~layer0_out[3213];
     layer1_out[773] <= ~layer0_out[7840] | layer0_out[7841];
     layer1_out[774] <= ~layer0_out[1709];
     layer1_out[775] <= ~(layer0_out[9360] & layer0_out[9361]);
     layer1_out[776] <= layer0_out[1985];
     layer1_out[777] <= layer0_out[2984];
     layer1_out[778] <= layer0_out[9691] | layer0_out[9692];
     layer1_out[779] <= layer0_out[10038] & ~layer0_out[10037];
     layer1_out[780] <= layer0_out[4087];
     layer1_out[781] <= layer0_out[10660];
     layer1_out[782] <= ~layer0_out[10832] | layer0_out[10833];
     layer1_out[783] <= layer0_out[2901] & ~layer0_out[2900];
     layer1_out[784] <= layer0_out[2915] & ~layer0_out[2916];
     layer1_out[785] <= layer0_out[4888] | layer0_out[4889];
     layer1_out[786] <= layer0_out[2970];
     layer1_out[787] <= 1'b1;
     layer1_out[788] <= layer0_out[1780];
     layer1_out[789] <= ~layer0_out[5804];
     layer1_out[790] <= layer0_out[5640];
     layer1_out[791] <= layer0_out[11191] & ~layer0_out[11192];
     layer1_out[792] <= ~layer0_out[3796];
     layer1_out[793] <= layer0_out[7237] & ~layer0_out[7238];
     layer1_out[794] <= ~(layer0_out[3865] & layer0_out[3866]);
     layer1_out[795] <= ~layer0_out[2736] | layer0_out[2737];
     layer1_out[796] <= layer0_out[4252] & layer0_out[4253];
     layer1_out[797] <= layer0_out[1547];
     layer1_out[798] <= layer0_out[2084] | layer0_out[2085];
     layer1_out[799] <= 1'b0;
     layer1_out[800] <= layer0_out[6200] & ~layer0_out[6201];
     layer1_out[801] <= ~layer0_out[5847] | layer0_out[5848];
     layer1_out[802] <= layer0_out[11218] & layer0_out[11219];
     layer1_out[803] <= layer0_out[2564] & ~layer0_out[2563];
     layer1_out[804] <= ~layer0_out[1934];
     layer1_out[805] <= layer0_out[5899];
     layer1_out[806] <= layer0_out[5584] & layer0_out[5585];
     layer1_out[807] <= ~layer0_out[6838] | layer0_out[6839];
     layer1_out[808] <= layer0_out[7535];
     layer1_out[809] <= layer0_out[7241];
     layer1_out[810] <= ~layer0_out[614];
     layer1_out[811] <= ~(layer0_out[1745] & layer0_out[1746]);
     layer1_out[812] <= layer0_out[6888];
     layer1_out[813] <= layer0_out[91] | layer0_out[92];
     layer1_out[814] <= layer0_out[10193] & ~layer0_out[10194];
     layer1_out[815] <= 1'b1;
     layer1_out[816] <= layer0_out[6663];
     layer1_out[817] <= 1'b0;
     layer1_out[818] <= ~layer0_out[8294] | layer0_out[8293];
     layer1_out[819] <= ~layer0_out[5634];
     layer1_out[820] <= layer0_out[7304];
     layer1_out[821] <= ~(layer0_out[11379] & layer0_out[11380]);
     layer1_out[822] <= ~(layer0_out[3792] | layer0_out[3793]);
     layer1_out[823] <= layer0_out[3714] | layer0_out[3715];
     layer1_out[824] <= layer0_out[10473] & layer0_out[10474];
     layer1_out[825] <= ~(layer0_out[1165] | layer0_out[1166]);
     layer1_out[826] <= ~layer0_out[1439];
     layer1_out[827] <= layer0_out[2363] & layer0_out[2364];
     layer1_out[828] <= ~layer0_out[3225] | layer0_out[3226];
     layer1_out[829] <= layer0_out[249];
     layer1_out[830] <= ~layer0_out[4532];
     layer1_out[831] <= ~layer0_out[10661] | layer0_out[10660];
     layer1_out[832] <= layer0_out[182];
     layer1_out[833] <= ~(layer0_out[8051] & layer0_out[8052]);
     layer1_out[834] <= ~(layer0_out[11096] | layer0_out[11097]);
     layer1_out[835] <= layer0_out[7190] & layer0_out[7191];
     layer1_out[836] <= layer0_out[5613] & ~layer0_out[5612];
     layer1_out[837] <= ~(layer0_out[9288] ^ layer0_out[9289]);
     layer1_out[838] <= ~layer0_out[8852];
     layer1_out[839] <= ~layer0_out[10210];
     layer1_out[840] <= layer0_out[635] & layer0_out[636];
     layer1_out[841] <= ~layer0_out[9614];
     layer1_out[842] <= layer0_out[216];
     layer1_out[843] <= layer0_out[11264];
     layer1_out[844] <= ~layer0_out[8036];
     layer1_out[845] <= layer0_out[6708] & layer0_out[6709];
     layer1_out[846] <= layer0_out[11450] ^ layer0_out[11451];
     layer1_out[847] <= layer0_out[9238];
     layer1_out[848] <= layer0_out[8296] & ~layer0_out[8295];
     layer1_out[849] <= ~layer0_out[4849] | layer0_out[4848];
     layer1_out[850] <= layer0_out[11455] & ~layer0_out[11454];
     layer1_out[851] <= ~layer0_out[6648];
     layer1_out[852] <= 1'b1;
     layer1_out[853] <= ~layer0_out[5658];
     layer1_out[854] <= layer0_out[10469];
     layer1_out[855] <= ~(layer0_out[637] | layer0_out[638]);
     layer1_out[856] <= layer0_out[9245] & layer0_out[9246];
     layer1_out[857] <= layer0_out[7543];
     layer1_out[858] <= layer0_out[9919] & layer0_out[9920];
     layer1_out[859] <= layer0_out[4083] & ~layer0_out[4084];
     layer1_out[860] <= layer0_out[6465] ^ layer0_out[6466];
     layer1_out[861] <= 1'b0;
     layer1_out[862] <= ~(layer0_out[2459] | layer0_out[2460]);
     layer1_out[863] <= ~layer0_out[1724];
     layer1_out[864] <= ~(layer0_out[1810] | layer0_out[1811]);
     layer1_out[865] <= layer0_out[6228];
     layer1_out[866] <= ~layer0_out[2323];
     layer1_out[867] <= ~layer0_out[3721];
     layer1_out[868] <= ~layer0_out[7161] | layer0_out[7160];
     layer1_out[869] <= 1'b1;
     layer1_out[870] <= layer0_out[8590];
     layer1_out[871] <= ~layer0_out[1705] | layer0_out[1704];
     layer1_out[872] <= ~layer0_out[4820];
     layer1_out[873] <= layer0_out[7100];
     layer1_out[874] <= ~layer0_out[9154];
     layer1_out[875] <= ~(layer0_out[3655] | layer0_out[3656]);
     layer1_out[876] <= ~layer0_out[10381] | layer0_out[10382];
     layer1_out[877] <= ~layer0_out[1175] | layer0_out[1176];
     layer1_out[878] <= ~(layer0_out[294] ^ layer0_out[295]);
     layer1_out[879] <= ~(layer0_out[7740] ^ layer0_out[7741]);
     layer1_out[880] <= layer0_out[3763];
     layer1_out[881] <= ~layer0_out[3090];
     layer1_out[882] <= ~layer0_out[5620] | layer0_out[5619];
     layer1_out[883] <= layer0_out[10891] & layer0_out[10892];
     layer1_out[884] <= layer0_out[3583] & ~layer0_out[3582];
     layer1_out[885] <= layer0_out[1639] & ~layer0_out[1640];
     layer1_out[886] <= layer0_out[5621];
     layer1_out[887] <= layer0_out[11050];
     layer1_out[888] <= ~(layer0_out[9562] | layer0_out[9563]);
     layer1_out[889] <= ~layer0_out[7294];
     layer1_out[890] <= ~layer0_out[7971];
     layer1_out[891] <= ~layer0_out[315];
     layer1_out[892] <= ~layer0_out[9794] | layer0_out[9795];
     layer1_out[893] <= ~layer0_out[1300];
     layer1_out[894] <= 1'b0;
     layer1_out[895] <= ~layer0_out[11834] | layer0_out[11835];
     layer1_out[896] <= layer0_out[10312];
     layer1_out[897] <= layer0_out[8533] | layer0_out[8534];
     layer1_out[898] <= ~layer0_out[5658] | layer0_out[5659];
     layer1_out[899] <= layer0_out[4579] & ~layer0_out[4580];
     layer1_out[900] <= ~(layer0_out[5973] | layer0_out[5974]);
     layer1_out[901] <= layer0_out[6950];
     layer1_out[902] <= layer0_out[2724] & layer0_out[2725];
     layer1_out[903] <= layer0_out[8916];
     layer1_out[904] <= layer0_out[8783] & layer0_out[8784];
     layer1_out[905] <= ~layer0_out[9065] | layer0_out[9066];
     layer1_out[906] <= layer0_out[5107] | layer0_out[5108];
     layer1_out[907] <= layer0_out[3621] & layer0_out[3622];
     layer1_out[908] <= ~layer0_out[1476] | layer0_out[1475];
     layer1_out[909] <= ~layer0_out[4945] | layer0_out[4944];
     layer1_out[910] <= ~layer0_out[8947];
     layer1_out[911] <= ~layer0_out[7990];
     layer1_out[912] <= layer0_out[904];
     layer1_out[913] <= ~(layer0_out[5719] | layer0_out[5720]);
     layer1_out[914] <= 1'b0;
     layer1_out[915] <= layer0_out[2299] & ~layer0_out[2300];
     layer1_out[916] <= layer0_out[8724];
     layer1_out[917] <= layer0_out[11742] & ~layer0_out[11741];
     layer1_out[918] <= layer0_out[7164] ^ layer0_out[7165];
     layer1_out[919] <= layer0_out[5885] & ~layer0_out[5886];
     layer1_out[920] <= ~(layer0_out[2288] ^ layer0_out[2289]);
     layer1_out[921] <= ~layer0_out[88];
     layer1_out[922] <= ~layer0_out[1398] | layer0_out[1399];
     layer1_out[923] <= layer0_out[4274] & ~layer0_out[4273];
     layer1_out[924] <= ~layer0_out[9740] | layer0_out[9741];
     layer1_out[925] <= ~(layer0_out[7783] & layer0_out[7784]);
     layer1_out[926] <= layer0_out[3912] | layer0_out[3913];
     layer1_out[927] <= ~(layer0_out[9981] | layer0_out[9982]);
     layer1_out[928] <= layer0_out[8265] & ~layer0_out[8266];
     layer1_out[929] <= ~layer0_out[6953];
     layer1_out[930] <= layer0_out[7036] & layer0_out[7037];
     layer1_out[931] <= ~layer0_out[7888];
     layer1_out[932] <= ~layer0_out[8983] | layer0_out[8984];
     layer1_out[933] <= layer0_out[3766];
     layer1_out[934] <= layer0_out[3238];
     layer1_out[935] <= layer0_out[9688] ^ layer0_out[9689];
     layer1_out[936] <= layer0_out[10058] & layer0_out[10059];
     layer1_out[937] <= ~layer0_out[7845] | layer0_out[7846];
     layer1_out[938] <= ~(layer0_out[7726] | layer0_out[7727]);
     layer1_out[939] <= ~layer0_out[7995] | layer0_out[7994];
     layer1_out[940] <= ~(layer0_out[121] & layer0_out[122]);
     layer1_out[941] <= ~layer0_out[1444] | layer0_out[1443];
     layer1_out[942] <= layer0_out[3195];
     layer1_out[943] <= layer0_out[5913] & layer0_out[5914];
     layer1_out[944] <= layer0_out[3876];
     layer1_out[945] <= layer0_out[10830] & ~layer0_out[10829];
     layer1_out[946] <= layer0_out[784] | layer0_out[785];
     layer1_out[947] <= layer0_out[9840];
     layer1_out[948] <= 1'b1;
     layer1_out[949] <= layer0_out[6297];
     layer1_out[950] <= ~layer0_out[3569];
     layer1_out[951] <= layer0_out[7654];
     layer1_out[952] <= ~(layer0_out[11629] & layer0_out[11630]);
     layer1_out[953] <= layer0_out[8100] | layer0_out[8101];
     layer1_out[954] <= ~layer0_out[7067] | layer0_out[7068];
     layer1_out[955] <= layer0_out[713] & ~layer0_out[714];
     layer1_out[956] <= ~layer0_out[3657];
     layer1_out[957] <= layer0_out[1969];
     layer1_out[958] <= ~layer0_out[1725] | layer0_out[1726];
     layer1_out[959] <= ~layer0_out[962];
     layer1_out[960] <= layer0_out[11229];
     layer1_out[961] <= layer0_out[6437];
     layer1_out[962] <= layer0_out[7263] | layer0_out[7264];
     layer1_out[963] <= layer0_out[9530] & layer0_out[9531];
     layer1_out[964] <= layer0_out[7860] & layer0_out[7861];
     layer1_out[965] <= ~layer0_out[11292] | layer0_out[11293];
     layer1_out[966] <= layer0_out[11121] | layer0_out[11122];
     layer1_out[967] <= ~layer0_out[8445];
     layer1_out[968] <= 1'b0;
     layer1_out[969] <= ~layer0_out[9742];
     layer1_out[970] <= layer0_out[10346] & ~layer0_out[10345];
     layer1_out[971] <= ~layer0_out[9864];
     layer1_out[972] <= ~(layer0_out[9772] ^ layer0_out[9773]);
     layer1_out[973] <= layer0_out[167];
     layer1_out[974] <= ~layer0_out[4603];
     layer1_out[975] <= layer0_out[2186] & ~layer0_out[2187];
     layer1_out[976] <= layer0_out[5736] & ~layer0_out[5735];
     layer1_out[977] <= layer0_out[10767];
     layer1_out[978] <= ~layer0_out[4731];
     layer1_out[979] <= ~layer0_out[5639];
     layer1_out[980] <= 1'b0;
     layer1_out[981] <= ~layer0_out[8729] | layer0_out[8730];
     layer1_out[982] <= ~(layer0_out[6175] & layer0_out[6176]);
     layer1_out[983] <= layer0_out[1843] ^ layer0_out[1844];
     layer1_out[984] <= ~layer0_out[11197];
     layer1_out[985] <= layer0_out[10360] | layer0_out[10361];
     layer1_out[986] <= layer0_out[11506] & ~layer0_out[11505];
     layer1_out[987] <= ~(layer0_out[1276] | layer0_out[1277]);
     layer1_out[988] <= layer0_out[3896] & layer0_out[3897];
     layer1_out[989] <= layer0_out[544] & ~layer0_out[545];
     layer1_out[990] <= layer0_out[610];
     layer1_out[991] <= ~layer0_out[2161] | layer0_out[2162];
     layer1_out[992] <= layer0_out[1280];
     layer1_out[993] <= layer0_out[3295] & ~layer0_out[3296];
     layer1_out[994] <= layer0_out[6032] & ~layer0_out[6031];
     layer1_out[995] <= layer0_out[11444];
     layer1_out[996] <= ~layer0_out[8546] | layer0_out[8547];
     layer1_out[997] <= layer0_out[6162] & layer0_out[6163];
     layer1_out[998] <= layer0_out[6102] & ~layer0_out[6101];
     layer1_out[999] <= ~(layer0_out[5193] & layer0_out[5194]);
     layer1_out[1000] <= layer0_out[11884];
     layer1_out[1001] <= layer0_out[8749];
     layer1_out[1002] <= 1'b1;
     layer1_out[1003] <= ~layer0_out[2614];
     layer1_out[1004] <= ~layer0_out[3005];
     layer1_out[1005] <= layer0_out[302] | layer0_out[303];
     layer1_out[1006] <= 1'b1;
     layer1_out[1007] <= layer0_out[7854] & layer0_out[7855];
     layer1_out[1008] <= ~(layer0_out[2683] & layer0_out[2684]);
     layer1_out[1009] <= ~(layer0_out[9722] | layer0_out[9723]);
     layer1_out[1010] <= layer0_out[718] ^ layer0_out[719];
     layer1_out[1011] <= layer0_out[6149] | layer0_out[6150];
     layer1_out[1012] <= ~layer0_out[11187] | layer0_out[11186];
     layer1_out[1013] <= layer0_out[2561] | layer0_out[2562];
     layer1_out[1014] <= ~(layer0_out[4190] ^ layer0_out[4191]);
     layer1_out[1015] <= ~(layer0_out[4914] | layer0_out[4915]);
     layer1_out[1016] <= 1'b1;
     layer1_out[1017] <= layer0_out[3054] & ~layer0_out[3053];
     layer1_out[1018] <= layer0_out[128];
     layer1_out[1019] <= layer0_out[5149] & layer0_out[5150];
     layer1_out[1020] <= layer0_out[11516];
     layer1_out[1021] <= ~(layer0_out[9024] & layer0_out[9025]);
     layer1_out[1022] <= layer0_out[5413] & ~layer0_out[5412];
     layer1_out[1023] <= layer0_out[6806] ^ layer0_out[6807];
     layer1_out[1024] <= layer0_out[2446] | layer0_out[2447];
     layer1_out[1025] <= ~(layer0_out[8879] | layer0_out[8880]);
     layer1_out[1026] <= layer0_out[7093];
     layer1_out[1027] <= layer0_out[8487] | layer0_out[8488];
     layer1_out[1028] <= layer0_out[4827];
     layer1_out[1029] <= ~(layer0_out[5291] & layer0_out[5292]);
     layer1_out[1030] <= ~(layer0_out[3623] | layer0_out[3624]);
     layer1_out[1031] <= layer0_out[355];
     layer1_out[1032] <= ~layer0_out[2217];
     layer1_out[1033] <= 1'b1;
     layer1_out[1034] <= layer0_out[11272] & ~layer0_out[11273];
     layer1_out[1035] <= layer0_out[4881] ^ layer0_out[4882];
     layer1_out[1036] <= ~layer0_out[3131] | layer0_out[3132];
     layer1_out[1037] <= ~layer0_out[9324];
     layer1_out[1038] <= ~(layer0_out[9630] & layer0_out[9631]);
     layer1_out[1039] <= layer0_out[4246] & layer0_out[4247];
     layer1_out[1040] <= ~layer0_out[9983] | layer0_out[9984];
     layer1_out[1041] <= layer0_out[2402];
     layer1_out[1042] <= ~(layer0_out[9881] | layer0_out[9882]);
     layer1_out[1043] <= layer0_out[6317];
     layer1_out[1044] <= ~layer0_out[3134];
     layer1_out[1045] <= layer0_out[3124];
     layer1_out[1046] <= layer0_out[5485];
     layer1_out[1047] <= layer0_out[9829];
     layer1_out[1048] <= layer0_out[10917] | layer0_out[10918];
     layer1_out[1049] <= ~layer0_out[1185];
     layer1_out[1050] <= ~layer0_out[6185] | layer0_out[6184];
     layer1_out[1051] <= layer0_out[4237];
     layer1_out[1052] <= ~layer0_out[990] | layer0_out[989];
     layer1_out[1053] <= layer0_out[10025] ^ layer0_out[10026];
     layer1_out[1054] <= ~(layer0_out[7166] ^ layer0_out[7167]);
     layer1_out[1055] <= 1'b0;
     layer1_out[1056] <= ~layer0_out[2126] | layer0_out[2125];
     layer1_out[1057] <= ~(layer0_out[9533] | layer0_out[9534]);
     layer1_out[1058] <= ~(layer0_out[1179] ^ layer0_out[1180]);
     layer1_out[1059] <= layer0_out[10074];
     layer1_out[1060] <= ~layer0_out[1322];
     layer1_out[1061] <= ~layer0_out[2247] | layer0_out[2246];
     layer1_out[1062] <= ~layer0_out[4116];
     layer1_out[1063] <= layer0_out[4232];
     layer1_out[1064] <= ~layer0_out[1815];
     layer1_out[1065] <= ~layer0_out[1908];
     layer1_out[1066] <= layer0_out[6272];
     layer1_out[1067] <= layer0_out[6244] ^ layer0_out[6245];
     layer1_out[1068] <= ~layer0_out[8462] | layer0_out[8461];
     layer1_out[1069] <= ~(layer0_out[9372] & layer0_out[9373]);
     layer1_out[1070] <= ~(layer0_out[1316] | layer0_out[1317]);
     layer1_out[1071] <= ~(layer0_out[8478] & layer0_out[8479]);
     layer1_out[1072] <= layer0_out[2696] ^ layer0_out[2697];
     layer1_out[1073] <= ~(layer0_out[10453] | layer0_out[10454]);
     layer1_out[1074] <= layer0_out[4437];
     layer1_out[1075] <= ~(layer0_out[1054] | layer0_out[1055]);
     layer1_out[1076] <= layer0_out[4151];
     layer1_out[1077] <= ~layer0_out[8965] | layer0_out[8964];
     layer1_out[1078] <= layer0_out[2726] & ~layer0_out[2727];
     layer1_out[1079] <= ~layer0_out[7536];
     layer1_out[1080] <= ~layer0_out[9671];
     layer1_out[1081] <= 1'b0;
     layer1_out[1082] <= 1'b1;
     layer1_out[1083] <= layer0_out[2265] & ~layer0_out[2266];
     layer1_out[1084] <= ~layer0_out[3621] | layer0_out[3620];
     layer1_out[1085] <= ~(layer0_out[11103] & layer0_out[11104]);
     layer1_out[1086] <= ~layer0_out[9010];
     layer1_out[1087] <= layer0_out[11180] | layer0_out[11181];
     layer1_out[1088] <= ~(layer0_out[6511] & layer0_out[6512]);
     layer1_out[1089] <= ~(layer0_out[4621] | layer0_out[4622]);
     layer1_out[1090] <= ~layer0_out[1723];
     layer1_out[1091] <= 1'b0;
     layer1_out[1092] <= 1'b0;
     layer1_out[1093] <= ~(layer0_out[6819] & layer0_out[6820]);
     layer1_out[1094] <= ~layer0_out[6255] | layer0_out[6254];
     layer1_out[1095] <= ~layer0_out[3239] | layer0_out[3240];
     layer1_out[1096] <= layer0_out[6567] & layer0_out[6568];
     layer1_out[1097] <= layer0_out[9698];
     layer1_out[1098] <= layer0_out[7001];
     layer1_out[1099] <= ~layer0_out[6146] | layer0_out[6145];
     layer1_out[1100] <= ~layer0_out[1961] | layer0_out[1960];
     layer1_out[1101] <= layer0_out[2747] ^ layer0_out[2748];
     layer1_out[1102] <= layer0_out[2946];
     layer1_out[1103] <= ~(layer0_out[6753] & layer0_out[6754]);
     layer1_out[1104] <= ~(layer0_out[1414] & layer0_out[1415]);
     layer1_out[1105] <= ~(layer0_out[1940] & layer0_out[1941]);
     layer1_out[1106] <= layer0_out[2793] & ~layer0_out[2792];
     layer1_out[1107] <= 1'b0;
     layer1_out[1108] <= ~layer0_out[7281] | layer0_out[7282];
     layer1_out[1109] <= layer0_out[10395] & layer0_out[10396];
     layer1_out[1110] <= 1'b0;
     layer1_out[1111] <= layer0_out[7884] & layer0_out[7885];
     layer1_out[1112] <= ~layer0_out[8488];
     layer1_out[1113] <= layer0_out[4911];
     layer1_out[1114] <= layer0_out[1646] & ~layer0_out[1647];
     layer1_out[1115] <= ~(layer0_out[7949] & layer0_out[7950]);
     layer1_out[1116] <= 1'b0;
     layer1_out[1117] <= layer0_out[8578] & layer0_out[8579];
     layer1_out[1118] <= ~(layer0_out[5960] | layer0_out[5961]);
     layer1_out[1119] <= layer0_out[6377];
     layer1_out[1120] <= layer0_out[9406] & layer0_out[9407];
     layer1_out[1121] <= ~layer0_out[4667];
     layer1_out[1122] <= ~(layer0_out[6431] & layer0_out[6432]);
     layer1_out[1123] <= layer0_out[10223];
     layer1_out[1124] <= layer0_out[10004];
     layer1_out[1125] <= layer0_out[5337] & layer0_out[5338];
     layer1_out[1126] <= ~layer0_out[8803];
     layer1_out[1127] <= ~(layer0_out[6561] & layer0_out[6562]);
     layer1_out[1128] <= layer0_out[7034];
     layer1_out[1129] <= ~(layer0_out[2137] & layer0_out[2138]);
     layer1_out[1130] <= layer0_out[2950];
     layer1_out[1131] <= layer0_out[894] & ~layer0_out[893];
     layer1_out[1132] <= ~(layer0_out[5545] ^ layer0_out[5546]);
     layer1_out[1133] <= ~(layer0_out[8371] & layer0_out[8372]);
     layer1_out[1134] <= ~layer0_out[8693] | layer0_out[8694];
     layer1_out[1135] <= layer0_out[4956];
     layer1_out[1136] <= layer0_out[6569];
     layer1_out[1137] <= layer0_out[1135] & ~layer0_out[1136];
     layer1_out[1138] <= layer0_out[9870];
     layer1_out[1139] <= ~layer0_out[1504];
     layer1_out[1140] <= layer0_out[475];
     layer1_out[1141] <= layer0_out[4236] ^ layer0_out[4237];
     layer1_out[1142] <= ~(layer0_out[6973] & layer0_out[6974]);
     layer1_out[1143] <= layer0_out[9335];
     layer1_out[1144] <= layer0_out[8769] | layer0_out[8770];
     layer1_out[1145] <= layer0_out[4251];
     layer1_out[1146] <= layer0_out[7454];
     layer1_out[1147] <= layer0_out[5269];
     layer1_out[1148] <= layer0_out[6641] & ~layer0_out[6642];
     layer1_out[1149] <= layer0_out[2765] & ~layer0_out[2764];
     layer1_out[1150] <= ~layer0_out[8658] | layer0_out[8657];
     layer1_out[1151] <= layer0_out[5388];
     layer1_out[1152] <= layer0_out[11908] & layer0_out[11909];
     layer1_out[1153] <= ~(layer0_out[5039] | layer0_out[5040]);
     layer1_out[1154] <= ~layer0_out[319] | layer0_out[318];
     layer1_out[1155] <= layer0_out[981] & ~layer0_out[982];
     layer1_out[1156] <= ~layer0_out[808] | layer0_out[809];
     layer1_out[1157] <= ~(layer0_out[6423] | layer0_out[6424]);
     layer1_out[1158] <= ~layer0_out[7269];
     layer1_out[1159] <= layer0_out[11620] | layer0_out[11621];
     layer1_out[1160] <= layer0_out[11772];
     layer1_out[1161] <= ~layer0_out[4597];
     layer1_out[1162] <= ~layer0_out[1740] | layer0_out[1741];
     layer1_out[1163] <= layer0_out[6986];
     layer1_out[1164] <= layer0_out[5808];
     layer1_out[1165] <= layer0_out[6137] & ~layer0_out[6138];
     layer1_out[1166] <= layer0_out[687] & layer0_out[688];
     layer1_out[1167] <= ~(layer0_out[5164] | layer0_out[5165]);
     layer1_out[1168] <= layer0_out[9822];
     layer1_out[1169] <= ~(layer0_out[8435] & layer0_out[8436]);
     layer1_out[1170] <= ~layer0_out[4595];
     layer1_out[1171] <= ~layer0_out[3152];
     layer1_out[1172] <= layer0_out[2707] & ~layer0_out[2706];
     layer1_out[1173] <= 1'b1;
     layer1_out[1174] <= ~layer0_out[1546] | layer0_out[1547];
     layer1_out[1175] <= ~layer0_out[1482] | layer0_out[1483];
     layer1_out[1176] <= layer0_out[3259] ^ layer0_out[3260];
     layer1_out[1177] <= 1'b0;
     layer1_out[1178] <= ~(layer0_out[7386] | layer0_out[7387]);
     layer1_out[1179] <= 1'b0;
     layer1_out[1180] <= ~layer0_out[705] | layer0_out[706];
     layer1_out[1181] <= layer0_out[6993];
     layer1_out[1182] <= ~layer0_out[9564] | layer0_out[9565];
     layer1_out[1183] <= layer0_out[1053] & layer0_out[1054];
     layer1_out[1184] <= layer0_out[665] & ~layer0_out[666];
     layer1_out[1185] <= layer0_out[11751] & ~layer0_out[11752];
     layer1_out[1186] <= layer0_out[6537];
     layer1_out[1187] <= layer0_out[6706];
     layer1_out[1188] <= layer0_out[8421] & ~layer0_out[8422];
     layer1_out[1189] <= ~layer0_out[7574];
     layer1_out[1190] <= 1'b1;
     layer1_out[1191] <= layer0_out[3994];
     layer1_out[1192] <= layer0_out[1407];
     layer1_out[1193] <= ~layer0_out[920] | layer0_out[919];
     layer1_out[1194] <= ~(layer0_out[10953] & layer0_out[10954]);
     layer1_out[1195] <= layer0_out[8768];
     layer1_out[1196] <= layer0_out[11422] & ~layer0_out[11421];
     layer1_out[1197] <= layer0_out[1197] & ~layer0_out[1198];
     layer1_out[1198] <= ~layer0_out[3844] | layer0_out[3845];
     layer1_out[1199] <= layer0_out[11813] | layer0_out[11814];
     layer1_out[1200] <= layer0_out[4005] & layer0_out[4006];
     layer1_out[1201] <= layer0_out[4187];
     layer1_out[1202] <= ~(layer0_out[10356] & layer0_out[10357]);
     layer1_out[1203] <= layer0_out[10608] & layer0_out[10609];
     layer1_out[1204] <= ~layer0_out[106];
     layer1_out[1205] <= ~layer0_out[2739];
     layer1_out[1206] <= ~layer0_out[9721];
     layer1_out[1207] <= ~(layer0_out[10979] & layer0_out[10980]);
     layer1_out[1208] <= layer0_out[624];
     layer1_out[1209] <= ~layer0_out[164];
     layer1_out[1210] <= layer0_out[7697] & layer0_out[7698];
     layer1_out[1211] <= layer0_out[8770];
     layer1_out[1212] <= ~layer0_out[9952];
     layer1_out[1213] <= layer0_out[3092] ^ layer0_out[3093];
     layer1_out[1214] <= ~(layer0_out[8049] & layer0_out[8050]);
     layer1_out[1215] <= 1'b1;
     layer1_out[1216] <= 1'b1;
     layer1_out[1217] <= ~(layer0_out[10452] | layer0_out[10453]);
     layer1_out[1218] <= layer0_out[3527] ^ layer0_out[3528];
     layer1_out[1219] <= layer0_out[7647] & ~layer0_out[7648];
     layer1_out[1220] <= ~layer0_out[2398];
     layer1_out[1221] <= ~(layer0_out[9991] & layer0_out[9992]);
     layer1_out[1222] <= ~layer0_out[8549];
     layer1_out[1223] <= ~(layer0_out[7271] ^ layer0_out[7272]);
     layer1_out[1224] <= ~layer0_out[9962];
     layer1_out[1225] <= 1'b1;
     layer1_out[1226] <= layer0_out[9147];
     layer1_out[1227] <= ~(layer0_out[7231] ^ layer0_out[7232]);
     layer1_out[1228] <= layer0_out[10772] & ~layer0_out[10771];
     layer1_out[1229] <= layer0_out[358] & ~layer0_out[357];
     layer1_out[1230] <= ~(layer0_out[1138] ^ layer0_out[1139]);
     layer1_out[1231] <= layer0_out[5325] | layer0_out[5326];
     layer1_out[1232] <= 1'b1;
     layer1_out[1233] <= ~layer0_out[8591];
     layer1_out[1234] <= ~layer0_out[8453];
     layer1_out[1235] <= layer0_out[8270] | layer0_out[8271];
     layer1_out[1236] <= ~(layer0_out[8967] | layer0_out[8968]);
     layer1_out[1237] <= layer0_out[4198];
     layer1_out[1238] <= layer0_out[11304] ^ layer0_out[11305];
     layer1_out[1239] <= ~layer0_out[1436];
     layer1_out[1240] <= ~layer0_out[7784];
     layer1_out[1241] <= ~(layer0_out[6290] | layer0_out[6291]);
     layer1_out[1242] <= ~layer0_out[6955] | layer0_out[6954];
     layer1_out[1243] <= ~(layer0_out[471] | layer0_out[472]);
     layer1_out[1244] <= layer0_out[11013] & ~layer0_out[11014];
     layer1_out[1245] <= layer0_out[1770] & ~layer0_out[1771];
     layer1_out[1246] <= ~layer0_out[2434];
     layer1_out[1247] <= ~layer0_out[3942];
     layer1_out[1248] <= layer0_out[5650] & ~layer0_out[5649];
     layer1_out[1249] <= layer0_out[1351];
     layer1_out[1250] <= layer0_out[1795] | layer0_out[1796];
     layer1_out[1251] <= ~(layer0_out[8929] | layer0_out[8930]);
     layer1_out[1252] <= ~layer0_out[10276];
     layer1_out[1253] <= layer0_out[1521];
     layer1_out[1254] <= 1'b0;
     layer1_out[1255] <= layer0_out[5785] & ~layer0_out[5786];
     layer1_out[1256] <= layer0_out[3977] & ~layer0_out[3976];
     layer1_out[1257] <= ~layer0_out[7537];
     layer1_out[1258] <= layer0_out[3071] & ~layer0_out[3070];
     layer1_out[1259] <= ~(layer0_out[11195] | layer0_out[11196]);
     layer1_out[1260] <= ~(layer0_out[5646] ^ layer0_out[5647]);
     layer1_out[1261] <= layer0_out[3664];
     layer1_out[1262] <= ~(layer0_out[2060] & layer0_out[2061]);
     layer1_out[1263] <= ~layer0_out[5169] | layer0_out[5170];
     layer1_out[1264] <= layer0_out[574];
     layer1_out[1265] <= ~layer0_out[4609] | layer0_out[4610];
     layer1_out[1266] <= 1'b1;
     layer1_out[1267] <= layer0_out[8040];
     layer1_out[1268] <= ~layer0_out[8025];
     layer1_out[1269] <= ~layer0_out[8380];
     layer1_out[1270] <= 1'b1;
     layer1_out[1271] <= layer0_out[6811];
     layer1_out[1272] <= layer0_out[10008] & ~layer0_out[10007];
     layer1_out[1273] <= ~layer0_out[1491];
     layer1_out[1274] <= layer0_out[518] & layer0_out[519];
     layer1_out[1275] <= ~(layer0_out[1188] | layer0_out[1189]);
     layer1_out[1276] <= ~layer0_out[2887];
     layer1_out[1277] <= layer0_out[6289] & ~layer0_out[6288];
     layer1_out[1278] <= layer0_out[10895] | layer0_out[10896];
     layer1_out[1279] <= layer0_out[8973];
     layer1_out[1280] <= layer0_out[579] & ~layer0_out[578];
     layer1_out[1281] <= ~layer0_out[2447];
     layer1_out[1282] <= ~layer0_out[1313] | layer0_out[1312];
     layer1_out[1283] <= ~(layer0_out[9035] ^ layer0_out[9036]);
     layer1_out[1284] <= ~layer0_out[8682];
     layer1_out[1285] <= layer0_out[11758];
     layer1_out[1286] <= layer0_out[3730];
     layer1_out[1287] <= ~layer0_out[7708] | layer0_out[7707];
     layer1_out[1288] <= layer0_out[8352] & ~layer0_out[8353];
     layer1_out[1289] <= layer0_out[2031];
     layer1_out[1290] <= layer0_out[11744] | layer0_out[11745];
     layer1_out[1291] <= ~layer0_out[9840];
     layer1_out[1292] <= layer0_out[7992];
     layer1_out[1293] <= ~(layer0_out[11152] | layer0_out[11153]);
     layer1_out[1294] <= layer0_out[3062] | layer0_out[3063];
     layer1_out[1295] <= layer0_out[8537] & layer0_out[8538];
     layer1_out[1296] <= ~layer0_out[10899];
     layer1_out[1297] <= ~layer0_out[363];
     layer1_out[1298] <= ~layer0_out[9158] | layer0_out[9159];
     layer1_out[1299] <= layer0_out[233] & ~layer0_out[232];
     layer1_out[1300] <= layer0_out[241] & ~layer0_out[242];
     layer1_out[1301] <= layer0_out[10584] & ~layer0_out[10583];
     layer1_out[1302] <= layer0_out[6827] ^ layer0_out[6828];
     layer1_out[1303] <= layer0_out[9436];
     layer1_out[1304] <= ~layer0_out[2769] | layer0_out[2768];
     layer1_out[1305] <= 1'b1;
     layer1_out[1306] <= layer0_out[90] & ~layer0_out[91];
     layer1_out[1307] <= ~layer0_out[11419];
     layer1_out[1308] <= layer0_out[11549] & ~layer0_out[11548];
     layer1_out[1309] <= ~layer0_out[3974];
     layer1_out[1310] <= layer0_out[901];
     layer1_out[1311] <= ~(layer0_out[9715] ^ layer0_out[9716]);
     layer1_out[1312] <= ~(layer0_out[1710] & layer0_out[1711]);
     layer1_out[1313] <= layer0_out[10528] & ~layer0_out[10527];
     layer1_out[1314] <= 1'b1;
     layer1_out[1315] <= layer0_out[8000];
     layer1_out[1316] <= ~layer0_out[3150];
     layer1_out[1317] <= layer0_out[9648] & layer0_out[9649];
     layer1_out[1318] <= layer0_out[10465];
     layer1_out[1319] <= layer0_out[5529] & layer0_out[5530];
     layer1_out[1320] <= ~(layer0_out[2587] ^ layer0_out[2588]);
     layer1_out[1321] <= layer0_out[9284] & ~layer0_out[9283];
     layer1_out[1322] <= ~layer0_out[306];
     layer1_out[1323] <= ~(layer0_out[4637] ^ layer0_out[4638]);
     layer1_out[1324] <= layer0_out[11042] | layer0_out[11043];
     layer1_out[1325] <= ~(layer0_out[7659] ^ layer0_out[7660]);
     layer1_out[1326] <= ~(layer0_out[7682] | layer0_out[7683]);
     layer1_out[1327] <= layer0_out[11260];
     layer1_out[1328] <= layer0_out[7371];
     layer1_out[1329] <= ~layer0_out[6473];
     layer1_out[1330] <= layer0_out[11324];
     layer1_out[1331] <= layer0_out[9154] | layer0_out[9155];
     layer1_out[1332] <= 1'b0;
     layer1_out[1333] <= ~layer0_out[2712];
     layer1_out[1334] <= ~(layer0_out[3106] ^ layer0_out[3107]);
     layer1_out[1335] <= 1'b0;
     layer1_out[1336] <= ~layer0_out[11711];
     layer1_out[1337] <= ~layer0_out[11463];
     layer1_out[1338] <= ~(layer0_out[5438] & layer0_out[5439]);
     layer1_out[1339] <= ~layer0_out[7676];
     layer1_out[1340] <= ~layer0_out[6888];
     layer1_out[1341] <= layer0_out[3975];
     layer1_out[1342] <= layer0_out[3358];
     layer1_out[1343] <= layer0_out[118];
     layer1_out[1344] <= ~layer0_out[3759] | layer0_out[3760];
     layer1_out[1345] <= ~(layer0_out[5102] & layer0_out[5103]);
     layer1_out[1346] <= ~(layer0_out[5138] ^ layer0_out[5139]);
     layer1_out[1347] <= layer0_out[3393];
     layer1_out[1348] <= ~layer0_out[7770] | layer0_out[7771];
     layer1_out[1349] <= layer0_out[2853] & layer0_out[2854];
     layer1_out[1350] <= ~(layer0_out[3161] | layer0_out[3162]);
     layer1_out[1351] <= ~layer0_out[5206];
     layer1_out[1352] <= ~layer0_out[1160];
     layer1_out[1353] <= ~layer0_out[2695];
     layer1_out[1354] <= layer0_out[359];
     layer1_out[1355] <= ~layer0_out[5860] | layer0_out[5861];
     layer1_out[1356] <= ~layer0_out[2921] | layer0_out[2920];
     layer1_out[1357] <= ~layer0_out[7447];
     layer1_out[1358] <= layer0_out[9184];
     layer1_out[1359] <= ~layer0_out[791];
     layer1_out[1360] <= layer0_out[6138] | layer0_out[6139];
     layer1_out[1361] <= layer0_out[1497];
     layer1_out[1362] <= layer0_out[3131];
     layer1_out[1363] <= layer0_out[6526];
     layer1_out[1364] <= layer0_out[7343];
     layer1_out[1365] <= layer0_out[11822];
     layer1_out[1366] <= layer0_out[8998] & layer0_out[8999];
     layer1_out[1367] <= layer0_out[4448] & ~layer0_out[4447];
     layer1_out[1368] <= ~(layer0_out[6592] | layer0_out[6593]);
     layer1_out[1369] <= 1'b1;
     layer1_out[1370] <= layer0_out[3];
     layer1_out[1371] <= layer0_out[3609] & ~layer0_out[3610];
     layer1_out[1372] <= ~layer0_out[10082] | layer0_out[10081];
     layer1_out[1373] <= ~(layer0_out[8080] & layer0_out[8081]);
     layer1_out[1374] <= layer0_out[4328] & layer0_out[4329];
     layer1_out[1375] <= layer0_out[10286] & layer0_out[10287];
     layer1_out[1376] <= ~layer0_out[11522];
     layer1_out[1377] <= ~(layer0_out[10616] | layer0_out[10617]);
     layer1_out[1378] <= layer0_out[839] & ~layer0_out[840];
     layer1_out[1379] <= ~layer0_out[3223];
     layer1_out[1380] <= layer0_out[1336];
     layer1_out[1381] <= ~layer0_out[3649];
     layer1_out[1382] <= ~layer0_out[8060] | layer0_out[8061];
     layer1_out[1383] <= layer0_out[3608] | layer0_out[3609];
     layer1_out[1384] <= ~layer0_out[5420] | layer0_out[5421];
     layer1_out[1385] <= ~layer0_out[10489];
     layer1_out[1386] <= layer0_out[2422];
     layer1_out[1387] <= layer0_out[7537] ^ layer0_out[7538];
     layer1_out[1388] <= ~(layer0_out[8493] ^ layer0_out[8494]);
     layer1_out[1389] <= layer0_out[3177] ^ layer0_out[3178];
     layer1_out[1390] <= ~(layer0_out[3238] & layer0_out[3239]);
     layer1_out[1391] <= 1'b0;
     layer1_out[1392] <= 1'b1;
     layer1_out[1393] <= layer0_out[5141] | layer0_out[5142];
     layer1_out[1394] <= ~layer0_out[6025] | layer0_out[6024];
     layer1_out[1395] <= ~(layer0_out[8712] & layer0_out[8713]);
     layer1_out[1396] <= layer0_out[10703];
     layer1_out[1397] <= ~(layer0_out[1327] & layer0_out[1328]);
     layer1_out[1398] <= layer0_out[7085];
     layer1_out[1399] <= 1'b1;
     layer1_out[1400] <= ~(layer0_out[10612] ^ layer0_out[10613]);
     layer1_out[1401] <= ~layer0_out[3190];
     layer1_out[1402] <= ~layer0_out[7632] | layer0_out[7633];
     layer1_out[1403] <= ~layer0_out[1128];
     layer1_out[1404] <= layer0_out[6] & ~layer0_out[5];
     layer1_out[1405] <= ~layer0_out[9202];
     layer1_out[1406] <= ~layer0_out[5031];
     layer1_out[1407] <= layer0_out[1654] & ~layer0_out[1653];
     layer1_out[1408] <= ~(layer0_out[5498] & layer0_out[5499]);
     layer1_out[1409] <= layer0_out[1865] | layer0_out[1866];
     layer1_out[1410] <= layer0_out[11543] & ~layer0_out[11542];
     layer1_out[1411] <= ~(layer0_out[7168] & layer0_out[7169]);
     layer1_out[1412] <= layer0_out[8983] & ~layer0_out[8982];
     layer1_out[1413] <= ~layer0_out[5680] | layer0_out[5679];
     layer1_out[1414] <= ~(layer0_out[5084] & layer0_out[5085]);
     layer1_out[1415] <= layer0_out[9788] | layer0_out[9789];
     layer1_out[1416] <= ~(layer0_out[3825] ^ layer0_out[3826]);
     layer1_out[1417] <= layer0_out[3227] & ~layer0_out[3228];
     layer1_out[1418] <= ~layer0_out[9389];
     layer1_out[1419] <= layer0_out[5925] & ~layer0_out[5926];
     layer1_out[1420] <= ~layer0_out[3689];
     layer1_out[1421] <= layer0_out[4334] & ~layer0_out[4335];
     layer1_out[1422] <= ~layer0_out[2197] | layer0_out[2196];
     layer1_out[1423] <= layer0_out[2316] & ~layer0_out[2315];
     layer1_out[1424] <= layer0_out[2646] | layer0_out[2647];
     layer1_out[1425] <= layer0_out[3518] & layer0_out[3519];
     layer1_out[1426] <= ~layer0_out[2];
     layer1_out[1427] <= ~layer0_out[7023];
     layer1_out[1428] <= ~(layer0_out[6292] & layer0_out[6293]);
     layer1_out[1429] <= ~(layer0_out[441] | layer0_out[442]);
     layer1_out[1430] <= ~layer0_out[6057];
     layer1_out[1431] <= layer0_out[8314] & ~layer0_out[8315];
     layer1_out[1432] <= layer0_out[3943] & ~layer0_out[3944];
     layer1_out[1433] <= ~(layer0_out[5082] & layer0_out[5083]);
     layer1_out[1434] <= ~layer0_out[9585] | layer0_out[9584];
     layer1_out[1435] <= layer0_out[68] & ~layer0_out[67];
     layer1_out[1436] <= ~(layer0_out[1692] | layer0_out[1693]);
     layer1_out[1437] <= layer0_out[10870];
     layer1_out[1438] <= layer0_out[8566] | layer0_out[8567];
     layer1_out[1439] <= ~layer0_out[3776] | layer0_out[3775];
     layer1_out[1440] <= layer0_out[1282] ^ layer0_out[1283];
     layer1_out[1441] <= layer0_out[5615] & ~layer0_out[5614];
     layer1_out[1442] <= ~(layer0_out[7706] & layer0_out[7707]);
     layer1_out[1443] <= layer0_out[322];
     layer1_out[1444] <= ~layer0_out[7690];
     layer1_out[1445] <= layer0_out[11166];
     layer1_out[1446] <= layer0_out[4326];
     layer1_out[1447] <= ~(layer0_out[7695] | layer0_out[7696]);
     layer1_out[1448] <= ~layer0_out[1325];
     layer1_out[1449] <= ~(layer0_out[438] & layer0_out[439]);
     layer1_out[1450] <= layer0_out[9113] & ~layer0_out[9114];
     layer1_out[1451] <= ~layer0_out[858] | layer0_out[857];
     layer1_out[1452] <= layer0_out[10976];
     layer1_out[1453] <= layer0_out[8766] & ~layer0_out[8767];
     layer1_out[1454] <= ~layer0_out[7675];
     layer1_out[1455] <= layer0_out[9620];
     layer1_out[1456] <= layer0_out[9615] & layer0_out[9616];
     layer1_out[1457] <= layer0_out[3406] & ~layer0_out[3405];
     layer1_out[1458] <= ~layer0_out[5921] | layer0_out[5920];
     layer1_out[1459] <= ~layer0_out[8898] | layer0_out[8899];
     layer1_out[1460] <= ~layer0_out[1115] | layer0_out[1116];
     layer1_out[1461] <= ~layer0_out[28];
     layer1_out[1462] <= ~(layer0_out[2264] | layer0_out[2265]);
     layer1_out[1463] <= layer0_out[2481];
     layer1_out[1464] <= layer0_out[3251];
     layer1_out[1465] <= layer0_out[6635];
     layer1_out[1466] <= ~layer0_out[1727] | layer0_out[1726];
     layer1_out[1467] <= layer0_out[3909] & ~layer0_out[3910];
     layer1_out[1468] <= ~layer0_out[1135] | layer0_out[1134];
     layer1_out[1469] <= ~(layer0_out[9717] | layer0_out[9718]);
     layer1_out[1470] <= layer0_out[4125] & ~layer0_out[4124];
     layer1_out[1471] <= ~layer0_out[8380] | layer0_out[8381];
     layer1_out[1472] <= layer0_out[8341];
     layer1_out[1473] <= ~layer0_out[4037];
     layer1_out[1474] <= ~(layer0_out[8795] ^ layer0_out[8796]);
     layer1_out[1475] <= layer0_out[5925];
     layer1_out[1476] <= ~layer0_out[5988] | layer0_out[5987];
     layer1_out[1477] <= ~layer0_out[9851];
     layer1_out[1478] <= layer0_out[1076] & ~layer0_out[1077];
     layer1_out[1479] <= layer0_out[7042];
     layer1_out[1480] <= layer0_out[669] ^ layer0_out[670];
     layer1_out[1481] <= ~(layer0_out[1799] ^ layer0_out[1800]);
     layer1_out[1482] <= layer0_out[7507] & ~layer0_out[7508];
     layer1_out[1483] <= ~layer0_out[11365] | layer0_out[11364];
     layer1_out[1484] <= ~(layer0_out[6046] & layer0_out[6047]);
     layer1_out[1485] <= layer0_out[10076] & layer0_out[10077];
     layer1_out[1486] <= layer0_out[4836];
     layer1_out[1487] <= layer0_out[2327] ^ layer0_out[2328];
     layer1_out[1488] <= layer0_out[2606] ^ layer0_out[2607];
     layer1_out[1489] <= layer0_out[6025] | layer0_out[6026];
     layer1_out[1490] <= layer0_out[7632] & ~layer0_out[7631];
     layer1_out[1491] <= layer0_out[5506] | layer0_out[5507];
     layer1_out[1492] <= layer0_out[3718];
     layer1_out[1493] <= ~layer0_out[10561];
     layer1_out[1494] <= ~layer0_out[6060] | layer0_out[6059];
     layer1_out[1495] <= layer0_out[4482] & ~layer0_out[4483];
     layer1_out[1496] <= layer0_out[4441];
     layer1_out[1497] <= ~layer0_out[10974] | layer0_out[10975];
     layer1_out[1498] <= ~layer0_out[883];
     layer1_out[1499] <= layer0_out[7298];
     layer1_out[1500] <= ~layer0_out[6418];
     layer1_out[1501] <= layer0_out[8020];
     layer1_out[1502] <= layer0_out[3882];
     layer1_out[1503] <= ~layer0_out[8555] | layer0_out[8556];
     layer1_out[1504] <= layer0_out[5184];
     layer1_out[1505] <= layer0_out[2009] & ~layer0_out[2010];
     layer1_out[1506] <= ~layer0_out[11571];
     layer1_out[1507] <= layer0_out[1159] & layer0_out[1160];
     layer1_out[1508] <= ~layer0_out[6657] | layer0_out[6658];
     layer1_out[1509] <= layer0_out[9097];
     layer1_out[1510] <= ~layer0_out[2997] | layer0_out[2996];
     layer1_out[1511] <= layer0_out[1753];
     layer1_out[1512] <= ~layer0_out[987];
     layer1_out[1513] <= ~layer0_out[1331];
     layer1_out[1514] <= ~layer0_out[6094];
     layer1_out[1515] <= layer0_out[421] ^ layer0_out[422];
     layer1_out[1516] <= ~(layer0_out[8756] ^ layer0_out[8757]);
     layer1_out[1517] <= 1'b1;
     layer1_out[1518] <= ~layer0_out[5706];
     layer1_out[1519] <= ~(layer0_out[5608] ^ layer0_out[5609]);
     layer1_out[1520] <= ~layer0_out[3717] | layer0_out[3716];
     layer1_out[1521] <= layer0_out[8974] & layer0_out[8975];
     layer1_out[1522] <= layer0_out[11041];
     layer1_out[1523] <= ~layer0_out[11838];
     layer1_out[1524] <= ~(layer0_out[6719] & layer0_out[6720]);
     layer1_out[1525] <= ~(layer0_out[5718] & layer0_out[5719]);
     layer1_out[1526] <= layer0_out[5798];
     layer1_out[1527] <= layer0_out[11143];
     layer1_out[1528] <= ~layer0_out[10444] | layer0_out[10443];
     layer1_out[1529] <= layer0_out[10581] & ~layer0_out[10582];
     layer1_out[1530] <= ~layer0_out[7869];
     layer1_out[1531] <= layer0_out[2024] & ~layer0_out[2025];
     layer1_out[1532] <= ~layer0_out[5333] | layer0_out[5334];
     layer1_out[1533] <= layer0_out[7388] & ~layer0_out[7389];
     layer1_out[1534] <= ~(layer0_out[10338] & layer0_out[10339]);
     layer1_out[1535] <= ~layer0_out[4495] | layer0_out[4496];
     layer1_out[1536] <= layer0_out[11618];
     layer1_out[1537] <= layer0_out[7992];
     layer1_out[1538] <= layer0_out[2159] ^ layer0_out[2160];
     layer1_out[1539] <= ~(layer0_out[5246] & layer0_out[5247]);
     layer1_out[1540] <= layer0_out[8608];
     layer1_out[1541] <= layer0_out[2662];
     layer1_out[1542] <= layer0_out[5898] & layer0_out[5899];
     layer1_out[1543] <= ~layer0_out[10780] | layer0_out[10779];
     layer1_out[1544] <= layer0_out[7960];
     layer1_out[1545] <= ~layer0_out[8311] | layer0_out[8312];
     layer1_out[1546] <= ~layer0_out[2374];
     layer1_out[1547] <= layer0_out[2534] | layer0_out[2535];
     layer1_out[1548] <= layer0_out[6454] & ~layer0_out[6455];
     layer1_out[1549] <= layer0_out[2558] & layer0_out[2559];
     layer1_out[1550] <= ~layer0_out[3740];
     layer1_out[1551] <= layer0_out[5762] | layer0_out[5763];
     layer1_out[1552] <= ~layer0_out[20];
     layer1_out[1553] <= ~layer0_out[4985];
     layer1_out[1554] <= layer0_out[11397] | layer0_out[11398];
     layer1_out[1555] <= ~(layer0_out[9848] | layer0_out[9849]);
     layer1_out[1556] <= ~(layer0_out[9990] & layer0_out[9991]);
     layer1_out[1557] <= 1'b0;
     layer1_out[1558] <= layer0_out[5376] & layer0_out[5377];
     layer1_out[1559] <= 1'b0;
     layer1_out[1560] <= layer0_out[3830] & ~layer0_out[3829];
     layer1_out[1561] <= layer0_out[4135] & layer0_out[4136];
     layer1_out[1562] <= layer0_out[10487] ^ layer0_out[10488];
     layer1_out[1563] <= layer0_out[6446] | layer0_out[6447];
     layer1_out[1564] <= layer0_out[4079];
     layer1_out[1565] <= ~layer0_out[9115] | layer0_out[9114];
     layer1_out[1566] <= 1'b1;
     layer1_out[1567] <= ~layer0_out[10304] | layer0_out[10303];
     layer1_out[1568] <= layer0_out[4714];
     layer1_out[1569] <= ~(layer0_out[6411] | layer0_out[6412]);
     layer1_out[1570] <= layer0_out[11603];
     layer1_out[1571] <= layer0_out[9664] & layer0_out[9665];
     layer1_out[1572] <= ~layer0_out[1967];
     layer1_out[1573] <= ~layer0_out[9829];
     layer1_out[1574] <= ~layer0_out[6398];
     layer1_out[1575] <= layer0_out[11422] & layer0_out[11423];
     layer1_out[1576] <= ~(layer0_out[6427] & layer0_out[6428]);
     layer1_out[1577] <= layer0_out[4712];
     layer1_out[1578] <= ~layer0_out[2581] | layer0_out[2580];
     layer1_out[1579] <= layer0_out[3769];
     layer1_out[1580] <= ~(layer0_out[10941] & layer0_out[10942]);
     layer1_out[1581] <= layer0_out[4059] & layer0_out[4060];
     layer1_out[1582] <= layer0_out[4433] | layer0_out[4434];
     layer1_out[1583] <= ~(layer0_out[11094] | layer0_out[11095]);
     layer1_out[1584] <= ~(layer0_out[3550] & layer0_out[3551]);
     layer1_out[1585] <= layer0_out[8267];
     layer1_out[1586] <= ~layer0_out[1629] | layer0_out[1630];
     layer1_out[1587] <= ~layer0_out[4669];
     layer1_out[1588] <= ~(layer0_out[4684] | layer0_out[4685]);
     layer1_out[1589] <= ~layer0_out[9272];
     layer1_out[1590] <= layer0_out[8881] | layer0_out[8882];
     layer1_out[1591] <= layer0_out[7225] ^ layer0_out[7226];
     layer1_out[1592] <= ~layer0_out[4435];
     layer1_out[1593] <= ~layer0_out[1461];
     layer1_out[1594] <= ~layer0_out[7255];
     layer1_out[1595] <= layer0_out[5139];
     layer1_out[1596] <= layer0_out[2032] | layer0_out[2033];
     layer1_out[1597] <= layer0_out[1260] & ~layer0_out[1259];
     layer1_out[1598] <= layer0_out[9979];
     layer1_out[1599] <= ~layer0_out[11912] | layer0_out[11913];
     layer1_out[1600] <= ~layer0_out[5255] | layer0_out[5256];
     layer1_out[1601] <= ~layer0_out[5062];
     layer1_out[1602] <= ~layer0_out[1586];
     layer1_out[1603] <= layer0_out[8910];
     layer1_out[1604] <= layer0_out[172] | layer0_out[173];
     layer1_out[1605] <= ~(layer0_out[4185] & layer0_out[4186]);
     layer1_out[1606] <= layer0_out[3870] & ~layer0_out[3871];
     layer1_out[1607] <= layer0_out[7443];
     layer1_out[1608] <= ~(layer0_out[2883] & layer0_out[2884]);
     layer1_out[1609] <= layer0_out[3209];
     layer1_out[1610] <= layer0_out[6873];
     layer1_out[1611] <= ~layer0_out[11542] | layer0_out[11541];
     layer1_out[1612] <= layer0_out[8103] & ~layer0_out[8102];
     layer1_out[1613] <= ~layer0_out[6984];
     layer1_out[1614] <= ~layer0_out[1790] | layer0_out[1791];
     layer1_out[1615] <= layer0_out[9985] & ~layer0_out[9986];
     layer1_out[1616] <= ~layer0_out[428] | layer0_out[429];
     layer1_out[1617] <= ~layer0_out[9162];
     layer1_out[1618] <= layer0_out[2591] & layer0_out[2592];
     layer1_out[1619] <= layer0_out[4669] & ~layer0_out[4668];
     layer1_out[1620] <= layer0_out[5655] & layer0_out[5656];
     layer1_out[1621] <= ~layer0_out[8474] | layer0_out[8473];
     layer1_out[1622] <= ~layer0_out[3125] | layer0_out[3126];
     layer1_out[1623] <= ~(layer0_out[3707] & layer0_out[3708]);
     layer1_out[1624] <= layer0_out[10693] & layer0_out[10694];
     layer1_out[1625] <= ~layer0_out[3471];
     layer1_out[1626] <= layer0_out[2293] ^ layer0_out[2294];
     layer1_out[1627] <= ~layer0_out[267];
     layer1_out[1628] <= layer0_out[2382] & ~layer0_out[2381];
     layer1_out[1629] <= layer0_out[8984] & ~layer0_out[8985];
     layer1_out[1630] <= layer0_out[3082] & layer0_out[3083];
     layer1_out[1631] <= ~layer0_out[10234] | layer0_out[10233];
     layer1_out[1632] <= layer0_out[1210];
     layer1_out[1633] <= ~layer0_out[10679];
     layer1_out[1634] <= ~layer0_out[9746];
     layer1_out[1635] <= ~layer0_out[6457] | layer0_out[6458];
     layer1_out[1636] <= layer0_out[6097] & ~layer0_out[6096];
     layer1_out[1637] <= layer0_out[11037] ^ layer0_out[11038];
     layer1_out[1638] <= 1'b0;
     layer1_out[1639] <= ~layer0_out[120] | layer0_out[119];
     layer1_out[1640] <= ~layer0_out[9067];
     layer1_out[1641] <= layer0_out[378];
     layer1_out[1642] <= layer0_out[7954] & ~layer0_out[7953];
     layer1_out[1643] <= layer0_out[4529] & ~layer0_out[4530];
     layer1_out[1644] <= ~layer0_out[4078] | layer0_out[4079];
     layer1_out[1645] <= ~(layer0_out[2652] ^ layer0_out[2653]);
     layer1_out[1646] <= layer0_out[3502];
     layer1_out[1647] <= 1'b0;
     layer1_out[1648] <= layer0_out[6896];
     layer1_out[1649] <= layer0_out[891];
     layer1_out[1650] <= layer0_out[10186];
     layer1_out[1651] <= layer0_out[3753];
     layer1_out[1652] <= layer0_out[7123] & layer0_out[7124];
     layer1_out[1653] <= layer0_out[8233];
     layer1_out[1654] <= ~layer0_out[6814] | layer0_out[6815];
     layer1_out[1655] <= layer0_out[11822];
     layer1_out[1656] <= layer0_out[3599];
     layer1_out[1657] <= ~layer0_out[8327] | layer0_out[8328];
     layer1_out[1658] <= ~(layer0_out[3491] & layer0_out[3492]);
     layer1_out[1659] <= 1'b1;
     layer1_out[1660] <= ~layer0_out[9608] | layer0_out[9607];
     layer1_out[1661] <= layer0_out[7901] & ~layer0_out[7902];
     layer1_out[1662] <= layer0_out[660];
     layer1_out[1663] <= ~layer0_out[10283] | layer0_out[10282];
     layer1_out[1664] <= 1'b1;
     layer1_out[1665] <= ~layer0_out[7378];
     layer1_out[1666] <= ~layer0_out[10170];
     layer1_out[1667] <= layer0_out[10235];
     layer1_out[1668] <= layer0_out[6678] & ~layer0_out[6679];
     layer1_out[1669] <= layer0_out[10995];
     layer1_out[1670] <= layer0_out[2776];
     layer1_out[1671] <= ~layer0_out[10239] | layer0_out[10238];
     layer1_out[1672] <= 1'b1;
     layer1_out[1673] <= layer0_out[315] | layer0_out[316];
     layer1_out[1674] <= 1'b0;
     layer1_out[1675] <= ~(layer0_out[991] | layer0_out[992]);
     layer1_out[1676] <= ~layer0_out[5523] | layer0_out[5524];
     layer1_out[1677] <= ~layer0_out[8089];
     layer1_out[1678] <= ~(layer0_out[7849] & layer0_out[7850]);
     layer1_out[1679] <= ~layer0_out[9729] | layer0_out[9728];
     layer1_out[1680] <= ~(layer0_out[1400] ^ layer0_out[1401]);
     layer1_out[1681] <= ~(layer0_out[9343] | layer0_out[9344]);
     layer1_out[1682] <= layer0_out[6880];
     layer1_out[1683] <= ~(layer0_out[670] ^ layer0_out[671]);
     layer1_out[1684] <= layer0_out[3530] & ~layer0_out[3531];
     layer1_out[1685] <= ~(layer0_out[9104] | layer0_out[9105]);
     layer1_out[1686] <= 1'b1;
     layer1_out[1687] <= ~(layer0_out[7083] | layer0_out[7084]);
     layer1_out[1688] <= layer0_out[7370] & ~layer0_out[7369];
     layer1_out[1689] <= 1'b1;
     layer1_out[1690] <= layer0_out[2093];
     layer1_out[1691] <= ~layer0_out[4911];
     layer1_out[1692] <= 1'b1;
     layer1_out[1693] <= ~(layer0_out[11200] ^ layer0_out[11201]);
     layer1_out[1694] <= ~layer0_out[5473];
     layer1_out[1695] <= 1'b1;
     layer1_out[1696] <= layer0_out[6160] | layer0_out[6161];
     layer1_out[1697] <= ~(layer0_out[4067] & layer0_out[4068]);
     layer1_out[1698] <= 1'b0;
     layer1_out[1699] <= layer0_out[6105];
     layer1_out[1700] <= layer0_out[140];
     layer1_out[1701] <= ~layer0_out[11947] | layer0_out[11948];
     layer1_out[1702] <= layer0_out[5934] & ~layer0_out[5935];
     layer1_out[1703] <= ~(layer0_out[9427] | layer0_out[9428]);
     layer1_out[1704] <= ~layer0_out[10708];
     layer1_out[1705] <= ~layer0_out[8423];
     layer1_out[1706] <= ~(layer0_out[6929] | layer0_out[6930]);
     layer1_out[1707] <= 1'b0;
     layer1_out[1708] <= ~layer0_out[9229];
     layer1_out[1709] <= layer0_out[2890] | layer0_out[2891];
     layer1_out[1710] <= ~layer0_out[8159];
     layer1_out[1711] <= layer0_out[5692] & layer0_out[5693];
     layer1_out[1712] <= layer0_out[581];
     layer1_out[1713] <= layer0_out[7367];
     layer1_out[1714] <= ~(layer0_out[3] | layer0_out[4]);
     layer1_out[1715] <= layer0_out[855] & ~layer0_out[856];
     layer1_out[1716] <= layer0_out[2660] & layer0_out[2661];
     layer1_out[1717] <= ~layer0_out[3851];
     layer1_out[1718] <= ~layer0_out[699] | layer0_out[700];
     layer1_out[1719] <= ~(layer0_out[10205] & layer0_out[10206]);
     layer1_out[1720] <= 1'b0;
     layer1_out[1721] <= ~(layer0_out[6835] | layer0_out[6836]);
     layer1_out[1722] <= ~layer0_out[9766] | layer0_out[9767];
     layer1_out[1723] <= layer0_out[5921];
     layer1_out[1724] <= layer0_out[1045];
     layer1_out[1725] <= layer0_out[5392] | layer0_out[5393];
     layer1_out[1726] <= layer0_out[5554] ^ layer0_out[5555];
     layer1_out[1727] <= layer0_out[3966];
     layer1_out[1728] <= layer0_out[9782] & ~layer0_out[9781];
     layer1_out[1729] <= ~(layer0_out[9371] & layer0_out[9372]);
     layer1_out[1730] <= layer0_out[825] & layer0_out[826];
     layer1_out[1731] <= layer0_out[5843] | layer0_out[5844];
     layer1_out[1732] <= ~layer0_out[2968];
     layer1_out[1733] <= ~(layer0_out[8234] ^ layer0_out[8235]);
     layer1_out[1734] <= ~layer0_out[10193];
     layer1_out[1735] <= ~layer0_out[3662] | layer0_out[3663];
     layer1_out[1736] <= layer0_out[6459] & ~layer0_out[6458];
     layer1_out[1737] <= layer0_out[2519];
     layer1_out[1738] <= ~layer0_out[7221];
     layer1_out[1739] <= layer0_out[3021] & layer0_out[3022];
     layer1_out[1740] <= layer0_out[9164];
     layer1_out[1741] <= ~(layer0_out[10462] | layer0_out[10463]);
     layer1_out[1742] <= layer0_out[7273];
     layer1_out[1743] <= layer0_out[2807] & ~layer0_out[2806];
     layer1_out[1744] <= ~(layer0_out[11321] & layer0_out[11322]);
     layer1_out[1745] <= ~(layer0_out[456] & layer0_out[457]);
     layer1_out[1746] <= ~layer0_out[9490];
     layer1_out[1747] <= layer0_out[4653];
     layer1_out[1748] <= layer0_out[216] & ~layer0_out[215];
     layer1_out[1749] <= layer0_out[11015] & ~layer0_out[11014];
     layer1_out[1750] <= layer0_out[654];
     layer1_out[1751] <= ~layer0_out[8403] | layer0_out[8402];
     layer1_out[1752] <= ~layer0_out[7163];
     layer1_out[1753] <= 1'b1;
     layer1_out[1754] <= layer0_out[2420] | layer0_out[2421];
     layer1_out[1755] <= ~layer0_out[2204] | layer0_out[2205];
     layer1_out[1756] <= layer0_out[3564] & ~layer0_out[3565];
     layer1_out[1757] <= layer0_out[8365] ^ layer0_out[8366];
     layer1_out[1758] <= ~layer0_out[2336];
     layer1_out[1759] <= 1'b1;
     layer1_out[1760] <= ~layer0_out[10992] | layer0_out[10993];
     layer1_out[1761] <= layer0_out[5500] & ~layer0_out[5501];
     layer1_out[1762] <= ~(layer0_out[11021] ^ layer0_out[11022]);
     layer1_out[1763] <= layer0_out[7985];
     layer1_out[1764] <= ~layer0_out[3371];
     layer1_out[1765] <= layer0_out[8833];
     layer1_out[1766] <= ~layer0_out[872];
     layer1_out[1767] <= layer0_out[9055];
     layer1_out[1768] <= layer0_out[550] & ~layer0_out[549];
     layer1_out[1769] <= layer0_out[6421] & ~layer0_out[6420];
     layer1_out[1770] <= layer0_out[6980];
     layer1_out[1771] <= layer0_out[4833];
     layer1_out[1772] <= ~layer0_out[9657];
     layer1_out[1773] <= ~layer0_out[7611];
     layer1_out[1774] <= layer0_out[4393];
     layer1_out[1775] <= layer0_out[7771] & ~layer0_out[7772];
     layer1_out[1776] <= layer0_out[3105] | layer0_out[3106];
     layer1_out[1777] <= ~(layer0_out[11818] & layer0_out[11819]);
     layer1_out[1778] <= layer0_out[9494] & ~layer0_out[9495];
     layer1_out[1779] <= layer0_out[3690] & layer0_out[3691];
     layer1_out[1780] <= ~layer0_out[3945];
     layer1_out[1781] <= layer0_out[11843] & layer0_out[11844];
     layer1_out[1782] <= ~layer0_out[4135];
     layer1_out[1783] <= ~layer0_out[1650] | layer0_out[1651];
     layer1_out[1784] <= layer0_out[6527] ^ layer0_out[6528];
     layer1_out[1785] <= layer0_out[6880] | layer0_out[6881];
     layer1_out[1786] <= layer0_out[10039];
     layer1_out[1787] <= layer0_out[6415];
     layer1_out[1788] <= layer0_out[10067] | layer0_out[10068];
     layer1_out[1789] <= ~layer0_out[11184] | layer0_out[11185];
     layer1_out[1790] <= ~layer0_out[3074] | layer0_out[3073];
     layer1_out[1791] <= layer0_out[53] & ~layer0_out[54];
     layer1_out[1792] <= layer0_out[7969];
     layer1_out[1793] <= layer0_out[11335] & ~layer0_out[11334];
     layer1_out[1794] <= 1'b0;
     layer1_out[1795] <= layer0_out[6864];
     layer1_out[1796] <= layer0_out[3758];
     layer1_out[1797] <= ~(layer0_out[8798] & layer0_out[8799]);
     layer1_out[1798] <= layer0_out[9843];
     layer1_out[1799] <= ~layer0_out[4005];
     layer1_out[1800] <= layer0_out[1447] | layer0_out[1448];
     layer1_out[1801] <= layer0_out[776] | layer0_out[777];
     layer1_out[1802] <= ~layer0_out[4140];
     layer1_out[1803] <= ~layer0_out[2066];
     layer1_out[1804] <= ~layer0_out[8038];
     layer1_out[1805] <= layer0_out[3452] & ~layer0_out[3453];
     layer1_out[1806] <= layer0_out[4470];
     layer1_out[1807] <= ~(layer0_out[6088] | layer0_out[6089]);
     layer1_out[1808] <= layer0_out[6988] & ~layer0_out[6989];
     layer1_out[1809] <= ~(layer0_out[1674] | layer0_out[1675]);
     layer1_out[1810] <= ~layer0_out[1559];
     layer1_out[1811] <= layer0_out[5548] & ~layer0_out[5547];
     layer1_out[1812] <= 1'b1;
     layer1_out[1813] <= ~layer0_out[11665] | layer0_out[11666];
     layer1_out[1814] <= ~layer0_out[7839] | layer0_out[7838];
     layer1_out[1815] <= ~layer0_out[8867] | layer0_out[8866];
     layer1_out[1816] <= 1'b1;
     layer1_out[1817] <= layer0_out[5251];
     layer1_out[1818] <= ~(layer0_out[8199] & layer0_out[8200]);
     layer1_out[1819] <= layer0_out[3358];
     layer1_out[1820] <= layer0_out[2645] ^ layer0_out[2646];
     layer1_out[1821] <= layer0_out[2690] & ~layer0_out[2691];
     layer1_out[1822] <= ~(layer0_out[2126] & layer0_out[2127]);
     layer1_out[1823] <= ~(layer0_out[3243] ^ layer0_out[3244]);
     layer1_out[1824] <= ~(layer0_out[6142] | layer0_out[6143]);
     layer1_out[1825] <= ~(layer0_out[5672] & layer0_out[5673]);
     layer1_out[1826] <= ~layer0_out[10186] | layer0_out[10185];
     layer1_out[1827] <= ~(layer0_out[479] & layer0_out[480]);
     layer1_out[1828] <= layer0_out[9171] & layer0_out[9172];
     layer1_out[1829] <= layer0_out[1558] ^ layer0_out[1559];
     layer1_out[1830] <= ~layer0_out[9151] | layer0_out[9150];
     layer1_out[1831] <= layer0_out[5802] | layer0_out[5803];
     layer1_out[1832] <= layer0_out[8115] & ~layer0_out[8116];
     layer1_out[1833] <= layer0_out[9095];
     layer1_out[1834] <= ~layer0_out[2272] | layer0_out[2271];
     layer1_out[1835] <= layer0_out[4578] & ~layer0_out[4577];
     layer1_out[1836] <= ~(layer0_out[9412] & layer0_out[9413]);
     layer1_out[1837] <= ~(layer0_out[8593] | layer0_out[8594]);
     layer1_out[1838] <= ~layer0_out[9129];
     layer1_out[1839] <= layer0_out[1902] ^ layer0_out[1903];
     layer1_out[1840] <= layer0_out[6283] & layer0_out[6284];
     layer1_out[1841] <= ~layer0_out[2264] | layer0_out[2263];
     layer1_out[1842] <= layer0_out[8231];
     layer1_out[1843] <= layer0_out[10731] | layer0_out[10732];
     layer1_out[1844] <= layer0_out[4282] & ~layer0_out[4281];
     layer1_out[1845] <= ~layer0_out[2904] | layer0_out[2903];
     layer1_out[1846] <= layer0_out[11294] ^ layer0_out[11295];
     layer1_out[1847] <= ~layer0_out[2236];
     layer1_out[1848] <= layer0_out[8526] ^ layer0_out[8527];
     layer1_out[1849] <= ~layer0_out[8502];
     layer1_out[1850] <= ~layer0_out[628];
     layer1_out[1851] <= ~layer0_out[4590] | layer0_out[4589];
     layer1_out[1852] <= ~layer0_out[1390];
     layer1_out[1853] <= ~layer0_out[9236];
     layer1_out[1854] <= ~layer0_out[8750];
     layer1_out[1855] <= layer0_out[7165] & ~layer0_out[7166];
     layer1_out[1856] <= layer0_out[1597] & layer0_out[1598];
     layer1_out[1857] <= ~layer0_out[2380] | layer0_out[2379];
     layer1_out[1858] <= layer0_out[11485] & ~layer0_out[11486];
     layer1_out[1859] <= layer0_out[5893];
     layer1_out[1860] <= layer0_out[1348];
     layer1_out[1861] <= 1'b1;
     layer1_out[1862] <= ~layer0_out[3124];
     layer1_out[1863] <= layer0_out[11234];
     layer1_out[1864] <= ~layer0_out[11916];
     layer1_out[1865] <= ~layer0_out[3480];
     layer1_out[1866] <= ~(layer0_out[7158] | layer0_out[7159]);
     layer1_out[1867] <= layer0_out[9447] & layer0_out[9448];
     layer1_out[1868] <= ~layer0_out[882];
     layer1_out[1869] <= layer0_out[3875];
     layer1_out[1870] <= ~layer0_out[6967] | layer0_out[6966];
     layer1_out[1871] <= layer0_out[908] & ~layer0_out[907];
     layer1_out[1872] <= layer0_out[87] & ~layer0_out[88];
     layer1_out[1873] <= ~(layer0_out[9330] & layer0_out[9331]);
     layer1_out[1874] <= 1'b1;
     layer1_out[1875] <= layer0_out[8741];
     layer1_out[1876] <= layer0_out[6022];
     layer1_out[1877] <= ~layer0_out[7554];
     layer1_out[1878] <= ~(layer0_out[5314] ^ layer0_out[5315]);
     layer1_out[1879] <= layer0_out[8158] & ~layer0_out[8157];
     layer1_out[1880] <= ~layer0_out[9164];
     layer1_out[1881] <= layer0_out[9964];
     layer1_out[1882] <= layer0_out[820];
     layer1_out[1883] <= ~(layer0_out[7938] | layer0_out[7939]);
     layer1_out[1884] <= ~layer0_out[11460];
     layer1_out[1885] <= ~layer0_out[5414] | layer0_out[5415];
     layer1_out[1886] <= layer0_out[11452] & ~layer0_out[11453];
     layer1_out[1887] <= layer0_out[3650] & layer0_out[3651];
     layer1_out[1888] <= layer0_out[11231] | layer0_out[11232];
     layer1_out[1889] <= layer0_out[2146];
     layer1_out[1890] <= ~layer0_out[4930] | layer0_out[4929];
     layer1_out[1891] <= ~layer0_out[11433];
     layer1_out[1892] <= layer0_out[2515];
     layer1_out[1893] <= ~(layer0_out[2548] | layer0_out[2549]);
     layer1_out[1894] <= ~layer0_out[7661];
     layer1_out[1895] <= ~(layer0_out[7819] ^ layer0_out[7820]);
     layer1_out[1896] <= layer0_out[149] & layer0_out[150];
     layer1_out[1897] <= ~(layer0_out[7097] | layer0_out[7098]);
     layer1_out[1898] <= ~layer0_out[6441];
     layer1_out[1899] <= layer0_out[1807] | layer0_out[1808];
     layer1_out[1900] <= ~layer0_out[1948];
     layer1_out[1901] <= layer0_out[329];
     layer1_out[1902] <= layer0_out[7212];
     layer1_out[1903] <= layer0_out[1946];
     layer1_out[1904] <= ~layer0_out[3550];
     layer1_out[1905] <= layer0_out[11155];
     layer1_out[1906] <= layer0_out[10618] & ~layer0_out[10617];
     layer1_out[1907] <= ~(layer0_out[4220] | layer0_out[4221]);
     layer1_out[1908] <= layer0_out[1024];
     layer1_out[1909] <= layer0_out[430] & ~layer0_out[429];
     layer1_out[1910] <= layer0_out[4129];
     layer1_out[1911] <= layer0_out[8354] & ~layer0_out[8355];
     layer1_out[1912] <= ~layer0_out[9282] | layer0_out[9281];
     layer1_out[1913] <= layer0_out[5416];
     layer1_out[1914] <= layer0_out[11446] & layer0_out[11447];
     layer1_out[1915] <= 1'b1;
     layer1_out[1916] <= ~layer0_out[10714] | layer0_out[10713];
     layer1_out[1917] <= layer0_out[6125];
     layer1_out[1918] <= ~(layer0_out[2106] & layer0_out[2107]);
     layer1_out[1919] <= layer0_out[9876] & ~layer0_out[9875];
     layer1_out[1920] <= layer0_out[7685] & ~layer0_out[7686];
     layer1_out[1921] <= layer0_out[8973];
     layer1_out[1922] <= 1'b1;
     layer1_out[1923] <= ~layer0_out[1629] | layer0_out[1628];
     layer1_out[1924] <= 1'b1;
     layer1_out[1925] <= ~layer0_out[4399];
     layer1_out[1926] <= ~(layer0_out[6382] ^ layer0_out[6383]);
     layer1_out[1927] <= layer0_out[8753];
     layer1_out[1928] <= layer0_out[11212] & ~layer0_out[11213];
     layer1_out[1929] <= ~layer0_out[536] | layer0_out[535];
     layer1_out[1930] <= layer0_out[7448] & ~layer0_out[7449];
     layer1_out[1931] <= layer0_out[9815] ^ layer0_out[9816];
     layer1_out[1932] <= ~(layer0_out[2802] ^ layer0_out[2803]);
     layer1_out[1933] <= ~(layer0_out[11582] & layer0_out[11583]);
     layer1_out[1934] <= layer0_out[11409] & layer0_out[11410];
     layer1_out[1935] <= layer0_out[4069] | layer0_out[4070];
     layer1_out[1936] <= ~layer0_out[10123] | layer0_out[10122];
     layer1_out[1937] <= layer0_out[5833] & ~layer0_out[5834];
     layer1_out[1938] <= layer0_out[9719] & ~layer0_out[9718];
     layer1_out[1939] <= ~(layer0_out[9434] & layer0_out[9435]);
     layer1_out[1940] <= ~(layer0_out[7410] & layer0_out[7411]);
     layer1_out[1941] <= ~layer0_out[6802] | layer0_out[6801];
     layer1_out[1942] <= layer0_out[2398];
     layer1_out[1943] <= ~(layer0_out[2642] & layer0_out[2643]);
     layer1_out[1944] <= ~layer0_out[1413];
     layer1_out[1945] <= ~(layer0_out[1285] ^ layer0_out[1286]);
     layer1_out[1946] <= layer0_out[4928] & ~layer0_out[4929];
     layer1_out[1947] <= ~(layer0_out[7744] & layer0_out[7745]);
     layer1_out[1948] <= ~layer0_out[5823];
     layer1_out[1949] <= ~(layer0_out[4034] | layer0_out[4035]);
     layer1_out[1950] <= layer0_out[11243] | layer0_out[11244];
     layer1_out[1951] <= layer0_out[7947] & ~layer0_out[7948];
     layer1_out[1952] <= layer0_out[7063];
     layer1_out[1953] <= layer0_out[494];
     layer1_out[1954] <= layer0_out[10396];
     layer1_out[1955] <= layer0_out[6759];
     layer1_out[1956] <= ~(layer0_out[1851] & layer0_out[1852]);
     layer1_out[1957] <= ~(layer0_out[483] & layer0_out[484]);
     layer1_out[1958] <= layer0_out[5014];
     layer1_out[1959] <= layer0_out[2690] & ~layer0_out[2689];
     layer1_out[1960] <= ~layer0_out[11502];
     layer1_out[1961] <= layer0_out[8103] & layer0_out[8104];
     layer1_out[1962] <= ~layer0_out[3600];
     layer1_out[1963] <= layer0_out[6379] | layer0_out[6380];
     layer1_out[1964] <= ~layer0_out[8732];
     layer1_out[1965] <= ~(layer0_out[9077] & layer0_out[9078]);
     layer1_out[1966] <= layer0_out[2473];
     layer1_out[1967] <= layer0_out[1959] & ~layer0_out[1958];
     layer1_out[1968] <= layer0_out[2838] & ~layer0_out[2839];
     layer1_out[1969] <= ~(layer0_out[3471] ^ layer0_out[3472]);
     layer1_out[1970] <= ~layer0_out[2312];
     layer1_out[1971] <= ~layer0_out[1517] | layer0_out[1518];
     layer1_out[1972] <= layer0_out[4174] & layer0_out[4175];
     layer1_out[1973] <= layer0_out[8027];
     layer1_out[1974] <= ~(layer0_out[786] | layer0_out[787]);
     layer1_out[1975] <= 1'b1;
     layer1_out[1976] <= ~layer0_out[4798] | layer0_out[4797];
     layer1_out[1977] <= ~layer0_out[5734] | layer0_out[5733];
     layer1_out[1978] <= 1'b0;
     layer1_out[1979] <= ~layer0_out[9990] | layer0_out[9989];
     layer1_out[1980] <= ~(layer0_out[7308] & layer0_out[7309]);
     layer1_out[1981] <= layer0_out[11612] | layer0_out[11613];
     layer1_out[1982] <= 1'b0;
     layer1_out[1983] <= layer0_out[5674] & ~layer0_out[5673];
     layer1_out[1984] <= layer0_out[222];
     layer1_out[1985] <= layer0_out[1994] & ~layer0_out[1993];
     layer1_out[1986] <= layer0_out[3907];
     layer1_out[1987] <= layer0_out[1250] & ~layer0_out[1249];
     layer1_out[1988] <= layer0_out[5325];
     layer1_out[1989] <= layer0_out[73] & ~layer0_out[74];
     layer1_out[1990] <= layer0_out[7412] & layer0_out[7413];
     layer1_out[1991] <= ~(layer0_out[9942] | layer0_out[9943]);
     layer1_out[1992] <= ~layer0_out[6479];
     layer1_out[1993] <= layer0_out[6106] & ~layer0_out[6107];
     layer1_out[1994] <= ~layer0_out[10201] | layer0_out[10202];
     layer1_out[1995] <= ~layer0_out[11059];
     layer1_out[1996] <= ~(layer0_out[8165] & layer0_out[8166]);
     layer1_out[1997] <= ~layer0_out[10668] | layer0_out[10669];
     layer1_out[1998] <= layer0_out[2207] & ~layer0_out[2206];
     layer1_out[1999] <= 1'b0;
     layer1_out[2000] <= 1'b0;
     layer1_out[2001] <= ~(layer0_out[10835] & layer0_out[10836]);
     layer1_out[2002] <= ~(layer0_out[729] ^ layer0_out[730]);
     layer1_out[2003] <= ~layer0_out[10945];
     layer1_out[2004] <= layer0_out[9460] & layer0_out[9461];
     layer1_out[2005] <= layer0_out[3934] & layer0_out[3935];
     layer1_out[2006] <= layer0_out[9168] | layer0_out[9169];
     layer1_out[2007] <= layer0_out[4476] & ~layer0_out[4475];
     layer1_out[2008] <= ~(layer0_out[8446] & layer0_out[8447]);
     layer1_out[2009] <= ~(layer0_out[365] & layer0_out[366]);
     layer1_out[2010] <= ~layer0_out[1798];
     layer1_out[2011] <= ~layer0_out[2719];
     layer1_out[2012] <= layer0_out[11118];
     layer1_out[2013] <= ~layer0_out[4188];
     layer1_out[2014] <= ~(layer0_out[9475] ^ layer0_out[9476]);
     layer1_out[2015] <= layer0_out[9215] ^ layer0_out[9216];
     layer1_out[2016] <= ~(layer0_out[5550] | layer0_out[5551]);
     layer1_out[2017] <= layer0_out[9216] | layer0_out[9217];
     layer1_out[2018] <= layer0_out[6832] & layer0_out[6833];
     layer1_out[2019] <= ~layer0_out[1545] | layer0_out[1544];
     layer1_out[2020] <= layer0_out[6990];
     layer1_out[2021] <= ~layer0_out[6405] | layer0_out[6406];
     layer1_out[2022] <= layer0_out[9923] & layer0_out[9924];
     layer1_out[2023] <= layer0_out[6768] & ~layer0_out[6767];
     layer1_out[2024] <= layer0_out[10824];
     layer1_out[2025] <= layer0_out[9142];
     layer1_out[2026] <= 1'b0;
     layer1_out[2027] <= ~layer0_out[2039];
     layer1_out[2028] <= layer0_out[11239];
     layer1_out[2029] <= layer0_out[9655] & ~layer0_out[9656];
     layer1_out[2030] <= ~layer0_out[2352];
     layer1_out[2031] <= layer0_out[6501] & ~layer0_out[6500];
     layer1_out[2032] <= layer0_out[3258];
     layer1_out[2033] <= ~(layer0_out[9506] | layer0_out[9507]);
     layer1_out[2034] <= ~layer0_out[3898] | layer0_out[3899];
     layer1_out[2035] <= layer0_out[371] & ~layer0_out[370];
     layer1_out[2036] <= layer0_out[8111] & ~layer0_out[8110];
     layer1_out[2037] <= ~(layer0_out[2880] | layer0_out[2881]);
     layer1_out[2038] <= 1'b1;
     layer1_out[2039] <= layer0_out[6904] & layer0_out[6905];
     layer1_out[2040] <= layer0_out[10531];
     layer1_out[2041] <= layer0_out[1996] & layer0_out[1997];
     layer1_out[2042] <= ~layer0_out[7243];
     layer1_out[2043] <= 1'b0;
     layer1_out[2044] <= layer0_out[10223] | layer0_out[10224];
     layer1_out[2045] <= layer0_out[3996];
     layer1_out[2046] <= layer0_out[7612] & ~layer0_out[7613];
     layer1_out[2047] <= ~layer0_out[5570];
     layer1_out[2048] <= layer0_out[1609] ^ layer0_out[1610];
     layer1_out[2049] <= layer0_out[605] & ~layer0_out[604];
     layer1_out[2050] <= ~layer0_out[725];
     layer1_out[2051] <= ~(layer0_out[9712] & layer0_out[9713]);
     layer1_out[2052] <= layer0_out[2119] & layer0_out[2120];
     layer1_out[2053] <= ~(layer0_out[6484] & layer0_out[6485]);
     layer1_out[2054] <= layer0_out[11401] | layer0_out[11402];
     layer1_out[2055] <= ~(layer0_out[2214] | layer0_out[2215]);
     layer1_out[2056] <= 1'b1;
     layer1_out[2057] <= layer0_out[4833];
     layer1_out[2058] <= layer0_out[811] & layer0_out[812];
     layer1_out[2059] <= layer0_out[2872] & layer0_out[2873];
     layer1_out[2060] <= ~(layer0_out[6649] | layer0_out[6650]);
     layer1_out[2061] <= layer0_out[2633];
     layer1_out[2062] <= layer0_out[8138];
     layer1_out[2063] <= ~layer0_out[3863];
     layer1_out[2064] <= layer0_out[11733] ^ layer0_out[11734];
     layer1_out[2065] <= layer0_out[11447] & layer0_out[11448];
     layer1_out[2066] <= layer0_out[10867] ^ layer0_out[10868];
     layer1_out[2067] <= 1'b0;
     layer1_out[2068] <= ~layer0_out[11380];
     layer1_out[2069] <= ~layer0_out[4346] | layer0_out[4345];
     layer1_out[2070] <= layer0_out[5708] & ~layer0_out[5707];
     layer1_out[2071] <= ~layer0_out[10701];
     layer1_out[2072] <= ~(layer0_out[5931] ^ layer0_out[5932]);
     layer1_out[2073] <= ~layer0_out[1051];
     layer1_out[2074] <= layer0_out[9062];
     layer1_out[2075] <= layer0_out[3320] & layer0_out[3321];
     layer1_out[2076] <= ~layer0_out[5461];
     layer1_out[2077] <= ~layer0_out[11368];
     layer1_out[2078] <= ~layer0_out[3772];
     layer1_out[2079] <= ~layer0_out[696];
     layer1_out[2080] <= ~(layer0_out[4152] | layer0_out[4153]);
     layer1_out[2081] <= ~(layer0_out[4749] ^ layer0_out[4750]);
     layer1_out[2082] <= ~(layer0_out[3490] & layer0_out[3491]);
     layer1_out[2083] <= ~(layer0_out[8896] | layer0_out[8897]);
     layer1_out[2084] <= layer0_out[4586] & layer0_out[4587];
     layer1_out[2085] <= 1'b0;
     layer1_out[2086] <= layer0_out[191];
     layer1_out[2087] <= layer0_out[8104] & layer0_out[8105];
     layer1_out[2088] <= ~layer0_out[9773];
     layer1_out[2089] <= layer0_out[4854] & ~layer0_out[4853];
     layer1_out[2090] <= ~layer0_out[532];
     layer1_out[2091] <= ~(layer0_out[8204] | layer0_out[8205]);
     layer1_out[2092] <= ~layer0_out[8828];
     layer1_out[2093] <= layer0_out[179];
     layer1_out[2094] <= layer0_out[10834];
     layer1_out[2095] <= layer0_out[3472] | layer0_out[3473];
     layer1_out[2096] <= ~(layer0_out[1987] ^ layer0_out[1988]);
     layer1_out[2097] <= ~(layer0_out[3805] & layer0_out[3806]);
     layer1_out[2098] <= ~(layer0_out[4570] ^ layer0_out[4571]);
     layer1_out[2099] <= ~layer0_out[5289];
     layer1_out[2100] <= layer0_out[5467];
     layer1_out[2101] <= layer0_out[9270];
     layer1_out[2102] <= ~layer0_out[4171];
     layer1_out[2103] <= ~(layer0_out[1623] & layer0_out[1624]);
     layer1_out[2104] <= layer0_out[1947] & ~layer0_out[1948];
     layer1_out[2105] <= ~layer0_out[1208] | layer0_out[1209];
     layer1_out[2106] <= layer0_out[1118] & ~layer0_out[1117];
     layer1_out[2107] <= ~layer0_out[6931];
     layer1_out[2108] <= ~layer0_out[644];
     layer1_out[2109] <= ~(layer0_out[4159] | layer0_out[4160]);
     layer1_out[2110] <= layer0_out[5396];
     layer1_out[2111] <= ~layer0_out[8687] | layer0_out[8686];
     layer1_out[2112] <= ~(layer0_out[10669] | layer0_out[10670]);
     layer1_out[2113] <= layer0_out[1853];
     layer1_out[2114] <= ~(layer0_out[157] | layer0_out[158]);
     layer1_out[2115] <= layer0_out[5529] & ~layer0_out[5528];
     layer1_out[2116] <= layer0_out[3960] & layer0_out[3961];
     layer1_out[2117] <= layer0_out[10948] & layer0_out[10949];
     layer1_out[2118] <= layer0_out[1522] | layer0_out[1523];
     layer1_out[2119] <= layer0_out[9083];
     layer1_out[2120] <= ~layer0_out[10108] | layer0_out[10109];
     layer1_out[2121] <= ~(layer0_out[1739] & layer0_out[1740]);
     layer1_out[2122] <= layer0_out[1593] & ~layer0_out[1592];
     layer1_out[2123] <= ~layer0_out[11599] | layer0_out[11600];
     layer1_out[2124] <= layer0_out[1108] & layer0_out[1109];
     layer1_out[2125] <= ~layer0_out[10756] | layer0_out[10755];
     layer1_out[2126] <= ~layer0_out[1804];
     layer1_out[2127] <= 1'b1;
     layer1_out[2128] <= ~layer0_out[3185];
     layer1_out[2129] <= ~(layer0_out[2487] ^ layer0_out[2488]);
     layer1_out[2130] <= layer0_out[9018];
     layer1_out[2131] <= layer0_out[8014] & layer0_out[8015];
     layer1_out[2132] <= ~(layer0_out[4703] ^ layer0_out[4704]);
     layer1_out[2133] <= ~layer0_out[8510] | layer0_out[8511];
     layer1_out[2134] <= layer0_out[4269] & layer0_out[4270];
     layer1_out[2135] <= layer0_out[8426];
     layer1_out[2136] <= layer0_out[9954] ^ layer0_out[9955];
     layer1_out[2137] <= layer0_out[5237];
     layer1_out[2138] <= ~layer0_out[11482];
     layer1_out[2139] <= ~layer0_out[5836] | layer0_out[5835];
     layer1_out[2140] <= 1'b1;
     layer1_out[2141] <= layer0_out[3988];
     layer1_out[2142] <= ~layer0_out[8787];
     layer1_out[2143] <= ~layer0_out[8846];
     layer1_out[2144] <= layer0_out[1385] | layer0_out[1386];
     layer1_out[2145] <= layer0_out[6946];
     layer1_out[2146] <= ~layer0_out[2675];
     layer1_out[2147] <= layer0_out[11755] | layer0_out[11756];
     layer1_out[2148] <= layer0_out[8951];
     layer1_out[2149] <= ~layer0_out[8945];
     layer1_out[2150] <= 1'b1;
     layer1_out[2151] <= ~layer0_out[1343];
     layer1_out[2152] <= layer0_out[5876] & layer0_out[5877];
     layer1_out[2153] <= 1'b0;
     layer1_out[2154] <= ~layer0_out[7187] | layer0_out[7186];
     layer1_out[2155] <= ~layer0_out[11257];
     layer1_out[2156] <= layer0_out[9386];
     layer1_out[2157] <= layer0_out[11352] & layer0_out[11353];
     layer1_out[2158] <= layer0_out[8272] & layer0_out[8273];
     layer1_out[2159] <= ~layer0_out[6980] | layer0_out[6979];
     layer1_out[2160] <= layer0_out[11420] & layer0_out[11421];
     layer1_out[2161] <= ~layer0_out[6005];
     layer1_out[2162] <= layer0_out[4926] & ~layer0_out[4927];
     layer1_out[2163] <= layer0_out[4690] & ~layer0_out[4689];
     layer1_out[2164] <= ~layer0_out[3284];
     layer1_out[2165] <= ~layer0_out[8827] | layer0_out[8826];
     layer1_out[2166] <= layer0_out[1341];
     layer1_out[2167] <= ~(layer0_out[11329] ^ layer0_out[11330]);
     layer1_out[2168] <= ~layer0_out[11723] | layer0_out[11722];
     layer1_out[2169] <= ~(layer0_out[10740] | layer0_out[10741]);
     layer1_out[2170] <= layer0_out[2626] & layer0_out[2627];
     layer1_out[2171] <= layer0_out[5916] & layer0_out[5917];
     layer1_out[2172] <= ~(layer0_out[2013] ^ layer0_out[2014]);
     layer1_out[2173] <= 1'b0;
     layer1_out[2174] <= ~layer0_out[11828];
     layer1_out[2175] <= ~(layer0_out[9389] ^ layer0_out[9390]);
     layer1_out[2176] <= ~(layer0_out[5503] | layer0_out[5504]);
     layer1_out[2177] <= layer0_out[5820] & ~layer0_out[5819];
     layer1_out[2178] <= ~layer0_out[6083] | layer0_out[6084];
     layer1_out[2179] <= ~(layer0_out[3590] | layer0_out[3591]);
     layer1_out[2180] <= ~layer0_out[4382];
     layer1_out[2181] <= ~layer0_out[2302] | layer0_out[2301];
     layer1_out[2182] <= ~(layer0_out[9111] & layer0_out[9112]);
     layer1_out[2183] <= layer0_out[6970] & ~layer0_out[6969];
     layer1_out[2184] <= ~layer0_out[11632];
     layer1_out[2185] <= ~(layer0_out[11475] | layer0_out[11476]);
     layer1_out[2186] <= layer0_out[11587] & ~layer0_out[11588];
     layer1_out[2187] <= 1'b0;
     layer1_out[2188] <= layer0_out[873];
     layer1_out[2189] <= ~(layer0_out[909] ^ layer0_out[910]);
     layer1_out[2190] <= ~layer0_out[10228];
     layer1_out[2191] <= ~(layer0_out[5220] & layer0_out[5221]);
     layer1_out[2192] <= layer0_out[2045] & ~layer0_out[2044];
     layer1_out[2193] <= ~(layer0_out[4239] | layer0_out[4240]);
     layer1_out[2194] <= ~layer0_out[6853] | layer0_out[6854];
     layer1_out[2195] <= layer0_out[4210] & layer0_out[4211];
     layer1_out[2196] <= layer0_out[4411] & layer0_out[4412];
     layer1_out[2197] <= ~(layer0_out[5571] | layer0_out[5572]);
     layer1_out[2198] <= layer0_out[2408] & ~layer0_out[2407];
     layer1_out[2199] <= layer0_out[2756] | layer0_out[2757];
     layer1_out[2200] <= ~layer0_out[4877];
     layer1_out[2201] <= ~(layer0_out[8653] & layer0_out[8654]);
     layer1_out[2202] <= 1'b0;
     layer1_out[2203] <= ~(layer0_out[7108] | layer0_out[7109]);
     layer1_out[2204] <= ~(layer0_out[9682] | layer0_out[9683]);
     layer1_out[2205] <= ~(layer0_out[10157] & layer0_out[10158]);
     layer1_out[2206] <= layer0_out[8098] & ~layer0_out[8099];
     layer1_out[2207] <= ~layer0_out[2923];
     layer1_out[2208] <= layer0_out[6575] & ~layer0_out[6576];
     layer1_out[2209] <= layer0_out[5380] | layer0_out[5381];
     layer1_out[2210] <= layer0_out[8101] & layer0_out[8102];
     layer1_out[2211] <= layer0_out[9269];
     layer1_out[2212] <= layer0_out[3378] ^ layer0_out[3379];
     layer1_out[2213] <= layer0_out[7396];
     layer1_out[2214] <= layer0_out[5746] | layer0_out[5747];
     layer1_out[2215] <= 1'b0;
     layer1_out[2216] <= ~layer0_out[10809] | layer0_out[10810];
     layer1_out[2217] <= 1'b1;
     layer1_out[2218] <= ~layer0_out[4048];
     layer1_out[2219] <= ~(layer0_out[3339] & layer0_out[3340]);
     layer1_out[2220] <= layer0_out[11926];
     layer1_out[2221] <= ~layer0_out[9345] | layer0_out[9346];
     layer1_out[2222] <= layer0_out[9421];
     layer1_out[2223] <= ~layer0_out[4099];
     layer1_out[2224] <= ~layer0_out[9938];
     layer1_out[2225] <= layer0_out[8958] | layer0_out[8959];
     layer1_out[2226] <= ~layer0_out[1432];
     layer1_out[2227] <= layer0_out[3607] ^ layer0_out[3608];
     layer1_out[2228] <= ~(layer0_out[1732] | layer0_out[1733]);
     layer1_out[2229] <= ~(layer0_out[960] ^ layer0_out[961]);
     layer1_out[2230] <= layer0_out[8734] & ~layer0_out[8733];
     layer1_out[2231] <= ~layer0_out[6682] | layer0_out[6681];
     layer1_out[2232] <= layer0_out[2258];
     layer1_out[2233] <= ~layer0_out[2429];
     layer1_out[2234] <= ~layer0_out[8370];
     layer1_out[2235] <= layer0_out[929] | layer0_out[930];
     layer1_out[2236] <= layer0_out[7144] ^ layer0_out[7145];
     layer1_out[2237] <= ~layer0_out[7258];
     layer1_out[2238] <= ~layer0_out[290];
     layer1_out[2239] <= ~layer0_out[4727];
     layer1_out[2240] <= layer0_out[653];
     layer1_out[2241] <= layer0_out[7283];
     layer1_out[2242] <= ~(layer0_out[9987] & layer0_out[9988]);
     layer1_out[2243] <= layer0_out[985];
     layer1_out[2244] <= layer0_out[6630];
     layer1_out[2245] <= ~(layer0_out[6270] | layer0_out[6271]);
     layer1_out[2246] <= ~(layer0_out[9117] | layer0_out[9118]);
     layer1_out[2247] <= layer0_out[8194] & ~layer0_out[8195];
     layer1_out[2248] <= ~(layer0_out[9377] & layer0_out[9378]);
     layer1_out[2249] <= ~layer0_out[4278] | layer0_out[4277];
     layer1_out[2250] <= layer0_out[6756];
     layer1_out[2251] <= ~layer0_out[1105];
     layer1_out[2252] <= ~layer0_out[1780];
     layer1_out[2253] <= layer0_out[10504] | layer0_out[10505];
     layer1_out[2254] <= layer0_out[7314] ^ layer0_out[7315];
     layer1_out[2255] <= layer0_out[10969] & layer0_out[10970];
     layer1_out[2256] <= layer0_out[4810] & ~layer0_out[4811];
     layer1_out[2257] <= layer0_out[4354] & layer0_out[4355];
     layer1_out[2258] <= ~(layer0_out[11657] & layer0_out[11658]);
     layer1_out[2259] <= ~(layer0_out[9573] & layer0_out[9574]);
     layer1_out[2260] <= layer0_out[9217];
     layer1_out[2261] <= ~layer0_out[7700];
     layer1_out[2262] <= layer0_out[4840] & ~layer0_out[4841];
     layer1_out[2263] <= layer0_out[7161];
     layer1_out[2264] <= layer0_out[7621] | layer0_out[7622];
     layer1_out[2265] <= layer0_out[1474];
     layer1_out[2266] <= ~layer0_out[9218];
     layer1_out[2267] <= layer0_out[10318];
     layer1_out[2268] <= layer0_out[11278];
     layer1_out[2269] <= layer0_out[5026] | layer0_out[5027];
     layer1_out[2270] <= layer0_out[9472] & layer0_out[9473];
     layer1_out[2271] <= ~layer0_out[11025] | layer0_out[11024];
     layer1_out[2272] <= layer0_out[7479];
     layer1_out[2273] <= layer0_out[5316] | layer0_out[5317];
     layer1_out[2274] <= ~layer0_out[3767] | layer0_out[3768];
     layer1_out[2275] <= 1'b1;
     layer1_out[2276] <= ~(layer0_out[7529] ^ layer0_out[7530]);
     layer1_out[2277] <= layer0_out[5057];
     layer1_out[2278] <= layer0_out[6948] & ~layer0_out[6947];
     layer1_out[2279] <= layer0_out[5530];
     layer1_out[2280] <= layer0_out[10376];
     layer1_out[2281] <= layer0_out[7015];
     layer1_out[2282] <= layer0_out[3317] & layer0_out[3318];
     layer1_out[2283] <= layer0_out[9562];
     layer1_out[2284] <= ~layer0_out[744];
     layer1_out[2285] <= layer0_out[8288] | layer0_out[8289];
     layer1_out[2286] <= layer0_out[896];
     layer1_out[2287] <= ~layer0_out[8511];
     layer1_out[2288] <= layer0_out[9819] & ~layer0_out[9818];
     layer1_out[2289] <= ~layer0_out[7383];
     layer1_out[2290] <= layer0_out[4966];
     layer1_out[2291] <= ~layer0_out[3273] | layer0_out[3272];
     layer1_out[2292] <= ~layer0_out[9558] | layer0_out[9557];
     layer1_out[2293] <= ~layer0_out[1827];
     layer1_out[2294] <= ~layer0_out[11824];
     layer1_out[2295] <= layer0_out[412];
     layer1_out[2296] <= ~layer0_out[2208];
     layer1_out[2297] <= ~(layer0_out[6550] | layer0_out[6551]);
     layer1_out[2298] <= ~layer0_out[3032];
     layer1_out[2299] <= ~layer0_out[5172] | layer0_out[5171];
     layer1_out[2300] <= layer0_out[2422] & layer0_out[2423];
     layer1_out[2301] <= ~(layer0_out[8324] | layer0_out[8325]);
     layer1_out[2302] <= layer0_out[5909] ^ layer0_out[5910];
     layer1_out[2303] <= ~(layer0_out[4598] ^ layer0_out[4599]);
     layer1_out[2304] <= layer0_out[10164] & ~layer0_out[10163];
     layer1_out[2305] <= layer0_out[3166];
     layer1_out[2306] <= layer0_out[4895] & layer0_out[4896];
     layer1_out[2307] <= layer0_out[2220];
     layer1_out[2308] <= ~layer0_out[10719] | layer0_out[10718];
     layer1_out[2309] <= 1'b0;
     layer1_out[2310] <= ~layer0_out[233];
     layer1_out[2311] <= layer0_out[2673];
     layer1_out[2312] <= 1'b1;
     layer1_out[2313] <= ~layer0_out[5880];
     layer1_out[2314] <= ~(layer0_out[1079] ^ layer0_out[1080]);
     layer1_out[2315] <= layer0_out[7320] | layer0_out[7321];
     layer1_out[2316] <= layer0_out[8887] & layer0_out[8888];
     layer1_out[2317] <= layer0_out[3597] | layer0_out[3598];
     layer1_out[2318] <= ~(layer0_out[7379] & layer0_out[7380]);
     layer1_out[2319] <= ~layer0_out[10039];
     layer1_out[2320] <= 1'b1;
     layer1_out[2321] <= ~layer0_out[6109] | layer0_out[6110];
     layer1_out[2322] <= ~layer0_out[8573] | layer0_out[8574];
     layer1_out[2323] <= layer0_out[1481] & ~layer0_out[1480];
     layer1_out[2324] <= ~layer0_out[3443] | layer0_out[3444];
     layer1_out[2325] <= ~(layer0_out[2955] & layer0_out[2956]);
     layer1_out[2326] <= layer0_out[9237];
     layer1_out[2327] <= ~layer0_out[7347];
     layer1_out[2328] <= ~layer0_out[7588] | layer0_out[7587];
     layer1_out[2329] <= ~(layer0_out[2253] ^ layer0_out[2254]);
     layer1_out[2330] <= ~layer0_out[1049];
     layer1_out[2331] <= layer0_out[1819] & ~layer0_out[1818];
     layer1_out[2332] <= ~layer0_out[4344];
     layer1_out[2333] <= layer0_out[6747] & ~layer0_out[6748];
     layer1_out[2334] <= layer0_out[3731] | layer0_out[3732];
     layer1_out[2335] <= ~layer0_out[1530];
     layer1_out[2336] <= ~layer0_out[9362];
     layer1_out[2337] <= layer0_out[9069];
     layer1_out[2338] <= layer0_out[10397] & layer0_out[10398];
     layer1_out[2339] <= layer0_out[416] & ~layer0_out[415];
     layer1_out[2340] <= layer0_out[3263] & ~layer0_out[3264];
     layer1_out[2341] <= layer0_out[4941] & layer0_out[4942];
     layer1_out[2342] <= layer0_out[10634] & layer0_out[10635];
     layer1_out[2343] <= 1'b1;
     layer1_out[2344] <= ~layer0_out[11652];
     layer1_out[2345] <= 1'b0;
     layer1_out[2346] <= ~layer0_out[5950];
     layer1_out[2347] <= layer0_out[9599];
     layer1_out[2348] <= ~layer0_out[9579];
     layer1_out[2349] <= ~(layer0_out[1055] | layer0_out[1056]);
     layer1_out[2350] <= ~(layer0_out[4626] ^ layer0_out[4627]);
     layer1_out[2351] <= layer0_out[2376] & ~layer0_out[2375];
     layer1_out[2352] <= ~(layer0_out[1318] ^ layer0_out[1319]);
     layer1_out[2353] <= layer0_out[1906];
     layer1_out[2354] <= ~(layer0_out[4247] & layer0_out[4248]);
     layer1_out[2355] <= 1'b0;
     layer1_out[2356] <= ~(layer0_out[10447] | layer0_out[10448]);
     layer1_out[2357] <= ~layer0_out[8451];
     layer1_out[2358] <= ~layer0_out[10202];
     layer1_out[2359] <= ~layer0_out[9855] | layer0_out[9854];
     layer1_out[2360] <= layer0_out[7749] & ~layer0_out[7750];
     layer1_out[2361] <= ~layer0_out[10470] | layer0_out[10471];
     layer1_out[2362] <= ~layer0_out[9020];
     layer1_out[2363] <= 1'b0;
     layer1_out[2364] <= ~layer0_out[675];
     layer1_out[2365] <= layer0_out[7049];
     layer1_out[2366] <= ~(layer0_out[5344] ^ layer0_out[5345]);
     layer1_out[2367] <= ~layer0_out[1802] | layer0_out[1801];
     layer1_out[2368] <= layer0_out[5300] & ~layer0_out[5299];
     layer1_out[2369] <= layer0_out[11775] & ~layer0_out[11774];
     layer1_out[2370] <= ~(layer0_out[3635] | layer0_out[3636]);
     layer1_out[2371] <= layer0_out[4678] & ~layer0_out[4677];
     layer1_out[2372] <= ~layer0_out[6534];
     layer1_out[2373] <= ~layer0_out[5831];
     layer1_out[2374] <= layer0_out[5728] | layer0_out[5729];
     layer1_out[2375] <= ~layer0_out[8377];
     layer1_out[2376] <= 1'b1;
     layer1_out[2377] <= ~layer0_out[3109];
     layer1_out[2378] <= layer0_out[7427] | layer0_out[7428];
     layer1_out[2379] <= ~(layer0_out[7282] | layer0_out[7283]);
     layer1_out[2380] <= ~layer0_out[9207];
     layer1_out[2381] <= ~layer0_out[9649];
     layer1_out[2382] <= layer0_out[5590] & ~layer0_out[5589];
     layer1_out[2383] <= ~(layer0_out[3576] ^ layer0_out[3577]);
     layer1_out[2384] <= ~layer0_out[7694] | layer0_out[7695];
     layer1_out[2385] <= ~layer0_out[7419] | layer0_out[7420];
     layer1_out[2386] <= ~layer0_out[2130];
     layer1_out[2387] <= layer0_out[1595] | layer0_out[1596];
     layer1_out[2388] <= 1'b1;
     layer1_out[2389] <= ~layer0_out[5348];
     layer1_out[2390] <= layer0_out[9776] & layer0_out[9777];
     layer1_out[2391] <= ~layer0_out[3276] | layer0_out[3277];
     layer1_out[2392] <= layer0_out[3485];
     layer1_out[2393] <= layer0_out[1101] & ~layer0_out[1100];
     layer1_out[2394] <= ~layer0_out[5875];
     layer1_out[2395] <= layer0_out[9745];
     layer1_out[2396] <= 1'b0;
     layer1_out[2397] <= ~(layer0_out[592] & layer0_out[593]);
     layer1_out[2398] <= ~(layer0_out[2502] | layer0_out[2503]);
     layer1_out[2399] <= layer0_out[2913] & layer0_out[2914];
     layer1_out[2400] <= layer0_out[11689] | layer0_out[11690];
     layer1_out[2401] <= layer0_out[10319] & ~layer0_out[10318];
     layer1_out[2402] <= layer0_out[2959] ^ layer0_out[2960];
     layer1_out[2403] <= layer0_out[9135] & layer0_out[9136];
     layer1_out[2404] <= ~(layer0_out[8333] | layer0_out[8334]);
     layer1_out[2405] <= layer0_out[2123] & layer0_out[2124];
     layer1_out[2406] <= layer0_out[794];
     layer1_out[2407] <= layer0_out[11393] ^ layer0_out[11394];
     layer1_out[2408] <= layer0_out[23] | layer0_out[24];
     layer1_out[2409] <= 1'b1;
     layer1_out[2410] <= 1'b1;
     layer1_out[2411] <= layer0_out[7500] & layer0_out[7501];
     layer1_out[2412] <= ~layer0_out[3824];
     layer1_out[2413] <= layer0_out[2449] & ~layer0_out[2448];
     layer1_out[2414] <= layer0_out[9663] & layer0_out[9664];
     layer1_out[2415] <= ~layer0_out[3205];
     layer1_out[2416] <= layer0_out[7622];
     layer1_out[2417] <= layer0_out[9948] & ~layer0_out[9947];
     layer1_out[2418] <= ~(layer0_out[3757] & layer0_out[3758]);
     layer1_out[2419] <= ~layer0_out[4077];
     layer1_out[2420] <= layer0_out[11085] & layer0_out[11086];
     layer1_out[2421] <= layer0_out[6416] & ~layer0_out[6417];
     layer1_out[2422] <= ~(layer0_out[2665] ^ layer0_out[2666]);
     layer1_out[2423] <= ~(layer0_out[8467] | layer0_out[8468]);
     layer1_out[2424] <= layer0_out[1281] & ~layer0_out[1282];
     layer1_out[2425] <= ~layer0_out[8571] | layer0_out[8572];
     layer1_out[2426] <= ~(layer0_out[1778] | layer0_out[1779]);
     layer1_out[2427] <= layer0_out[7428] | layer0_out[7429];
     layer1_out[2428] <= ~layer0_out[11361] | layer0_out[11360];
     layer1_out[2429] <= ~layer0_out[6571] | layer0_out[6570];
     layer1_out[2430] <= ~layer0_out[1366];
     layer1_out[2431] <= ~layer0_out[7424];
     layer1_out[2432] <= ~layer0_out[11545];
     layer1_out[2433] <= ~layer0_out[3199];
     layer1_out[2434] <= ~(layer0_out[9102] ^ layer0_out[9103]);
     layer1_out[2435] <= layer0_out[9514] ^ layer0_out[9515];
     layer1_out[2436] <= layer0_out[302] & ~layer0_out[301];
     layer1_out[2437] <= layer0_out[3883];
     layer1_out[2438] <= layer0_out[5580];
     layer1_out[2439] <= ~(layer0_out[4472] | layer0_out[4473]);
     layer1_out[2440] <= layer0_out[6306] & ~layer0_out[6305];
     layer1_out[2441] <= layer0_out[1962] ^ layer0_out[1963];
     layer1_out[2442] <= layer0_out[3577] & ~layer0_out[3578];
     layer1_out[2443] <= ~layer0_out[9152] | layer0_out[9151];
     layer1_out[2444] <= ~layer0_out[9238];
     layer1_out[2445] <= ~layer0_out[8140] | layer0_out[8139];
     layer1_out[2446] <= layer0_out[2787];
     layer1_out[2447] <= layer0_out[1952] & layer0_out[1953];
     layer1_out[2448] <= layer0_out[1410];
     layer1_out[2449] <= layer0_out[7941] & layer0_out[7942];
     layer1_out[2450] <= ~layer0_out[4829] | layer0_out[4828];
     layer1_out[2451] <= ~layer0_out[8839] | layer0_out[8838];
     layer1_out[2452] <= layer0_out[6721];
     layer1_out[2453] <= ~layer0_out[934];
     layer1_out[2454] <= layer0_out[8580];
     layer1_out[2455] <= layer0_out[11286] & ~layer0_out[11285];
     layer1_out[2456] <= ~layer0_out[1915];
     layer1_out[2457] <= layer0_out[830] & ~layer0_out[831];
     layer1_out[2458] <= layer0_out[11217];
     layer1_out[2459] <= 1'b0;
     layer1_out[2460] <= layer0_out[11869] & ~layer0_out[11870];
     layer1_out[2461] <= layer0_out[11699];
     layer1_out[2462] <= 1'b1;
     layer1_out[2463] <= layer0_out[4211] & layer0_out[4212];
     layer1_out[2464] <= layer0_out[11806] & ~layer0_out[11807];
     layer1_out[2465] <= ~layer0_out[11608];
     layer1_out[2466] <= layer0_out[9128];
     layer1_out[2467] <= 1'b1;
     layer1_out[2468] <= ~layer0_out[10427];
     layer1_out[2469] <= ~layer0_out[4856] | layer0_out[4857];
     layer1_out[2470] <= ~layer0_out[8801];
     layer1_out[2471] <= ~layer0_out[10439];
     layer1_out[2472] <= layer0_out[9069] & ~layer0_out[9068];
     layer1_out[2473] <= 1'b1;
     layer1_out[2474] <= layer0_out[5728];
     layer1_out[2475] <= ~(layer0_out[3546] ^ layer0_out[3547]);
     layer1_out[2476] <= layer0_out[9790];
     layer1_out[2477] <= layer0_out[5094] | layer0_out[5095];
     layer1_out[2478] <= layer0_out[8248] | layer0_out[8249];
     layer1_out[2479] <= layer0_out[7668];
     layer1_out[2480] <= layer0_out[8490] & ~layer0_out[8489];
     layer1_out[2481] <= layer0_out[4060] | layer0_out[4061];
     layer1_out[2482] <= 1'b1;
     layer1_out[2483] <= layer0_out[11771];
     layer1_out[2484] <= layer0_out[8844];
     layer1_out[2485] <= ~(layer0_out[10011] & layer0_out[10012]);
     layer1_out[2486] <= ~layer0_out[11318] | layer0_out[11317];
     layer1_out[2487] <= ~(layer0_out[171] ^ layer0_out[172]);
     layer1_out[2488] <= ~layer0_out[4218];
     layer1_out[2489] <= layer0_out[8544];
     layer1_out[2490] <= ~layer0_out[7095];
     layer1_out[2491] <= ~layer0_out[3219];
     layer1_out[2492] <= layer0_out[1161];
     layer1_out[2493] <= ~(layer0_out[1976] | layer0_out[1977]);
     layer1_out[2494] <= layer0_out[2028];
     layer1_out[2495] <= layer0_out[7931] & ~layer0_out[7932];
     layer1_out[2496] <= ~(layer0_out[1271] & layer0_out[1272]);
     layer1_out[2497] <= ~layer0_out[5514] | layer0_out[5513];
     layer1_out[2498] <= layer0_out[197] & ~layer0_out[196];
     layer1_out[2499] <= ~(layer0_out[10908] & layer0_out[10909]);
     layer1_out[2500] <= ~(layer0_out[4736] ^ layer0_out[4737]);
     layer1_out[2501] <= ~(layer0_out[5315] ^ layer0_out[5316]);
     layer1_out[2502] <= layer0_out[770] | layer0_out[771];
     layer1_out[2503] <= ~layer0_out[6216];
     layer1_out[2504] <= layer0_out[3590];
     layer1_out[2505] <= layer0_out[5144] & layer0_out[5145];
     layer1_out[2506] <= ~layer0_out[3213];
     layer1_out[2507] <= layer0_out[7038];
     layer1_out[2508] <= layer0_out[7271];
     layer1_out[2509] <= layer0_out[6886] & layer0_out[6887];
     layer1_out[2510] <= layer0_out[10708];
     layer1_out[2511] <= layer0_out[2136];
     layer1_out[2512] <= layer0_out[11472];
     layer1_out[2513] <= 1'b1;
     layer1_out[2514] <= ~layer0_out[2792];
     layer1_out[2515] <= ~layer0_out[5165];
     layer1_out[2516] <= ~layer0_out[10135] | layer0_out[10134];
     layer1_out[2517] <= ~layer0_out[9519];
     layer1_out[2518] <= layer0_out[2734];
     layer1_out[2519] <= ~(layer0_out[7521] | layer0_out[7522]);
     layer1_out[2520] <= layer0_out[6662] | layer0_out[6663];
     layer1_out[2521] <= layer0_out[2356] & layer0_out[2357];
     layer1_out[2522] <= ~(layer0_out[1260] & layer0_out[1261]);
     layer1_out[2523] <= layer0_out[2589] & layer0_out[2590];
     layer1_out[2524] <= layer0_out[6757] & ~layer0_out[6758];
     layer1_out[2525] <= ~layer0_out[4066];
     layer1_out[2526] <= ~layer0_out[8738] | layer0_out[8739];
     layer1_out[2527] <= layer0_out[3391];
     layer1_out[2528] <= layer0_out[704] ^ layer0_out[705];
     layer1_out[2529] <= ~layer0_out[8168];
     layer1_out[2530] <= ~layer0_out[11646] | layer0_out[11645];
     layer1_out[2531] <= ~(layer0_out[1187] & layer0_out[1188]);
     layer1_out[2532] <= ~layer0_out[10327] | layer0_out[10326];
     layer1_out[2533] <= ~(layer0_out[4036] | layer0_out[4037]);
     layer1_out[2534] <= ~layer0_out[4928];
     layer1_out[2535] <= layer0_out[1255] | layer0_out[1256];
     layer1_out[2536] <= ~(layer0_out[9754] | layer0_out[9755]);
     layer1_out[2537] <= layer0_out[10704] ^ layer0_out[10705];
     layer1_out[2538] <= 1'b0;
     layer1_out[2539] <= ~layer0_out[5696];
     layer1_out[2540] <= ~layer0_out[142] | layer0_out[141];
     layer1_out[2541] <= ~(layer0_out[6176] | layer0_out[6177]);
     layer1_out[2542] <= ~layer0_out[9731];
     layer1_out[2543] <= layer0_out[4243] | layer0_out[4244];
     layer1_out[2544] <= layer0_out[4016];
     layer1_out[2545] <= layer0_out[11264];
     layer1_out[2546] <= layer0_out[3419] ^ layer0_out[3420];
     layer1_out[2547] <= layer0_out[8438];
     layer1_out[2548] <= layer0_out[8929] & ~layer0_out[8928];
     layer1_out[2549] <= ~layer0_out[4296] | layer0_out[4295];
     layer1_out[2550] <= ~layer0_out[1590] | layer0_out[1591];
     layer1_out[2551] <= ~layer0_out[8976];
     layer1_out[2552] <= layer0_out[4951] ^ layer0_out[4952];
     layer1_out[2553] <= ~layer0_out[5988] | layer0_out[5989];
     layer1_out[2554] <= layer0_out[10309] | layer0_out[10310];
     layer1_out[2555] <= layer0_out[1829];
     layer1_out[2556] <= ~(layer0_out[3628] & layer0_out[3629]);
     layer1_out[2557] <= layer0_out[9092] | layer0_out[9093];
     layer1_out[2558] <= layer0_out[2944];
     layer1_out[2559] <= ~(layer0_out[2409] ^ layer0_out[2410]);
     layer1_out[2560] <= layer0_out[10724] & ~layer0_out[10725];
     layer1_out[2561] <= ~layer0_out[448] | layer0_out[447];
     layer1_out[2562] <= layer0_out[2549] | layer0_out[2550];
     layer1_out[2563] <= layer0_out[11107];
     layer1_out[2564] <= layer0_out[8295] & ~layer0_out[8294];
     layer1_out[2565] <= layer0_out[1831];
     layer1_out[2566] <= layer0_out[11799] & layer0_out[11800];
     layer1_out[2567] <= ~layer0_out[7327];
     layer1_out[2568] <= layer0_out[11675] | layer0_out[11676];
     layer1_out[2569] <= ~layer0_out[11457] | layer0_out[11458];
     layer1_out[2570] <= layer0_out[9214] & ~layer0_out[9215];
     layer1_out[2571] <= layer0_out[218];
     layer1_out[2572] <= layer0_out[60];
     layer1_out[2573] <= layer0_out[10015] & ~layer0_out[10014];
     layer1_out[2574] <= ~layer0_out[2532] | layer0_out[2531];
     layer1_out[2575] <= ~layer0_out[286] | layer0_out[287];
     layer1_out[2576] <= ~layer0_out[6482];
     layer1_out[2577] <= layer0_out[11802] & ~layer0_out[11803];
     layer1_out[2578] <= layer0_out[11281];
     layer1_out[2579] <= layer0_out[8817] & ~layer0_out[8816];
     layer1_out[2580] <= ~(layer0_out[2190] | layer0_out[2191]);
     layer1_out[2581] <= ~layer0_out[5698] | layer0_out[5697];
     layer1_out[2582] <= layer0_out[5630];
     layer1_out[2583] <= layer0_out[1707] | layer0_out[1708];
     layer1_out[2584] <= ~layer0_out[4093];
     layer1_out[2585] <= ~layer0_out[5645] | layer0_out[5646];
     layer1_out[2586] <= ~(layer0_out[5217] | layer0_out[5218]);
     layer1_out[2587] <= ~(layer0_out[8535] ^ layer0_out[8536]);
     layer1_out[2588] <= ~layer0_out[5475] | layer0_out[5474];
     layer1_out[2589] <= ~layer0_out[3820];
     layer1_out[2590] <= layer0_out[6115] ^ layer0_out[6116];
     layer1_out[2591] <= ~layer0_out[4540];
     layer1_out[2592] <= ~layer0_out[2961];
     layer1_out[2593] <= layer0_out[9904] & layer0_out[9905];
     layer1_out[2594] <= ~layer0_out[10639];
     layer1_out[2595] <= layer0_out[10529] | layer0_out[10530];
     layer1_out[2596] <= ~(layer0_out[736] | layer0_out[737]);
     layer1_out[2597] <= layer0_out[4389];
     layer1_out[2598] <= ~(layer0_out[11815] | layer0_out[11816]);
     layer1_out[2599] <= layer0_out[3957] & ~layer0_out[3956];
     layer1_out[2600] <= ~(layer0_out[8330] | layer0_out[8331]);
     layer1_out[2601] <= layer0_out[1172] ^ layer0_out[1173];
     layer1_out[2602] <= layer0_out[7796] & ~layer0_out[7797];
     layer1_out[2603] <= layer0_out[11075] & ~layer0_out[11076];
     layer1_out[2604] <= ~(layer0_out[342] | layer0_out[343]);
     layer1_out[2605] <= layer0_out[7148] & layer0_out[7149];
     layer1_out[2606] <= layer0_out[10101];
     layer1_out[2607] <= layer0_out[9225];
     layer1_out[2608] <= layer0_out[4560] & ~layer0_out[4559];
     layer1_out[2609] <= layer0_out[5394] & layer0_out[5395];
     layer1_out[2610] <= layer0_out[1141] & layer0_out[1142];
     layer1_out[2611] <= layer0_out[7954] & layer0_out[7955];
     layer1_out[2612] <= ~(layer0_out[2507] ^ layer0_out[2508]);
     layer1_out[2613] <= layer0_out[312];
     layer1_out[2614] <= layer0_out[6311] & ~layer0_out[6312];
     layer1_out[2615] <= layer0_out[6139] & ~layer0_out[6140];
     layer1_out[2616] <= layer0_out[3851] | layer0_out[3852];
     layer1_out[2617] <= ~layer0_out[1515] | layer0_out[1516];
     layer1_out[2618] <= layer0_out[6917] ^ layer0_out[6918];
     layer1_out[2619] <= ~layer0_out[4737];
     layer1_out[2620] <= layer0_out[1448] & ~layer0_out[1449];
     layer1_out[2621] <= ~layer0_out[4481] | layer0_out[4482];
     layer1_out[2622] <= layer0_out[9631] & layer0_out[9632];
     layer1_out[2623] <= layer0_out[2327];
     layer1_out[2624] <= ~layer0_out[1961] | layer0_out[1962];
     layer1_out[2625] <= 1'b1;
     layer1_out[2626] <= ~layer0_out[3502] | layer0_out[3503];
     layer1_out[2627] <= ~layer0_out[814];
     layer1_out[2628] <= layer0_out[9365];
     layer1_out[2629] <= ~(layer0_out[10346] & layer0_out[10347]);
     layer1_out[2630] <= ~layer0_out[1425];
     layer1_out[2631] <= layer0_out[8581] | layer0_out[8582];
     layer1_out[2632] <= ~layer0_out[1654] | layer0_out[1655];
     layer1_out[2633] <= ~layer0_out[2973];
     layer1_out[2634] <= layer0_out[5021] & ~layer0_out[5022];
     layer1_out[2635] <= ~layer0_out[2733];
     layer1_out[2636] <= layer0_out[6236] & ~layer0_out[6235];
     layer1_out[2637] <= layer0_out[8373] & ~layer0_out[8374];
     layer1_out[2638] <= ~layer0_out[2984];
     layer1_out[2639] <= layer0_out[11985];
     layer1_out[2640] <= ~(layer0_out[8304] & layer0_out[8305]);
     layer1_out[2641] <= ~layer0_out[8229] | layer0_out[8230];
     layer1_out[2642] <= ~(layer0_out[8687] & layer0_out[8688]);
     layer1_out[2643] <= ~layer0_out[4174] | layer0_out[4173];
     layer1_out[2644] <= ~layer0_out[3781] | layer0_out[3780];
     layer1_out[2645] <= layer0_out[10637] | layer0_out[10638];
     layer1_out[2646] <= layer0_out[7260] ^ layer0_out[7261];
     layer1_out[2647] <= ~layer0_out[540] | layer0_out[541];
     layer1_out[2648] <= ~layer0_out[1539] | layer0_out[1540];
     layer1_out[2649] <= layer0_out[11782] & ~layer0_out[11783];
     layer1_out[2650] <= layer0_out[5551] | layer0_out[5552];
     layer1_out[2651] <= ~layer0_out[1567] | layer0_out[1568];
     layer1_out[2652] <= layer0_out[5840] | layer0_out[5841];
     layer1_out[2653] <= ~layer0_out[3347] | layer0_out[3348];
     layer1_out[2654] <= layer0_out[4744] | layer0_out[4745];
     layer1_out[2655] <= layer0_out[8727] ^ layer0_out[8728];
     layer1_out[2656] <= ~(layer0_out[1819] & layer0_out[1820]);
     layer1_out[2657] <= ~(layer0_out[9765] & layer0_out[9766]);
     layer1_out[2658] <= ~(layer0_out[8331] & layer0_out[8332]);
     layer1_out[2659] <= ~(layer0_out[8762] | layer0_out[8763]);
     layer1_out[2660] <= ~layer0_out[10477];
     layer1_out[2661] <= ~(layer0_out[9348] | layer0_out[9349]);
     layer1_out[2662] <= ~(layer0_out[10706] & layer0_out[10707]);
     layer1_out[2663] <= layer0_out[2135] & ~layer0_out[2136];
     layer1_out[2664] <= ~layer0_out[6119] | layer0_out[6120];
     layer1_out[2665] <= ~layer0_out[6653];
     layer1_out[2666] <= ~layer0_out[9748] | layer0_out[9747];
     layer1_out[2667] <= ~(layer0_out[6074] & layer0_out[6075]);
     layer1_out[2668] <= layer0_out[6868];
     layer1_out[2669] <= ~layer0_out[634] | layer0_out[633];
     layer1_out[2670] <= layer0_out[10688] | layer0_out[10689];
     layer1_out[2671] <= layer0_out[7307];
     layer1_out[2672] <= layer0_out[5848] & ~layer0_out[5849];
     layer1_out[2673] <= layer0_out[6540] & ~layer0_out[6541];
     layer1_out[2674] <= ~layer0_out[3129];
     layer1_out[2675] <= layer0_out[7756];
     layer1_out[2676] <= layer0_out[10261] & layer0_out[10262];
     layer1_out[2677] <= layer0_out[10208] & ~layer0_out[10209];
     layer1_out[2678] <= layer0_out[10644];
     layer1_out[2679] <= layer0_out[859] | layer0_out[860];
     layer1_out[2680] <= layer0_out[11911] & ~layer0_out[11910];
     layer1_out[2681] <= ~(layer0_out[8315] & layer0_out[8316]);
     layer1_out[2682] <= layer0_out[9943] | layer0_out[9944];
     layer1_out[2683] <= layer0_out[11054] & ~layer0_out[11053];
     layer1_out[2684] <= ~(layer0_out[5378] & layer0_out[5379]);
     layer1_out[2685] <= ~(layer0_out[7822] ^ layer0_out[7823]);
     layer1_out[2686] <= ~(layer0_out[6364] ^ layer0_out[6365]);
     layer1_out[2687] <= ~layer0_out[226];
     layer1_out[2688] <= layer0_out[3703];
     layer1_out[2689] <= layer0_out[4957] & layer0_out[4958];
     layer1_out[2690] <= ~layer0_out[6665] | layer0_out[6666];
     layer1_out[2691] <= ~layer0_out[5197] | layer0_out[5196];
     layer1_out[2692] <= 1'b0;
     layer1_out[2693] <= ~layer0_out[9126] | layer0_out[9125];
     layer1_out[2694] <= layer0_out[10355] & ~layer0_out[10354];
     layer1_out[2695] <= ~layer0_out[10304];
     layer1_out[2696] <= ~layer0_out[7479];
     layer1_out[2697] <= layer0_out[5190] ^ layer0_out[5191];
     layer1_out[2698] <= ~layer0_out[6310];
     layer1_out[2699] <= layer0_out[3249] | layer0_out[3250];
     layer1_out[2700] <= ~layer0_out[10241] | layer0_out[10242];
     layer1_out[2701] <= layer0_out[9968] & layer0_out[9969];
     layer1_out[2702] <= ~layer0_out[2999];
     layer1_out[2703] <= ~(layer0_out[6151] & layer0_out[6152]);
     layer1_out[2704] <= layer0_out[5428] & layer0_out[5429];
     layer1_out[2705] <= ~(layer0_out[3270] | layer0_out[3271]);
     layer1_out[2706] <= layer0_out[6981] | layer0_out[6982];
     layer1_out[2707] <= ~layer0_out[8521] | layer0_out[8520];
     layer1_out[2708] <= ~layer0_out[10944];
     layer1_out[2709] <= ~(layer0_out[751] | layer0_out[752]);
     layer1_out[2710] <= layer0_out[3805];
     layer1_out[2711] <= 1'b0;
     layer1_out[2712] <= ~layer0_out[4322];
     layer1_out[2713] <= ~layer0_out[5489] | layer0_out[5490];
     layer1_out[2714] <= ~layer0_out[8299] | layer0_out[8300];
     layer1_out[2715] <= layer0_out[7199];
     layer1_out[2716] <= layer0_out[4029] & layer0_out[4030];
     layer1_out[2717] <= layer0_out[4168] & ~layer0_out[4169];
     layer1_out[2718] <= ~layer0_out[2596];
     layer1_out[2719] <= layer0_out[9474] & ~layer0_out[9473];
     layer1_out[2720] <= ~layer0_out[5454];
     layer1_out[2721] <= ~layer0_out[8608] | layer0_out[8607];
     layer1_out[2722] <= ~(layer0_out[3914] | layer0_out[3915]);
     layer1_out[2723] <= ~layer0_out[9446] | layer0_out[9445];
     layer1_out[2724] <= layer0_out[10265] & ~layer0_out[10266];
     layer1_out[2725] <= ~layer0_out[674];
     layer1_out[2726] <= ~layer0_out[11560] | layer0_out[11559];
     layer1_out[2727] <= ~layer0_out[5257];
     layer1_out[2728] <= layer0_out[11962] & layer0_out[11963];
     layer1_out[2729] <= layer0_out[11021];
     layer1_out[2730] <= ~layer0_out[7962] | layer0_out[7963];
     layer1_out[2731] <= ~(layer0_out[5363] & layer0_out[5364]);
     layer1_out[2732] <= ~layer0_out[8478];
     layer1_out[2733] <= layer0_out[8949];
     layer1_out[2734] <= layer0_out[6010];
     layer1_out[2735] <= layer0_out[8420] & ~layer0_out[8419];
     layer1_out[2736] <= layer0_out[9246] | layer0_out[9247];
     layer1_out[2737] <= layer0_out[5871] & layer0_out[5872];
     layer1_out[2738] <= layer0_out[1791] & ~layer0_out[1792];
     layer1_out[2739] <= ~layer0_out[9263] | layer0_out[9264];
     layer1_out[2740] <= ~layer0_out[8413] | layer0_out[8412];
     layer1_out[2741] <= ~layer0_out[3159] | layer0_out[3160];
     layer1_out[2742] <= layer0_out[9043] & layer0_out[9044];
     layer1_out[2743] <= layer0_out[3852];
     layer1_out[2744] <= ~(layer0_out[11004] | layer0_out[11005]);
     layer1_out[2745] <= ~(layer0_out[8180] & layer0_out[8181]);
     layer1_out[2746] <= ~layer0_out[4262] | layer0_out[4261];
     layer1_out[2747] <= layer0_out[7633] & ~layer0_out[7634];
     layer1_out[2748] <= ~(layer0_out[1681] ^ layer0_out[1682]);
     layer1_out[2749] <= ~layer0_out[5602];
     layer1_out[2750] <= ~(layer0_out[1594] | layer0_out[1595]);
     layer1_out[2751] <= layer0_out[1136] & ~layer0_out[1137];
     layer1_out[2752] <= layer0_out[6428] & layer0_out[6429];
     layer1_out[2753] <= layer0_out[8882] ^ layer0_out[8883];
     layer1_out[2754] <= ~layer0_out[1827] | layer0_out[1828];
     layer1_out[2755] <= ~layer0_out[1020];
     layer1_out[2756] <= layer0_out[6273] & layer0_out[6274];
     layer1_out[2757] <= ~layer0_out[9470];
     layer1_out[2758] <= layer0_out[9709];
     layer1_out[2759] <= layer0_out[6928] & ~layer0_out[6927];
     layer1_out[2760] <= layer0_out[1316];
     layer1_out[2761] <= ~layer0_out[11759] | layer0_out[11758];
     layer1_out[2762] <= ~layer0_out[7558] | layer0_out[7557];
     layer1_out[2763] <= ~layer0_out[3050];
     layer1_out[2764] <= ~(layer0_out[6419] ^ layer0_out[6420]);
     layer1_out[2765] <= ~layer0_out[1410];
     layer1_out[2766] <= ~layer0_out[6867];
     layer1_out[2767] <= ~layer0_out[1678];
     layer1_out[2768] <= ~layer0_out[4057];
     layer1_out[2769] <= ~layer0_out[5644];
     layer1_out[2770] <= ~layer0_out[2639];
     layer1_out[2771] <= layer0_out[7835] ^ layer0_out[7836];
     layer1_out[2772] <= layer0_out[4631];
     layer1_out[2773] <= ~(layer0_out[8718] & layer0_out[8719]);
     layer1_out[2774] <= layer0_out[7107] & ~layer0_out[7108];
     layer1_out[2775] <= ~layer0_out[3531];
     layer1_out[2776] <= layer0_out[2200] & layer0_out[2201];
     layer1_out[2777] <= layer0_out[9672] & layer0_out[9673];
     layer1_out[2778] <= layer0_out[10407] & ~layer0_out[10406];
     layer1_out[2779] <= ~layer0_out[11767];
     layer1_out[2780] <= layer0_out[5442] | layer0_out[5443];
     layer1_out[2781] <= layer0_out[2035] & layer0_out[2036];
     layer1_out[2782] <= layer0_out[6204] & ~layer0_out[6203];
     layer1_out[2783] <= ~layer0_out[6142];
     layer1_out[2784] <= layer0_out[2763] | layer0_out[2764];
     layer1_out[2785] <= layer0_out[10564];
     layer1_out[2786] <= layer0_out[37];
     layer1_out[2787] <= layer0_out[8610];
     layer1_out[2788] <= ~layer0_out[6198];
     layer1_out[2789] <= ~(layer0_out[11993] | layer0_out[11994]);
     layer1_out[2790] <= layer0_out[258] ^ layer0_out[259];
     layer1_out[2791] <= ~layer0_out[11208] | layer0_out[11209];
     layer1_out[2792] <= 1'b0;
     layer1_out[2793] <= layer0_out[412];
     layer1_out[2794] <= ~layer0_out[2590] | layer0_out[2591];
     layer1_out[2795] <= ~layer0_out[11287] | layer0_out[11288];
     layer1_out[2796] <= ~layer0_out[4291] | layer0_out[4290];
     layer1_out[2797] <= ~layer0_out[8308] | layer0_out[8307];
     layer1_out[2798] <= layer0_out[11817];
     layer1_out[2799] <= ~(layer0_out[6389] & layer0_out[6390]);
     layer1_out[2800] <= ~layer0_out[3528] | layer0_out[3529];
     layer1_out[2801] <= layer0_out[3352] | layer0_out[3353];
     layer1_out[2802] <= ~(layer0_out[9570] | layer0_out[9571]);
     layer1_out[2803] <= ~(layer0_out[6052] | layer0_out[6053]);
     layer1_out[2804] <= layer0_out[7192];
     layer1_out[2805] <= layer0_out[738] ^ layer0_out[739];
     layer1_out[2806] <= ~layer0_out[4906] | layer0_out[4907];
     layer1_out[2807] <= layer0_out[8774];
     layer1_out[2808] <= layer0_out[10413] & ~layer0_out[10412];
     layer1_out[2809] <= layer0_out[1373];
     layer1_out[2810] <= layer0_out[11106] & ~layer0_out[11105];
     layer1_out[2811] <= layer0_out[6024] & ~layer0_out[6023];
     layer1_out[2812] <= layer0_out[4281];
     layer1_out[2813] <= ~(layer0_out[2380] ^ layer0_out[2381]);
     layer1_out[2814] <= ~layer0_out[3019] | layer0_out[3018];
     layer1_out[2815] <= layer0_out[600] ^ layer0_out[601];
     layer1_out[2816] <= layer0_out[7921];
     layer1_out[2817] <= ~layer0_out[7025];
     layer1_out[2818] <= layer0_out[8884] ^ layer0_out[8885];
     layer1_out[2819] <= 1'b1;
     layer1_out[2820] <= layer0_out[916];
     layer1_out[2821] <= layer0_out[9498] & ~layer0_out[9497];
     layer1_out[2822] <= layer0_out[4267] | layer0_out[4268];
     layer1_out[2823] <= ~layer0_out[7662];
     layer1_out[2824] <= layer0_out[2898];
     layer1_out[2825] <= layer0_out[6837] & ~layer0_out[6838];
     layer1_out[2826] <= 1'b1;
     layer1_out[2827] <= ~layer0_out[4429];
     layer1_out[2828] <= layer0_out[4992] ^ layer0_out[4993];
     layer1_out[2829] <= ~layer0_out[8074];
     layer1_out[2830] <= layer0_out[1484] & layer0_out[1485];
     layer1_out[2831] <= ~(layer0_out[7376] ^ layer0_out[7377]);
     layer1_out[2832] <= layer0_out[11971] ^ layer0_out[11972];
     layer1_out[2833] <= layer0_out[7718] | layer0_out[7719];
     layer1_out[2834] <= ~layer0_out[3898];
     layer1_out[2835] <= layer0_out[8695] & ~layer0_out[8694];
     layer1_out[2836] <= layer0_out[5063];
     layer1_out[2837] <= layer0_out[8164] ^ layer0_out[8165];
     layer1_out[2838] <= ~layer0_out[9746];
     layer1_out[2839] <= ~(layer0_out[861] | layer0_out[862]);
     layer1_out[2840] <= 1'b1;
     layer1_out[2841] <= ~layer0_out[7151];
     layer1_out[2842] <= ~(layer0_out[4492] | layer0_out[4493]);
     layer1_out[2843] <= ~(layer0_out[10104] | layer0_out[10105]);
     layer1_out[2844] <= ~layer0_out[2897] | layer0_out[2896];
     layer1_out[2845] <= ~layer0_out[3989];
     layer1_out[2846] <= ~layer0_out[994] | layer0_out[993];
     layer1_out[2847] <= layer0_out[5243] | layer0_out[5244];
     layer1_out[2848] <= ~layer0_out[5479];
     layer1_out[2849] <= layer0_out[6794] ^ layer0_out[6795];
     layer1_out[2850] <= ~(layer0_out[7492] & layer0_out[7493]);
     layer1_out[2851] <= layer0_out[7915] & ~layer0_out[7916];
     layer1_out[2852] <= ~layer0_out[8515];
     layer1_out[2853] <= layer0_out[4544] & layer0_out[4545];
     layer1_out[2854] <= layer0_out[1922] & layer0_out[1923];
     layer1_out[2855] <= ~layer0_out[9700] | layer0_out[9701];
     layer1_out[2856] <= ~(layer0_out[6172] & layer0_out[6173]);
     layer1_out[2857] <= layer0_out[4886] & layer0_out[4887];
     layer1_out[2858] <= ~(layer0_out[4850] ^ layer0_out[4851]);
     layer1_out[2859] <= layer0_out[6085] & ~layer0_out[6086];
     layer1_out[2860] <= ~(layer0_out[446] & layer0_out[447]);
     layer1_out[2861] <= layer0_out[6029];
     layer1_out[2862] <= ~layer0_out[5873] | layer0_out[5872];
     layer1_out[2863] <= layer0_out[701] & ~layer0_out[700];
     layer1_out[2864] <= layer0_out[11719];
     layer1_out[2865] <= layer0_out[3040] & ~layer0_out[3039];
     layer1_out[2866] <= layer0_out[6327] & layer0_out[6328];
     layer1_out[2867] <= ~(layer0_out[1293] | layer0_out[1294]);
     layer1_out[2868] <= layer0_out[10293];
     layer1_out[2869] <= ~(layer0_out[6907] & layer0_out[6908]);
     layer1_out[2870] <= ~layer0_out[10322];
     layer1_out[2871] <= ~(layer0_out[10765] & layer0_out[10766]);
     layer1_out[2872] <= ~layer0_out[12];
     layer1_out[2873] <= ~layer0_out[6609] | layer0_out[6608];
     layer1_out[2874] <= layer0_out[5515] | layer0_out[5516];
     layer1_out[2875] <= layer0_out[11007] ^ layer0_out[11008];
     layer1_out[2876] <= layer0_out[2623] & layer0_out[2624];
     layer1_out[2877] <= ~layer0_out[3551];
     layer1_out[2878] <= ~layer0_out[9497] | layer0_out[9496];
     layer1_out[2879] <= layer0_out[2680];
     layer1_out[2880] <= layer0_out[4655] | layer0_out[4656];
     layer1_out[2881] <= ~layer0_out[8902];
     layer1_out[2882] <= ~layer0_out[1997] | layer0_out[1998];
     layer1_out[2883] <= ~layer0_out[11945] | layer0_out[11946];
     layer1_out[2884] <= layer0_out[8275] & ~layer0_out[8274];
     layer1_out[2885] <= layer0_out[7324];
     layer1_out[2886] <= 1'b1;
     layer1_out[2887] <= layer0_out[5405] ^ layer0_out[5406];
     layer1_out[2888] <= ~layer0_out[2521];
     layer1_out[2889] <= ~layer0_out[3515];
     layer1_out[2890] <= ~layer0_out[48] | layer0_out[49];
     layer1_out[2891] <= layer0_out[8717] ^ layer0_out[8718];
     layer1_out[2892] <= ~layer0_out[9024];
     layer1_out[2893] <= layer0_out[2337] & ~layer0_out[2338];
     layer1_out[2894] <= layer0_out[4341] & ~layer0_out[4342];
     layer1_out[2895] <= layer0_out[10352];
     layer1_out[2896] <= layer0_out[2085] & layer0_out[2086];
     layer1_out[2897] <= layer0_out[7349] | layer0_out[7350];
     layer1_out[2898] <= ~layer0_out[7872] | layer0_out[7873];
     layer1_out[2899] <= 1'b0;
     layer1_out[2900] <= ~layer0_out[7584];
     layer1_out[2901] <= ~layer0_out[9484];
     layer1_out[2902] <= ~layer0_out[3859];
     layer1_out[2903] <= layer0_out[9194] | layer0_out[9195];
     layer1_out[2904] <= layer0_out[7656];
     layer1_out[2905] <= layer0_out[4980];
     layer1_out[2906] <= layer0_out[7787] & ~layer0_out[7788];
     layer1_out[2907] <= layer0_out[10363];
     layer1_out[2908] <= ~layer0_out[10921];
     layer1_out[2909] <= layer0_out[5322] & ~layer0_out[5321];
     layer1_out[2910] <= layer0_out[8088];
     layer1_out[2911] <= layer0_out[4606] & ~layer0_out[4605];
     layer1_out[2912] <= layer0_out[5072];
     layer1_out[2913] <= ~layer0_out[2493] | layer0_out[2492];
     layer1_out[2914] <= ~layer0_out[1573];
     layer1_out[2915] <= ~(layer0_out[9837] | layer0_out[9838]);
     layer1_out[2916] <= layer0_out[3283] & ~layer0_out[3284];
     layer1_out[2917] <= layer0_out[11510] & layer0_out[11511];
     layer1_out[2918] <= ~(layer0_out[5561] & layer0_out[5562]);
     layer1_out[2919] <= layer0_out[6504] | layer0_out[6505];
     layer1_out[2920] <= ~layer0_out[5965];
     layer1_out[2921] <= layer0_out[11819] & layer0_out[11820];
     layer1_out[2922] <= ~(layer0_out[1604] & layer0_out[1605]);
     layer1_out[2923] <= ~layer0_out[985];
     layer1_out[2924] <= layer0_out[6515] & ~layer0_out[6514];
     layer1_out[2925] <= layer0_out[10592] & ~layer0_out[10591];
     layer1_out[2926] <= layer0_out[4650];
     layer1_out[2927] <= ~layer0_out[3838];
     layer1_out[2928] <= layer0_out[6539] & layer0_out[6540];
     layer1_out[2929] <= layer0_out[2576] ^ layer0_out[2577];
     layer1_out[2930] <= layer0_out[9198] & ~layer0_out[9199];
     layer1_out[2931] <= ~(layer0_out[11907] | layer0_out[11908]);
     layer1_out[2932] <= ~layer0_out[5777] | layer0_out[5778];
     layer1_out[2933] <= ~layer0_out[10651];
     layer1_out[2934] <= layer0_out[951];
     layer1_out[2935] <= layer0_out[11473];
     layer1_out[2936] <= layer0_out[7029];
     layer1_out[2937] <= layer0_out[2128];
     layer1_out[2938] <= ~(layer0_out[7087] & layer0_out[7088]);
     layer1_out[2939] <= ~layer0_out[7064];
     layer1_out[2940] <= layer0_out[351];
     layer1_out[2941] <= ~layer0_out[3922] | layer0_out[3923];
     layer1_out[2942] <= layer0_out[2203] & ~layer0_out[2202];
     layer1_out[2943] <= ~(layer0_out[513] & layer0_out[514]);
     layer1_out[2944] <= layer0_out[6745] & ~layer0_out[6746];
     layer1_out[2945] <= ~layer0_out[9464] | layer0_out[9465];
     layer1_out[2946] <= ~layer0_out[11934];
     layer1_out[2947] <= ~layer0_out[5067];
     layer1_out[2948] <= ~layer0_out[3411] | layer0_out[3412];
     layer1_out[2949] <= layer0_out[7441];
     layer1_out[2950] <= ~(layer0_out[11514] & layer0_out[11515]);
     layer1_out[2951] <= layer0_out[727] | layer0_out[728];
     layer1_out[2952] <= ~layer0_out[3383];
     layer1_out[2953] <= layer0_out[2335];
     layer1_out[2954] <= ~layer0_out[2349];
     layer1_out[2955] <= ~(layer0_out[7839] & layer0_out[7840]);
     layer1_out[2956] <= 1'b0;
     layer1_out[2957] <= layer0_out[5178] ^ layer0_out[5179];
     layer1_out[2958] <= layer0_out[4594] | layer0_out[4595];
     layer1_out[2959] <= layer0_out[6847] | layer0_out[6848];
     layer1_out[2960] <= ~layer0_out[530] | layer0_out[531];
     layer1_out[2961] <= ~layer0_out[11534];
     layer1_out[2962] <= ~layer0_out[9588];
     layer1_out[2963] <= ~layer0_out[8743];
     layer1_out[2964] <= ~layer0_out[11199] | layer0_out[11198];
     layer1_out[2965] <= ~layer0_out[4147] | layer0_out[4148];
     layer1_out[2966] <= layer0_out[10772] | layer0_out[10773];
     layer1_out[2967] <= ~layer0_out[8834] | layer0_out[8835];
     layer1_out[2968] <= ~layer0_out[6489];
     layer1_out[2969] <= ~layer0_out[957] | layer0_out[958];
     layer1_out[2970] <= layer0_out[383] & layer0_out[384];
     layer1_out[2971] <= ~layer0_out[2019] | layer0_out[2018];
     layer1_out[2972] <= ~(layer0_out[2342] & layer0_out[2343]);
     layer1_out[2973] <= ~layer0_out[2109] | layer0_out[2108];
     layer1_out[2974] <= layer0_out[437];
     layer1_out[2975] <= 1'b1;
     layer1_out[2976] <= 1'b0;
     layer1_out[2977] <= layer0_out[8584];
     layer1_out[2978] <= layer0_out[4782] & ~layer0_out[4781];
     layer1_out[2979] <= layer0_out[8553] & layer0_out[8554];
     layer1_out[2980] <= layer0_out[7637] & ~layer0_out[7636];
     layer1_out[2981] <= ~layer0_out[8941];
     layer1_out[2982] <= layer0_out[93] & ~layer0_out[94];
     layer1_out[2983] <= ~(layer0_out[10245] | layer0_out[10246]);
     layer1_out[2984] <= ~(layer0_out[9272] ^ layer0_out[9273]);
     layer1_out[2985] <= layer0_out[1064];
     layer1_out[2986] <= ~layer0_out[8090] | layer0_out[8091];
     layer1_out[2987] <= layer0_out[1302];
     layer1_out[2988] <= ~layer0_out[8568];
     layer1_out[2989] <= layer0_out[7936] & layer0_out[7937];
     layer1_out[2990] <= layer0_out[11205] & ~layer0_out[11206];
     layer1_out[2991] <= 1'b0;
     layer1_out[2992] <= layer0_out[6500];
     layer1_out[2993] <= ~layer0_out[7554] | layer0_out[7553];
     layer1_out[2994] <= layer0_out[2099] | layer0_out[2100];
     layer1_out[2995] <= ~layer0_out[8878] | layer0_out[8879];
     layer1_out[2996] <= ~layer0_out[2798] | layer0_out[2797];
     layer1_out[2997] <= ~(layer0_out[8859] & layer0_out[8860]);
     layer1_out[2998] <= layer0_out[4120] & layer0_out[4121];
     layer1_out[2999] <= ~layer0_out[9882] | layer0_out[9883];
     layer1_out[3000] <= ~layer0_out[2572] | layer0_out[2571];
     layer1_out[3001] <= ~layer0_out[11939] | layer0_out[11940];
     layer1_out[3002] <= layer0_out[5125];
     layer1_out[3003] <= layer0_out[5970] & layer0_out[5971];
     layer1_out[3004] <= layer0_out[8836];
     layer1_out[3005] <= ~layer0_out[7967] | layer0_out[7968];
     layer1_out[3006] <= layer0_out[8786] & layer0_out[8787];
     layer1_out[3007] <= layer0_out[6464] & ~layer0_out[6465];
     layer1_out[3008] <= layer0_out[9689] & layer0_out[9690];
     layer1_out[3009] <= ~layer0_out[8439] | layer0_out[8438];
     layer1_out[3010] <= layer0_out[1878];
     layer1_out[3011] <= ~(layer0_out[11005] | layer0_out[11006]);
     layer1_out[3012] <= ~(layer0_out[10433] ^ layer0_out[10434]);
     layer1_out[3013] <= layer0_out[8349] | layer0_out[8350];
     layer1_out[3014] <= ~(layer0_out[3950] & layer0_out[3951]);
     layer1_out[3015] <= 1'b0;
     layer1_out[3016] <= layer0_out[1977];
     layer1_out[3017] <= layer0_out[11739] | layer0_out[11740];
     layer1_out[3018] <= ~layer0_out[167] | layer0_out[166];
     layer1_out[3019] <= ~(layer0_out[5409] & layer0_out[5410]);
     layer1_out[3020] <= ~layer0_out[11399] | layer0_out[11400];
     layer1_out[3021] <= layer0_out[4145] & ~layer0_out[4146];
     layer1_out[3022] <= layer0_out[200];
     layer1_out[3023] <= ~(layer0_out[4329] | layer0_out[4330]);
     layer1_out[3024] <= layer0_out[2055] & layer0_out[2056];
     layer1_out[3025] <= layer0_out[9188] | layer0_out[9189];
     layer1_out[3026] <= layer0_out[11857] & layer0_out[11858];
     layer1_out[3027] <= ~(layer0_out[3052] | layer0_out[3053]);
     layer1_out[3028] <= ~(layer0_out[11532] & layer0_out[11533]);
     layer1_out[3029] <= ~(layer0_out[6680] | layer0_out[6681]);
     layer1_out[3030] <= layer0_out[2877] & layer0_out[2878];
     layer1_out[3031] <= layer0_out[5526];
     layer1_out[3032] <= layer0_out[6914] ^ layer0_out[6915];
     layer1_out[3033] <= ~(layer0_out[2739] | layer0_out[2740]);
     layer1_out[3034] <= layer0_out[10253] & ~layer0_out[10254];
     layer1_out[3035] <= ~layer0_out[3439];
     layer1_out[3036] <= layer0_out[3692] & layer0_out[3693];
     layer1_out[3037] <= layer0_out[8912] ^ layer0_out[8913];
     layer1_out[3038] <= 1'b0;
     layer1_out[3039] <= ~layer0_out[318];
     layer1_out[3040] <= 1'b1;
     layer1_out[3041] <= layer0_out[10497] & ~layer0_out[10496];
     layer1_out[3042] <= ~(layer0_out[4845] ^ layer0_out[4846]);
     layer1_out[3043] <= ~layer0_out[9127];
     layer1_out[3044] <= layer0_out[10313];
     layer1_out[3045] <= ~(layer0_out[6233] ^ layer0_out[6234]);
     layer1_out[3046] <= 1'b0;
     layer1_out[3047] <= layer0_out[1001] & ~layer0_out[1000];
     layer1_out[3048] <= layer0_out[3066] | layer0_out[3067];
     layer1_out[3049] <= 1'b0;
     layer1_out[3050] <= layer0_out[3798];
     layer1_out[3051] <= layer0_out[9993] | layer0_out[9994];
     layer1_out[3052] <= ~layer0_out[4710] | layer0_out[4711];
     layer1_out[3053] <= layer0_out[6808] | layer0_out[6809];
     layer1_out[3054] <= layer0_out[5979];
     layer1_out[3055] <= ~(layer0_out[3539] & layer0_out[3540]);
     layer1_out[3056] <= ~layer0_out[1631];
     layer1_out[3057] <= ~(layer0_out[489] | layer0_out[490]);
     layer1_out[3058] <= layer0_out[4208] & ~layer0_out[4207];
     layer1_out[3059] <= ~(layer0_out[4296] & layer0_out[4297]);
     layer1_out[3060] <= layer0_out[6972] & ~layer0_out[6971];
     layer1_out[3061] <= layer0_out[3549] & ~layer0_out[3548];
     layer1_out[3062] <= layer0_out[4525];
     layer1_out[3063] <= layer0_out[6438] ^ layer0_out[6439];
     layer1_out[3064] <= 1'b1;
     layer1_out[3065] <= ~(layer0_out[5650] ^ layer0_out[5651]);
     layer1_out[3066] <= layer0_out[2169] & layer0_out[2170];
     layer1_out[3067] <= layer0_out[1111] & layer0_out[1112];
     layer1_out[3068] <= layer0_out[6875];
     layer1_out[3069] <= ~layer0_out[4989];
     layer1_out[3070] <= layer0_out[10732];
     layer1_out[3071] <= layer0_out[1533];
     layer1_out[3072] <= layer0_out[4003] ^ layer0_out[4004];
     layer1_out[3073] <= layer0_out[7353];
     layer1_out[3074] <= layer0_out[2471];
     layer1_out[3075] <= 1'b0;
     layer1_out[3076] <= layer0_out[7865];
     layer1_out[3077] <= ~layer0_out[4725];
     layer1_out[3078] <= layer0_out[9567] & ~layer0_out[9568];
     layer1_out[3079] <= layer0_out[11576] & ~layer0_out[11575];
     layer1_out[3080] <= ~layer0_out[1917];
     layer1_out[3081] <= layer0_out[2505] | layer0_out[2506];
     layer1_out[3082] <= layer0_out[4933];
     layer1_out[3083] <= layer0_out[5476] ^ layer0_out[5477];
     layer1_out[3084] <= ~layer0_out[3333];
     layer1_out[3085] <= ~(layer0_out[1242] & layer0_out[1243]);
     layer1_out[3086] <= ~layer0_out[9633] | layer0_out[9634];
     layer1_out[3087] <= layer0_out[10906] ^ layer0_out[10907];
     layer1_out[3088] <= layer0_out[5502];
     layer1_out[3089] <= layer0_out[2953] ^ layer0_out[2954];
     layer1_out[3090] <= layer0_out[7265];
     layer1_out[3091] <= layer0_out[1259] & ~layer0_out[1258];
     layer1_out[3092] <= layer0_out[7815] & ~layer0_out[7814];
     layer1_out[3093] <= ~(layer0_out[7061] ^ layer0_out[7062]);
     layer1_out[3094] <= ~(layer0_out[484] | layer0_out[485]);
     layer1_out[3095] <= layer0_out[9337] & layer0_out[9338];
     layer1_out[3096] <= ~layer0_out[4480] | layer0_out[4479];
     layer1_out[3097] <= ~layer0_out[9103] | layer0_out[9104];
     layer1_out[3098] <= layer0_out[7313] ^ layer0_out[7314];
     layer1_out[3099] <= ~layer0_out[10759];
     layer1_out[3100] <= ~layer0_out[851] | layer0_out[850];
     layer1_out[3101] <= ~layer0_out[8185];
     layer1_out[3102] <= ~(layer0_out[9392] | layer0_out[9393]);
     layer1_out[3103] <= layer0_out[418];
     layer1_out[3104] <= ~layer0_out[5188];
     layer1_out[3105] <= 1'b1;
     layer1_out[3106] <= layer0_out[1364] & ~layer0_out[1365];
     layer1_out[3107] <= layer0_out[5301] & ~layer0_out[5300];
     layer1_out[3108] <= ~(layer0_out[9286] ^ layer0_out[9287]);
     layer1_out[3109] <= layer0_out[2453] & ~layer0_out[2454];
     layer1_out[3110] <= ~layer0_out[3972];
     layer1_out[3111] <= ~(layer0_out[11453] ^ layer0_out[11454]);
     layer1_out[3112] <= layer0_out[5048];
     layer1_out[3113] <= ~layer0_out[9049];
     layer1_out[3114] <= ~(layer0_out[11551] | layer0_out[11552]);
     layer1_out[3115] <= ~(layer0_out[5407] ^ layer0_out[5408]);
     layer1_out[3116] <= layer0_out[1329] & ~layer0_out[1330];
     layer1_out[3117] <= layer0_out[11987] | layer0_out[11988];
     layer1_out[3118] <= layer0_out[10331] & layer0_out[10332];
     layer1_out[3119] <= layer0_out[11171];
     layer1_out[3120] <= ~layer0_out[11913] | layer0_out[11914];
     layer1_out[3121] <= layer0_out[7930] & ~layer0_out[7929];
     layer1_out[3122] <= layer0_out[2248] | layer0_out[2249];
     layer1_out[3123] <= ~layer0_out[7549];
     layer1_out[3124] <= layer0_out[9660] | layer0_out[9661];
     layer1_out[3125] <= layer0_out[10371] ^ layer0_out[10372];
     layer1_out[3126] <= ~(layer0_out[6569] | layer0_out[6570]);
     layer1_out[3127] <= ~(layer0_out[10075] | layer0_out[10076]);
     layer1_out[3128] <= layer0_out[4813] & layer0_out[4814];
     layer1_out[3129] <= 1'b0;
     layer1_out[3130] <= ~layer0_out[11578] | layer0_out[11577];
     layer1_out[3131] <= layer0_out[5578];
     layer1_out[3132] <= layer0_out[6461] | layer0_out[6462];
     layer1_out[3133] <= layer0_out[8901] | layer0_out[8902];
     layer1_out[3134] <= ~(layer0_out[9110] & layer0_out[9111]);
     layer1_out[3135] <= layer0_out[11350];
     layer1_out[3136] <= ~layer0_out[2522];
     layer1_out[3137] <= ~(layer0_out[1010] & layer0_out[1011]);
     layer1_out[3138] <= ~layer0_out[5279];
     layer1_out[3139] <= ~(layer0_out[10638] | layer0_out[10639]);
     layer1_out[3140] <= layer0_out[9856];
     layer1_out[3141] <= layer0_out[1497] | layer0_out[1498];
     layer1_out[3142] <= ~layer0_out[1606] | layer0_out[1607];
     layer1_out[3143] <= layer0_out[11805];
     layer1_out[3144] <= ~(layer0_out[11070] & layer0_out[11071]);
     layer1_out[3145] <= layer0_out[4730] & ~layer0_out[4729];
     layer1_out[3146] <= ~(layer0_out[3199] ^ layer0_out[3200]);
     layer1_out[3147] <= layer0_out[2945];
     layer1_out[3148] <= layer0_out[9118];
     layer1_out[3149] <= layer0_out[575] | layer0_out[576];
     layer1_out[3150] <= layer0_out[8544] & ~layer0_out[8543];
     layer1_out[3151] <= layer0_out[4094] & ~layer0_out[4095];
     layer1_out[3152] <= layer0_out[6317] ^ layer0_out[6318];
     layer1_out[3153] <= layer0_out[8497] | layer0_out[8498];
     layer1_out[3154] <= layer0_out[8955] & ~layer0_out[8956];
     layer1_out[3155] <= layer0_out[8226];
     layer1_out[3156] <= layer0_out[10932] & layer0_out[10933];
     layer1_out[3157] <= 1'b1;
     layer1_out[3158] <= ~(layer0_out[3188] | layer0_out[3189]);
     layer1_out[3159] <= layer0_out[7723];
     layer1_out[3160] <= layer0_out[389];
     layer1_out[3161] <= layer0_out[6403] ^ layer0_out[6404];
     layer1_out[3162] <= 1'b1;
     layer1_out[3163] <= ~layer0_out[7055] | layer0_out[7054];
     layer1_out[3164] <= layer0_out[1769] & ~layer0_out[1770];
     layer1_out[3165] <= 1'b1;
     layer1_out[3166] <= ~layer0_out[6557];
     layer1_out[3167] <= ~layer0_out[7434] | layer0_out[7433];
     layer1_out[3168] <= layer0_out[3855];
     layer1_out[3169] <= layer0_out[9255];
     layer1_out[3170] <= ~layer0_out[4162] | layer0_out[4161];
     layer1_out[3171] <= ~layer0_out[11431] | layer0_out[11432];
     layer1_out[3172] <= ~layer0_out[8155];
     layer1_out[3173] <= ~(layer0_out[6848] & layer0_out[6849]);
     layer1_out[3174] <= layer0_out[6086] & ~layer0_out[6087];
     layer1_out[3175] <= ~layer0_out[2798] | layer0_out[2799];
     layer1_out[3176] <= layer0_out[7793] & layer0_out[7794];
     layer1_out[3177] <= ~layer0_out[10404] | layer0_out[10403];
     layer1_out[3178] <= layer0_out[8720];
     layer1_out[3179] <= ~layer0_out[7643] | layer0_out[7644];
     layer1_out[3180] <= layer0_out[8283] & ~layer0_out[8282];
     layer1_out[3181] <= ~layer0_out[9003];
     layer1_out[3182] <= ~layer0_out[6518] | layer0_out[6519];
     layer1_out[3183] <= layer0_out[3402];
     layer1_out[3184] <= ~layer0_out[879];
     layer1_out[3185] <= ~layer0_out[10560];
     layer1_out[3186] <= layer0_out[1048] & ~layer0_out[1049];
     layer1_out[3187] <= layer0_out[446];
     layer1_out[3188] <= ~(layer0_out[10062] ^ layer0_out[10063]);
     layer1_out[3189] <= ~(layer0_out[8600] | layer0_out[8601]);
     layer1_out[3190] <= ~layer0_out[404];
     layer1_out[3191] <= layer0_out[7352] | layer0_out[7353];
     layer1_out[3192] <= layer0_out[7853] & ~layer0_out[7854];
     layer1_out[3193] <= ~layer0_out[3236] | layer0_out[3237];
     layer1_out[3194] <= ~layer0_out[3584];
     layer1_out[3195] <= layer0_out[4325];
     layer1_out[3196] <= ~(layer0_out[6377] & layer0_out[6378]);
     layer1_out[3197] <= ~(layer0_out[4338] ^ layer0_out[4339]);
     layer1_out[3198] <= layer0_out[488];
     layer1_out[3199] <= layer0_out[11876] & layer0_out[11877];
     layer1_out[3200] <= layer0_out[10429];
     layer1_out[3201] <= layer0_out[8763];
     layer1_out[3202] <= ~(layer0_out[4465] ^ layer0_out[4466]);
     layer1_out[3203] <= layer0_out[11874] ^ layer0_out[11875];
     layer1_out[3204] <= ~(layer0_out[10191] | layer0_out[10192]);
     layer1_out[3205] <= layer0_out[4547] & layer0_out[4548];
     layer1_out[3206] <= ~layer0_out[2113];
     layer1_out[3207] <= ~layer0_out[2747];
     layer1_out[3208] <= layer0_out[2843] & layer0_out[2844];
     layer1_out[3209] <= layer0_out[6216] & ~layer0_out[6217];
     layer1_out[3210] <= layer0_out[7646] ^ layer0_out[7647];
     layer1_out[3211] <= layer0_out[6053];
     layer1_out[3212] <= ~layer0_out[1702];
     layer1_out[3213] <= layer0_out[5222];
     layer1_out[3214] <= ~layer0_out[2587] | layer0_out[2586];
     layer1_out[3215] <= ~(layer0_out[7355] | layer0_out[7356]);
     layer1_out[3216] <= layer0_out[11795] & ~layer0_out[11794];
     layer1_out[3217] <= ~layer0_out[9910];
     layer1_out[3218] <= ~(layer0_out[1254] | layer0_out[1255]);
     layer1_out[3219] <= layer0_out[1014] & ~layer0_out[1013];
     layer1_out[3220] <= layer0_out[5083] | layer0_out[5084];
     layer1_out[3221] <= layer0_out[3492];
     layer1_out[3222] <= layer0_out[4137] ^ layer0_out[4138];
     layer1_out[3223] <= ~layer0_out[7722];
     layer1_out[3224] <= layer0_out[1495] & ~layer0_out[1494];
     layer1_out[3225] <= ~layer0_out[7349];
     layer1_out[3226] <= layer0_out[1019];
     layer1_out[3227] <= layer0_out[8612] & ~layer0_out[8611];
     layer1_out[3228] <= ~layer0_out[11506];
     layer1_out[3229] <= ~(layer0_out[4399] ^ layer0_out[4400]);
     layer1_out[3230] <= layer0_out[9000];
     layer1_out[3231] <= layer0_out[11309];
     layer1_out[3232] <= layer0_out[1005];
     layer1_out[3233] <= layer0_out[2947] & ~layer0_out[2948];
     layer1_out[3234] <= ~layer0_out[549] | layer0_out[548];
     layer1_out[3235] <= layer0_out[7056] & layer0_out[7057];
     layer1_out[3236] <= layer0_out[11369] & layer0_out[11370];
     layer1_out[3237] <= layer0_out[9170];
     layer1_out[3238] <= ~layer0_out[995] | layer0_out[996];
     layer1_out[3239] <= ~(layer0_out[406] | layer0_out[407]);
     layer1_out[3240] <= ~layer0_out[8558];
     layer1_out[3241] <= layer0_out[257] & ~layer0_out[256];
     layer1_out[3242] <= layer0_out[8068];
     layer1_out[3243] <= 1'b1;
     layer1_out[3244] <= layer0_out[2862] | layer0_out[2863];
     layer1_out[3245] <= ~layer0_out[7478];
     layer1_out[3246] <= layer0_out[1935];
     layer1_out[3247] <= layer0_out[5546];
     layer1_out[3248] <= layer0_out[4490] & layer0_out[4491];
     layer1_out[3249] <= 1'b0;
     layer1_out[3250] <= layer0_out[8053] | layer0_out[8054];
     layer1_out[3251] <= layer0_out[11610] & ~layer0_out[11611];
     layer1_out[3252] <= layer0_out[955] & ~layer0_out[956];
     layer1_out[3253] <= layer0_out[11339] | layer0_out[11340];
     layer1_out[3254] <= 1'b1;
     layer1_out[3255] <= layer0_out[1041];
     layer1_out[3256] <= ~layer0_out[1013];
     layer1_out[3257] <= ~layer0_out[7895];
     layer1_out[3258] <= layer0_out[9031] & ~layer0_out[9030];
     layer1_out[3259] <= ~layer0_out[9231];
     layer1_out[3260] <= ~layer0_out[4117];
     layer1_out[3261] <= ~layer0_out[904] | layer0_out[903];
     layer1_out[3262] <= layer0_out[2358];
     layer1_out[3263] <= layer0_out[11578] ^ layer0_out[11579];
     layer1_out[3264] <= ~layer0_out[11801];
     layer1_out[3265] <= ~layer0_out[7844] | layer0_out[7845];
     layer1_out[3266] <= layer0_out[3068] | layer0_out[3069];
     layer1_out[3267] <= ~(layer0_out[1214] & layer0_out[1215]);
     layer1_out[3268] <= ~(layer0_out[9645] | layer0_out[9646]);
     layer1_out[3269] <= ~layer0_out[8767] | layer0_out[8768];
     layer1_out[3270] <= layer0_out[276] | layer0_out[277];
     layer1_out[3271] <= layer0_out[45] & ~layer0_out[46];
     layer1_out[3272] <= layer0_out[283] & layer0_out[284];
     layer1_out[3273] <= ~layer0_out[1071];
     layer1_out[3274] <= ~layer0_out[2834];
     layer1_out[3275] <= ~(layer0_out[7470] & layer0_out[7471]);
     layer1_out[3276] <= ~layer0_out[4636];
     layer1_out[3277] <= layer0_out[8262] & ~layer0_out[8263];
     layer1_out[3278] <= ~layer0_out[9583];
     layer1_out[3279] <= layer0_out[8336] | layer0_out[8337];
     layer1_out[3280] <= layer0_out[4286];
     layer1_out[3281] <= 1'b0;
     layer1_out[3282] <= ~layer0_out[8059] | layer0_out[8058];
     layer1_out[3283] <= layer0_out[4772] & layer0_out[4773];
     layer1_out[3284] <= ~layer0_out[5026] | layer0_out[5025];
     layer1_out[3285] <= layer0_out[143];
     layer1_out[3286] <= layer0_out[4483] & layer0_out[4484];
     layer1_out[3287] <= layer0_out[4662];
     layer1_out[3288] <= 1'b0;
     layer1_out[3289] <= layer0_out[6394] & ~layer0_out[6395];
     layer1_out[3290] <= layer0_out[4075] & layer0_out[4076];
     layer1_out[3291] <= ~layer0_out[2628] | layer0_out[2629];
     layer1_out[3292] <= ~layer0_out[5262];
     layer1_out[3293] <= layer0_out[4162] & ~layer0_out[4163];
     layer1_out[3294] <= ~(layer0_out[10468] ^ layer0_out[10469]);
     layer1_out[3295] <= layer0_out[2439];
     layer1_out[3296] <= layer0_out[2877];
     layer1_out[3297] <= layer0_out[6340];
     layer1_out[3298] <= ~(layer0_out[3700] & layer0_out[3701]);
     layer1_out[3299] <= layer0_out[3536] ^ layer0_out[3537];
     layer1_out[3300] <= ~layer0_out[2083] | layer0_out[2082];
     layer1_out[3301] <= layer0_out[5050];
     layer1_out[3302] <= ~layer0_out[2207] | layer0_out[2208];
     layer1_out[3303] <= layer0_out[2373] & ~layer0_out[2372];
     layer1_out[3304] <= layer0_out[4560] & layer0_out[4561];
     layer1_out[3305] <= ~layer0_out[4921];
     layer1_out[3306] <= ~layer0_out[1304] | layer0_out[1303];
     layer1_out[3307] <= ~layer0_out[10024] | layer0_out[10023];
     layer1_out[3308] <= layer0_out[2062] | layer0_out[2063];
     layer1_out[3309] <= ~layer0_out[6579];
     layer1_out[3310] <= layer0_out[6100] & ~layer0_out[6101];
     layer1_out[3311] <= layer0_out[2173];
     layer1_out[3312] <= ~(layer0_out[730] & layer0_out[731]);
     layer1_out[3313] <= layer0_out[10700] | layer0_out[10701];
     layer1_out[3314] <= layer0_out[11687] & layer0_out[11688];
     layer1_out[3315] <= layer0_out[1370];
     layer1_out[3316] <= layer0_out[8872] & ~layer0_out[8871];
     layer1_out[3317] <= layer0_out[11597];
     layer1_out[3318] <= layer0_out[8979] & layer0_out[8980];
     layer1_out[3319] <= ~layer0_out[5199];
     layer1_out[3320] <= layer0_out[10625] | layer0_out[10626];
     layer1_out[3321] <= ~(layer0_out[4716] | layer0_out[4717]);
     layer1_out[3322] <= layer0_out[7099] & layer0_out[7100];
     layer1_out[3323] <= ~layer0_out[9286];
     layer1_out[3324] <= ~(layer0_out[6687] & layer0_out[6688]);
     layer1_out[3325] <= layer0_out[1737] & ~layer0_out[1736];
     layer1_out[3326] <= 1'b1;
     layer1_out[3327] <= ~(layer0_out[9042] | layer0_out[9043]);
     layer1_out[3328] <= ~(layer0_out[6604] ^ layer0_out[6605]);
     layer1_out[3329] <= ~layer0_out[3859] | layer0_out[3858];
     layer1_out[3330] <= layer0_out[8572];
     layer1_out[3331] <= ~layer0_out[7205] | layer0_out[7206];
     layer1_out[3332] <= layer0_out[8400] & ~layer0_out[8399];
     layer1_out[3333] <= layer0_out[8278];
     layer1_out[3334] <= layer0_out[6435] ^ layer0_out[6436];
     layer1_out[3335] <= layer0_out[7477] & ~layer0_out[7476];
     layer1_out[3336] <= ~(layer0_out[2272] & layer0_out[2273]);
     layer1_out[3337] <= 1'b1;
     layer1_out[3338] <= ~layer0_out[830];
     layer1_out[3339] <= layer0_out[337];
     layer1_out[3340] <= ~(layer0_out[2151] ^ layer0_out[2152]);
     layer1_out[3341] <= layer0_out[8232];
     layer1_out[3342] <= ~layer0_out[4664];
     layer1_out[3343] <= layer0_out[5553] & ~layer0_out[5554];
     layer1_out[3344] <= layer0_out[11626];
     layer1_out[3345] <= ~layer0_out[2860] | layer0_out[2861];
     layer1_out[3346] <= ~(layer0_out[9196] | layer0_out[9197]);
     layer1_out[3347] <= layer0_out[3246];
     layer1_out[3348] <= ~layer0_out[3456] | layer0_out[3457];
     layer1_out[3349] <= 1'b0;
     layer1_out[3350] <= ~layer0_out[9639];
     layer1_out[3351] <= layer0_out[1034] & ~layer0_out[1035];
     layer1_out[3352] <= ~(layer0_out[10055] & layer0_out[10056]);
     layer1_out[3353] <= layer0_out[2760] & ~layer0_out[2759];
     layer1_out[3354] <= ~(layer0_out[9866] ^ layer0_out[9867]);
     layer1_out[3355] <= ~(layer0_out[2821] | layer0_out[2822]);
     layer1_out[3356] <= layer0_out[10977];
     layer1_out[3357] <= layer0_out[1105] & layer0_out[1106];
     layer1_out[3358] <= ~(layer0_out[4826] & layer0_out[4827]);
     layer1_out[3359] <= layer0_out[6925] ^ layer0_out[6926];
     layer1_out[3360] <= ~(layer0_out[8075] | layer0_out[8076]);
     layer1_out[3361] <= layer0_out[1817];
     layer1_out[3362] <= layer0_out[10940];
     layer1_out[3363] <= layer0_out[9002];
     layer1_out[3364] <= ~(layer0_out[2006] & layer0_out[2007]);
     layer1_out[3365] <= layer0_out[9834];
     layer1_out[3366] <= layer0_out[6262];
     layer1_out[3367] <= 1'b1;
     layer1_out[3368] <= ~(layer0_out[10167] | layer0_out[10168]);
     layer1_out[3369] <= ~layer0_out[6135];
     layer1_out[3370] <= ~layer0_out[9025] | layer0_out[9026];
     layer1_out[3371] <= layer0_out[9537] ^ layer0_out[9538];
     layer1_out[3372] <= ~(layer0_out[5856] | layer0_out[5857]);
     layer1_out[3373] <= layer0_out[607] & ~layer0_out[606];
     layer1_out[3374] <= ~layer0_out[10361];
     layer1_out[3375] <= 1'b0;
     layer1_out[3376] <= ~(layer0_out[1476] | layer0_out[1477]);
     layer1_out[3377] <= layer0_out[2153] | layer0_out[2154];
     layer1_out[3378] <= 1'b1;
     layer1_out[3379] <= ~(layer0_out[11322] | layer0_out[11323]);
     layer1_out[3380] <= ~layer0_out[6775];
     layer1_out[3381] <= ~layer0_out[10875];
     layer1_out[3382] <= layer0_out[10998] ^ layer0_out[10999];
     layer1_out[3383] <= layer0_out[5623] | layer0_out[5624];
     layer1_out[3384] <= ~(layer0_out[789] | layer0_out[790]);
     layer1_out[3385] <= layer0_out[10030] & layer0_out[10031];
     layer1_out[3386] <= layer0_out[3661];
     layer1_out[3387] <= layer0_out[1119] | layer0_out[1120];
     layer1_out[3388] <= ~layer0_out[4885] | layer0_out[4884];
     layer1_out[3389] <= layer0_out[1823];
     layer1_out[3390] <= ~layer0_out[11031];
     layer1_out[3391] <= layer0_out[10419] & layer0_out[10420];
     layer1_out[3392] <= layer0_out[10445];
     layer1_out[3393] <= ~layer0_out[906] | layer0_out[907];
     layer1_out[3394] <= ~layer0_out[76] | layer0_out[77];
     layer1_out[3395] <= layer0_out[7082];
     layer1_out[3396] <= ~layer0_out[11928] | layer0_out[11929];
     layer1_out[3397] <= layer0_out[1696];
     layer1_out[3398] <= layer0_out[5012] & layer0_out[5013];
     layer1_out[3399] <= layer0_out[9382] | layer0_out[9383];
     layer1_out[3400] <= layer0_out[9296];
     layer1_out[3401] <= ~layer0_out[7776] | layer0_out[7777];
     layer1_out[3402] <= ~layer0_out[9770];
     layer1_out[3403] <= layer0_out[6773] & ~layer0_out[6772];
     layer1_out[3404] <= layer0_out[321];
     layer1_out[3405] <= layer0_out[6674];
     layer1_out[3406] <= layer0_out[3814];
     layer1_out[3407] <= layer0_out[7742] & ~layer0_out[7743];
     layer1_out[3408] <= layer0_out[4364] ^ layer0_out[4365];
     layer1_out[3409] <= ~layer0_out[9444] | layer0_out[9445];
     layer1_out[3410] <= ~(layer0_out[2400] | layer0_out[2401]);
     layer1_out[3411] <= layer0_out[6783] & ~layer0_out[6782];
     layer1_out[3412] <= ~(layer0_out[8264] | layer0_out[8265]);
     layer1_out[3413] <= ~(layer0_out[4829] | layer0_out[4830]);
     layer1_out[3414] <= layer0_out[9331] | layer0_out[9332];
     layer1_out[3415] <= ~layer0_out[911] | layer0_out[910];
     layer1_out[3416] <= ~layer0_out[8530] | layer0_out[8529];
     layer1_out[3417] <= ~layer0_out[5893];
     layer1_out[3418] <= layer0_out[2489] | layer0_out[2490];
     layer1_out[3419] <= layer0_out[2008] & layer0_out[2009];
     layer1_out[3420] <= 1'b0;
     layer1_out[3421] <= ~layer0_out[9542];
     layer1_out[3422] <= layer0_out[6007] ^ layer0_out[6008];
     layer1_out[3423] <= ~layer0_out[1694];
     layer1_out[3424] <= layer0_out[6816] & ~layer0_out[6817];
     layer1_out[3425] <= ~layer0_out[6595] | layer0_out[6594];
     layer1_out[3426] <= layer0_out[2052] & ~layer0_out[2051];
     layer1_out[3427] <= layer0_out[10982];
     layer1_out[3428] <= layer0_out[3687] & layer0_out[3688];
     layer1_out[3429] <= layer0_out[6829];
     layer1_out[3430] <= layer0_out[496] & ~layer0_out[497];
     layer1_out[3431] <= ~layer0_out[938];
     layer1_out[3432] <= ~layer0_out[9250] | layer0_out[9249];
     layer1_out[3433] <= 1'b0;
     layer1_out[3434] <= ~(layer0_out[2931] & layer0_out[2932]);
     layer1_out[3435] <= layer0_out[8606] & layer0_out[8607];
     layer1_out[3436] <= layer0_out[8034] | layer0_out[8035];
     layer1_out[3437] <= layer0_out[5878];
     layer1_out[3438] <= ~layer0_out[9241];
     layer1_out[3439] <= layer0_out[1712];
     layer1_out[3440] <= ~(layer0_out[7902] | layer0_out[7903]);
     layer1_out[3441] <= layer0_out[7961] & layer0_out[7962];
     layer1_out[3442] <= layer0_out[641];
     layer1_out[3443] <= ~(layer0_out[8138] & layer0_out[8139]);
     layer1_out[3444] <= layer0_out[4785] | layer0_out[4786];
     layer1_out[3445] <= ~layer0_out[2854];
     layer1_out[3446] <= ~(layer0_out[11701] | layer0_out[11702]);
     layer1_out[3447] <= ~layer0_out[8318];
     layer1_out[3448] <= layer0_out[6983] & ~layer0_out[6984];
     layer1_out[3449] <= layer0_out[10766] & layer0_out[10767];
     layer1_out[3450] <= ~(layer0_out[5557] & layer0_out[5558]);
     layer1_out[3451] <= layer0_out[1190] & ~layer0_out[1191];
     layer1_out[3452] <= layer0_out[3683] & ~layer0_out[3684];
     layer1_out[3453] <= ~(layer0_out[250] & layer0_out[251]);
     layer1_out[3454] <= layer0_out[2504];
     layer1_out[3455] <= layer0_out[1214];
     layer1_out[3456] <= ~layer0_out[8729];
     layer1_out[3457] <= layer0_out[4445];
     layer1_out[3458] <= layer0_out[2429];
     layer1_out[3459] <= layer0_out[10312];
     layer1_out[3460] <= ~layer0_out[5700];
     layer1_out[3461] <= layer0_out[11952] & ~layer0_out[11951];
     layer1_out[3462] <= ~(layer0_out[2981] | layer0_out[2982]);
     layer1_out[3463] <= layer0_out[8777] ^ layer0_out[8778];
     layer1_out[3464] <= ~layer0_out[10684] | layer0_out[10683];
     layer1_out[3465] <= 1'b0;
     layer1_out[3466] <= ~layer0_out[3266];
     layer1_out[3467] <= layer0_out[3025];
     layer1_out[3468] <= ~(layer0_out[4825] & layer0_out[4826]);
     layer1_out[3469] <= ~(layer0_out[7852] ^ layer0_out[7853]);
     layer1_out[3470] <= ~layer0_out[664];
     layer1_out[3471] <= ~layer0_out[5201] | layer0_out[5200];
     layer1_out[3472] <= layer0_out[3194] & ~layer0_out[3193];
     layer1_out[3473] <= ~layer0_out[10570] | layer0_out[10571];
     layer1_out[3474] <= layer0_out[4012] & ~layer0_out[4013];
     layer1_out[3475] <= layer0_out[9253];
     layer1_out[3476] <= layer0_out[9654];
     layer1_out[3477] <= ~layer0_out[11376] | layer0_out[11375];
     layer1_out[3478] <= ~layer0_out[2905];
     layer1_out[3479] <= ~layer0_out[1750] | layer0_out[1751];
     layer1_out[3480] <= layer0_out[4538] & layer0_out[4539];
     layer1_out[3481] <= layer0_out[2529];
     layer1_out[3482] <= layer0_out[6020] ^ layer0_out[6021];
     layer1_out[3483] <= layer0_out[7810];
     layer1_out[3484] <= ~layer0_out[2935];
     layer1_out[3485] <= ~layer0_out[3523] | layer0_out[3524];
     layer1_out[3486] <= ~layer0_out[583] | layer0_out[584];
     layer1_out[3487] <= layer0_out[7274] | layer0_out[7275];
     layer1_out[3488] <= layer0_out[8192] & ~layer0_out[8191];
     layer1_out[3489] <= ~layer0_out[724] | layer0_out[723];
     layer1_out[3490] <= ~layer0_out[2040] | layer0_out[2039];
     layer1_out[3491] <= ~layer0_out[6833];
     layer1_out[3492] <= ~(layer0_out[6314] | layer0_out[6315]);
     layer1_out[3493] <= ~layer0_out[9059] | layer0_out[9058];
     layer1_out[3494] <= ~layer0_out[10675] | layer0_out[10676];
     layer1_out[3495] <= ~layer0_out[10597] | layer0_out[10596];
     layer1_out[3496] <= layer0_out[10691] | layer0_out[10692];
     layer1_out[3497] <= layer0_out[8223] & layer0_out[8224];
     layer1_out[3498] <= ~(layer0_out[2187] | layer0_out[2188]);
     layer1_out[3499] <= ~layer0_out[9011];
     layer1_out[3500] <= ~layer0_out[5702] | layer0_out[5703];
     layer1_out[3501] <= layer0_out[1453];
     layer1_out[3502] <= layer0_out[3953] ^ layer0_out[3954];
     layer1_out[3503] <= ~layer0_out[4761];
     layer1_out[3504] <= ~layer0_out[1140] | layer0_out[1141];
     layer1_out[3505] <= layer0_out[5461] & ~layer0_out[5460];
     layer1_out[3506] <= layer0_out[11284] & layer0_out[11285];
     layer1_out[3507] <= ~(layer0_out[1613] ^ layer0_out[1614]);
     layer1_out[3508] <= layer0_out[813] & ~layer0_out[812];
     layer1_out[3509] <= ~layer0_out[1311];
     layer1_out[3510] <= layer0_out[10697] & ~layer0_out[10698];
     layer1_out[3511] <= layer0_out[8661] & layer0_out[8662];
     layer1_out[3512] <= ~(layer0_out[3306] ^ layer0_out[3307]);
     layer1_out[3513] <= ~layer0_out[9900] | layer0_out[9899];
     layer1_out[3514] <= ~(layer0_out[194] & layer0_out[195]);
     layer1_out[3515] <= layer0_out[2180];
     layer1_out[3516] <= ~(layer0_out[702] & layer0_out[703]);
     layer1_out[3517] <= layer0_out[2822] | layer0_out[2823];
     layer1_out[3518] <= layer0_out[10800] & ~layer0_out[10799];
     layer1_out[3519] <= 1'b0;
     layer1_out[3520] <= layer0_out[3885] & ~layer0_out[3884];
     layer1_out[3521] <= layer0_out[6938];
     layer1_out[3522] <= ~(layer0_out[2522] & layer0_out[2523]);
     layer1_out[3523] <= ~(layer0_out[3141] & layer0_out[3142]);
     layer1_out[3524] <= layer0_out[4995] & layer0_out[4996];
     layer1_out[3525] <= ~(layer0_out[2158] & layer0_out[2159]);
     layer1_out[3526] <= layer0_out[543] & ~layer0_out[542];
     layer1_out[3527] <= layer0_out[4660];
     layer1_out[3528] <= ~layer0_out[5033];
     layer1_out[3529] <= ~(layer0_out[9309] ^ layer0_out[9310]);
     layer1_out[3530] <= ~layer0_out[10141];
     layer1_out[3531] <= ~layer0_out[7234] | layer0_out[7233];
     layer1_out[3532] <= ~layer0_out[169];
     layer1_out[3533] <= ~(layer0_out[10632] | layer0_out[10633]);
     layer1_out[3534] <= ~layer0_out[5170];
     layer1_out[3535] <= layer0_out[10024];
     layer1_out[3536] <= layer0_out[2978] & ~layer0_out[2977];
     layer1_out[3537] <= ~layer0_out[1274];
     layer1_out[3538] <= ~layer0_out[2669];
     layer1_out[3539] <= layer0_out[8564] | layer0_out[8565];
     layer1_out[3540] <= layer0_out[11312];
     layer1_out[3541] <= 1'b0;
     layer1_out[3542] <= ~layer0_out[5150] | layer0_out[5151];
     layer1_out[3543] <= ~layer0_out[8118];
     layer1_out[3544] <= ~(layer0_out[10278] | layer0_out[10279]);
     layer1_out[3545] <= layer0_out[8684] | layer0_out[8685];
     layer1_out[3546] <= layer0_out[7332] & ~layer0_out[7331];
     layer1_out[3547] <= ~(layer0_out[5814] | layer0_out[5815]);
     layer1_out[3548] <= layer0_out[3770];
     layer1_out[3549] <= layer0_out[9441] & layer0_out[9442];
     layer1_out[3550] <= ~layer0_out[5637];
     layer1_out[3551] <= layer0_out[2912];
     layer1_out[3552] <= layer0_out[9636] & layer0_out[9637];
     layer1_out[3553] <= layer0_out[8206] & ~layer0_out[8207];
     layer1_out[3554] <= layer0_out[2935] & ~layer0_out[2936];
     layer1_out[3555] <= ~layer0_out[4263] | layer0_out[4264];
     layer1_out[3556] <= layer0_out[9054] & ~layer0_out[9055];
     layer1_out[3557] <= ~layer0_out[10126];
     layer1_out[3558] <= ~(layer0_out[271] | layer0_out[272]);
     layer1_out[3559] <= ~(layer0_out[6501] | layer0_out[6502]);
     layer1_out[3560] <= layer0_out[4411] & ~layer0_out[4410];
     layer1_out[3561] <= ~layer0_out[10517];
     layer1_out[3562] <= layer0_out[8296] | layer0_out[8297];
     layer1_out[3563] <= ~(layer0_out[4896] & layer0_out[4897]);
     layer1_out[3564] <= ~layer0_out[4202] | layer0_out[4201];
     layer1_out[3565] <= 1'b1;
     layer1_out[3566] <= layer0_out[6752] & ~layer0_out[6753];
     layer1_out[3567] <= ~(layer0_out[7295] | layer0_out[7296]);
     layer1_out[3568] <= layer0_out[5745];
     layer1_out[3569] <= layer0_out[5147];
     layer1_out[3570] <= ~(layer0_out[4451] | layer0_out[4452]);
     layer1_out[3571] <= ~(layer0_out[6061] | layer0_out[6062]);
     layer1_out[3572] <= layer0_out[534];
     layer1_out[3573] <= layer0_out[10757];
     layer1_out[3574] <= ~layer0_out[11528] | layer0_out[11529];
     layer1_out[3575] <= ~layer0_out[29];
     layer1_out[3576] <= ~layer0_out[2656] | layer0_out[2655];
     layer1_out[3577] <= layer0_out[6754] & layer0_out[6755];
     layer1_out[3578] <= ~(layer0_out[2087] & layer0_out[2088]);
     layer1_out[3579] <= layer0_out[1525];
     layer1_out[3580] <= layer0_out[7057] | layer0_out[7058];
     layer1_out[3581] <= ~layer0_out[5580];
     layer1_out[3582] <= layer0_out[7421] | layer0_out[7422];
     layer1_out[3583] <= layer0_out[2663] ^ layer0_out[2664];
     layer1_out[3584] <= layer0_out[4442] & ~layer0_out[4443];
     layer1_out[3585] <= layer0_out[10848] & ~layer0_out[10849];
     layer1_out[3586] <= layer0_out[8989] & ~layer0_out[8990];
     layer1_out[3587] <= layer0_out[8627] & ~layer0_out[8626];
     layer1_out[3588] <= layer0_out[1166];
     layer1_out[3589] <= ~(layer0_out[9997] | layer0_out[9998]);
     layer1_out[3590] <= ~layer0_out[9132] | layer0_out[9133];
     layer1_out[3591] <= layer0_out[8519] | layer0_out[8520];
     layer1_out[3592] <= ~layer0_out[3891] | layer0_out[3892];
     layer1_out[3593] <= ~(layer0_out[3480] | layer0_out[3481]);
     layer1_out[3594] <= layer0_out[1397] ^ layer0_out[1398];
     layer1_out[3595] <= layer0_out[5318] ^ layer0_out[5319];
     layer1_out[3596] <= layer0_out[4956] | layer0_out[4957];
     layer1_out[3597] <= ~layer0_out[4950];
     layer1_out[3598] <= ~(layer0_out[8858] ^ layer0_out[8859]);
     layer1_out[3599] <= layer0_out[4623];
     layer1_out[3600] <= ~(layer0_out[603] | layer0_out[604]);
     layer1_out[3601] <= layer0_out[693] & layer0_out[694];
     layer1_out[3602] <= ~(layer0_out[7865] | layer0_out[7866]);
     layer1_out[3603] <= ~layer0_out[10718] | layer0_out[10717];
     layer1_out[3604] <= ~(layer0_out[2147] ^ layer0_out[2148]);
     layer1_out[3605] <= layer0_out[2098];
     layer1_out[3606] <= layer0_out[9079] & layer0_out[9080];
     layer1_out[3607] <= layer0_out[8183];
     layer1_out[3608] <= layer0_out[1123] & ~layer0_out[1122];
     layer1_out[3609] <= layer0_out[7082] & ~layer0_out[7083];
     layer1_out[3610] <= layer0_out[10217];
     layer1_out[3611] <= layer0_out[7752] & ~layer0_out[7753];
     layer1_out[3612] <= ~(layer0_out[4249] & layer0_out[4250]);
     layer1_out[3613] <= ~layer0_out[4404];
     layer1_out[3614] <= layer0_out[2753] & ~layer0_out[2754];
     layer1_out[3615] <= layer0_out[2790];
     layer1_out[3616] <= ~layer0_out[8068];
     layer1_out[3617] <= 1'b0;
     layer1_out[3618] <= layer0_out[6973] & ~layer0_out[6972];
     layer1_out[3619] <= layer0_out[11351] & ~layer0_out[11352];
     layer1_out[3620] <= ~(layer0_out[2928] & layer0_out[2929]);
     layer1_out[3621] <= ~layer0_out[8673] | layer0_out[8672];
     layer1_out[3622] <= layer0_out[10943];
     layer1_out[3623] <= layer0_out[298];
     layer1_out[3624] <= layer0_out[5914];
     layer1_out[3625] <= ~(layer0_out[4478] | layer0_out[4479]);
     layer1_out[3626] <= ~layer0_out[3940];
     layer1_out[3627] <= ~layer0_out[2179];
     layer1_out[3628] <= layer0_out[3842] & ~layer0_out[3843];
     layer1_out[3629] <= 1'b0;
     layer1_out[3630] <= ~layer0_out[2759];
     layer1_out[3631] <= layer0_out[4883] & ~layer0_out[4884];
     layer1_out[3632] <= layer0_out[399];
     layer1_out[3633] <= ~(layer0_out[4556] | layer0_out[4557]);
     layer1_out[3634] <= ~layer0_out[1044];
     layer1_out[3635] <= layer0_out[3399] | layer0_out[3400];
     layer1_out[3636] <= layer0_out[3359] & ~layer0_out[3360];
     layer1_out[3637] <= ~layer0_out[7051] | layer0_out[7050];
     layer1_out[3638] <= ~layer0_out[10429];
     layer1_out[3639] <= ~layer0_out[11170];
     layer1_out[3640] <= ~layer0_out[5826] | layer0_out[5827];
     layer1_out[3641] <= 1'b1;
     layer1_out[3642] <= ~layer0_out[4040];
     layer1_out[3643] <= layer0_out[4327] & ~layer0_out[4328];
     layer1_out[3644] <= ~layer0_out[8689] | layer0_out[8690];
     layer1_out[3645] <= ~layer0_out[5775] | layer0_out[5776];
     layer1_out[3646] <= ~(layer0_out[4033] ^ layer0_out[4034]);
     layer1_out[3647] <= ~layer0_out[7651] | layer0_out[7650];
     layer1_out[3648] <= ~layer0_out[8910];
     layer1_out[3649] <= ~layer0_out[1328] | layer0_out[1329];
     layer1_out[3650] <= layer0_out[6037] & layer0_out[6038];
     layer1_out[3651] <= ~layer0_out[8275];
     layer1_out[3652] <= ~(layer0_out[9384] ^ layer0_out[9385]);
     layer1_out[3653] <= layer0_out[1929];
     layer1_out[3654] <= layer0_out[4614] | layer0_out[4615];
     layer1_out[3655] <= layer0_out[2523] & ~layer0_out[2524];
     layer1_out[3656] <= ~layer0_out[10873] | layer0_out[10872];
     layer1_out[3657] <= layer0_out[11033];
     layer1_out[3658] <= layer0_out[7439] | layer0_out[7440];
     layer1_out[3659] <= layer0_out[8358];
     layer1_out[3660] <= layer0_out[8400] | layer0_out[8401];
     layer1_out[3661] <= ~layer0_out[4006] | layer0_out[4007];
     layer1_out[3662] <= layer0_out[10646] ^ layer0_out[10647];
     layer1_out[3663] <= layer0_out[2678] & layer0_out[2679];
     layer1_out[3664] <= layer0_out[368] & ~layer0_out[367];
     layer1_out[3665] <= ~layer0_out[9885];
     layer1_out[3666] <= ~layer0_out[10179] | layer0_out[10178];
     layer1_out[3667] <= layer0_out[2355];
     layer1_out[3668] <= layer0_out[3241] & ~layer0_out[3240];
     layer1_out[3669] <= layer0_out[11601];
     layer1_out[3670] <= ~(layer0_out[4557] ^ layer0_out[4558]);
     layer1_out[3671] <= layer0_out[11163] & layer0_out[11164];
     layer1_out[3672] <= layer0_out[1234] & ~layer0_out[1233];
     layer1_out[3673] <= ~(layer0_out[7829] | layer0_out[7830]);
     layer1_out[3674] <= layer0_out[11172] ^ layer0_out[11173];
     layer1_out[3675] <= ~layer0_out[1692];
     layer1_out[3676] <= ~(layer0_out[9244] ^ layer0_out[9245]);
     layer1_out[3677] <= ~(layer0_out[5173] & layer0_out[5174]);
     layer1_out[3678] <= layer0_out[3751];
     layer1_out[3679] <= layer0_out[1430] & ~layer0_out[1431];
     layer1_out[3680] <= ~layer0_out[3627];
     layer1_out[3681] <= ~(layer0_out[9187] & layer0_out[9188]);
     layer1_out[3682] <= ~layer0_out[9782];
     layer1_out[3683] <= ~layer0_out[8564];
     layer1_out[3684] <= layer0_out[729] & ~layer0_out[728];
     layer1_out[3685] <= ~layer0_out[11878] | layer0_out[11877];
     layer1_out[3686] <= ~layer0_out[11149] | layer0_out[11148];
     layer1_out[3687] <= ~(layer0_out[3005] & layer0_out[3006]);
     layer1_out[3688] <= layer0_out[8308];
     layer1_out[3689] <= ~(layer0_out[9819] & layer0_out[9820]);
     layer1_out[3690] <= layer0_out[4938];
     layer1_out[3691] <= ~layer0_out[9848];
     layer1_out[3692] <= 1'b0;
     layer1_out[3693] <= ~layer0_out[9760] | layer0_out[9759];
     layer1_out[3694] <= layer0_out[3211];
     layer1_out[3695] <= layer0_out[9289] | layer0_out[9290];
     layer1_out[3696] <= layer0_out[558] & layer0_out[559];
     layer1_out[3697] <= layer0_out[6128] & ~layer0_out[6127];
     layer1_out[3698] <= ~(layer0_out[10552] & layer0_out[10553]);
     layer1_out[3699] <= ~layer0_out[4654] | layer0_out[4655];
     layer1_out[3700] <= layer0_out[2873] ^ layer0_out[2874];
     layer1_out[3701] <= layer0_out[655];
     layer1_out[3702] <= ~layer0_out[8621];
     layer1_out[3703] <= 1'b0;
     layer1_out[3704] <= ~layer0_out[6665] | layer0_out[6664];
     layer1_out[3705] <= ~(layer0_out[4869] & layer0_out[4870]);
     layer1_out[3706] <= layer0_out[9162];
     layer1_out[3707] <= ~(layer0_out[4376] ^ layer0_out[4377]);
     layer1_out[3708] <= layer0_out[5568] ^ layer0_out[5569];
     layer1_out[3709] <= layer0_out[938];
     layer1_out[3710] <= ~layer0_out[967];
     layer1_out[3711] <= ~(layer0_out[6242] & layer0_out[6243]);
     layer1_out[3712] <= ~(layer0_out[11072] | layer0_out[11073]);
     layer1_out[3713] <= layer0_out[7125] & ~layer0_out[7124];
     layer1_out[3714] <= ~layer0_out[4260];
     layer1_out[3715] <= layer0_out[3087] ^ layer0_out[3088];
     layer1_out[3716] <= ~(layer0_out[10965] | layer0_out[10966]);
     layer1_out[3717] <= ~(layer0_out[9031] | layer0_out[9032]);
     layer1_out[3718] <= layer0_out[763];
     layer1_out[3719] <= ~(layer0_out[2439] | layer0_out[2440]);
     layer1_out[3720] <= ~layer0_out[2688];
     layer1_out[3721] <= ~layer0_out[2472];
     layer1_out[3722] <= layer0_out[11673] ^ layer0_out[11674];
     layer1_out[3723] <= layer0_out[1387] | layer0_out[1388];
     layer1_out[3724] <= layer0_out[1428] | layer0_out[1429];
     layer1_out[3725] <= layer0_out[7625] & ~layer0_out[7626];
     layer1_out[3726] <= layer0_out[2927];
     layer1_out[3727] <= layer0_out[8310] & layer0_out[8311];
     layer1_out[3728] <= ~layer0_out[4839];
     layer1_out[3729] <= ~layer0_out[10922] | layer0_out[10923];
     layer1_out[3730] <= layer0_out[160] & ~layer0_out[159];
     layer1_out[3731] <= layer0_out[10096];
     layer1_out[3732] <= ~(layer0_out[7460] & layer0_out[7461]);
     layer1_out[3733] <= ~layer0_out[1155] | layer0_out[1156];
     layer1_out[3734] <= layer0_out[1821] & layer0_out[1822];
     layer1_out[3735] <= ~layer0_out[11709] | layer0_out[11708];
     layer1_out[3736] <= 1'b0;
     layer1_out[3737] <= ~layer0_out[1605] | layer0_out[1606];
     layer1_out[3738] <= layer0_out[11980] & layer0_out[11981];
     layer1_out[3739] <= layer0_out[5773];
     layer1_out[3740] <= ~layer0_out[7146] | layer0_out[7145];
     layer1_out[3741] <= 1'b1;
     layer1_out[3742] <= layer0_out[9149] ^ layer0_out[9150];
     layer1_out[3743] <= layer0_out[11408] & ~layer0_out[11407];
     layer1_out[3744] <= layer0_out[7964] & ~layer0_out[7963];
     layer1_out[3745] <= ~(layer0_out[4732] ^ layer0_out[4733]);
     layer1_out[3746] <= layer0_out[2800] & ~layer0_out[2799];
     layer1_out[3747] <= layer0_out[2023] & ~layer0_out[2022];
     layer1_out[3748] <= ~layer0_out[9767] | layer0_out[9768];
     layer1_out[3749] <= layer0_out[3375];
     layer1_out[3750] <= ~(layer0_out[51] ^ layer0_out[52]);
     layer1_out[3751] <= layer0_out[11425];
     layer1_out[3752] <= layer0_out[7618] & layer0_out[7619];
     layer1_out[3753] <= layer0_out[10406] & ~layer0_out[10405];
     layer1_out[3754] <= layer0_out[4477];
     layer1_out[3755] <= layer0_out[10893] & ~layer0_out[10892];
     layer1_out[3756] <= layer0_out[8587] | layer0_out[8588];
     layer1_out[3757] <= layer0_out[3989];
     layer1_out[3758] <= layer0_out[5224] & ~layer0_out[5225];
     layer1_out[3759] <= layer0_out[1467];
     layer1_out[3760] <= layer0_out[5393];
     layer1_out[3761] <= ~(layer0_out[7299] | layer0_out[7300]);
     layer1_out[3762] <= ~layer0_out[9930];
     layer1_out[3763] <= ~layer0_out[5607];
     layer1_out[3764] <= layer0_out[5121] & layer0_out[5122];
     layer1_out[3765] <= layer0_out[8754];
     layer1_out[3766] <= layer0_out[11044] & ~layer0_out[11043];
     layer1_out[3767] <= layer0_out[360] & layer0_out[361];
     layer1_out[3768] <= layer0_out[3927] & layer0_out[3928];
     layer1_out[3769] <= layer0_out[4924] & layer0_out[4925];
     layer1_out[3770] <= layer0_out[3429] & ~layer0_out[3428];
     layer1_out[3771] <= ~layer0_out[11713] | layer0_out[11712];
     layer1_out[3772] <= ~(layer0_out[7218] ^ layer0_out[7219]);
     layer1_out[3773] <= ~layer0_out[9710];
     layer1_out[3774] <= ~layer0_out[3221];
     layer1_out[3775] <= ~layer0_out[5904];
     layer1_out[3776] <= ~layer0_out[11952];
     layer1_out[3777] <= 1'b0;
     layer1_out[3778] <= layer0_out[5402] | layer0_out[5403];
     layer1_out[3779] <= ~(layer0_out[7177] ^ layer0_out[7178]);
     layer1_out[3780] <= layer0_out[2195];
     layer1_out[3781] <= layer0_out[964];
     layer1_out[3782] <= layer0_out[2138] | layer0_out[2139];
     layer1_out[3783] <= layer0_out[4657];
     layer1_out[3784] <= ~(layer0_out[5665] & layer0_out[5666]);
     layer1_out[3785] <= ~layer0_out[6756];
     layer1_out[3786] <= layer0_out[2097] & ~layer0_out[2096];
     layer1_out[3787] <= layer0_out[9805] & ~layer0_out[9806];
     layer1_out[3788] <= layer0_out[8775] & layer0_out[8776];
     layer1_out[3789] <= ~(layer0_out[6122] ^ layer0_out[6123]);
     layer1_out[3790] <= 1'b0;
     layer1_out[3791] <= ~(layer0_out[1338] ^ layer0_out[1339]);
     layer1_out[3792] <= 1'b1;
     layer1_out[3793] <= layer0_out[4904] ^ layer0_out[4905];
     layer1_out[3794] <= ~(layer0_out[4940] ^ layer0_out[4941]);
     layer1_out[3795] <= layer0_out[10648];
     layer1_out[3796] <= layer0_out[4582];
     layer1_out[3797] <= ~layer0_out[7590];
     layer1_out[3798] <= ~layer0_out[10605];
     layer1_out[3799] <= layer0_out[6276] & ~layer0_out[6277];
     layer1_out[3800] <= ~layer0_out[5883];
     layer1_out[3801] <= layer0_out[2469] & layer0_out[2470];
     layer1_out[3802] <= layer0_out[10691];
     layer1_out[3803] <= ~layer0_out[11864];
     layer1_out[3804] <= ~layer0_out[11942] | layer0_out[11943];
     layer1_out[3805] <= ~layer0_out[8541];
     layer1_out[3806] <= ~layer0_out[1797] | layer0_out[1796];
     layer1_out[3807] <= ~layer0_out[7453];
     layer1_out[3808] <= ~layer0_out[9426] | layer0_out[9427];
     layer1_out[3809] <= layer0_out[7618];
     layer1_out[3810] <= ~layer0_out[3933] | layer0_out[3934];
     layer1_out[3811] <= ~(layer0_out[2195] & layer0_out[2196]);
     layer1_out[3812] <= ~layer0_out[7430];
     layer1_out[3813] <= layer0_out[5369] ^ layer0_out[5370];
     layer1_out[3814] <= layer0_out[3248] & ~layer0_out[3247];
     layer1_out[3815] <= ~layer0_out[3811] | layer0_out[3812];
     layer1_out[3816] <= layer0_out[3278] & ~layer0_out[3277];
     layer1_out[3817] <= ~(layer0_out[11927] & layer0_out[11928]);
     layer1_out[3818] <= ~layer0_out[8042] | layer0_out[8041];
     layer1_out[3819] <= layer0_out[9109];
     layer1_out[3820] <= layer0_out[9316] | layer0_out[9317];
     layer1_out[3821] <= ~layer0_out[5575];
     layer1_out[3822] <= layer0_out[11403] ^ layer0_out[11404];
     layer1_out[3823] <= ~layer0_out[1265] | layer0_out[1266];
     layer1_out[3824] <= ~layer0_out[4589];
     layer1_out[3825] <= layer0_out[2499];
     layer1_out[3826] <= ~(layer0_out[6802] | layer0_out[6803]);
     layer1_out[3827] <= ~(layer0_out[10455] & layer0_out[10456]);
     layer1_out[3828] <= ~layer0_out[6940] | layer0_out[6939];
     layer1_out[3829] <= layer0_out[89] & layer0_out[90];
     layer1_out[3830] <= layer0_out[7751] | layer0_out[7752];
     layer1_out[3831] <= ~(layer0_out[11084] | layer0_out[11085]);
     layer1_out[3832] <= ~layer0_out[9007];
     layer1_out[3833] <= 1'b1;
     layer1_out[3834] <= layer0_out[7329] ^ layer0_out[7330];
     layer1_out[3835] <= layer0_out[3542] & ~layer0_out[3543];
     layer1_out[3836] <= ~(layer0_out[3596] | layer0_out[3597]);
     layer1_out[3837] <= layer0_out[9954] & ~layer0_out[9953];
     layer1_out[3838] <= layer0_out[61];
     layer1_out[3839] <= 1'b0;
     layer1_out[3840] <= layer0_out[7956];
     layer1_out[3841] <= layer0_out[5669];
     layer1_out[3842] <= ~(layer0_out[11213] & layer0_out[11214]);
     layer1_out[3843] <= ~layer0_out[6553] | layer0_out[6552];
     layer1_out[3844] <= ~layer0_out[520] | layer0_out[521];
     layer1_out[3845] <= ~(layer0_out[11618] & layer0_out[11619]);
     layer1_out[3846] <= ~layer0_out[10713] | layer0_out[10712];
     layer1_out[3847] <= ~(layer0_out[11320] ^ layer0_out[11321]);
     layer1_out[3848] <= layer0_out[8723] ^ layer0_out[8724];
     layer1_out[3849] <= layer0_out[3695] & layer0_out[3696];
     layer1_out[3850] <= ~layer0_out[5423];
     layer1_out[3851] <= layer0_out[2180] & layer0_out[2181];
     layer1_out[3852] <= ~layer0_out[8989];
     layer1_out[3853] <= layer0_out[8190] ^ layer0_out[8191];
     layer1_out[3854] <= layer0_out[3013] & layer0_out[3014];
     layer1_out[3855] <= ~layer0_out[6493] | layer0_out[6494];
     layer1_out[3856] <= layer0_out[3140];
     layer1_out[3857] <= layer0_out[4321] & layer0_out[4322];
     layer1_out[3858] <= layer0_out[414] & layer0_out[415];
     layer1_out[3859] <= layer0_out[9479] ^ layer0_out[9480];
     layer1_out[3860] <= ~(layer0_out[2676] & layer0_out[2677]);
     layer1_out[3861] <= ~(layer0_out[11539] & layer0_out[11540]);
     layer1_out[3862] <= ~layer0_out[1307];
     layer1_out[3863] <= ~(layer0_out[5729] ^ layer0_out[5730]);
     layer1_out[3864] <= layer0_out[6158];
     layer1_out[3865] <= 1'b0;
     layer1_out[3866] <= layer0_out[5867] & ~layer0_out[5868];
     layer1_out[3867] <= layer0_out[3774];
     layer1_out[3868] <= layer0_out[5113];
     layer1_out[3869] <= layer0_out[11419];
     layer1_out[3870] <= layer0_out[1812] & ~layer0_out[1811];
     layer1_out[3871] <= ~layer0_out[2093] | layer0_out[2092];
     layer1_out[3872] <= layer0_out[8499];
     layer1_out[3873] <= ~layer0_out[3925] | layer0_out[3926];
     layer1_out[3874] <= layer0_out[6188] & layer0_out[6189];
     layer1_out[3875] <= ~layer0_out[2976];
     layer1_out[3876] <= ~layer0_out[6175] | layer0_out[6174];
     layer1_out[3877] <= ~(layer0_out[2440] & layer0_out[2441]);
     layer1_out[3878] <= layer0_out[3473];
     layer1_out[3879] <= ~layer0_out[11775];
     layer1_out[3880] <= ~layer0_out[5128];
     layer1_out[3881] <= layer0_out[5951] & ~layer0_out[5950];
     layer1_out[3882] <= ~layer0_out[11084];
     layer1_out[3883] <= ~(layer0_out[7359] ^ layer0_out[7360]);
     layer1_out[3884] <= layer0_out[1359] & layer0_out[1360];
     layer1_out[3885] <= ~layer0_out[695];
     layer1_out[3886] <= layer0_out[536];
     layer1_out[3887] <= ~layer0_out[35] | layer0_out[36];
     layer1_out[3888] <= layer0_out[5038] & ~layer0_out[5037];
     layer1_out[3889] <= 1'b1;
     layer1_out[3890] <= 1'b0;
     layer1_out[3891] <= layer0_out[9663];
     layer1_out[3892] <= 1'b0;
     layer1_out[3893] <= layer0_out[4738] | layer0_out[4739];
     layer1_out[3894] <= layer0_out[11732];
     layer1_out[3895] <= ~(layer0_out[11101] ^ layer0_out[11102]);
     layer1_out[3896] <= 1'b0;
     layer1_out[3897] <= ~(layer0_out[5759] & layer0_out[5760]);
     layer1_out[3898] <= ~layer0_out[3269] | layer0_out[3268];
     layer1_out[3899] <= layer0_out[9059];
     layer1_out[3900] <= layer0_out[10649] & ~layer0_out[10650];
     layer1_out[3901] <= ~layer0_out[10433] | layer0_out[10432];
     layer1_out[3902] <= ~layer0_out[2365];
     layer1_out[3903] <= ~layer0_out[1838] | layer0_out[1839];
     layer1_out[3904] <= layer0_out[11184] & ~layer0_out[11183];
     layer1_out[3905] <= layer0_out[6653];
     layer1_out[3906] <= ~layer0_out[10938];
     layer1_out[3907] <= layer0_out[6530] ^ layer0_out[6531];
     layer1_out[3908] <= layer0_out[8141] & ~layer0_out[8140];
     layer1_out[3909] <= 1'b0;
     layer1_out[3910] <= ~layer0_out[1060] | layer0_out[1061];
     layer1_out[3911] <= layer0_out[2104];
     layer1_out[3912] <= layer0_out[9012] ^ layer0_out[9013];
     layer1_out[3913] <= ~layer0_out[8481] | layer0_out[8480];
     layer1_out[3914] <= layer0_out[6480];
     layer1_out[3915] <= layer0_out[976] & ~layer0_out[975];
     layer1_out[3916] <= ~layer0_out[5576];
     layer1_out[3917] <= ~layer0_out[4974];
     layer1_out[3918] <= layer0_out[9260];
     layer1_out[3919] <= ~(layer0_out[6626] & layer0_out[6627]);
     layer1_out[3920] <= layer0_out[240];
     layer1_out[3921] <= ~layer0_out[395] | layer0_out[394];
     layer1_out[3922] <= layer0_out[10464] & ~layer0_out[10463];
     layer1_out[3923] <= layer0_out[8353] | layer0_out[8354];
     layer1_out[3924] <= layer0_out[5583] & layer0_out[5584];
     layer1_out[3925] <= layer0_out[1493] | layer0_out[1494];
     layer1_out[3926] <= layer0_out[2091] & layer0_out[2092];
     layer1_out[3927] <= ~layer0_out[11204] | layer0_out[11203];
     layer1_out[3928] <= layer0_out[11792] & layer0_out[11793];
     layer1_out[3929] <= layer0_out[6045] & layer0_out[6046];
     layer1_out[3930] <= layer0_out[7754];
     layer1_out[3931] <= ~layer0_out[5586] | layer0_out[5587];
     layer1_out[3932] <= ~layer0_out[2496] | layer0_out[2497];
     layer1_out[3933] <= layer0_out[11847];
     layer1_out[3934] <= layer0_out[876] & ~layer0_out[877];
     layer1_out[3935] <= layer0_out[2368] & layer0_out[2369];
     layer1_out[3936] <= layer0_out[948];
     layer1_out[3937] <= ~(layer0_out[9651] ^ layer0_out[9652]);
     layer1_out[3938] <= layer0_out[10410];
     layer1_out[3939] <= ~layer0_out[4413];
     layer1_out[3940] <= layer0_out[6714] & layer0_out[6715];
     layer1_out[3941] <= ~(layer0_out[8071] | layer0_out[8072]);
     layer1_out[3942] <= ~(layer0_out[5298] | layer0_out[5299]);
     layer1_out[3943] <= layer0_out[6788] & layer0_out[6789];
     layer1_out[3944] <= layer0_out[8471] | layer0_out[8472];
     layer1_out[3945] <= ~layer0_out[5778];
     layer1_out[3946] <= layer0_out[5079];
     layer1_out[3947] <= ~layer0_out[5865];
     layer1_out[3948] <= ~(layer0_out[10915] ^ layer0_out[10916]);
     layer1_out[3949] <= layer0_out[6927];
     layer1_out[3950] <= ~(layer0_out[4020] & layer0_out[4021]);
     layer1_out[3951] <= 1'b0;
     layer1_out[3952] <= ~layer0_out[534];
     layer1_out[3953] <= ~(layer0_out[5758] & layer0_out[5759]);
     layer1_out[3954] <= 1'b0;
     layer1_out[3955] <= 1'b0;
     layer1_out[3956] <= layer0_out[5397] & ~layer0_out[5398];
     layer1_out[3957] <= ~(layer0_out[275] ^ layer0_out[276]);
     layer1_out[3958] <= ~layer0_out[63];
     layer1_out[3959] <= ~layer0_out[11955];
     layer1_out[3960] <= ~(layer0_out[5257] | layer0_out[5258]);
     layer1_out[3961] <= layer0_out[9305];
     layer1_out[3962] <= ~layer0_out[3667];
     layer1_out[3963] <= layer0_out[9108] & ~layer0_out[9109];
     layer1_out[3964] <= ~(layer0_out[10642] | layer0_out[10643]);
     layer1_out[3965] <= layer0_out[802];
     layer1_out[3966] <= layer0_out[1107];
     layer1_out[3967] <= layer0_out[8121];
     layer1_out[3968] <= ~layer0_out[6196];
     layer1_out[3969] <= layer0_out[514] ^ layer0_out[515];
     layer1_out[3970] <= ~(layer0_out[5662] | layer0_out[5663]);
     layer1_out[3971] <= ~(layer0_out[2490] ^ layer0_out[2491]);
     layer1_out[3972] <= ~layer0_out[10872] | layer0_out[10871];
     layer1_out[3973] <= layer0_out[3816];
     layer1_out[3974] <= layer0_out[6865];
     layer1_out[3975] <= ~(layer0_out[1237] & layer0_out[1238]);
     layer1_out[3976] <= layer0_out[10739];
     layer1_out[3977] <= layer0_out[3393];
     layer1_out[3978] <= ~layer0_out[5163] | layer0_out[5162];
     layer1_out[3979] <= ~(layer0_out[5241] & layer0_out[5242]);
     layer1_out[3980] <= ~layer0_out[10531];
     layer1_out[3981] <= layer0_out[658] & layer0_out[659];
     layer1_out[3982] <= ~(layer0_out[7333] | layer0_out[7334]);
     layer1_out[3983] <= ~layer0_out[6123];
     layer1_out[3984] <= 1'b1;
     layer1_out[3985] <= ~layer0_out[7964];
     layer1_out[3986] <= ~layer0_out[2410];
     layer1_out[3987] <= 1'b0;
     layer1_out[3988] <= layer0_out[6613] & ~layer0_out[6614];
     layer1_out[3989] <= ~layer0_out[9587];
     layer1_out[3990] <= 1'b1;
     layer1_out[3991] <= layer0_out[9400] & layer0_out[9401];
     layer1_out[3992] <= layer0_out[6616] & ~layer0_out[6615];
     layer1_out[3993] <= layer0_out[4670];
     layer1_out[3994] <= ~layer0_out[8777];
     layer1_out[3995] <= ~layer0_out[4464];
     layer1_out[3996] <= layer0_out[567] ^ layer0_out[568];
     layer1_out[3997] <= ~layer0_out[10085];
     layer1_out[3998] <= layer0_out[11536] & layer0_out[11537];
     layer1_out[3999] <= ~layer0_out[1833] | layer0_out[1834];
     layer1_out[4000] <= layer0_out[3136] & layer0_out[3137];
     layer1_out[4001] <= layer0_out[6790] & layer0_out[6791];
     layer1_out[4002] <= layer0_out[1558] & ~layer0_out[1557];
     layer1_out[4003] <= ~(layer0_out[6781] & layer0_out[6782]);
     layer1_out[4004] <= layer0_out[4125];
     layer1_out[4005] <= layer0_out[6148];
     layer1_out[4006] <= layer0_out[9098] | layer0_out[9099];
     layer1_out[4007] <= ~layer0_out[689];
     layer1_out[4008] <= layer0_out[3792] & ~layer0_out[3791];
     layer1_out[4009] <= layer0_out[230] | layer0_out[231];
     layer1_out[4010] <= ~layer0_out[1155] | layer0_out[1154];
     layer1_out[4011] <= ~layer0_out[5226] | layer0_out[5225];
     layer1_out[4012] <= ~layer0_out[4996] | layer0_out[4997];
     layer1_out[4013] <= 1'b1;
     layer1_out[4014] <= ~layer0_out[8594];
     layer1_out[4015] <= ~layer0_out[4923];
     layer1_out[4016] <= layer0_out[11436];
     layer1_out[4017] <= layer0_out[2465] & ~layer0_out[2464];
     layer1_out[4018] <= layer0_out[6520];
     layer1_out[4019] <= ~layer0_out[11790] | layer0_out[11791];
     layer1_out[4020] <= ~(layer0_out[8965] | layer0_out[8966]);
     layer1_out[4021] <= 1'b0;
     layer1_out[4022] <= ~layer0_out[2339];
     layer1_out[4023] <= layer0_out[170];
     layer1_out[4024] <= ~layer0_out[6358] | layer0_out[6357];
     layer1_out[4025] <= ~layer0_out[235] | layer0_out[236];
     layer1_out[4026] <= ~layer0_out[7163];
     layer1_out[4027] <= layer0_out[3200] & ~layer0_out[3201];
     layer1_out[4028] <= ~layer0_out[5408];
     layer1_out[4029] <= layer0_out[3380];
     layer1_out[4030] <= layer0_out[2089];
     layer1_out[4031] <= 1'b1;
     layer1_out[4032] <= ~(layer0_out[356] | layer0_out[357]);
     layer1_out[4033] <= ~layer0_out[1570] | layer0_out[1569];
     layer1_out[4034] <= layer0_out[9433] & ~layer0_out[9432];
     layer1_out[4035] <= layer0_out[3071] | layer0_out[3072];
     layer1_out[4036] <= layer0_out[7550] | layer0_out[7551];
     layer1_out[4037] <= layer0_out[8228] & layer0_out[8229];
     layer1_out[4038] <= ~layer0_out[6205];
     layer1_out[4039] <= ~layer0_out[8648] | layer0_out[8647];
     layer1_out[4040] <= ~layer0_out[2031] | layer0_out[2030];
     layer1_out[4041] <= ~layer0_out[290];
     layer1_out[4042] <= layer0_out[1181] & layer0_out[1182];
     layer1_out[4043] <= layer0_out[1489];
     layer1_out[4044] <= ~layer0_out[758];
     layer1_out[4045] <= layer0_out[7738] | layer0_out[7739];
     layer1_out[4046] <= layer0_out[7410] & ~layer0_out[7409];
     layer1_out[4047] <= layer0_out[11700];
     layer1_out[4048] <= 1'b0;
     layer1_out[4049] <= ~layer0_out[4184] | layer0_out[4183];
     layer1_out[4050] <= layer0_out[6617] | layer0_out[6618];
     layer1_out[4051] <= ~layer0_out[5264] | layer0_out[5265];
     layer1_out[4052] <= ~layer0_out[1368];
     layer1_out[4053] <= layer0_out[977] ^ layer0_out[978];
     layer1_out[4054] <= layer0_out[646] & ~layer0_out[645];
     layer1_out[4055] <= ~(layer0_out[9850] | layer0_out[9851]);
     layer1_out[4056] <= layer0_out[7501];
     layer1_out[4057] <= layer0_out[2830] & ~layer0_out[2831];
     layer1_out[4058] <= ~layer0_out[11174];
     layer1_out[4059] <= ~layer0_out[11848];
     layer1_out[4060] <= ~layer0_out[7375];
     layer1_out[4061] <= ~layer0_out[8863] | layer0_out[8862];
     layer1_out[4062] <= ~(layer0_out[1762] & layer0_out[1763]);
     layer1_out[4063] <= layer0_out[865] & ~layer0_out[864];
     layer1_out[4064] <= layer0_out[6760] ^ layer0_out[6761];
     layer1_out[4065] <= ~layer0_out[4844];
     layer1_out[4066] <= layer0_out[2691] & ~layer0_out[2692];
     layer1_out[4067] <= layer0_out[11863] & layer0_out[11864];
     layer1_out[4068] <= layer0_out[10000];
     layer1_out[4069] <= layer0_out[6013];
     layer1_out[4070] <= ~layer0_out[2289];
     layer1_out[4071] <= layer0_out[7003];
     layer1_out[4072] <= ~(layer0_out[8848] | layer0_out[8849]);
     layer1_out[4073] <= layer0_out[5044];
     layer1_out[4074] <= ~(layer0_out[9541] | layer0_out[9542]);
     layer1_out[4075] <= 1'b1;
     layer1_out[4076] <= layer0_out[2456] & layer0_out[2457];
     layer1_out[4077] <= ~layer0_out[1405];
     layer1_out[4078] <= ~(layer0_out[1450] | layer0_out[1451]);
     layer1_out[4079] <= ~layer0_out[5188] | layer0_out[5189];
     layer1_out[4080] <= layer0_out[6082];
     layer1_out[4081] <= layer0_out[4831];
     layer1_out[4082] <= ~layer0_out[326] | layer0_out[327];
     layer1_out[4083] <= layer0_out[6464] & ~layer0_out[6463];
     layer1_out[4084] <= ~layer0_out[1691] | layer0_out[1690];
     layer1_out[4085] <= layer0_out[9513] & ~layer0_out[9512];
     layer1_out[4086] <= layer0_out[10856] ^ layer0_out[10857];
     layer1_out[4087] <= ~(layer0_out[4113] | layer0_out[4114]);
     layer1_out[4088] <= layer0_out[7851];
     layer1_out[4089] <= ~(layer0_out[5431] & layer0_out[5432]);
     layer1_out[4090] <= layer0_out[7711] & ~layer0_out[7710];
     layer1_out[4091] <= ~layer0_out[2634];
     layer1_out[4092] <= ~(layer0_out[7121] ^ layer0_out[7122]);
     layer1_out[4093] <= 1'b0;
     layer1_out[4094] <= ~(layer0_out[841] & layer0_out[842]);
     layer1_out[4095] <= ~layer0_out[10523];
     layer1_out[4096] <= ~layer0_out[10909] | layer0_out[10910];
     layer1_out[4097] <= ~layer0_out[7390];
     layer1_out[4098] <= layer0_out[11093] | layer0_out[11094];
     layer1_out[4099] <= layer0_out[3088];
     layer1_out[4100] <= ~layer0_out[9553] | layer0_out[9552];
     layer1_out[4101] <= ~(layer0_out[8987] | layer0_out[8988]);
     layer1_out[4102] <= layer0_out[8343];
     layer1_out[4103] <= 1'b1;
     layer1_out[4104] <= layer0_out[7263];
     layer1_out[4105] <= layer0_out[9240] ^ layer0_out[9241];
     layer1_out[4106] <= ~layer0_out[10004];
     layer1_out[4107] <= ~layer0_out[11057];
     layer1_out[4108] <= layer0_out[6820] & layer0_out[6821];
     layer1_out[4109] <= ~(layer0_out[10111] | layer0_out[10112]);
     layer1_out[4110] <= ~layer0_out[10344] | layer0_out[10343];
     layer1_out[4111] <= ~(layer0_out[706] & layer0_out[707]);
     layer1_out[4112] <= layer0_out[9038] | layer0_out[9039];
     layer1_out[4113] <= ~(layer0_out[8637] & layer0_out[8638]);
     layer1_out[4114] <= layer0_out[4962] & ~layer0_out[4961];
     layer1_out[4115] <= ~layer0_out[8854] | layer0_out[8853];
     layer1_out[4116] <= ~layer0_out[11544];
     layer1_out[4117] <= ~layer0_out[3979] | layer0_out[3978];
     layer1_out[4118] <= layer0_out[11269] ^ layer0_out[11270];
     layer1_out[4119] <= layer0_out[10219] & ~layer0_out[10220];
     layer1_out[4120] <= layer0_out[5888];
     layer1_out[4121] <= layer0_out[4801];
     layer1_out[4122] <= layer0_out[932];
     layer1_out[4123] <= 1'b0;
     layer1_out[4124] <= ~layer0_out[2755] | layer0_out[2754];
     layer1_out[4125] <= layer0_out[6954];
     layer1_out[4126] <= layer0_out[7114] | layer0_out[7115];
     layer1_out[4127] <= ~(layer0_out[6732] | layer0_out[6733]);
     layer1_out[4128] <= layer0_out[3143] & layer0_out[3144];
     layer1_out[4129] <= ~layer0_out[5309];
     layer1_out[4130] <= ~layer0_out[9434] | layer0_out[9433];
     layer1_out[4131] <= ~(layer0_out[4783] ^ layer0_out[4784]);
     layer1_out[4132] <= ~layer0_out[10007];
     layer1_out[4133] <= layer0_out[8904] & ~layer0_out[8903];
     layer1_out[4134] <= 1'b1;
     layer1_out[4135] <= ~layer0_out[5907] | layer0_out[5906];
     layer1_out[4136] <= layer0_out[7944];
     layer1_out[4137] <= ~(layer0_out[6486] ^ layer0_out[6487]);
     layer1_out[4138] <= layer0_out[9076] & ~layer0_out[9075];
     layer1_out[4139] <= ~(layer0_out[8688] & layer0_out[8689]);
     layer1_out[4140] <= ~(layer0_out[9610] ^ layer0_out[9611]);
     layer1_out[4141] <= ~layer0_out[4624] | layer0_out[4625];
     layer1_out[4142] <= ~(layer0_out[11865] | layer0_out[11866]);
     layer1_out[4143] <= ~layer0_out[6977];
     layer1_out[4144] <= layer0_out[4963] & layer0_out[4964];
     layer1_out[4145] <= layer0_out[8582] & ~layer0_out[8583];
     layer1_out[4146] <= ~layer0_out[9902] | layer0_out[9901];
     layer1_out[4147] <= layer0_out[6967] & layer0_out[6968];
     layer1_out[4148] <= ~layer0_out[6784] | layer0_out[6783];
     layer1_out[4149] <= 1'b1;
     layer1_out[4150] <= ~(layer0_out[1744] ^ layer0_out[1745]);
     layer1_out[4151] <= ~layer0_out[648] | layer0_out[649];
     layer1_out[4152] <= layer0_out[2615] | layer0_out[2616];
     layer1_out[4153] <= ~layer0_out[2354];
     layer1_out[4154] <= layer0_out[9284] & layer0_out[9285];
     layer1_out[4155] <= layer0_out[4487] | layer0_out[4488];
     layer1_out[4156] <= ~layer0_out[5718] | layer0_out[5717];
     layer1_out[4157] <= layer0_out[7391];
     layer1_out[4158] <= layer0_out[6360];
     layer1_out[4159] <= layer0_out[3894];
     layer1_out[4160] <= layer0_out[2767] ^ layer0_out[2768];
     layer1_out[4161] <= ~layer0_out[4014];
     layer1_out[4162] <= layer0_out[8994] & ~layer0_out[8993];
     layer1_out[4163] <= layer0_out[3207];
     layer1_out[4164] <= layer0_out[3417];
     layer1_out[4165] <= layer0_out[9046];
     layer1_out[4166] <= 1'b1;
     layer1_out[4167] <= ~(layer0_out[4242] ^ layer0_out[4243]);
     layer1_out[4168] <= layer0_out[5198] & layer0_out[5199];
     layer1_out[4169] <= layer0_out[6661];
     layer1_out[4170] <= ~layer0_out[1284] | layer0_out[1285];
     layer1_out[4171] <= 1'b0;
     layer1_out[4172] <= layer0_out[9313];
     layer1_out[4173] <= layer0_out[8618] | layer0_out[8619];
     layer1_out[4174] <= 1'b0;
     layer1_out[4175] <= layer0_out[6805] & ~layer0_out[6806];
     layer1_out[4176] <= ~layer0_out[3808];
     layer1_out[4177] <= layer0_out[10493];
     layer1_out[4178] <= ~layer0_out[5052] | layer0_out[5051];
     layer1_out[4179] <= layer0_out[10143];
     layer1_out[4180] <= ~layer0_out[6456];
     layer1_out[4181] <= ~(layer0_out[7937] ^ layer0_out[7938]);
     layer1_out[4182] <= layer0_out[528] & layer0_out[529];
     layer1_out[4183] <= layer0_out[10736];
     layer1_out[4184] <= layer0_out[5278];
     layer1_out[4185] <= layer0_out[1936] ^ layer0_out[1937];
     layer1_out[4186] <= ~layer0_out[2191] | layer0_out[2192];
     layer1_out[4187] <= ~layer0_out[5342];
     layer1_out[4188] <= layer0_out[5894] & layer0_out[5895];
     layer1_out[4189] <= ~(layer0_out[4782] ^ layer0_out[4783]);
     layer1_out[4190] <= ~layer0_out[3668] | layer0_out[3669];
     layer1_out[4191] <= ~(layer0_out[11730] | layer0_out[11731]);
     layer1_out[4192] <= layer0_out[9868] & layer0_out[9869];
     layer1_out[4193] <= ~layer0_out[8713] | layer0_out[8714];
     layer1_out[4194] <= layer0_out[260];
     layer1_out[4195] <= layer0_out[2958];
     layer1_out[4196] <= layer0_out[11051] & layer0_out[11052];
     layer1_out[4197] <= layer0_out[2719] & layer0_out[2720];
     layer1_out[4198] <= layer0_out[2012];
     layer1_out[4199] <= ~layer0_out[6143] | layer0_out[6144];
     layer1_out[4200] <= ~layer0_out[7228] | layer0_out[7227];
     layer1_out[4201] <= layer0_out[5698] ^ layer0_out[5699];
     layer1_out[4202] <= ~(layer0_out[1682] ^ layer0_out[1683]);
     layer1_out[4203] <= ~layer0_out[10125] | layer0_out[10124];
     layer1_out[4204] <= layer0_out[11416] & ~layer0_out[11417];
     layer1_out[4205] <= ~layer0_out[7289];
     layer1_out[4206] <= ~layer0_out[8056] | layer0_out[8055];
     layer1_out[4207] <= layer0_out[7122];
     layer1_out[4208] <= layer0_out[2222] & ~layer0_out[2223];
     layer1_out[4209] <= ~layer0_out[7644] | layer0_out[7645];
     layer1_out[4210] <= ~layer0_out[1468];
     layer1_out[4211] <= layer0_out[5569] | layer0_out[5570];
     layer1_out[4212] <= layer0_out[7458];
     layer1_out[4213] <= ~layer0_out[5678] | layer0_out[5679];
     layer1_out[4214] <= ~layer0_out[2864] | layer0_out[2863];
     layer1_out[4215] <= ~layer0_out[11639] | layer0_out[11640];
     layer1_out[4216] <= ~layer0_out[6485];
     layer1_out[4217] <= ~layer0_out[10408] | layer0_out[10407];
     layer1_out[4218] <= ~layer0_out[8261] | layer0_out[8260];
     layer1_out[4219] <= layer0_out[2665] & ~layer0_out[2664];
     layer1_out[4220] <= layer0_out[11963] | layer0_out[11964];
     layer1_out[4221] <= layer0_out[6010];
     layer1_out[4222] <= ~layer0_out[9849];
     layer1_out[4223] <= ~(layer0_out[11914] & layer0_out[11915]);
     layer1_out[4224] <= ~layer0_out[11130] | layer0_out[11131];
     layer1_out[4225] <= 1'b1;
     layer1_out[4226] <= layer0_out[9168];
     layer1_out[4227] <= layer0_out[11826];
     layer1_out[4228] <= layer0_out[1667] & layer0_out[1668];
     layer1_out[4229] <= layer0_out[9983] & ~layer0_out[9982];
     layer1_out[4230] <= layer0_out[6546] & ~layer0_out[6545];
     layer1_out[4231] <= layer0_out[3069];
     layer1_out[4232] <= 1'b0;
     layer1_out[4233] <= ~layer0_out[7335];
     layer1_out[4234] <= ~(layer0_out[1943] ^ layer0_out[1944]);
     layer1_out[4235] <= ~(layer0_out[457] & layer0_out[458]);
     layer1_out[4236] <= ~layer0_out[6056] | layer0_out[6055];
     layer1_out[4237] <= 1'b0;
     layer1_out[4238] <= layer0_out[7945];
     layer1_out[4239] <= ~(layer0_out[8906] ^ layer0_out[8907]);
     layer1_out[4240] <= ~layer0_out[8449];
     layer1_out[4241] <= layer0_out[6414];
     layer1_out[4242] <= layer0_out[182];
     layer1_out[4243] <= ~layer0_out[5823];
     layer1_out[4244] <= ~layer0_out[5140] | layer0_out[5141];
     layer1_out[4245] <= layer0_out[4485] & layer0_out[4486];
     layer1_out[4246] <= 1'b0;
     layer1_out[4247] <= layer0_out[6795] ^ layer0_out[6796];
     layer1_out[4248] <= ~(layer0_out[6744] ^ layer0_out[6745]);
     layer1_out[4249] <= layer0_out[396];
     layer1_out[4250] <= layer0_out[2545] & ~layer0_out[2546];
     layer1_out[4251] <= layer0_out[9074] & layer0_out[9075];
     layer1_out[4252] <= ~layer0_out[9919];
     layer1_out[4253] <= ~(layer0_out[782] ^ layer0_out[783]);
     layer1_out[4254] <= layer0_out[10540] & layer0_out[10541];
     layer1_out[4255] <= layer0_out[7575];
     layer1_out[4256] <= layer0_out[8450];
     layer1_out[4257] <= layer0_out[6403];
     layer1_out[4258] <= layer0_out[849] | layer0_out[850];
     layer1_out[4259] <= layer0_out[2402];
     layer1_out[4260] <= layer0_out[2982] ^ layer0_out[2983];
     layer1_out[4261] <= layer0_out[7285] & ~layer0_out[7284];
     layer1_out[4262] <= ~layer0_out[4139];
     layer1_out[4263] <= ~layer0_out[3136] | layer0_out[3135];
     layer1_out[4264] <= layer0_out[5287];
     layer1_out[4265] <= ~(layer0_out[4045] | layer0_out[4046]);
     layer1_out[4266] <= ~layer0_out[4332];
     layer1_out[4267] <= ~layer0_out[10815] | layer0_out[10814];
     layer1_out[4268] <= layer0_out[10219];
     layer1_out[4269] <= ~(layer0_out[9278] ^ layer0_out[9279]);
     layer1_out[4270] <= layer0_out[2561];
     layer1_out[4271] <= layer0_out[11201] ^ layer0_out[11202];
     layer1_out[4272] <= ~(layer0_out[1719] ^ layer0_out[1720]);
     layer1_out[4273] <= ~layer0_out[768] | layer0_out[767];
     layer1_out[4274] <= layer0_out[8993];
     layer1_out[4275] <= ~layer0_out[9836];
     layer1_out[4276] <= ~layer0_out[11510];
     layer1_out[4277] <= layer0_out[9374];
     layer1_out[4278] <= layer0_out[829];
     layer1_out[4279] <= layer0_out[3505] & ~layer0_out[3504];
     layer1_out[4280] <= ~(layer0_out[3094] | layer0_out[3095]);
     layer1_out[4281] <= 1'b0;
     layer1_out[4282] <= layer0_out[9204] & ~layer0_out[9203];
     layer1_out[4283] <= layer0_out[11438] & ~layer0_out[11439];
     layer1_out[4284] <= ~(layer0_out[9099] & layer0_out[9100]);
     layer1_out[4285] <= layer0_out[8044] | layer0_out[8045];
     layer1_out[4286] <= layer0_out[7300];
     layer1_out[4287] <= ~layer0_out[983];
     layer1_out[4288] <= layer0_out[5642];
     layer1_out[4289] <= ~(layer0_out[3078] & layer0_out[3079]);
     layer1_out[4290] <= layer0_out[1624];
     layer1_out[4291] <= ~layer0_out[8851];
     layer1_out[4292] <= layer0_out[9931] | layer0_out[9932];
     layer1_out[4293] <= ~layer0_out[3838] | layer0_out[3837];
     layer1_out[4294] <= ~layer0_out[3810];
     layer1_out[4295] <= ~(layer0_out[765] & layer0_out[766]);
     layer1_out[4296] <= ~layer0_out[6560];
     layer1_out[4297] <= layer0_out[6911];
     layer1_out[4298] <= 1'b1;
     layer1_out[4299] <= layer0_out[10273] & ~layer0_out[10274];
     layer1_out[4300] <= ~layer0_out[5386];
     layer1_out[4301] <= layer0_out[9941];
     layer1_out[4302] <= ~layer0_out[3665] | layer0_out[3666];
     layer1_out[4303] <= layer0_out[11468] | layer0_out[11469];
     layer1_out[4304] <= ~(layer0_out[11683] & layer0_out[11684]);
     layer1_out[4305] <= ~layer0_out[2767] | layer0_out[2766];
     layer1_out[4306] <= layer0_out[5928] & layer0_out[5929];
     layer1_out[4307] <= layer0_out[135] & ~layer0_out[134];
     layer1_out[4308] <= ~layer0_out[5385];
     layer1_out[4309] <= ~(layer0_out[6923] | layer0_out[6924]);
     layer1_out[4310] <= ~layer0_out[8496] | layer0_out[8497];
     layer1_out[4311] <= layer0_out[4090];
     layer1_out[4312] <= layer0_out[4008];
     layer1_out[4313] <= ~layer0_out[5512];
     layer1_out[4314] <= layer0_out[9035] & ~layer0_out[9034];
     layer1_out[4315] <= ~layer0_out[8126];
     layer1_out[4316] <= layer0_out[8408];
     layer1_out[4317] <= ~layer0_out[8247];
     layer1_out[4318] <= ~layer0_out[966];
     layer1_out[4319] <= ~(layer0_out[4734] | layer0_out[4735]);
     layer1_out[4320] <= ~(layer0_out[6958] ^ layer0_out[6959]);
     layer1_out[4321] <= ~layer0_out[2715] | layer0_out[2714];
     layer1_out[4322] <= ~layer0_out[10590];
     layer1_out[4323] <= ~layer0_out[11633] | layer0_out[11632];
     layer1_out[4324] <= layer0_out[9762] & ~layer0_out[9763];
     layer1_out[4325] <= ~(layer0_out[8635] & layer0_out[8636]);
     layer1_out[4326] <= ~(layer0_out[58] ^ layer0_out[59]);
     layer1_out[4327] <= layer0_out[1657];
     layer1_out[4328] <= 1'b1;
     layer1_out[4329] <= ~layer0_out[4368] | layer0_out[4367];
     layer1_out[4330] <= layer0_out[81];
     layer1_out[4331] <= ~layer0_out[715];
     layer1_out[4332] <= ~(layer0_out[2320] & layer0_out[2321]);
     layer1_out[4333] <= layer0_out[6240] & layer0_out[6241];
     layer1_out[4334] <= ~(layer0_out[9906] ^ layer0_out[9907]);
     layer1_out[4335] <= layer0_out[972] & ~layer0_out[971];
     layer1_out[4336] <= layer0_out[1754] & ~layer0_out[1753];
     layer1_out[4337] <= layer0_out[2769] & layer0_out[2770];
     layer1_out[4338] <= layer0_out[1981] & layer0_out[1982];
     layer1_out[4339] <= layer0_out[6012];
     layer1_out[4340] <= layer0_out[3537] & ~layer0_out[3538];
     layer1_out[4341] <= ~layer0_out[6895] | layer0_out[6894];
     layer1_out[4342] <= layer0_out[5962] & layer0_out[5963];
     layer1_out[4343] <= layer0_out[4567];
     layer1_out[4344] <= layer0_out[7566] & ~layer0_out[7565];
     layer1_out[4345] <= ~layer0_out[11345];
     layer1_out[4346] <= ~(layer0_out[591] | layer0_out[592]);
     layer1_out[4347] <= layer0_out[11055] & ~layer0_out[11056];
     layer1_out[4348] <= layer0_out[3680] & ~layer0_out[3679];
     layer1_out[4349] <= layer0_out[6278] & layer0_out[6279];
     layer1_out[4350] <= ~(layer0_out[2870] | layer0_out[2871]);
     layer1_out[4351] <= ~layer0_out[10084];
     layer1_out[4352] <= ~layer0_out[9817];
     layer1_out[4353] <= ~layer0_out[425];
     layer1_out[4354] <= ~(layer0_out[5927] & layer0_out[5928]);
     layer1_out[4355] <= ~(layer0_out[5266] & layer0_out[5267]);
     layer1_out[4356] <= layer0_out[7512] & ~layer0_out[7513];
     layer1_out[4357] <= layer0_out[9801] & ~layer0_out[9800];
     layer1_out[4358] <= layer0_out[6886];
     layer1_out[4359] <= layer0_out[3921];
     layer1_out[4360] <= 1'b1;
     layer1_out[4361] <= ~layer0_out[5132] | layer0_out[5133];
     layer1_out[4362] <= layer0_out[5587];
     layer1_out[4363] <= layer0_out[6779] | layer0_out[6780];
     layer1_out[4364] <= ~(layer0_out[10698] | layer0_out[10699]);
     layer1_out[4365] <= layer0_out[9877] ^ layer0_out[9878];
     layer1_out[4366] <= ~layer0_out[3977];
     layer1_out[4367] <= layer0_out[10578] ^ layer0_out[10579];
     layer1_out[4368] <= layer0_out[7775];
     layer1_out[4369] <= layer0_out[2974] & ~layer0_out[2975];
     layer1_out[4370] <= ~layer0_out[9498] | layer0_out[9499];
     layer1_out[4371] <= ~(layer0_out[7799] ^ layer0_out[7800]);
     layer1_out[4372] <= layer0_out[8782] & layer0_out[8783];
     layer1_out[4373] <= ~layer0_out[4958];
     layer1_out[4374] <= layer0_out[2245] | layer0_out[2246];
     layer1_out[4375] <= layer0_out[10314];
     layer1_out[4376] <= ~(layer0_out[6320] | layer0_out[6321]);
     layer1_out[4377] <= ~(layer0_out[10930] & layer0_out[10931]);
     layer1_out[4378] <= layer0_out[4339] & ~layer0_out[4340];
     layer1_out[4379] <= layer0_out[11810] & ~layer0_out[11811];
     layer1_out[4380] <= layer0_out[3888];
     layer1_out[4381] <= layer0_out[9477] | layer0_out[9478];
     layer1_out[4382] <= ~(layer0_out[10327] & layer0_out[10328]);
     layer1_out[4383] <= layer0_out[8240] | layer0_out[8241];
     layer1_out[4384] <= layer0_out[9590];
     layer1_out[4385] <= layer0_out[331] & layer0_out[332];
     layer1_out[4386] <= layer0_out[11194] & layer0_out[11195];
     layer1_out[4387] <= ~layer0_out[2389] | layer0_out[2388];
     layer1_out[4388] <= ~layer0_out[10794] | layer0_out[10793];
     layer1_out[4389] <= ~layer0_out[2533];
     layer1_out[4390] <= layer0_out[5771] | layer0_out[5772];
     layer1_out[4391] <= layer0_out[767];
     layer1_out[4392] <= layer0_out[8907] | layer0_out[8908];
     layer1_out[4393] <= layer0_out[2848];
     layer1_out[4394] <= layer0_out[11710] & ~layer0_out[11711];
     layer1_out[4395] <= ~layer0_out[5366];
     layer1_out[4396] <= ~layer0_out[3574] | layer0_out[3575];
     layer1_out[4397] <= layer0_out[11706];
     layer1_out[4398] <= layer0_out[7192];
     layer1_out[4399] <= layer0_out[4723];
     layer1_out[4400] <= layer0_out[4183];
     layer1_out[4401] <= ~layer0_out[4841];
     layer1_out[4402] <= ~(layer0_out[3565] ^ layer0_out[3566]);
     layer1_out[4403] <= ~(layer0_out[8736] & layer0_out[8737]);
     layer1_out[4404] <= layer0_out[4530] & layer0_out[4531];
     layer1_out[4405] <= layer0_out[9460] & ~layer0_out[9459];
     layer1_out[4406] <= layer0_out[9780] & ~layer0_out[9779];
     layer1_out[4407] <= ~layer0_out[504] | layer0_out[505];
     layer1_out[4408] <= layer0_out[2412] | layer0_out[2413];
     layer1_out[4409] <= layer0_out[10294] | layer0_out[10295];
     layer1_out[4410] <= ~(layer0_out[3138] | layer0_out[3139]);
     layer1_out[4411] <= layer0_out[5784] & ~layer0_out[5783];
     layer1_out[4412] <= layer0_out[73] & ~layer0_out[72];
     layer1_out[4413] <= ~(layer0_out[6291] & layer0_out[6292]);
     layer1_out[4414] <= layer0_out[9907] | layer0_out[9908];
     layer1_out[4415] <= ~layer0_out[1151] | layer0_out[1152];
     layer1_out[4416] <= layer0_out[4511] & ~layer0_out[4512];
     layer1_out[4417] <= ~(layer0_out[7363] & layer0_out[7364]);
     layer1_out[4418] <= layer0_out[7761] & layer0_out[7762];
     layer1_out[4419] <= ~(layer0_out[8091] | layer0_out[8092]);
     layer1_out[4420] <= ~layer0_out[11136];
     layer1_out[4421] <= layer0_out[2511] & layer0_out[2512];
     layer1_out[4422] <= layer0_out[1578];
     layer1_out[4423] <= layer0_out[11010];
     layer1_out[4424] <= ~(layer0_out[462] & layer0_out[463]);
     layer1_out[4425] <= ~(layer0_out[7580] | layer0_out[7581]);
     layer1_out[4426] <= ~layer0_out[6367] | layer0_out[6366];
     layer1_out[4427] <= layer0_out[9777];
     layer1_out[4428] <= ~layer0_out[6296];
     layer1_out[4429] <= layer0_out[6121];
     layer1_out[4430] <= layer0_out[6690] & ~layer0_out[6689];
     layer1_out[4431] <= ~layer0_out[3783];
     layer1_out[4432] <= layer0_out[516] & layer0_out[517];
     layer1_out[4433] <= ~layer0_out[7290];
     layer1_out[4434] <= layer0_out[4792];
     layer1_out[4435] <= layer0_out[11754];
     layer1_out[4436] <= layer0_out[3025] ^ layer0_out[3026];
     layer1_out[4437] <= ~layer0_out[6921] | layer0_out[6920];
     layer1_out[4438] <= ~(layer0_out[9624] & layer0_out[9625]);
     layer1_out[4439] <= 1'b0;
     layer1_out[4440] <= layer0_out[10244] | layer0_out[10245];
     layer1_out[4441] <= ~(layer0_out[3448] ^ layer0_out[3449]);
     layer1_out[4442] <= ~(layer0_out[10802] | layer0_out[10803]);
     layer1_out[4443] <= layer0_out[3857];
     layer1_out[4444] <= layer0_out[4573] | layer0_out[4574];
     layer1_out[4445] <= ~layer0_out[3592] | layer0_out[3593];
     layer1_out[4446] <= ~(layer0_out[7576] & layer0_out[7577]);
     layer1_out[4447] <= ~layer0_out[1503];
     layer1_out[4448] <= ~layer0_out[2952];
     layer1_out[4449] <= ~layer0_out[5089] | layer0_out[5088];
     layer1_out[4450] <= ~(layer0_out[9527] | layer0_out[9528]);
     layer1_out[4451] <= layer0_out[9539] & ~layer0_out[9538];
     layer1_out[4452] <= ~layer0_out[6337];
     layer1_out[4453] <= ~(layer0_out[176] ^ layer0_out[177]);
     layer1_out[4454] <= ~layer0_out[3254];
     layer1_out[4455] <= 1'b1;
     layer1_out[4456] <= layer0_out[10148] & ~layer0_out[10147];
     layer1_out[4457] <= ~(layer0_out[5413] & layer0_out[5414]);
     layer1_out[4458] <= 1'b0;
     layer1_out[4459] <= layer0_out[923] & ~layer0_out[924];
     layer1_out[4460] <= ~layer0_out[3445];
     layer1_out[4461] <= ~layer0_out[2964] | layer0_out[2963];
     layer1_out[4462] <= layer0_out[5471] ^ layer0_out[5472];
     layer1_out[4463] <= layer0_out[11241];
     layer1_out[4464] <= layer0_out[8087] ^ layer0_out[8088];
     layer1_out[4465] <= layer0_out[2461] & ~layer0_out[2460];
     layer1_out[4466] <= ~layer0_out[5703] | layer0_out[5704];
     layer1_out[4467] <= ~layer0_out[5177];
     layer1_out[4468] <= ~layer0_out[3784];
     layer1_out[4469] <= 1'b1;
     layer1_out[4470] <= ~layer0_out[5613] | layer0_out[5614];
     layer1_out[4471] <= layer0_out[7996];
     layer1_out[4472] <= layer0_out[2491];
     layer1_out[4473] <= layer0_out[1717] ^ layer0_out[1718];
     layer1_out[4474] <= ~layer0_out[5977];
     layer1_out[4475] <= ~(layer0_out[740] | layer0_out[741]);
     layer1_out[4476] <= ~layer0_out[3463];
     layer1_out[4477] <= ~layer0_out[5090] | layer0_out[5089];
     layer1_out[4478] <= ~layer0_out[2952];
     layer1_out[4479] <= ~layer0_out[8962] | layer0_out[8961];
     layer1_out[4480] <= layer0_out[7511] | layer0_out[7512];
     layer1_out[4481] <= ~layer0_out[4256];
     layer1_out[4482] <= ~(layer0_out[3262] & layer0_out[3263]);
     layer1_out[4483] <= ~(layer0_out[8922] | layer0_out[8923]);
     layer1_out[4484] <= ~layer0_out[4645];
     layer1_out[4485] <= layer0_out[7972] & layer0_out[7973];
     layer1_out[4486] <= layer0_out[4430] & ~layer0_out[4431];
     layer1_out[4487] <= ~layer0_out[1117];
     layer1_out[4488] <= ~(layer0_out[11588] & layer0_out[11589]);
     layer1_out[4489] <= ~(layer0_out[7434] & layer0_out[7435]);
     layer1_out[4490] <= ~layer0_out[9219] | layer0_out[9220];
     layer1_out[4491] <= ~layer0_out[987];
     layer1_out[4492] <= layer0_out[10576] & layer0_out[10577];
     layer1_out[4493] <= layer0_out[6307] & layer0_out[6308];
     layer1_out[4494] <= layer0_out[8626];
     layer1_out[4495] <= layer0_out[2385];
     layer1_out[4496] <= ~(layer0_out[7748] & layer0_out[7749]);
     layer1_out[4497] <= layer0_out[1767] & layer0_out[1768];
     layer1_out[4498] <= ~layer0_out[11893] | layer0_out[11892];
     layer1_out[4499] <= ~layer0_out[5055];
     layer1_out[4500] <= 1'b1;
     layer1_out[4501] <= ~layer0_out[6962];
     layer1_out[4502] <= layer0_out[4740];
     layer1_out[4503] <= ~(layer0_out[10595] ^ layer0_out[10596]);
     layer1_out[4504] <= ~layer0_out[11564] | layer0_out[11563];
     layer1_out[4505] <= ~layer0_out[4335] | layer0_out[4336];
     layer1_out[4506] <= layer0_out[2045] & ~layer0_out[2046];
     layer1_out[4507] <= layer0_out[2117];
     layer1_out[4508] <= layer0_out[1616] & ~layer0_out[1615];
     layer1_out[4509] <= ~(layer0_out[8811] ^ layer0_out[8812]);
     layer1_out[4510] <= layer0_out[8663] ^ layer0_out[8664];
     layer1_out[4511] <= layer0_out[5573] & ~layer0_out[5574];
     layer1_out[4512] <= layer0_out[9551] & layer0_out[9552];
     layer1_out[4513] <= ~layer0_out[5294];
     layer1_out[4514] <= layer0_out[10689];
     layer1_out[4515] <= ~layer0_out[6877] | layer0_out[6878];
     layer1_out[4516] <= ~layer0_out[8149] | layer0_out[8148];
     layer1_out[4517] <= ~layer0_out[6394];
     layer1_out[4518] <= ~(layer0_out[2650] ^ layer0_out[2651]);
     layer1_out[4519] <= ~layer0_out[10101];
     layer1_out[4520] <= ~(layer0_out[120] & layer0_out[121]);
     layer1_out[4521] <= layer0_out[4794];
     layer1_out[4522] <= layer0_out[9531] ^ layer0_out[9532];
     layer1_out[4523] <= layer0_out[9914];
     layer1_out[4524] <= layer0_out[9306];
     layer1_out[4525] <= ~layer0_out[6590];
     layer1_out[4526] <= 1'b0;
     layer1_out[4527] <= ~(layer0_out[10306] | layer0_out[10307]);
     layer1_out[4528] <= layer0_out[7546] | layer0_out[7547];
     layer1_out[4529] <= ~(layer0_out[6161] ^ layer0_out[6162]);
     layer1_out[4530] <= layer0_out[509];
     layer1_out[4531] <= ~(layer0_out[2300] ^ layer0_out[2301]);
     layer1_out[4532] <= ~layer0_out[6898] | layer0_out[6897];
     layer1_out[4533] <= ~(layer0_out[1294] ^ layer0_out[1295]);
     layer1_out[4534] <= layer0_out[6185] | layer0_out[6186];
     layer1_out[4535] <= layer0_out[1357];
     layer1_out[4536] <= layer0_out[1664] | layer0_out[1665];
     layer1_out[4537] <= layer0_out[5008];
     layer1_out[4538] <= layer0_out[1729] | layer0_out[1730];
     layer1_out[4539] <= ~layer0_out[2771];
     layer1_out[4540] <= ~(layer0_out[2276] | layer0_out[2277]);
     layer1_out[4541] <= ~layer0_out[3462];
     layer1_out[4542] <= layer0_out[4149] & layer0_out[4150];
     layer1_out[4543] <= ~layer0_out[9974];
     layer1_out[4544] <= layer0_out[5595];
     layer1_out[4545] <= layer0_out[3061];
     layer1_out[4546] <= ~(layer0_out[8830] | layer0_out[8831]);
     layer1_out[4547] <= layer0_out[2314] | layer0_out[2315];
     layer1_out[4548] <= ~layer0_out[9762];
     layer1_out[4549] <= ~layer0_out[7088];
     layer1_out[4550] <= ~layer0_out[2378] | layer0_out[2379];
     layer1_out[4551] <= ~layer0_out[9894] | layer0_out[9895];
     layer1_out[4552] <= layer0_out[1631];
     layer1_out[4553] <= ~(layer0_out[3047] | layer0_out[3048]);
     layer1_out[4554] <= 1'b1;
     layer1_out[4555] <= ~layer0_out[10227] | layer0_out[10226];
     layer1_out[4556] <= ~layer0_out[1009];
     layer1_out[4557] <= ~layer0_out[55];
     layer1_out[4558] <= layer0_out[8711] & layer0_out[8712];
     layer1_out[4559] <= ~layer0_out[2080];
     layer1_out[4560] <= layer0_out[4287] ^ layer0_out[4288];
     layer1_out[4561] <= ~(layer0_out[8328] & layer0_out[8329]);
     layer1_out[4562] <= ~layer0_out[8215] | layer0_out[8216];
     layer1_out[4563] <= ~layer0_out[4672] | layer0_out[4673];
     layer1_out[4564] <= ~(layer0_out[2779] & layer0_out[2780]);
     layer1_out[4565] <= layer0_out[5999] & ~layer0_out[6000];
     layer1_out[4566] <= layer0_out[9797] & ~layer0_out[9796];
     layer1_out[4567] <= layer0_out[925];
     layer1_out[4568] <= layer0_out[11655];
     layer1_out[4569] <= ~layer0_out[2840];
     layer1_out[4570] <= ~layer0_out[1790] | layer0_out[1789];
     layer1_out[4571] <= layer0_out[8528];
     layer1_out[4572] <= layer0_out[7916] & layer0_out[7917];
     layer1_out[4573] <= ~layer0_out[7137] | layer0_out[7136];
     layer1_out[4574] <= ~layer0_out[1087] | layer0_out[1086];
     layer1_out[4575] <= ~(layer0_out[3823] & layer0_out[3824]);
     layer1_out[4576] <= 1'b1;
     layer1_out[4577] <= layer0_out[2537] & layer0_out[2538];
     layer1_out[4578] <= ~layer0_out[7795] | layer0_out[7794];
     layer1_out[4579] <= ~layer0_out[9994];
     layer1_out[4580] <= layer0_out[988];
     layer1_out[4581] <= layer0_out[4309] & ~layer0_out[4310];
     layer1_out[4582] <= ~layer0_out[3877];
     layer1_out[4583] <= layer0_out[7748] & ~layer0_out[7747];
     layer1_out[4584] <= ~layer0_out[8947] | layer0_out[8946];
     layer1_out[4585] <= ~layer0_out[2189] | layer0_out[2188];
     layer1_out[4586] <= layer0_out[3835] & ~layer0_out[3836];
     layer1_out[4587] <= ~layer0_out[2700];
     layer1_out[4588] <= ~(layer0_out[7960] & layer0_out[7961]);
     layer1_out[4589] <= layer0_out[4503] & ~layer0_out[4504];
     layer1_out[4590] <= ~layer0_out[8615] | layer0_out[8616];
     layer1_out[4591] <= layer0_out[5329] & ~layer0_out[5330];
     layer1_out[4592] <= ~layer0_out[3928];
     layer1_out[4593] <= layer0_out[5813] & ~layer0_out[5812];
     layer1_out[4594] <= 1'b1;
     layer1_out[4595] <= ~layer0_out[7247] | layer0_out[7246];
     layer1_out[4596] <= layer0_out[5945] & layer0_out[5946];
     layer1_out[4597] <= layer0_out[1258];
     layer1_out[4598] <= layer0_out[11155] & layer0_out[11156];
     layer1_out[4599] <= layer0_out[11614] ^ layer0_out[11615];
     layer1_out[4600] <= layer0_out[8485];
     layer1_out[4601] <= layer0_out[2543] & ~layer0_out[2542];
     layer1_out[4602] <= layer0_out[6706] & layer0_out[6707];
     layer1_out[4603] <= layer0_out[5078] ^ layer0_out[5079];
     layer1_out[4604] <= layer0_out[1536] & ~layer0_out[1535];
     layer1_out[4605] <= layer0_out[10769];
     layer1_out[4606] <= ~layer0_out[5063] | layer0_out[5062];
     layer1_out[4607] <= ~layer0_out[3254];
     layer1_out[4608] <= ~(layer0_out[4943] & layer0_out[4944]);
     layer1_out[4609] <= ~layer0_out[8801] | layer0_out[8802];
     layer1_out[4610] <= ~layer0_out[8218];
     layer1_out[4611] <= ~(layer0_out[5596] & layer0_out[5597]);
     layer1_out[4612] <= layer0_out[3043] & layer0_out[3044];
     layer1_out[4613] <= ~layer0_out[1335] | layer0_out[1336];
     layer1_out[4614] <= layer0_out[1584] & layer0_out[1585];
     layer1_out[4615] <= layer0_out[2886] & ~layer0_out[2885];
     layer1_out[4616] <= ~(layer0_out[249] & layer0_out[250]);
     layer1_out[4617] <= layer0_out[6224] & ~layer0_out[6225];
     layer1_out[4618] <= layer0_out[10045] & ~layer0_out[10046];
     layer1_out[4619] <= layer0_out[5360] & ~layer0_out[5361];
     layer1_out[4620] <= ~layer0_out[9940] | layer0_out[9939];
     layer1_out[4621] <= layer0_out[1491];
     layer1_out[4622] <= layer0_out[10285] & ~layer0_out[10284];
     layer1_out[4623] <= layer0_out[585];
     layer1_out[4624] <= ~layer0_out[5862] | layer0_out[5861];
     layer1_out[4625] <= layer0_out[1816];
     layer1_out[4626] <= ~layer0_out[4748];
     layer1_out[4627] <= ~layer0_out[6081] | layer0_out[6080];
     layer1_out[4628] <= ~layer0_out[6986] | layer0_out[6985];
     layer1_out[4629] <= ~layer0_out[10371] | layer0_out[10370];
     layer1_out[4630] <= ~layer0_out[5254];
     layer1_out[4631] <= 1'b1;
     layer1_out[4632] <= ~layer0_out[2078];
     layer1_out[4633] <= layer0_out[9965] | layer0_out[9966];
     layer1_out[4634] <= ~layer0_out[8749];
     layer1_out[4635] <= ~(layer0_out[7137] & layer0_out[7138]);
     layer1_out[4636] <= layer0_out[2330] & layer0_out[2331];
     layer1_out[4637] <= layer0_out[1276];
     layer1_out[4638] <= ~layer0_out[9838] | layer0_out[9839];
     layer1_out[4639] <= ~layer0_out[10818] | layer0_out[10819];
     layer1_out[4640] <= ~layer0_out[6498] | layer0_out[6499];
     layer1_out[4641] <= ~layer0_out[2678];
     layer1_out[4642] <= ~layer0_out[7791];
     layer1_out[4643] <= ~layer0_out[539];
     layer1_out[4644] <= layer0_out[9705] | layer0_out[9706];
     layer1_out[4645] <= layer0_out[4728] & layer0_out[4729];
     layer1_out[4646] <= layer0_out[8460] & layer0_out[8461];
     layer1_out[4647] <= ~(layer0_out[2425] | layer0_out[2426]);
     layer1_out[4648] <= layer0_out[607];
     layer1_out[4649] <= ~(layer0_out[4073] & layer0_out[4074]);
     layer1_out[4650] <= layer0_out[352] & ~layer0_out[353];
     layer1_out[4651] <= layer0_out[8804];
     layer1_out[4652] <= layer0_out[7292];
     layer1_out[4653] <= layer0_out[9033] & ~layer0_out[9034];
     layer1_out[4654] <= layer0_out[5531] & ~layer0_out[5532];
     layer1_out[4655] <= ~layer0_out[10261];
     layer1_out[4656] <= ~(layer0_out[6738] & layer0_out[6739]);
     layer1_out[4657] <= ~layer0_out[1552];
     layer1_out[4658] <= ~layer0_out[11412];
     layer1_out[4659] <= layer0_out[9352];
     layer1_out[4660] <= ~layer0_out[6959] | layer0_out[6960];
     layer1_out[4661] <= ~layer0_out[7824] | layer0_out[7825];
     layer1_out[4662] <= ~layer0_out[1438];
     layer1_out[4663] <= layer0_out[3999] & ~layer0_out[4000];
     layer1_out[4664] <= ~layer0_out[4121] | layer0_out[4122];
     layer1_out[4665] <= layer0_out[199] ^ layer0_out[200];
     layer1_out[4666] <= ~layer0_out[846];
     layer1_out[4667] <= ~(layer0_out[1487] & layer0_out[1488]);
     layer1_out[4668] <= layer0_out[7206];
     layer1_out[4669] <= layer0_out[6898];
     layer1_out[4670] <= layer0_out[3075] & ~layer0_out[3076];
     layer1_out[4671] <= ~layer0_out[8914];
     layer1_out[4672] <= ~(layer0_out[4141] | layer0_out[4142]);
     layer1_out[4673] <= ~layer0_out[954] | layer0_out[953];
     layer1_out[4674] <= ~(layer0_out[10543] | layer0_out[10544]);
     layer1_out[4675] <= ~(layer0_out[6344] ^ layer0_out[6345]);
     layer1_out[4676] <= layer0_out[4258];
     layer1_out[4677] <= layer0_out[426];
     layer1_out[4678] <= layer0_out[6072] ^ layer0_out[6073];
     layer1_out[4679] <= 1'b1;
     layer1_out[4680] <= layer0_out[4642] & ~layer0_out[4643];
     layer1_out[4681] <= ~layer0_out[5489] | layer0_out[5488];
     layer1_out[4682] <= 1'b0;
     layer1_out[4683] <= ~layer0_out[1600];
     layer1_out[4684] <= ~(layer0_out[11793] & layer0_out[11794]);
     layer1_out[4685] <= layer0_out[9905];
     layer1_out[4686] <= ~(layer0_out[2443] ^ layer0_out[2444]);
     layer1_out[4687] <= ~(layer0_out[11814] | layer0_out[11815]);
     layer1_out[4688] <= layer0_out[7922] | layer0_out[7923];
     layer1_out[4689] <= layer0_out[11562] & ~layer0_out[11561];
     layer1_out[4690] <= layer0_out[1092] & layer0_out[1093];
     layer1_out[4691] <= layer0_out[8996] & ~layer0_out[8997];
     layer1_out[4692] <= layer0_out[2938] & layer0_out[2939];
     layer1_out[4693] <= layer0_out[3267] | layer0_out[3268];
     layer1_out[4694] <= ~layer0_out[278];
     layer1_out[4695] <= ~layer0_out[6919] | layer0_out[6920];
     layer1_out[4696] <= ~layer0_out[4314];
     layer1_out[4697] <= ~layer0_out[9230] | layer0_out[9229];
     layer1_out[4698] <= layer0_out[5019] & layer0_out[5020];
     layer1_out[4699] <= layer0_out[529];
     layer1_out[4700] <= layer0_out[7789] | layer0_out[7790];
     layer1_out[4701] <= layer0_out[8490];
     layer1_out[4702] <= 1'b0;
     layer1_out[4703] <= ~layer0_out[8285] | layer0_out[8284];
     layer1_out[4704] <= ~layer0_out[1586];
     layer1_out[4705] <= layer0_out[7386];
     layer1_out[4706] <= ~(layer0_out[3697] & layer0_out[3698]);
     layer1_out[4707] <= ~(layer0_out[905] & layer0_out[906]);
     layer1_out[4708] <= ~(layer0_out[5896] & layer0_out[5897]);
     layer1_out[4709] <= 1'b0;
     layer1_out[4710] <= ~layer0_out[3448];
     layer1_out[4711] <= layer0_out[7672];
     layer1_out[4712] <= layer0_out[3333];
     layer1_out[4713] <= ~(layer0_out[1910] | layer0_out[1911]);
     layer1_out[4714] <= 1'b0;
     layer1_out[4715] <= ~layer0_out[11720];
     layer1_out[4716] <= ~(layer0_out[1420] ^ layer0_out[1421]);
     layer1_out[4717] <= ~(layer0_out[4330] ^ layer0_out[4331]);
     layer1_out[4718] <= ~layer0_out[86];
     layer1_out[4719] <= layer0_out[1461];
     layer1_out[4720] <= ~layer0_out[3425];
     layer1_out[4721] <= layer0_out[11098] & ~layer0_out[11099];
     layer1_out[4722] <= ~layer0_out[158] | layer0_out[159];
     layer1_out[4723] <= ~(layer0_out[1504] ^ layer0_out[1505]);
     layer1_out[4724] <= layer0_out[9091];
     layer1_out[4725] <= ~layer0_out[9798];
     layer1_out[4726] <= ~layer0_out[7603] | layer0_out[7604];
     layer1_out[4727] <= ~layer0_out[8073] | layer0_out[8074];
     layer1_out[4728] <= layer0_out[10296] & layer0_out[10297];
     layer1_out[4729] <= ~(layer0_out[5836] ^ layer0_out[5837]);
     layer1_out[4730] <= layer0_out[6303];
     layer1_out[4731] <= ~(layer0_out[11260] & layer0_out[11261]);
     layer1_out[4732] <= ~layer0_out[6977];
     layer1_out[4733] <= ~layer0_out[2564] | layer0_out[2565];
     layer1_out[4734] <= layer0_out[7023];
     layer1_out[4735] <= layer0_out[1995] & ~layer0_out[1994];
     layer1_out[4736] <= layer0_out[10342] ^ layer0_out[10343];
     layer1_out[4737] <= ~(layer0_out[8656] | layer0_out[8657]);
     layer1_out[4738] <= layer0_out[3288];
     layer1_out[4739] <= layer0_out[2735];
     layer1_out[4740] <= ~(layer0_out[11495] | layer0_out[11496]);
     layer1_out[4741] <= 1'b0;
     layer1_out[4742] <= ~(layer0_out[3453] & layer0_out[3454]);
     layer1_out[4743] <= ~layer0_out[11120];
     layer1_out[4744] <= layer0_out[1298];
     layer1_out[4745] <= ~layer0_out[10817];
     layer1_out[4746] <= ~layer0_out[4644];
     layer1_out[4747] <= layer0_out[3305] & ~layer0_out[3306];
     layer1_out[4748] <= 1'b1;
     layer1_out[4749] <= layer0_out[9383];
     layer1_out[4750] <= layer0_out[7092] & ~layer0_out[7093];
     layer1_out[4751] <= layer0_out[4497] & ~layer0_out[4498];
     layer1_out[4752] <= ~layer0_out[7092];
     layer1_out[4753] <= layer0_out[4101] | layer0_out[4102];
     layer1_out[4754] <= ~layer0_out[1832];
     layer1_out[4755] <= ~layer0_out[5169] | layer0_out[5168];
     layer1_out[4756] <= layer0_out[10618];
     layer1_out[4757] <= layer0_out[9067] | layer0_out[9068];
     layer1_out[4758] <= layer0_out[7235] & ~layer0_out[7236];
     layer1_out[4759] <= layer0_out[7026];
     layer1_out[4760] <= ~layer0_out[8508];
     layer1_out[4761] <= ~(layer0_out[11932] & layer0_out[11933]);
     layer1_out[4762] <= layer0_out[11362] & ~layer0_out[11363];
     layer1_out[4763] <= layer0_out[2377] & ~layer0_out[2376];
     layer1_out[4764] <= layer0_out[11151] & ~layer0_out[11152];
     layer1_out[4765] <= ~(layer0_out[6089] | layer0_out[6090]);
     layer1_out[4766] <= ~layer0_out[4003];
     layer1_out[4767] <= ~(layer0_out[5770] | layer0_out[5771]);
     layer1_out[4768] <= 1'b0;
     layer1_out[4769] <= ~(layer0_out[7973] ^ layer0_out[7974]);
     layer1_out[4770] <= layer0_out[6044] | layer0_out[6045];
     layer1_out[4771] <= ~layer0_out[7822];
     layer1_out[4772] <= ~layer0_out[10726];
     layer1_out[4773] <= ~layer0_out[5219] | layer0_out[5220];
     layer1_out[4774] <= layer0_out[11872] ^ layer0_out[11873];
     layer1_out[4775] <= ~(layer0_out[8936] | layer0_out[8937]);
     layer1_out[4776] <= ~layer0_out[9320];
     layer1_out[4777] <= layer0_out[7774] & ~layer0_out[7775];
     layer1_out[4778] <= layer0_out[5280] | layer0_out[5281];
     layer1_out[4779] <= layer0_out[3356] | layer0_out[3357];
     layer1_out[4780] <= ~layer0_out[10041];
     layer1_out[4781] <= ~layer0_out[165];
     layer1_out[4782] <= layer0_out[11525] & layer0_out[11526];
     layer1_out[4783] <= layer0_out[1573];
     layer1_out[4784] <= ~(layer0_out[6301] & layer0_out[6302]);
     layer1_out[4785] <= ~layer0_out[5706];
     layer1_out[4786] <= layer0_out[8114] & layer0_out[8115];
     layer1_out[4787] <= layer0_out[2287] & ~layer0_out[2288];
     layer1_out[4788] <= ~layer0_out[6211];
     layer1_out[4789] <= ~(layer0_out[8313] & layer0_out[8314]);
     layer1_out[4790] <= ~(layer0_out[281] | layer0_out[282]);
     layer1_out[4791] <= 1'b0;
     layer1_out[4792] <= ~(layer0_out[8633] | layer0_out[8634]);
     layer1_out[4793] <= layer0_out[5262] & ~layer0_out[5261];
     layer1_out[4794] <= layer0_out[8584] & ~layer0_out[8585];
     layer1_out[4795] <= layer0_out[716] | layer0_out[717];
     layer1_out[4796] <= layer0_out[7194] & ~layer0_out[7193];
     layer1_out[4797] <= ~layer0_out[11941] | layer0_out[11940];
     layer1_out[4798] <= layer0_out[6392] & ~layer0_out[6391];
     layer1_out[4799] <= ~layer0_out[7394] | layer0_out[7393];
     layer1_out[4800] <= layer0_out[1841];
     layer1_out[4801] <= ~(layer0_out[10152] | layer0_out[10153]);
     layer1_out[4802] <= layer0_out[11398] | layer0_out[11399];
     layer1_out[4803] <= ~layer0_out[8538];
     layer1_out[4804] <= ~layer0_out[8150] | layer0_out[8151];
     layer1_out[4805] <= 1'b0;
     layer1_out[4806] <= ~(layer0_out[9182] & layer0_out[9183]);
     layer1_out[4807] <= layer0_out[3041];
     layer1_out[4808] <= layer0_out[10489] & layer0_out[10490];
     layer1_out[4809] <= ~layer0_out[10676];
     layer1_out[4810] <= layer0_out[264] & ~layer0_out[263];
     layer1_out[4811] <= ~(layer0_out[9355] ^ layer0_out[9356]);
     layer1_out[4812] <= ~(layer0_out[6862] & layer0_out[6863]);
     layer1_out[4813] <= layer0_out[9052] & layer0_out[9053];
     layer1_out[4814] <= layer0_out[11859];
     layer1_out[4815] <= ~layer0_out[7798] | layer0_out[7799];
     layer1_out[4816] <= layer0_out[10021];
     layer1_out[4817] <= layer0_out[8483] & ~layer0_out[8484];
     layer1_out[4818] <= layer0_out[8356];
     layer1_out[4819] <= ~(layer0_out[668] | layer0_out[669]);
     layer1_out[4820] <= ~layer0_out[7198] | layer0_out[7197];
     layer1_out[4821] <= ~(layer0_out[10846] | layer0_out[10847]);
     layer1_out[4822] <= ~layer0_out[4285];
     layer1_out[4823] <= layer0_out[11306];
     layer1_out[4824] <= ~layer0_out[9417];
     layer1_out[4825] <= ~layer0_out[6922];
     layer1_out[4826] <= ~layer0_out[3914] | layer0_out[3913];
     layer1_out[4827] <= layer0_out[5543];
     layer1_out[4828] <= ~(layer0_out[1417] | layer0_out[1418]);
     layer1_out[4829] <= ~layer0_out[10922] | layer0_out[10921];
     layer1_out[4830] <= layer0_out[10795] & ~layer0_out[10794];
     layer1_out[4831] <= layer0_out[5245] ^ layer0_out[5246];
     layer1_out[4832] <= layer0_out[11805] & ~layer0_out[11806];
     layer1_out[4833] <= ~(layer0_out[1800] | layer0_out[1801]);
     layer1_out[4834] <= layer0_out[4266];
     layer1_out[4835] <= layer0_out[10053] | layer0_out[10054];
     layer1_out[4836] <= layer0_out[5910] & ~layer0_out[5911];
     layer1_out[4837] <= ~(layer0_out[9493] ^ layer0_out[9494]);
     layer1_out[4838] <= layer0_out[1671] & layer0_out[1672];
     layer1_out[4839] <= layer0_out[3643];
     layer1_out[4840] <= layer0_out[2517];
     layer1_out[4841] <= layer0_out[11253] ^ layer0_out[11254];
     layer1_out[4842] <= layer0_out[4513] & layer0_out[4514];
     layer1_out[4843] <= ~(layer0_out[242] ^ layer0_out[243]);
     layer1_out[4844] <= layer0_out[8439] & ~layer0_out[8440];
     layer1_out[4845] <= ~layer0_out[9738] | layer0_out[9737];
     layer1_out[4846] <= layer0_out[2507];
     layer1_out[4847] <= layer0_out[7009];
     layer1_out[4848] <= layer0_out[9212] & layer0_out[9213];
     layer1_out[4849] <= ~layer0_out[1747] | layer0_out[1746];
     layer1_out[4850] <= ~(layer0_out[2403] & layer0_out[2404]);
     layer1_out[4851] <= layer0_out[4222] | layer0_out[4223];
     layer1_out[4852] <= layer0_out[5350] & ~layer0_out[5351];
     layer1_out[4853] <= 1'b0;
     layer1_out[4854] <= layer0_out[3677] & ~layer0_out[3678];
     layer1_out[4855] <= layer0_out[3831] & ~layer0_out[3832];
     layer1_out[4856] <= layer0_out[2991] & ~layer0_out[2992];
     layer1_out[4857] <= ~layer0_out[1555] | layer0_out[1556];
     layer1_out[4858] <= layer0_out[3465] ^ layer0_out[3466];
     layer1_out[4859] <= ~layer0_out[1799];
     layer1_out[4860] <= ~(layer0_out[10072] & layer0_out[10073]);
     layer1_out[4861] <= layer0_out[5627] & layer0_out[5628];
     layer1_out[4862] <= layer0_out[10800] & layer0_out[10801];
     layer1_out[4863] <= layer0_out[2941];
     layer1_out[4864] <= ~(layer0_out[10860] & layer0_out[10861]);
     layer1_out[4865] <= ~layer0_out[6497] | layer0_out[6498];
     layer1_out[4866] <= layer0_out[5756] & layer0_out[5757];
     layer1_out[4867] <= ~layer0_out[1200];
     layer1_out[4868] <= ~layer0_out[2236];
     layer1_out[4869] <= layer0_out[8193] & layer0_out[8194];
     layer1_out[4870] <= ~layer0_out[3401];
     layer1_out[4871] <= layer0_out[2918] & ~layer0_out[2919];
     layer1_out[4872] <= ~layer0_out[4875] | layer0_out[4876];
     layer1_out[4873] <= layer0_out[10168] & ~layer0_out[10169];
     layer1_out[4874] <= layer0_out[8905] & ~layer0_out[8906];
     layer1_out[4875] <= layer0_out[10086] & layer0_out[10087];
     layer1_out[4876] <= ~layer0_out[1641];
     layer1_out[4877] <= ~layer0_out[10788];
     layer1_out[4878] <= layer0_out[1875];
     layer1_out[4879] <= ~layer0_out[5123] | layer0_out[5124];
     layer1_out[4880] <= ~layer0_out[9301] | layer0_out[9302];
     layer1_out[4881] <= ~layer0_out[10851];
     layer1_out[4882] <= ~(layer0_out[8781] & layer0_out[8782]);
     layer1_out[4883] <= layer0_out[7438];
     layer1_out[4884] <= layer0_out[7194];
     layer1_out[4885] <= layer0_out[8562] | layer0_out[8563];
     layer1_out[4886] <= layer0_out[2340] & ~layer0_out[2341];
     layer1_out[4887] <= 1'b1;
     layer1_out[4888] <= layer0_out[8159] & ~layer0_out[8158];
     layer1_out[4889] <= layer0_out[466] ^ layer0_out[467];
     layer1_out[4890] <= ~layer0_out[6227];
     layer1_out[4891] <= layer0_out[9652];
     layer1_out[4892] <= ~layer0_out[10614] | layer0_out[10615];
     layer1_out[4893] <= layer0_out[5163] ^ layer0_out[5164];
     layer1_out[4894] <= layer0_out[5432] & ~layer0_out[5433];
     layer1_out[4895] <= ~layer0_out[1168] | layer0_out[1169];
     layer1_out[4896] <= ~(layer0_out[3691] & layer0_out[3692]);
     layer1_out[4897] <= layer0_out[10512];
     layer1_out[4898] <= layer0_out[4614] & ~layer0_out[4613];
     layer1_out[4899] <= layer0_out[3279] & ~layer0_out[3278];
     layer1_out[4900] <= ~layer0_out[5798];
     layer1_out[4901] <= ~layer0_out[11251];
     layer1_out[4902] <= layer0_out[8414] | layer0_out[8415];
     layer1_out[4903] <= layer0_out[5040];
     layer1_out[4904] <= ~layer0_out[4517];
     layer1_out[4905] <= ~layer0_out[8789];
     layer1_out[4906] <= layer0_out[8202] & ~layer0_out[8203];
     layer1_out[4907] <= layer0_out[10468];
     layer1_out[4908] <= layer0_out[1812] | layer0_out[1813];
     layer1_out[4909] <= layer0_out[11333];
     layer1_out[4910] <= layer0_out[3821];
     layer1_out[4911] <= ~layer0_out[11922];
     layer1_out[4912] <= ~layer0_out[901];
     layer1_out[4913] <= layer0_out[1737];
     layer1_out[4914] <= ~layer0_out[5792] | layer0_out[5791];
     layer1_out[4915] <= layer0_out[7948] & layer0_out[7949];
     layer1_out[4916] <= ~(layer0_out[5956] | layer0_out[5957]);
     layer1_out[4917] <= ~layer0_out[10434];
     layer1_out[4918] <= layer0_out[1577];
     layer1_out[4919] <= ~layer0_out[3316];
     layer1_out[4920] <= ~layer0_out[2183] | layer0_out[2184];
     layer1_out[4921] <= layer0_out[439];
     layer1_out[4922] <= layer0_out[8980];
     layer1_out[4923] <= layer0_out[198];
     layer1_out[4924] <= layer0_out[11611];
     layer1_out[4925] <= ~layer0_out[752];
     layer1_out[4926] <= layer0_out[573];
     layer1_out[4927] <= layer0_out[6387] & ~layer0_out[6388];
     layer1_out[4928] <= ~layer0_out[11713];
     layer1_out[4929] <= layer0_out[1923] ^ layer0_out[1924];
     layer1_out[4930] <= layer0_out[9891] & ~layer0_out[9892];
     layer1_out[4931] <= layer0_out[10593] & layer0_out[10594];
     layer1_out[4932] <= 1'b1;
     layer1_out[4933] <= layer0_out[6324] & ~layer0_out[6325];
     layer1_out[4934] <= ~(layer0_out[7028] ^ layer0_out[7029]);
     layer1_out[4935] <= ~(layer0_out[3122] & layer0_out[3123]);
     layer1_out[4936] <= layer0_out[10221];
     layer1_out[4937] <= layer0_out[4930];
     layer1_out[4938] <= ~layer0_out[7222];
     layer1_out[4939] <= ~(layer0_out[1599] | layer0_out[1600]);
     layer1_out[4940] <= ~layer0_out[3517];
     layer1_out[4941] <= layer0_out[6744];
     layer1_out[4942] <= layer0_out[7563] | layer0_out[7564];
     layer1_out[4943] <= layer0_out[3786] & ~layer0_out[3787];
     layer1_out[4944] <= ~layer0_out[3507] | layer0_out[3506];
     layer1_out[4945] <= layer0_out[10621] & ~layer0_out[10620];
     layer1_out[4946] <= ~(layer0_out[9015] ^ layer0_out[9016]);
     layer1_out[4947] <= ~layer0_out[6906];
     layer1_out[4948] <= ~layer0_out[5859];
     layer1_out[4949] <= ~(layer0_out[10150] & layer0_out[10151]);
     layer1_out[4950] <= ~layer0_out[6255];
     layer1_out[4951] <= layer0_out[4535] & ~layer0_out[4534];
     layer1_out[4952] <= layer0_out[2884] & ~layer0_out[2885];
     layer1_out[4953] <= ~(layer0_out[10240] | layer0_out[10241]);
     layer1_out[4954] <= layer0_out[3579];
     layer1_out[4955] <= layer0_out[11396] | layer0_out[11397];
     layer1_out[4956] <= ~layer0_out[4284] | layer0_out[4283];
     layer1_out[4957] <= ~layer0_out[11250] | layer0_out[11249];
     layer1_out[4958] <= layer0_out[2199] & ~layer0_out[2200];
     layer1_out[4959] <= layer0_out[274] ^ layer0_out[275];
     layer1_out[4960] <= ~layer0_out[2152];
     layer1_out[4961] <= ~layer0_out[65];
     layer1_out[4962] <= layer0_out[5035] & ~layer0_out[5036];
     layer1_out[4963] <= ~(layer0_out[2233] & layer0_out[2234]);
     layer1_out[4964] <= ~layer0_out[2786] | layer0_out[2785];
     layer1_out[4965] <= 1'b0;
     layer1_out[4966] <= layer0_out[4192] | layer0_out[4193];
     layer1_out[4967] <= ~(layer0_out[9967] & layer0_out[9968]);
     layer1_out[4968] <= ~layer0_out[4473] | layer0_out[4474];
     layer1_out[4969] <= layer0_out[4032] & ~layer0_out[4031];
     layer1_out[4970] <= ~layer0_out[1103] | layer0_out[1102];
     layer1_out[4971] <= ~(layer0_out[11158] | layer0_out[11159]);
     layer1_out[4972] <= layer0_out[10276] & ~layer0_out[10277];
     layer1_out[4973] <= ~layer0_out[8846] | layer0_out[8847];
     layer1_out[4974] <= layer0_out[8007];
     layer1_out[4975] <= ~layer0_out[1196];
     layer1_out[4976] <= ~layer0_out[1942];
     layer1_out[4977] <= layer0_out[16] ^ layer0_out[17];
     layer1_out[4978] <= layer0_out[9277] | layer0_out[9278];
     layer1_out[4979] <= ~(layer0_out[5429] | layer0_out[5430]);
     layer1_out[4980] <= layer0_out[10670] | layer0_out[10671];
     layer1_out[4981] <= ~layer0_out[7091] | layer0_out[7090];
     layer1_out[4982] <= layer0_out[9191] & ~layer0_out[9192];
     layer1_out[4983] <= layer0_out[6812] | layer0_out[6813];
     layer1_out[4984] <= ~layer0_out[3289];
     layer1_out[4985] <= ~(layer0_out[10077] & layer0_out[10078]);
     layer1_out[4986] <= layer0_out[3646] & layer0_out[3647];
     layer1_out[4987] <= ~layer0_out[3575];
     layer1_out[4988] <= layer0_out[6915];
     layer1_out[4989] <= layer0_out[4610];
     layer1_out[4990] <= ~(layer0_out[7934] | layer0_out[7935]);
     layer1_out[4991] <= 1'b1;
     layer1_out[4992] <= layer0_out[4967] & ~layer0_out[4968];
     layer1_out[4993] <= ~layer0_out[2437];
     layer1_out[4994] <= ~(layer0_out[4704] ^ layer0_out[4705]);
     layer1_out[4995] <= ~layer0_out[2756];
     layer1_out[4996] <= layer0_out[3704] & ~layer0_out[3705];
     layer1_out[4997] <= ~layer0_out[11735] | layer0_out[11734];
     layer1_out[4998] <= layer0_out[9894];
     layer1_out[4999] <= layer0_out[2965];
     layer1_out[5000] <= layer0_out[8876];
     layer1_out[5001] <= layer0_out[5980] & ~layer0_out[5981];
     layer1_out[5002] <= ~layer0_out[1568] | layer0_out[1569];
     layer1_out[5003] <= layer0_out[7646] & ~layer0_out[7645];
     layer1_out[5004] <= layer0_out[1032] & ~layer0_out[1033];
     layer1_out[5005] <= ~(layer0_out[3431] ^ layer0_out[3432]);
     layer1_out[5006] <= layer0_out[1868] | layer0_out[1869];
     layer1_out[5007] <= ~layer0_out[8083] | layer0_out[8082];
     layer1_out[5008] <= ~(layer0_out[5815] | layer0_out[5816]);
     layer1_out[5009] <= ~(layer0_out[1880] ^ layer0_out[1881]);
     layer1_out[5010] <= ~(layer0_out[9723] ^ layer0_out[9724]);
     layer1_out[5011] <= layer0_out[6796] | layer0_out[6797];
     layer1_out[5012] <= ~layer0_out[210];
     layer1_out[5013] <= layer0_out[6525];
     layer1_out[5014] <= ~(layer0_out[3801] & layer0_out[3802]);
     layer1_out[5015] <= layer0_out[3037];
     layer1_out[5016] <= ~(layer0_out[858] | layer0_out[859]);
     layer1_out[5017] <= layer0_out[1408];
     layer1_out[5018] <= layer0_out[10988] & layer0_out[10989];
     layer1_out[5019] <= ~layer0_out[1641] | layer0_out[1642];
     layer1_out[5020] <= ~layer0_out[7882];
     layer1_out[5021] <= 1'b1;
     layer1_out[5022] <= ~layer0_out[5731] | layer0_out[5730];
     layer1_out[5023] <= layer0_out[6333] & layer0_out[6334];
     layer1_out[5024] <= ~(layer0_out[3915] | layer0_out[3916]);
     layer1_out[5025] <= 1'b0;
     layer1_out[5026] <= layer0_out[3660];
     layer1_out[5027] <= ~layer0_out[7210] | layer0_out[7209];
     layer1_out[5028] <= ~layer0_out[2049];
     layer1_out[5029] <= layer0_out[5153] & ~layer0_out[5152];
     layer1_out[5030] <= layer0_out[3168];
     layer1_out[5031] <= ~(layer0_out[10557] | layer0_out[10558]);
     layer1_out[5032] <= ~layer0_out[556];
     layer1_out[5033] <= ~layer0_out[10331];
     layer1_out[5034] <= layer0_out[11892];
     layer1_out[5035] <= ~layer0_out[6867];
     layer1_out[5036] <= ~(layer0_out[2707] ^ layer0_out[2708]);
     layer1_out[5037] <= 1'b0;
     layer1_out[5038] <= layer0_out[10299] & ~layer0_out[10300];
     layer1_out[5039] <= layer0_out[5688] & ~layer0_out[5689];
     layer1_out[5040] <= layer0_out[1240] & ~layer0_out[1241];
     layer1_out[5041] <= layer0_out[10630] & ~layer0_out[10629];
     layer1_out[5042] <= layer0_out[9282];
     layer1_out[5043] <= ~layer0_out[11369];
     layer1_out[5044] <= layer0_out[10462];
     layer1_out[5045] <= ~(layer0_out[3313] & layer0_out[3314]);
     layer1_out[5046] <= ~(layer0_out[650] & layer0_out[651]);
     layer1_out[5047] <= layer0_out[5440] | layer0_out[5441];
     layer1_out[5048] <= layer0_out[5284];
     layer1_out[5049] <= layer0_out[347] | layer0_out[348];
     layer1_out[5050] <= layer0_out[8548] & ~layer0_out[8547];
     layer1_out[5051] <= layer0_out[11281] ^ layer0_out[11282];
     layer1_out[5052] <= ~(layer0_out[1080] | layer0_out[1081]);
     layer1_out[5053] <= ~(layer0_out[5750] | layer0_out[5751]);
     layer1_out[5054] <= ~(layer0_out[1514] | layer0_out[1515]);
     layer1_out[5055] <= ~(layer0_out[10199] ^ layer0_out[10200]);
     layer1_out[5056] <= ~(layer0_out[11534] | layer0_out[11535]);
     layer1_out[5057] <= ~(layer0_out[11265] & layer0_out[11266]);
     layer1_out[5058] <= ~(layer0_out[3315] ^ layer0_out[3316]);
     layer1_out[5059] <= layer0_out[6000];
     layer1_out[5060] <= layer0_out[6787] ^ layer0_out[6788];
     layer1_out[5061] <= layer0_out[3155] | layer0_out[3156];
     layer1_out[5062] <= ~layer0_out[661] | layer0_out[662];
     layer1_out[5063] <= ~layer0_out[7235];
     layer1_out[5064] <= ~(layer0_out[4730] ^ layer0_out[4731]);
     layer1_out[5065] <= ~(layer0_out[8970] ^ layer0_out[8971]);
     layer1_out[5066] <= ~layer0_out[589];
     layer1_out[5067] <= layer0_out[9714] & ~layer0_out[9713];
     layer1_out[5068] <= ~(layer0_out[8397] ^ layer0_out[8398]);
     layer1_out[5069] <= ~(layer0_out[1634] & layer0_out[1635]);
     layer1_out[5070] <= ~layer0_out[9993];
     layer1_out[5071] <= ~(layer0_out[3573] | layer0_out[3574]);
     layer1_out[5072] <= layer0_out[10189] & layer0_out[10190];
     layer1_out[5073] <= 1'b0;
     layer1_out[5074] <= ~(layer0_out[8652] | layer0_out[8653]);
     layer1_out[5075] <= layer0_out[8057] & ~layer0_out[8056];
     layer1_out[5076] <= layer0_out[5880] & ~layer0_out[5879];
     layer1_out[5077] <= ~layer0_out[3482];
     layer1_out[5078] <= ~layer0_out[6901] | layer0_out[6900];
     layer1_out[5079] <= ~layer0_out[2643];
     layer1_out[5080] <= ~layer0_out[4021];
     layer1_out[5081] <= 1'b1;
     layer1_out[5082] <= layer0_out[11451] ^ layer0_out[11452];
     layer1_out[5083] <= ~(layer0_out[11011] | layer0_out[11012]);
     layer1_out[5084] <= ~layer0_out[7156];
     layer1_out[5085] <= layer0_out[4032] | layer0_out[4033];
     layer1_out[5086] <= layer0_out[2232];
     layer1_out[5087] <= layer0_out[5731];
     layer1_out[5088] <= ~(layer0_out[1957] | layer0_out[1958]);
     layer1_out[5089] <= ~layer0_out[7982] | layer0_out[7983];
     layer1_out[5090] <= ~(layer0_out[2783] | layer0_out[2784]);
     layer1_out[5091] <= ~(layer0_out[8731] | layer0_out[8732]);
     layer1_out[5092] <= layer0_out[7887] & ~layer0_out[7886];
     layer1_out[5093] <= ~layer0_out[10015] | layer0_out[10016];
     layer1_out[5094] <= ~layer0_out[6965] | layer0_out[6966];
     layer1_out[5095] <= ~layer0_out[5470];
     layer1_out[5096] <= layer0_out[5434] & ~layer0_out[5433];
     layer1_out[5097] <= ~(layer0_out[3244] ^ layer0_out[3245]);
     layer1_out[5098] <= ~(layer0_out[436] ^ layer0_out[437]);
     layer1_out[5099] <= ~layer0_out[10175] | layer0_out[10174];
     layer1_out[5100] <= layer0_out[9588] & layer0_out[9589];
     layer1_out[5101] <= layer0_out[66] & ~layer0_out[67];
     layer1_out[5102] <= layer0_out[11363] | layer0_out[11364];
     layer1_out[5103] <= ~layer0_out[1062] | layer0_out[1063];
     layer1_out[5104] <= ~layer0_out[6303] | layer0_out[6304];
     layer1_out[5105] <= layer0_out[11059] | layer0_out[11060];
     layer1_out[5106] <= layer0_out[155] & layer0_out[156];
     layer1_out[5107] <= layer0_out[9404] & ~layer0_out[9405];
     layer1_out[5108] <= ~layer0_out[11295] | layer0_out[11296];
     layer1_out[5109] <= layer0_out[5195] | layer0_out[5196];
     layer1_out[5110] <= layer0_out[3488] & ~layer0_out[3489];
     layer1_out[5111] <= layer0_out[5981] | layer0_out[5982];
     layer1_out[5112] <= layer0_out[9872];
     layer1_out[5113] <= 1'b0;
     layer1_out[5114] <= ~layer0_out[7944] | layer0_out[7943];
     layer1_out[5115] <= layer0_out[6107] & layer0_out[6108];
     layer1_out[5116] <= ~(layer0_out[6614] | layer0_out[6615]);
     layer1_out[5117] <= ~(layer0_out[5881] | layer0_out[5882]);
     layer1_out[5118] <= layer0_out[11757];
     layer1_out[5119] <= ~layer0_out[810];
     layer1_out[5120] <= layer0_out[3167] | layer0_out[3168];
     layer1_out[5121] <= layer0_out[1565] & layer0_out[1566];
     layer1_out[5122] <= ~layer0_out[2933];
     layer1_out[5123] <= 1'b0;
     layer1_out[5124] <= ~layer0_out[11223];
     layer1_out[5125] <= ~layer0_out[10248] | layer0_out[10247];
     layer1_out[5126] <= layer0_out[7321];
     layer1_out[5127] <= layer0_out[1489] & ~layer0_out[1490];
     layer1_out[5128] <= ~(layer0_out[3083] ^ layer0_out[3084]);
     layer1_out[5129] <= ~layer0_out[9708];
     layer1_out[5130] <= layer0_out[11851] | layer0_out[11852];
     layer1_out[5131] <= ~(layer0_out[9632] ^ layer0_out[9633]);
     layer1_out[5132] <= ~(layer0_out[922] | layer0_out[923]);
     layer1_out[5133] <= layer0_out[4723];
     layer1_out[5134] <= ~(layer0_out[9807] | layer0_out[9808]);
     layer1_out[5135] <= ~(layer0_out[11823] | layer0_out[11824]);
     layer1_out[5136] <= layer0_out[8855] & layer0_out[8856];
     layer1_out[5137] <= layer0_out[6589] & ~layer0_out[6588];
     layer1_out[5138] <= ~layer0_out[11035];
     layer1_out[5139] <= ~(layer0_out[11232] | layer0_out[11233]);
     layer1_out[5140] <= ~layer0_out[690] | layer0_out[691];
     layer1_out[5141] <= ~layer0_out[6503] | layer0_out[6504];
     layer1_out[5142] <= ~(layer0_out[4788] & layer0_out[4789]);
     layer1_out[5143] <= layer0_out[1036] ^ layer0_out[1037];
     layer1_out[5144] <= ~layer0_out[2328];
     layer1_out[5145] <= layer0_out[9638];
     layer1_out[5146] <= ~(layer0_out[9540] ^ layer0_out[9541]);
     layer1_out[5147] <= layer0_out[8933] & layer0_out[8934];
     layer1_out[5148] <= layer0_out[8513] ^ layer0_out[8514];
     layer1_out[5149] <= ~layer0_out[7420];
     layer1_out[5150] <= layer0_out[11361] | layer0_out[11362];
     layer1_out[5151] <= ~(layer0_out[122] ^ layer0_out[123]);
     layer1_out[5152] <= ~layer0_out[9956];
     layer1_out[5153] <= 1'b0;
     layer1_out[5154] <= ~(layer0_out[322] | layer0_out[323]);
     layer1_out[5155] <= layer0_out[6709];
     layer1_out[5156] <= ~(layer0_out[3512] ^ layer0_out[3513]);
     layer1_out[5157] <= layer0_out[1319] & ~layer0_out[1320];
     layer1_out[5158] <= layer0_out[153] & layer0_out[154];
     layer1_out[5159] <= ~layer0_out[11270] | layer0_out[11271];
     layer1_out[5160] <= layer0_out[6443];
     layer1_out[5161] <= ~(layer0_out[490] | layer0_out[491]);
     layer1_out[5162] <= layer0_out[11743] ^ layer0_out[11744];
     layer1_out[5163] <= layer0_out[8794];
     layer1_out[5164] <= ~(layer0_out[3503] & layer0_out[3504]);
     layer1_out[5165] <= ~layer0_out[6028] | layer0_out[6027];
     layer1_out[5166] <= layer0_out[5855];
     layer1_out[5167] <= ~layer0_out[1360] | layer0_out[1361];
     layer1_out[5168] <= layer0_out[5232] & layer0_out[5233];
     layer1_out[5169] <= ~(layer0_out[461] & layer0_out[462]);
     layer1_out[5170] <= layer0_out[7451] & ~layer0_out[7450];
     layer1_out[5171] <= layer0_out[2867];
     layer1_out[5172] <= layer0_out[6437];
     layer1_out[5173] <= layer0_out[11854];
     layer1_out[5174] <= ~(layer0_out[6334] | layer0_out[6335]);
     layer1_out[5175] <= ~(layer0_out[8043] ^ layer0_out[8044]);
     layer1_out[5176] <= ~(layer0_out[1446] | layer0_out[1447]);
     layer1_out[5177] <= layer0_out[4099] ^ layer0_out[4100];
     layer1_out[5178] <= layer0_out[208];
     layer1_out[5179] <= layer0_out[3497] | layer0_out[3498];
     layer1_out[5180] <= ~layer0_out[9628] | layer0_out[9627];
     layer1_out[5181] <= layer0_out[11569] & ~layer0_out[11568];
     layer1_out[5182] <= layer0_out[2682];
     layer1_out[5183] <= layer0_out[4092] & ~layer0_out[4093];
     layer1_out[5184] <= ~layer0_out[7114] | layer0_out[7113];
     layer1_out[5185] <= layer0_out[4867] & layer0_out[4868];
     layer1_out[5186] <= layer0_out[6686];
     layer1_out[5187] <= ~layer0_out[11991];
     layer1_out[5188] <= layer0_out[9635] | layer0_out[9636];
     layer1_out[5189] <= layer0_out[5230] ^ layer0_out[5231];
     layer1_out[5190] <= ~layer0_out[7253];
     layer1_out[5191] <= layer0_out[4824] | layer0_out[4825];
     layer1_out[5192] <= ~(layer0_out[6282] & layer0_out[6283]);
     layer1_out[5193] <= layer0_out[5401] & ~layer0_out[5402];
     layer1_out[5194] <= ~layer0_out[832] | layer0_out[833];
     layer1_out[5195] <= ~layer0_out[1339];
     layer1_out[5196] <= layer0_out[1005] ^ layer0_out[1006];
     layer1_out[5197] <= layer0_out[11518] & ~layer0_out[11517];
     layer1_out[5198] <= layer0_out[5626] & layer0_out[5627];
     layer1_out[5199] <= layer0_out[7065] & ~layer0_out[7066];
     layer1_out[5200] <= ~layer0_out[6865] | layer0_out[6866];
     layer1_out[5201] <= layer0_out[11839] ^ layer0_out[11840];
     layer1_out[5202] <= ~layer0_out[5961] | layer0_out[5962];
     layer1_out[5203] <= layer0_out[3234];
     layer1_out[5204] <= ~layer0_out[2697] | layer0_out[2698];
     layer1_out[5205] <= layer0_out[10131] & layer0_out[10132];
     layer1_out[5206] <= layer0_out[7636] & ~layer0_out[7635];
     layer1_out[5207] <= layer0_out[11899];
     layer1_out[5208] <= ~(layer0_out[9270] & layer0_out[9271]);
     layer1_out[5209] <= ~layer0_out[880];
     layer1_out[5210] <= ~layer0_out[5884];
     layer1_out[5211] <= 1'b0;
     layer1_out[5212] <= layer0_out[11018] & layer0_out[11019];
     layer1_out[5213] <= ~layer0_out[207];
     layer1_out[5214] <= ~layer0_out[6723];
     layer1_out[5215] <= ~(layer0_out[288] & layer0_out[289]);
     layer1_out[5216] <= ~layer0_out[3177];
     layer1_out[5217] <= 1'b1;
     layer1_out[5218] <= ~layer0_out[387] | layer0_out[386];
     layer1_out[5219] <= layer0_out[3081] | layer0_out[3082];
     layer1_out[5220] <= ~(layer0_out[10500] & layer0_out[10501]);
     layer1_out[5221] <= ~layer0_out[4375] | layer0_out[4376];
     layer1_out[5222] <= ~layer0_out[10257];
     layer1_out[5223] <= layer0_out[3076] & layer0_out[3077];
     layer1_out[5224] <= ~(layer0_out[1862] | layer0_out[1863]);
     layer1_out[5225] <= ~layer0_out[11835];
     layer1_out[5226] <= layer0_out[11132];
     layer1_out[5227] <= ~layer0_out[5072] | layer0_out[5071];
     layer1_out[5228] <= layer0_out[11809] & ~layer0_out[11808];
     layer1_out[5229] <= 1'b0;
     layer1_out[5230] <= layer0_out[2029] | layer0_out[2030];
     layer1_out[5231] <= ~(layer0_out[8900] ^ layer0_out[8901]);
     layer1_out[5232] <= layer0_out[566] & ~layer0_out[565];
     layer1_out[5233] <= ~layer0_out[5723] | layer0_out[5722];
     layer1_out[5234] <= layer0_out[4672] & ~layer0_out[4671];
     layer1_out[5235] <= layer0_out[11411];
     layer1_out[5236] <= ~layer0_out[7090];
     layer1_out[5237] <= layer0_out[10056] ^ layer0_out[10057];
     layer1_out[5238] <= layer0_out[253] ^ layer0_out[254];
     layer1_out[5239] <= ~layer0_out[3207];
     layer1_out[5240] <= layer0_out[2286] | layer0_out[2287];
     layer1_out[5241] <= ~(layer0_out[4558] | layer0_out[4559]);
     layer1_out[5242] <= ~layer0_out[1096];
     layer1_out[5243] <= ~layer0_out[2887];
     layer1_out[5244] <= ~layer0_out[1416] | layer0_out[1417];
     layer1_out[5245] <= ~(layer0_out[3534] ^ layer0_out[3535]);
     layer1_out[5246] <= ~(layer0_out[4454] ^ layer0_out[4455]);
     layer1_out[5247] <= layer0_out[2242] | layer0_out[2243];
     layer1_out[5248] <= layer0_out[1033] & ~layer0_out[1034];
     layer1_out[5249] <= ~layer0_out[7542] | layer0_out[7543];
     layer1_out[5250] <= layer0_out[3935];
     layer1_out[5251] <= ~layer0_out[755];
     layer1_out[5252] <= layer0_out[11233];
     layer1_out[5253] <= ~layer0_out[11246];
     layer1_out[5254] <= layer0_out[844] & layer0_out[845];
     layer1_out[5255] <= layer0_out[1377] & layer0_out[1378];
     layer1_out[5256] <= ~layer0_out[7110];
     layer1_out[5257] <= ~layer0_out[2094] | layer0_out[2095];
     layer1_out[5258] <= ~layer0_out[9828] | layer0_out[9827];
     layer1_out[5259] <= layer0_out[7244] & layer0_out[7245];
     layer1_out[5260] <= 1'b0;
     layer1_out[5261] <= layer0_out[3242];
     layer1_out[5262] <= layer0_out[4504] ^ layer0_out[4505];
     layer1_out[5263] <= ~(layer0_out[6313] | layer0_out[6314]);
     layer1_out[5264] <= ~(layer0_out[8079] & layer0_out[8080]);
     layer1_out[5265] <= layer0_out[10520];
     layer1_out[5266] <= layer0_out[3410];
     layer1_out[5267] <= layer0_out[3562];
     layer1_out[5268] <= ~layer0_out[6471];
     layer1_out[5269] <= layer0_out[3908] & layer0_out[3909];
     layer1_out[5270] <= layer0_out[2383] & layer0_out[2384];
     layer1_out[5271] <= ~layer0_out[562];
     layer1_out[5272] <= layer0_out[7482] ^ layer0_out[7483];
     layer1_out[5273] <= ~(layer0_out[6872] | layer0_out[6873]);
     layer1_out[5274] <= layer0_out[10170];
     layer1_out[5275] <= layer0_out[3096] & ~layer0_out[3097];
     layer1_out[5276] <= ~layer0_out[7160];
     layer1_out[5277] <= layer0_out[3126] & layer0_out[3127];
     layer1_out[5278] <= ~(layer0_out[9354] | layer0_out[9355]);
     layer1_out[5279] <= ~layer0_out[2177];
     layer1_out[5280] <= layer0_out[3798] & layer0_out[3799];
     layer1_out[5281] <= ~layer0_out[760] | layer0_out[759];
     layer1_out[5282] <= layer0_out[4662];
     layer1_out[5283] <= layer0_out[8705] ^ layer0_out[8706];
     layer1_out[5284] <= layer0_out[7737] & ~layer0_out[7736];
     layer1_out[5285] <= layer0_out[11176] & layer0_out[11177];
     layer1_out[5286] <= layer0_out[11023] ^ layer0_out[11024];
     layer1_out[5287] <= layer0_out[8880] | layer0_out[8881];
     layer1_out[5288] <= layer0_out[1989] & layer0_out[1990];
     layer1_out[5289] <= layer0_out[3160] & layer0_out[3161];
     layer1_out[5290] <= layer0_out[10109] ^ layer0_out[10110];
     layer1_out[5291] <= ~layer0_out[10963];
     layer1_out[5292] <= layer0_out[432] & layer0_out[433];
     layer1_out[5293] <= layer0_out[9616] & ~layer0_out[9617];
     layer1_out[5294] <= ~layer0_out[3920] | layer0_out[3921];
     layer1_out[5295] <= ~(layer0_out[8303] & layer0_out[8304]);
     layer1_out[5296] <= ~layer0_out[10580];
     layer1_out[5297] <= ~(layer0_out[5625] ^ layer0_out[5626]);
     layer1_out[5298] <= layer0_out[10499];
     layer1_out[5299] <= layer0_out[7199] & ~layer0_out[7200];
     layer1_out[5300] <= layer0_out[2386];
     layer1_out[5301] <= ~(layer0_out[742] | layer0_out[743]);
     layer1_out[5302] <= ~layer0_out[478] | layer0_out[477];
     layer1_out[5303] <= ~layer0_out[3885];
     layer1_out[5304] <= layer0_out[2575];
     layer1_out[5305] <= ~(layer0_out[8895] ^ layer0_out[8896]);
     layer1_out[5306] <= ~layer0_out[11717];
     layer1_out[5307] <= ~layer0_out[1750];
     layer1_out[5308] <= layer0_out[3031] ^ layer0_out[3032];
     layer1_out[5309] <= ~layer0_out[5923];
     layer1_out[5310] <= layer0_out[5944] & ~layer0_out[5943];
     layer1_out[5311] <= layer0_out[4816] & layer0_out[4817];
     layer1_out[5312] <= layer0_out[7041] | layer0_out[7042];
     layer1_out[5313] <= layer0_out[3603];
     layer1_out[5314] <= ~layer0_out[11899] | layer0_out[11900];
     layer1_out[5315] <= layer0_out[10894];
     layer1_out[5316] <= layer0_out[5454] | layer0_out[5455];
     layer1_out[5317] <= ~layer0_out[10840] | layer0_out[10841];
     layer1_out[5318] <= layer0_out[10873] & ~layer0_out[10874];
     layer1_out[5319] <= ~layer0_out[11728];
     layer1_out[5320] <= layer0_out[3634] & layer0_out[3635];
     layer1_out[5321] <= ~layer0_out[6557] | layer0_out[6558];
     layer1_out[5322] <= ~layer0_out[2875];
     layer1_out[5323] <= ~layer0_out[11698];
     layer1_out[5324] <= layer0_out[7201];
     layer1_out[5325] <= ~(layer0_out[967] ^ layer0_out[968]);
     layer1_out[5326] <= ~layer0_out[11931];
     layer1_out[5327] <= ~layer0_out[8640];
     layer1_out[5328] <= layer0_out[7700] & ~layer0_out[7701];
     layer1_out[5329] <= ~layer0_out[6735];
     layer1_out[5330] <= 1'b0;
     layer1_out[5331] <= ~layer0_out[10379];
     layer1_out[5332] <= layer0_out[3361] & ~layer0_out[3360];
     layer1_out[5333] <= ~layer0_out[1302];
     layer1_out[5334] <= layer0_out[9376] & layer0_out[9377];
     layer1_out[5335] <= layer0_out[11681];
     layer1_out[5336] <= layer0_out[5153];
     layer1_out[5337] <= ~(layer0_out[10236] | layer0_out[10237]);
     layer1_out[5338] <= layer0_out[2295];
     layer1_out[5339] <= ~layer0_out[10866] | layer0_out[10865];
     layer1_out[5340] <= ~layer0_out[2536] | layer0_out[2535];
     layer1_out[5341] <= ~layer0_out[848];
     layer1_out[5342] <= layer0_out[8812];
     layer1_out[5343] <= layer0_out[9951];
     layer1_out[5344] <= layer0_out[9051];
     layer1_out[5345] <= layer0_out[4969];
     layer1_out[5346] <= layer0_out[6353];
     layer1_out[5347] <= ~(layer0_out[3591] | layer0_out[3592]);
     layer1_out[5348] <= layer0_out[3256] & ~layer0_out[3257];
     layer1_out[5349] <= ~(layer0_out[9072] & layer0_out[9073]);
     layer1_out[5350] <= ~layer0_out[11961] | layer0_out[11962];
     layer1_out[5351] <= ~(layer0_out[2197] ^ layer0_out[2198]);
     layer1_out[5352] <= ~layer0_out[1880];
     layer1_out[5353] <= layer0_out[800] & layer0_out[801];
     layer1_out[5354] <= layer0_out[6067];
     layer1_out[5355] <= ~layer0_out[8152] | layer0_out[8153];
     layer1_out[5356] <= ~(layer0_out[2710] | layer0_out[2711]);
     layer1_out[5357] <= ~layer0_out[6401] | layer0_out[6402];
     layer1_out[5358] <= ~layer0_out[744];
     layer1_out[5359] <= layer0_out[7909];
     layer1_out[5360] <= layer0_out[6063] & ~layer0_out[6062];
     layer1_out[5361] <= layer0_out[11366];
     layer1_out[5362] <= ~layer0_out[3013] | layer0_out[3012];
     layer1_out[5363] <= ~layer0_out[7720];
     layer1_out[5364] <= layer0_out[1955];
     layer1_out[5365] <= ~layer0_out[4164];
     layer1_out[5366] <= ~layer0_out[978];
     layer1_out[5367] <= layer0_out[10090];
     layer1_out[5368] <= layer0_out[10332];
     layer1_out[5369] <= layer0_out[2573] | layer0_out[2574];
     layer1_out[5370] <= ~layer0_out[1501];
     layer1_out[5371] <= layer0_out[7619];
     layer1_out[5372] <= layer0_out[11664];
     layer1_out[5373] <= ~(layer0_out[2127] ^ layer0_out[2128]);
     layer1_out[5374] <= layer0_out[251] | layer0_out[252];
     layer1_out[5375] <= ~layer0_out[2500];
     layer1_out[5376] <= ~layer0_out[4960] | layer0_out[4961];
     layer1_out[5377] <= ~layer0_out[10601];
     layer1_out[5378] <= ~layer0_out[8772] | layer0_out[8771];
     layer1_out[5379] <= layer0_out[11030] & ~layer0_out[11029];
     layer1_out[5380] <= layer0_out[4863] | layer0_out[4864];
     layer1_out[5381] <= layer0_out[11254] | layer0_out[11255];
     layer1_out[5382] <= layer0_out[37];
     layer1_out[5383] <= layer0_out[8658] ^ layer0_out[8659];
     layer1_out[5384] <= ~layer0_out[2793] | layer0_out[2794];
     layer1_out[5385] <= layer0_out[4164];
     layer1_out[5386] <= layer0_out[3689] & ~layer0_out[3690];
     layer1_out[5387] <= layer0_out[5270] & ~layer0_out[5271];
     layer1_out[5388] <= 1'b1;
     layer1_out[5389] <= ~layer0_out[629];
     layer1_out[5390] <= layer0_out[10437];
     layer1_out[5391] <= layer0_out[1297];
     layer1_out[5392] <= ~(layer0_out[10896] & layer0_out[10897]);
     layer1_out[5393] <= layer0_out[11635] & layer0_out[11636];
     layer1_out[5394] <= layer0_out[6294] ^ layer0_out[6295];
     layer1_out[5395] <= layer0_out[2223] & layer0_out[2224];
     layer1_out[5396] <= 1'b0;
     layer1_out[5397] <= layer0_out[3889] ^ layer0_out[3890];
     layer1_out[5398] <= 1'b1;
     layer1_out[5399] <= ~(layer0_out[10705] & layer0_out[10706]);
     layer1_out[5400] <= ~layer0_out[2221];
     layer1_out[5401] <= 1'b0;
     layer1_out[5402] <= layer0_out[6909];
     layer1_out[5403] <= layer0_out[1345];
     layer1_out[5404] <= ~layer0_out[2483];
     layer1_out[5405] <= layer0_out[8971] & ~layer0_out[8972];
     layer1_out[5406] <= ~layer0_out[10291] | layer0_out[10292];
     layer1_out[5407] <= ~(layer0_out[5536] | layer0_out[5537]);
     layer1_out[5408] <= ~layer0_out[2313];
     layer1_out[5409] <= layer0_out[10177] & layer0_out[10178];
     layer1_out[5410] <= layer0_out[11108] | layer0_out[11109];
     layer1_out[5411] <= layer0_out[1223];
     layer1_out[5412] <= ~layer0_out[3967] | layer0_out[3968];
     layer1_out[5413] <= layer0_out[3166] & layer0_out[3167];
     layer1_out[5414] <= ~layer0_out[9005];
     layer1_out[5415] <= layer0_out[9300] & layer0_out[9301];
     layer1_out[5416] <= layer0_out[2124] & ~layer0_out[2125];
     layer1_out[5417] <= layer0_out[10935];
     layer1_out[5418] <= ~(layer0_out[4983] ^ layer0_out[4984]);
     layer1_out[5419] <= layer0_out[7798] & ~layer0_out[7797];
     layer1_out[5420] <= ~(layer0_out[7679] & layer0_out[7680]);
     layer1_out[5421] <= layer0_out[5187] & ~layer0_out[5186];
     layer1_out[5422] <= layer0_out[4426] & ~layer0_out[4427];
     layer1_out[5423] <= ~layer0_out[10421] | layer0_out[10420];
     layer1_out[5424] <= layer0_out[10904];
     layer1_out[5425] <= 1'b0;
     layer1_out[5426] <= layer0_out[4484] ^ layer0_out[4485];
     layer1_out[5427] <= ~layer0_out[2552];
     layer1_out[5428] <= ~(layer0_out[4491] | layer0_out[4492]);
     layer1_out[5429] <= layer0_out[11236];
     layer1_out[5430] <= ~(layer0_out[11789] & layer0_out[11790]);
     layer1_out[5431] <= layer0_out[2027];
     layer1_out[5432] <= layer0_out[6707];
     layer1_out[5433] <= layer0_out[7345];
     layer1_out[5434] <= ~layer0_out[2466];
     layer1_out[5435] <= layer0_out[7143];
     layer1_out[5436] <= ~(layer0_out[2906] & layer0_out[2907]);
     layer1_out[5437] <= ~layer0_out[9856] | layer0_out[9855];
     layer1_out[5438] <= ~(layer0_out[10271] ^ layer0_out[10272]);
     layer1_out[5439] <= ~layer0_out[11768];
     layer1_out[5440] <= layer0_out[156];
     layer1_out[5441] <= ~layer0_out[10051];
     layer1_out[5442] <= ~layer0_out[3345];
     layer1_out[5443] <= ~layer0_out[3826];
     layer1_out[5444] <= ~layer0_out[3150];
     layer1_out[5445] <= layer0_out[6844] | layer0_out[6845];
     layer1_out[5446] <= layer0_out[2005];
     layer1_out[5447] <= ~(layer0_out[8216] | layer0_out[8217]);
     layer1_out[5448] <= ~layer0_out[3086];
     layer1_out[5449] <= ~(layer0_out[8865] | layer0_out[8866]);
     layer1_out[5450] <= layer0_out[7143] | layer0_out[7144];
     layer1_out[5451] <= layer0_out[2771] | layer0_out[2772];
     layer1_out[5452] <= ~(layer0_out[1355] ^ layer0_out[1356]);
     layer1_out[5453] <= layer0_out[10549] ^ layer0_out[10550];
     layer1_out[5454] <= layer0_out[2988];
     layer1_out[5455] <= layer0_out[6906];
     layer1_out[5456] <= layer0_out[8620] & ~layer0_out[8619];
     layer1_out[5457] <= layer0_out[261];
     layer1_out[5458] <= ~(layer0_out[3414] & layer0_out[3415]);
     layer1_out[5459] <= layer0_out[8668] | layer0_out[8669];
     layer1_out[5460] <= layer0_out[6449];
     layer1_out[5461] <= ~(layer0_out[5883] ^ layer0_out[5884]);
     layer1_out[5462] <= layer0_out[9946] & ~layer0_out[9947];
     layer1_out[5463] <= layer0_out[7953] & ~layer0_out[7952];
     layer1_out[5464] <= layer0_out[9673] ^ layer0_out[9674];
     layer1_out[5465] <= layer0_out[8121];
     layer1_out[5466] <= layer0_out[40] & ~layer0_out[41];
     layer1_out[5467] <= ~layer0_out[11696] | layer0_out[11695];
     layer1_out[5468] <= ~(layer0_out[10138] | layer0_out[10139]);
     layer1_out[5469] <= ~layer0_out[11249];
     layer1_out[5470] <= ~layer0_out[597] | layer0_out[598];
     layer1_out[5471] <= ~layer0_out[9537] | layer0_out[9536];
     layer1_out[5472] <= layer0_out[1454];
     layer1_out[5473] <= layer0_out[8211] & layer0_out[8212];
     layer1_out[5474] <= 1'b1;
     layer1_out[5475] <= layer0_out[11832] & layer0_out[11833];
     layer1_out[5476] <= layer0_out[452];
     layer1_out[5477] <= ~layer0_out[7216];
     layer1_out[5478] <= layer0_out[8362];
     layer1_out[5479] <= layer0_out[6700] | layer0_out[6701];
     layer1_out[5480] <= ~layer0_out[150];
     layer1_out[5481] <= layer0_out[2735] & ~layer0_out[2734];
     layer1_out[5482] <= ~(layer0_out[1017] & layer0_out[1018]);
     layer1_out[5483] <= layer0_out[10384];
     layer1_out[5484] <= layer0_out[7150];
     layer1_out[5485] <= layer0_out[6882] & ~layer0_out[6881];
     layer1_out[5486] <= ~(layer0_out[4804] ^ layer0_out[4805]);
     layer1_out[5487] <= layer0_out[8641] ^ layer0_out[8642];
     layer1_out[5488] <= ~(layer0_out[8765] & layer0_out[8766]);
     layer1_out[5489] <= ~(layer0_out[9826] | layer0_out[9827]);
     layer1_out[5490] <= layer0_out[5873] | layer0_out[5874];
     layer1_out[5491] <= layer0_out[3438] & ~layer0_out[3437];
     layer1_out[5492] <= layer0_out[1172];
     layer1_out[5493] <= ~layer0_out[5070];
     layer1_out[5494] <= ~layer0_out[8147];
     layer1_out[5495] <= 1'b0;
     layer1_out[5496] <= ~(layer0_out[1059] & layer0_out[1060]);
     layer1_out[5497] <= layer0_out[3304] & ~layer0_out[3303];
     layer1_out[5498] <= layer0_out[1659] | layer0_out[1660];
     layer1_out[5499] <= ~layer0_out[822];
     layer1_out[5500] <= ~layer0_out[6365] | layer0_out[6366];
     layer1_out[5501] <= layer0_out[6875];
     layer1_out[5502] <= layer0_out[11428];
     layer1_out[5503] <= layer0_out[8253];
     layer1_out[5504] <= ~layer0_out[6338];
     layer1_out[5505] <= layer0_out[4601];
     layer1_out[5506] <= layer0_out[7696];
     layer1_out[5507] <= layer0_out[10532] ^ layer0_out[10533];
     layer1_out[5508] <= ~(layer0_out[11493] | layer0_out[11494]);
     layer1_out[5509] <= layer0_out[2514] & ~layer0_out[2515];
     layer1_out[5510] <= ~layer0_out[1356];
     layer1_out[5511] <= ~(layer0_out[9578] | layer0_out[9579]);
     layer1_out[5512] <= layer0_out[552] & layer0_out[553];
     layer1_out[5513] <= layer0_out[3686];
     layer1_out[5514] <= ~layer0_out[4695] | layer0_out[4696];
     layer1_out[5515] <= layer0_out[6849];
     layer1_out[5516] <= layer0_out[7422] & layer0_out[7423];
     layer1_out[5517] <= layer0_out[1008] & layer0_out[1009];
     layer1_out[5518] <= 1'b1;
     layer1_out[5519] <= layer0_out[10129];
     layer1_out[5520] <= ~layer0_out[2659];
     layer1_out[5521] <= layer0_out[6414] & ~layer0_out[6413];
     layer1_out[5522] <= ~(layer0_out[4091] | layer0_out[4092]);
     layer1_out[5523] <= layer0_out[10574];
     layer1_out[5524] <= layer0_out[3337];
     layer1_out[5525] <= layer0_out[4531] & ~layer0_out[4532];
     layer1_out[5526] <= layer0_out[3501];
     layer1_out[5527] <= ~layer0_out[410] | layer0_out[411];
     layer1_out[5528] <= layer0_out[10881] & ~layer0_out[10880];
     layer1_out[5529] <= ~layer0_out[3999] | layer0_out[3998];
     layer1_out[5530] <= layer0_out[5598];
     layer1_out[5531] <= ~layer0_out[8706];
     layer1_out[5532] <= ~layer0_out[8018];
     layer1_out[5533] <= layer0_out[10913] & layer0_out[10914];
     layer1_out[5534] <= layer0_out[5632];
     layer1_out[5535] <= ~layer0_out[8458];
     layer1_out[5536] <= ~layer0_out[9859] | layer0_out[9858];
     layer1_out[5537] <= layer0_out[9841] & layer0_out[9842];
     layer1_out[5538] <= layer0_out[131];
     layer1_out[5539] <= layer0_out[6167] & layer0_out[6168];
     layer1_out[5540] <= layer0_out[10521] & ~layer0_out[10522];
     layer1_out[5541] <= ~layer0_out[6184] | layer0_out[6183];
     layer1_out[5542] <= ~(layer0_out[4550] & layer0_out[4551]);
     layer1_out[5543] <= layer0_out[5765] & ~layer0_out[5764];
     layer1_out[5544] <= layer0_out[10017];
     layer1_out[5545] <= ~(layer0_out[7171] & layer0_out[7172]);
     layer1_out[5546] <= 1'b1;
     layer1_out[5547] <= ~layer0_out[2252];
     layer1_out[5548] <= ~(layer0_out[7440] | layer0_out[7441]);
     layer1_out[5549] <= ~layer0_out[740] | layer0_out[739];
     layer1_out[5550] <= ~layer0_out[778];
     layer1_out[5551] <= layer0_out[3042] & layer0_out[3043];
     layer1_out[5552] <= ~layer0_out[11223] | layer0_out[11222];
     layer1_out[5553] <= layer0_out[6066];
     layer1_out[5554] <= ~(layer0_out[9853] | layer0_out[9854]);
     layer1_out[5555] <= layer0_out[381];
     layer1_out[5556] <= layer0_out[657];
     layer1_out[5557] <= layer0_out[5213] | layer0_out[5214];
     layer1_out[5558] <= ~layer0_out[10687] | layer0_out[10686];
     layer1_out[5559] <= ~(layer0_out[10344] ^ layer0_out[10345]);
     layer1_out[5560] <= 1'b1;
     layer1_out[5561] <= ~layer0_out[11521];
     layer1_out[5562] <= layer0_out[3232] & layer0_out[3233];
     layer1_out[5563] <= ~layer0_out[3456] | layer0_out[3455];
     layer1_out[5564] <= layer0_out[5119];
     layer1_out[5565] <= layer0_out[9469] & ~layer0_out[9468];
     layer1_out[5566] <= ~(layer0_out[2557] & layer0_out[2558]);
     layer1_out[5567] <= layer0_out[1493] & ~layer0_out[1492];
     layer1_out[5568] <= ~layer0_out[2467];
     layer1_out[5569] <= layer0_out[3141];
     layer1_out[5570] <= ~layer0_out[5827];
     layer1_out[5571] <= 1'b0;
     layer1_out[5572] <= ~(layer0_out[6549] ^ layer0_out[6550]);
     layer1_out[5573] <= ~(layer0_out[6618] | layer0_out[6619]);
     layer1_out[5574] <= ~layer0_out[6075];
     layer1_out[5575] <= ~layer0_out[407] | layer0_out[408];
     layer1_out[5576] <= ~layer0_out[5604] | layer0_out[5603];
     layer1_out[5577] <= layer0_out[9173];
     layer1_out[5578] <= ~layer0_out[11644] | layer0_out[11643];
     layer1_out[5579] <= ~layer0_out[7754];
     layer1_out[5580] <= ~layer0_out[8129] | layer0_out[8130];
     layer1_out[5581] <= ~(layer0_out[5254] & layer0_out[5255]);
     layer1_out[5582] <= ~layer0_out[9836];
     layer1_out[5583] <= layer0_out[7492];
     layer1_out[5584] <= layer0_out[7605] & ~layer0_out[7606];
     layer1_out[5585] <= layer0_out[4607] & layer0_out[4608];
     layer1_out[5586] <= layer0_out[5008];
     layer1_out[5587] <= ~layer0_out[9748];
     layer1_out[5588] <= layer0_out[9696] & ~layer0_out[9697];
     layer1_out[5589] <= ~layer0_out[7882];
     layer1_out[5590] <= layer0_out[1757];
     layer1_out[5591] <= ~layer0_out[10731];
     layer1_out[5592] <= layer0_out[7951];
     layer1_out[5593] <= layer0_out[4347] & layer0_out[4348];
     layer1_out[5594] <= ~layer0_out[1648];
     layer1_out[5595] <= layer0_out[1145] | layer0_out[1146];
     layer1_out[5596] <= layer0_out[6388];
     layer1_out[5597] <= ~layer0_out[4970] | layer0_out[4971];
     layer1_out[5598] <= ~layer0_out[3869];
     layer1_out[5599] <= ~(layer0_out[5058] ^ layer0_out[5059]);
     layer1_out[5600] <= ~(layer0_out[9157] & layer0_out[9158]);
     layer1_out[5601] <= layer0_out[5362] & ~layer0_out[5361];
     layer1_out[5602] <= layer0_out[721];
     layer1_out[5603] <= ~layer0_out[6692];
     layer1_out[5604] <= layer0_out[5286] & ~layer0_out[5285];
     layer1_out[5605] <= layer0_out[10359] & layer0_out[10360];
     layer1_out[5606] <= layer0_out[1239] & layer0_out[1240];
     layer1_out[5607] <= layer0_out[1519] & layer0_out[1520];
     layer1_out[5608] <= layer0_out[10980] & ~layer0_out[10981];
     layer1_out[5609] <= layer0_out[6463];
     layer1_out[5610] <= ~layer0_out[3280];
     layer1_out[5611] <= 1'b0;
     layer1_out[5612] <= layer0_out[5367];
     layer1_out[5613] <= layer0_out[9327] & layer0_out[9328];
     layer1_out[5614] <= ~layer0_out[1940];
     layer1_out[5615] <= layer0_out[1716];
     layer1_out[5616] <= 1'b0;
     layer1_out[5617] <= ~layer0_out[6656];
     layer1_out[5618] <= 1'b1;
     layer1_out[5619] <= layer0_out[3006] ^ layer0_out[3007];
     layer1_out[5620] <= layer0_out[4439] & layer0_out[4440];
     layer1_out[5621] <= layer0_out[5951];
     layer1_out[5622] <= ~(layer0_out[2582] & layer0_out[2583]);
     layer1_out[5623] <= ~layer0_out[1346];
     layer1_out[5624] <= ~layer0_out[4842];
     layer1_out[5625] <= layer0_out[7640] & ~layer0_out[7641];
     layer1_out[5626] <= layer0_out[9056];
     layer1_out[5627] <= ~layer0_out[6822] | layer0_out[6823];
     layer1_out[5628] <= layer0_out[3261] & ~layer0_out[3260];
     layer1_out[5629] <= ~layer0_out[1814];
     layer1_out[5630] <= layer0_out[747];
     layer1_out[5631] <= ~(layer0_out[10744] | layer0_out[10745]);
     layer1_out[5632] <= layer0_out[1915] & ~layer0_out[1916];
     layer1_out[5633] <= layer0_out[5724];
     layer1_out[5634] <= ~(layer0_out[9825] & layer0_out[9826]);
     layer1_out[5635] <= ~layer0_out[11489] | layer0_out[11490];
     layer1_out[5636] <= ~layer0_out[3365];
     layer1_out[5637] <= layer0_out[3149] & ~layer0_out[3148];
     layer1_out[5638] <= ~layer0_out[9097];
     layer1_out[5639] <= layer0_out[7377];
     layer1_out[5640] <= ~(layer0_out[4404] & layer0_out[4405]);
     layer1_out[5641] <= layer0_out[3940] & ~layer0_out[3939];
     layer1_out[5642] <= 1'b1;
     layer1_out[5643] <= ~(layer0_out[9018] & layer0_out[9019]);
     layer1_out[5644] <= layer0_out[5382];
     layer1_out[5645] <= ~layer0_out[4199] | layer0_out[4200];
     layer1_out[5646] <= ~(layer0_out[7842] | layer0_out[7843]);
     layer1_out[5647] <= ~layer0_out[11575] | layer0_out[11574];
     layer1_out[5648] <= layer0_out[4556] & ~layer0_out[4555];
     layer1_out[5649] <= layer0_out[204] & ~layer0_out[205];
     layer1_out[5650] <= ~(layer0_out[6655] & layer0_out[6656]);
     layer1_out[5651] <= layer0_out[3349];
     layer1_out[5652] <= ~layer0_out[9501];
     layer1_out[5653] <= ~layer0_out[7075];
     layer1_out[5654] <= layer0_out[9516];
     layer1_out[5655] <= layer0_out[4278] ^ layer0_out[4279];
     layer1_out[5656] <= 1'b1;
     layer1_out[5657] <= ~(layer0_out[3394] | layer0_out[3395]);
     layer1_out[5658] <= ~layer0_out[902];
     layer1_out[5659] <= ~layer0_out[3534] | layer0_out[3533];
     layer1_out[5660] <= layer0_out[11886] & layer0_out[11887];
     layer1_out[5661] <= ~layer0_out[1267];
     layer1_out[5662] <= 1'b1;
     layer1_out[5663] <= layer0_out[553] & layer0_out[554];
     layer1_out[5664] <= ~layer0_out[7781];
     layer1_out[5665] <= ~layer0_out[93];
     layer1_out[5666] <= layer0_out[5003] & ~layer0_out[5002];
     layer1_out[5667] <= ~(layer0_out[10040] & layer0_out[10041]);
     layer1_out[5668] <= layer0_out[11593] | layer0_out[11594];
     layer1_out[5669] <= ~(layer0_out[3114] | layer0_out[3115]);
     layer1_out[5670] <= 1'b0;
     layer1_out[5671] <= ~layer0_out[6636];
     layer1_out[5672] <= ~layer0_out[4680] | layer0_out[4679];
     layer1_out[5673] <= ~layer0_out[5283] | layer0_out[5284];
     layer1_out[5674] <= layer0_out[4803] & ~layer0_out[4802];
     layer1_out[5675] <= layer0_out[5265];
     layer1_out[5676] <= ~layer0_out[11267] | layer0_out[11268];
     layer1_out[5677] <= layer0_out[708];
     layer1_out[5678] <= layer0_out[8427];
     layer1_out[5679] <= ~layer0_out[11304];
     layer1_out[5680] <= ~layer0_out[9934];
     layer1_out[5681] <= 1'b1;
     layer1_out[5682] <= layer0_out[605] & layer0_out[606];
     layer1_out[5683] <= ~(layer0_out[11370] & layer0_out[11371]);
     layer1_out[5684] <= ~layer0_out[10441] | layer0_out[10440];
     layer1_out[5685] <= layer0_out[2899] ^ layer0_out[2900];
     layer1_out[5686] <= ~(layer0_out[9349] & layer0_out[9350]);
     layer1_out[5687] <= ~layer0_out[8638];
     layer1_out[5688] <= layer0_out[4592] & layer0_out[4593];
     layer1_out[5689] <= layer0_out[207] & layer0_out[208];
     layer1_out[5690] <= layer0_out[2911] & layer0_out[2912];
     layer1_out[5691] <= layer0_out[14] | layer0_out[15];
     layer1_out[5692] <= ~layer0_out[1892] | layer0_out[1891];
     layer1_out[5693] <= ~layer0_out[8721] | layer0_out[8720];
     layer1_out[5694] <= layer0_out[1912] & ~layer0_out[1913];
     layer1_out[5695] <= layer0_out[3152] & ~layer0_out[3153];
     layer1_out[5696] <= ~layer0_out[4577];
     layer1_out[5697] <= layer0_out[4546] & ~layer0_out[4545];
     layer1_out[5698] <= ~layer0_out[8268];
     layer1_out[5699] <= layer0_out[3869] & layer0_out[3870];
     layer1_out[5700] <= layer0_out[6542] ^ layer0_out[6543];
     layer1_out[5701] <= layer0_out[8207];
     layer1_out[5702] <= layer0_out[10832] & ~layer0_out[10831];
     layer1_out[5703] <= layer0_out[3505];
     layer1_out[5704] <= layer0_out[1097] & layer0_out[1098];
     layer1_out[5705] <= ~(layer0_out[1189] ^ layer0_out[1190]);
     layer1_out[5706] <= ~layer0_out[8007];
     layer1_out[5707] <= ~layer0_out[8357] | layer0_out[8356];
     layer1_out[5708] <= layer0_out[6422] & ~layer0_out[6423];
     layer1_out[5709] <= ~(layer0_out[1384] | layer0_out[1385]);
     layer1_out[5710] <= layer0_out[6194];
     layer1_out[5711] <= ~(layer0_out[4767] ^ layer0_out[4768]);
     layer1_out[5712] <= layer0_out[933];
     layer1_out[5713] <= layer0_out[8824] ^ layer0_out[8825];
     layer1_out[5714] <= ~(layer0_out[2654] ^ layer0_out[2655]);
     layer1_out[5715] <= ~layer0_out[5904];
     layer1_out[5716] <= ~layer0_out[2631] | layer0_out[2632];
     layer1_out[5717] <= layer0_out[7431];
     layer1_out[5718] <= layer0_out[2104];
     layer1_out[5719] <= ~layer0_out[869] | layer0_out[868];
     layer1_out[5720] <= layer0_out[10602] ^ layer0_out[10603];
     layer1_out[5721] <= layer0_out[1139] & layer0_out[1140];
     layer1_out[5722] <= ~(layer0_out[1858] | layer0_out[1859]);
     layer1_out[5723] <= 1'b0;
     layer1_out[5724] <= layer0_out[8759];
     layer1_out[5725] <= layer0_out[11330];
     layer1_out[5726] <= ~layer0_out[99] | layer0_out[100];
     layer1_out[5727] <= layer0_out[6691] & ~layer0_out[6690];
     layer1_out[5728] <= ~layer0_out[11748];
     layer1_out[5729] <= layer0_out[6766] | layer0_out[6767];
     layer1_out[5730] <= ~layer0_out[6770] | layer0_out[6771];
     layer1_out[5731] <= ~(layer0_out[4448] & layer0_out[4449]);
     layer1_out[5732] <= ~(layer0_out[6063] ^ layer0_out[6064]);
     layer1_out[5733] <= layer0_out[2084];
     layer1_out[5734] <= ~(layer0_out[2079] & layer0_out[2080]);
     layer1_out[5735] <= 1'b1;
     layer1_out[5736] <= ~layer0_out[6482];
     layer1_out[5737] <= layer0_out[5342];
     layer1_out[5738] <= layer0_out[8832];
     layer1_out[5739] <= layer0_out[6768] & layer0_out[6769];
     layer1_out[5740] <= ~layer0_out[197] | layer0_out[198];
     layer1_out[5741] <= layer0_out[10662];
     layer1_out[5742] <= layer0_out[643] & ~layer0_out[644];
     layer1_out[5743] <= layer0_out[10890] & ~layer0_out[10891];
     layer1_out[5744] <= layer0_out[9461] | layer0_out[9462];
     layer1_out[5745] <= ~layer0_out[1864] | layer0_out[1865];
     layer1_out[5746] <= layer0_out[8404] & ~layer0_out[8405];
     layer1_out[5747] <= ~(layer0_out[11123] & layer0_out[11124]);
     layer1_out[5748] <= ~(layer0_out[6426] & layer0_out[6427]);
     layer1_out[5749] <= layer0_out[9863] ^ layer0_out[9864];
     layer1_out[5750] <= 1'b0;
     layer1_out[5751] <= ~(layer0_out[5713] | layer0_out[5714]);
     layer1_out[5752] <= ~(layer0_out[6343] & layer0_out[6344]);
     layer1_out[5753] <= ~layer0_out[5522];
     layer1_out[5754] <= ~layer0_out[7820];
     layer1_out[5755] <= 1'b1;
     layer1_out[5756] <= ~(layer0_out[4870] | layer0_out[4871]);
     layer1_out[5757] <= ~layer0_out[8549];
     layer1_out[5758] <= ~layer0_out[8829] | layer0_out[8828];
     layer1_out[5759] <= layer0_out[3924] & ~layer0_out[3923];
     layer1_out[5760] <= ~(layer0_out[3204] | layer0_out[3205]);
     layer1_out[5761] <= ~layer0_out[9500] | layer0_out[9499];
     layer1_out[5762] <= layer0_out[2936] & layer0_out[2937];
     layer1_out[5763] <= ~layer0_out[758] | layer0_out[759];
     layer1_out[5764] <= 1'b1;
     layer1_out[5765] <= ~(layer0_out[7548] | layer0_out[7549]);
     layer1_out[5766] <= ~(layer0_out[11298] & layer0_out[11299]);
     layer1_out[5767] <= layer0_out[2268] ^ layer0_out[2269];
     layer1_out[5768] <= 1'b1;
     layer1_out[5769] <= layer0_out[1902] & ~layer0_out[1901];
     layer1_out[5770] <= layer0_out[9276] | layer0_out[9277];
     layer1_out[5771] <= ~layer0_out[8000] | layer0_out[7999];
     layer1_out[5772] <= layer0_out[9791] & ~layer0_out[9792];
     layer1_out[5773] <= ~layer0_out[6597] | layer0_out[6596];
     layer1_out[5774] <= ~layer0_out[1201] | layer0_out[1202];
     layer1_out[5775] <= layer0_out[8700] & ~layer0_out[8699];
     layer1_out[5776] <= layer0_out[9878] & ~layer0_out[9879];
     layer1_out[5777] <= layer0_out[1920];
     layer1_out[5778] <= ~(layer0_out[6531] & layer0_out[6532]);
     layer1_out[5779] <= ~(layer0_out[348] & layer0_out[349]);
     layer1_out[5780] <= 1'b1;
     layer1_out[5781] <= ~(layer0_out[5189] | layer0_out[5190]);
     layer1_out[5782] <= ~(layer0_out[7105] ^ layer0_out[7106]);
     layer1_out[5783] <= layer0_out[1983] & ~layer0_out[1984];
     layer1_out[5784] <= ~layer0_out[6250] | layer0_out[6249];
     layer1_out[5785] <= layer0_out[11377];
     layer1_out[5786] <= ~(layer0_out[3323] ^ layer0_out[3324]);
     layer1_out[5787] <= layer0_out[3104] & layer0_out[3105];
     layer1_out[5788] <= layer0_out[1281] & ~layer0_out[1280];
     layer1_out[5789] <= layer0_out[2393] & ~layer0_out[2392];
     layer1_out[5790] <= ~layer0_out[6859] | layer0_out[6860];
     layer1_out[5791] <= layer0_out[7484];
     layer1_out[5792] <= layer0_out[1332] & ~layer0_out[1333];
     layer1_out[5793] <= ~(layer0_out[7917] ^ layer0_out[7918]);
     layer1_out[5794] <= ~(layer0_out[4580] & layer0_out[4581]);
     layer1_out[5795] <= ~layer0_out[4450];
     layer1_out[5796] <= ~(layer0_out[9667] | layer0_out[9668]);
     layer1_out[5797] <= 1'b0;
     layer1_out[5798] <= ~(layer0_out[9424] & layer0_out[9425]);
     layer1_out[5799] <= ~layer0_out[5517] | layer0_out[5516];
     layer1_out[5800] <= ~layer0_out[5458];
     layer1_out[5801] <= layer0_out[4422];
     layer1_out[5802] <= ~layer0_out[3191];
     layer1_out[5803] <= ~layer0_out[11319];
     layer1_out[5804] <= ~layer0_out[3917];
     layer1_out[5805] <= layer0_out[3671] & ~layer0_out[3670];
     layer1_out[5806] <= ~layer0_out[7705] | layer0_out[7704];
     layer1_out[5807] <= ~layer0_out[10968] | layer0_out[10969];
     layer1_out[5808] <= layer0_out[11141] & ~layer0_out[11142];
     layer1_out[5809] <= ~(layer0_out[1388] ^ layer0_out[1389]);
     layer1_out[5810] <= 1'b0;
     layer1_out[5811] <= layer0_out[7592];
     layer1_out[5812] <= layer0_out[1167] & layer0_out[1168];
     layer1_out[5813] <= layer0_out[9390] & layer0_out[9391];
     layer1_out[5814] <= ~layer0_out[6780];
     layer1_out[5815] <= ~layer0_out[963];
     layer1_out[5816] <= layer0_out[7140] ^ layer0_out[7141];
     layer1_out[5817] <= layer0_out[9420] & layer0_out[9421];
     layer1_out[5818] <= ~(layer0_out[11373] & layer0_out[11374]);
     layer1_out[5819] <= ~(layer0_out[4118] | layer0_out[4119]);
     layer1_out[5820] <= ~layer0_out[8726] | layer0_out[8727];
     layer1_out[5821] <= layer0_out[6623] | layer0_out[6624];
     layer1_out[5822] <= ~layer0_out[11113];
     layer1_out[5823] <= ~layer0_out[3389];
     layer1_out[5824] <= 1'b1;
     layer1_out[5825] <= layer0_out[5011];
     layer1_out[5826] <= ~layer0_out[8543] | layer0_out[8542];
     layer1_out[5827] <= ~layer0_out[9600];
     layer1_out[5828] <= layer0_out[10822] | layer0_out[10823];
     layer1_out[5829] <= ~layer0_out[11718] | layer0_out[11719];
     layer1_out[5830] <= 1'b1;
     layer1_out[5831] <= layer0_out[11326] & layer0_out[11327];
     layer1_out[5832] <= ~(layer0_out[3446] | layer0_out[3447]);
     layer1_out[5833] <= ~(layer0_out[9786] & layer0_out[9787]);
     layer1_out[5834] <= ~(layer0_out[507] & layer0_out[508]);
     layer1_out[5835] <= ~layer0_out[2972];
     layer1_out[5836] <= layer0_out[7254] | layer0_out[7255];
     layer1_out[5837] <= ~(layer0_out[10837] & layer0_out[10838]);
     layer1_out[5838] <= layer0_out[3611] & ~layer0_out[3612];
     layer1_out[5839] <= ~(layer0_out[5212] & layer0_out[5213]);
     layer1_out[5840] <= ~(layer0_out[852] | layer0_out[853]);
     layer1_out[5841] <= layer0_out[3619];
     layer1_out[5842] <= 1'b1;
     layer1_out[5843] <= ~layer0_out[1747] | layer0_out[1748];
     layer1_out[5844] <= layer0_out[9073] & layer0_out[9074];
     layer1_out[5845] <= ~layer0_out[5295] | layer0_out[5296];
     layer1_out[5846] <= layer0_out[10476] & ~layer0_out[10477];
     layer1_out[5847] <= ~layer0_out[10476] | layer0_out[10475];
     layer1_out[5848] <= layer0_out[2648] & layer0_out[2649];
     layer1_out[5849] <= ~layer0_out[4276] | layer0_out[4275];
     layer1_out[5850] <= ~(layer0_out[1899] | layer0_out[1900]);
     layer1_out[5851] <= layer0_out[10392] & layer0_out[10393];
     layer1_out[5852] <= layer0_out[11206];
     layer1_out[5853] <= layer0_out[3641] & layer0_out[3642];
     layer1_out[5854] <= ~layer0_out[10195];
     layer1_out[5855] <= layer0_out[10081];
     layer1_out[5856] <= ~layer0_out[9733] | layer0_out[9734];
     layer1_out[5857] <= ~layer0_out[6612];
     layer1_out[5858] <= ~layer0_out[11598];
     layer1_out[5859] <= ~(layer0_out[6718] & layer0_out[6719]);
     layer1_out[5860] <= ~layer0_out[4987];
     layer1_out[5861] <= layer0_out[1871] & layer0_out[1872];
     layer1_out[5862] <= ~layer0_out[8894] | layer0_out[8895];
     layer1_out[5863] <= layer0_out[7008] & layer0_out[7009];
     layer1_out[5864] <= layer0_out[4193] ^ layer0_out[4194];
     layer1_out[5865] <= layer0_out[11090] ^ layer0_out[11091];
     layer1_out[5866] <= 1'b1;
     layer1_out[5867] <= layer0_out[10578] & ~layer0_out[10577];
     layer1_out[5868] <= ~layer0_out[11231];
     layer1_out[5869] <= ~layer0_out[392];
     layer1_out[5870] <= ~layer0_out[11348] | layer0_out[11347];
     layer1_out[5871] <= layer0_out[885];
     layer1_out[5872] <= layer0_out[10196] | layer0_out[10197];
     layer1_out[5873] <= ~(layer0_out[9211] ^ layer0_out[9212]);
     layer1_out[5874] <= ~layer0_out[11781];
     layer1_out[5875] <= layer0_out[8] | layer0_out[9];
     layer1_out[5876] <= ~layer0_out[6381] | layer0_out[6382];
     layer1_out[5877] <= ~layer0_out[1571] | layer0_out[1572];
     layer1_out[5878] <= ~layer0_out[5085];
     layer1_out[5879] <= layer0_out[8097] | layer0_out[8098];
     layer1_out[5880] <= layer0_out[2610];
     layer1_out[5881] <= ~(layer0_out[10783] & layer0_out[10784]);
     layer1_out[5882] <= ~(layer0_out[4527] ^ layer0_out[4528]);
     layer1_out[5883] <= 1'b0;
     layer1_out[5884] <= layer0_out[9934] & ~layer0_out[9935];
     layer1_out[5885] <= layer0_out[7230];
     layer1_out[5886] <= ~(layer0_out[7497] | layer0_out[7498]);
     layer1_out[5887] <= ~layer0_out[565];
     layer1_out[5888] <= layer0_out[7701] & layer0_out[7702];
     layer1_out[5889] <= layer0_out[898] & ~layer0_out[897];
     layer1_out[5890] <= ~layer0_out[5161];
     layer1_out[5891] <= ~layer0_out[9444] | layer0_out[9443];
     layer1_out[5892] <= layer0_out[590];
     layer1_out[5893] <= layer0_out[11852] ^ layer0_out[11853];
     layer1_out[5894] <= layer0_out[11277] & ~layer0_out[11276];
     layer1_out[5895] <= layer0_out[761] | layer0_out[762];
     layer1_out[5896] <= layer0_out[885];
     layer1_out[5897] <= ~(layer0_out[8384] & layer0_out[8385]);
     layer1_out[5898] <= ~layer0_out[2446];
     layer1_out[5899] <= ~layer0_out[945];
     layer1_out[5900] <= ~(layer0_out[870] & layer0_out[871]);
     layer1_out[5901] <= ~(layer0_out[5203] | layer0_out[5204]);
     layer1_out[5902] <= 1'b1;
     layer1_out[5903] <= layer0_out[5941];
     layer1_out[5904] <= ~(layer0_out[4316] | layer0_out[4317]);
     layer1_out[5905] <= ~layer0_out[625];
     layer1_out[5906] <= ~layer0_out[4908];
     layer1_out[5907] <= layer0_out[10410] ^ layer0_out[10411];
     layer1_out[5908] <= layer0_out[5532] & ~layer0_out[5533];
     layer1_out[5909] <= ~layer0_out[8935] | layer0_out[8936];
     layer1_out[5910] <= ~layer0_out[4490];
     layer1_out[5911] <= ~layer0_out[10997] | layer0_out[10996];
     layer1_out[5912] <= ~layer0_out[2766];
     layer1_out[5913] <= ~layer0_out[1088] | layer0_out[1089];
     layer1_out[5914] <= layer0_out[6187];
     layer1_out[5915] <= ~layer0_out[11792] | layer0_out[11791];
     layer1_out[5916] <= 1'b0;
     layer1_out[5917] <= layer0_out[7860];
     layer1_out[5918] <= layer0_out[3385] ^ layer0_out[3386];
     layer1_out[5919] <= ~layer0_out[1721] | layer0_out[1720];
     layer1_out[5920] <= layer0_out[2021] | layer0_out[2022];
     layer1_out[5921] <= layer0_out[11482];
     layer1_out[5922] <= ~layer0_out[9061] | layer0_out[9060];
     layer1_out[5923] <= ~layer0_out[8437];
     layer1_out[5924] <= ~layer0_out[2011] | layer0_out[2010];
     layer1_out[5925] <= 1'b1;
     layer1_out[5926] <= 1'b0;
     layer1_out[5927] <= ~layer0_out[6223];
     layer1_out[5928] <= ~layer0_out[10783];
     layer1_out[5929] <= ~layer0_out[9508];
     layer1_out[5930] <= layer0_out[1164] & layer0_out[1165];
     layer1_out[5931] <= layer0_out[1270] & ~layer0_out[1269];
     layer1_out[5932] <= layer0_out[454] & ~layer0_out[453];
     layer1_out[5933] <= layer0_out[7486] | layer0_out[7487];
     layer1_out[5934] <= ~(layer0_out[3387] | layer0_out[3388]);
     layer1_out[5935] <= ~layer0_out[400];
     layer1_out[5936] <= layer0_out[5994] & ~layer0_out[5993];
     layer1_out[5937] <= ~layer0_out[2484];
     layer1_out[5938] <= ~layer0_out[448] | layer0_out[449];
     layer1_out[5939] <= ~layer0_out[7096] | layer0_out[7095];
     layer1_out[5940] <= layer0_out[2036];
     layer1_out[5941] <= ~layer0_out[10998];
     layer1_out[5942] <= layer0_out[943] & ~layer0_out[944];
     layer1_out[5943] <= layer0_out[2818];
     layer1_out[5944] <= ~layer0_out[11373] | layer0_out[11372];
     layer1_out[5945] <= layer0_out[2965] ^ layer0_out[2966];
     layer1_out[5946] <= layer0_out[2608];
     layer1_out[5947] <= ~layer0_out[2071];
     layer1_out[5948] <= layer0_out[78] & ~layer0_out[77];
     layer1_out[5949] <= ~layer0_out[4300] | layer0_out[4299];
     layer1_out[5950] <= layer0_out[2286];
     layer1_out[5951] <= layer0_out[9310] ^ layer0_out[9311];
     layer1_out[5952] <= ~layer0_out[3901];
     layer1_out[5953] <= ~layer0_out[4561];
     layer1_out[5954] <= layer0_out[2291] & ~layer0_out[2290];
     layer1_out[5955] <= layer0_out[7017];
     layer1_out[5956] <= layer0_out[11070] & ~layer0_out[11069];
     layer1_out[5957] <= layer0_out[6262];
     layer1_out[5958] <= layer0_out[1130] & ~layer0_out[1131];
     layer1_out[5959] <= ~(layer0_out[10861] | layer0_out[10862]);
     layer1_out[5960] <= layer0_out[2226] & ~layer0_out[2225];
     layer1_out[5961] <= layer0_out[5209];
     layer1_out[5962] <= 1'b0;
     layer1_out[5963] <= layer0_out[8820] | layer0_out[8821];
     layer1_out[5964] <= layer0_out[10795] & layer0_out[10796];
     layer1_out[5965] <= ~layer0_out[4548];
     layer1_out[5966] <= ~layer0_out[2004];
     layer1_out[5967] <= ~layer0_out[1652] | layer0_out[1653];
     layer1_out[5968] <= ~layer0_out[6764] | layer0_out[6763];
     layer1_out[5969] <= layer0_out[2510] & layer0_out[2511];
     layer1_out[5970] <= layer0_out[9089] & ~layer0_out[9088];
     layer1_out[5971] <= layer0_out[8431] & ~layer0_out[8430];
     layer1_out[5972] <= 1'b1;
     layer1_out[5973] <= layer0_out[3390];
     layer1_out[5974] <= ~layer0_out[9311] | layer0_out[9312];
     layer1_out[5975] <= ~layer0_out[2369];
     layer1_out[5976] <= ~(layer0_out[7126] & layer0_out[7127]);
     layer1_out[5977] <= ~layer0_out[7768] | layer0_out[7769];
     layer1_out[5978] <= ~layer0_out[749];
     layer1_out[5979] <= ~(layer0_out[10878] | layer0_out[10879]);
     layer1_out[5980] <= ~(layer0_out[7777] ^ layer0_out[7778]);
     layer1_out[5981] <= ~(layer0_out[1038] | layer0_out[1039]);
     layer1_out[5982] <= ~(layer0_out[9169] | layer0_out[9170]);
     layer1_out[5983] <= ~(layer0_out[8516] & layer0_out[8517]);
     layer1_out[5984] <= layer0_out[9139];
     layer1_out[5985] <= layer0_out[5448];
     layer1_out[5986] <= ~(layer0_out[8026] | layer0_out[8027]);
     layer1_out[5987] <= ~layer0_out[1179];
     layer1_out[5988] <= layer0_out[5611] & ~layer0_out[5610];
     layer1_out[5989] <= ~(layer0_out[10586] | layer0_out[10587]);
     layer1_out[5990] <= 1'b0;
     layer1_out[5991] <= layer0_out[10253];
     layer1_out[5992] <= ~(layer0_out[9816] ^ layer0_out[9817]);
     layer1_out[5993] <= layer0_out[8186];
     layer1_out[5994] <= layer0_out[722] & layer0_out[723];
     layer1_out[5995] <= ~layer0_out[9926];
     layer1_out[5996] <= layer0_out[5724] & ~layer0_out[5723];
     layer1_out[5997] <= layer0_out[7174] & ~layer0_out[7175];
     layer1_out[5998] <= layer0_out[8124] & ~layer0_out[8125];
     layer1_out[5999] <= ~layer0_out[7457];
     layer1_out[6000] <= ~layer0_out[10060];
     layer1_out[6001] <= ~(layer0_out[7540] & layer0_out[7541]);
     layer1_out[6002] <= layer0_out[4465];
     layer1_out[6003] <= layer0_out[7292] & ~layer0_out[7293];
     layer1_out[6004] <= layer0_out[9474] & ~layer0_out[9475];
     layer1_out[6005] <= layer0_out[10645] ^ layer0_out[10646];
     layer1_out[6006] <= layer0_out[8459] | layer0_out[8460];
     layer1_out[6007] <= ~(layer0_out[5567] & layer0_out[5568]);
     layer1_out[6008] <= layer0_out[1183] & ~layer0_out[1184];
     layer1_out[6009] <= layer0_out[11125] | layer0_out[11126];
     layer1_out[6010] <= ~layer0_out[153];
     layer1_out[6011] <= ~(layer0_out[10323] ^ layer0_out[10324]);
     layer1_out[6012] <= layer0_out[2217];
     layer1_out[6013] <= layer0_out[1363];
     layer1_out[6014] <= ~layer0_out[4698] | layer0_out[4697];
     layer1_out[6015] <= ~layer0_out[9179];
     layer1_out[6016] <= ~layer0_out[7252] | layer0_out[7251];
     layer1_out[6017] <= ~layer0_out[75];
     layer1_out[6018] <= layer0_out[3992] & ~layer0_out[3993];
     layer1_out[6019] <= ~(layer0_out[6268] & layer0_out[6269]);
     layer1_out[6020] <= layer0_out[6822] & ~layer0_out[6821];
     layer1_out[6021] <= ~layer0_out[4899];
     layer1_out[6022] <= ~(layer0_out[750] | layer0_out[751]);
     layer1_out[6023] <= layer0_out[9437];
     layer1_out[6024] <= ~layer0_out[10326];
     layer1_out[6025] <= layer0_out[3475];
     layer1_out[6026] <= layer0_out[3086];
     layer1_out[6027] <= ~layer0_out[4554] | layer0_out[4553];
     layer1_out[6028] <= layer0_out[2827] & ~layer0_out[2826];
     layer1_out[6029] <= layer0_out[4234] & ~layer0_out[4235];
     layer1_out[6030] <= ~layer0_out[3642];
     layer1_out[6031] <= ~layer0_out[5242] | layer0_out[5243];
     layer1_out[6032] <= ~(layer0_out[6987] & layer0_out[6988]);
     layer1_out[6033] <= ~(layer0_out[1361] & layer0_out[1362]);
     layer1_out[6034] <= ~layer0_out[5441];
     layer1_out[6035] <= ~(layer0_out[1878] | layer0_out[1879]);
     layer1_out[6036] <= ~layer0_out[1529] | layer0_out[1528];
     layer1_out[6037] <= layer0_out[9292];
     layer1_out[6038] <= ~(layer0_out[2874] & layer0_out[2875]);
     layer1_out[6039] <= layer0_out[1577] | layer0_out[1578];
     layer1_out[6040] <= ~layer0_out[8685];
     layer1_out[6041] <= layer0_out[2193] & ~layer0_out[2194];
     layer1_out[6042] <= ~(layer0_out[8245] | layer0_out[8246]);
     layer1_out[6043] <= ~(layer0_out[2086] | layer0_out[2087]);
     layer1_out[6044] <= layer0_out[6042] & ~layer0_out[6043];
     layer1_out[6045] <= ~layer0_out[11625] | layer0_out[11624];
     layer1_out[6046] <= layer0_out[2508] & layer0_out[2509];
     layer1_out[6047] <= ~layer0_out[2731];
     layer1_out[6048] <= ~layer0_out[1062];
     layer1_out[6049] <= ~layer0_out[3701] | layer0_out[3702];
     layer1_out[6050] <= ~layer0_out[5671];
     layer1_out[6051] <= ~layer0_out[5553] | layer0_out[5552];
     layer1_out[6052] <= layer0_out[8877] ^ layer0_out[8878];
     layer1_out[6053] <= layer0_out[2475] & layer0_out[2476];
     layer1_out[6054] <= ~layer0_out[72];
     layer1_out[6055] <= ~(layer0_out[3926] ^ layer0_out[3927]);
     layer1_out[6056] <= ~layer0_out[2555];
     layer1_out[6057] <= ~(layer0_out[3740] & layer0_out[3741]);
     layer1_out[6058] <= ~layer0_out[1636];
     layer1_out[6059] <= layer0_out[3440] | layer0_out[3441];
     layer1_out[6060] <= layer0_out[7266];
     layer1_out[6061] <= ~layer0_out[7806] | layer0_out[7807];
     layer1_out[6062] <= ~layer0_out[1716];
     layer1_out[6063] <= layer0_out[11039];
     layer1_out[6064] <= layer0_out[8891] | layer0_out[8892];
     layer1_out[6065] <= ~layer0_out[7573];
     layer1_out[6066] <= ~layer0_out[5969] | layer0_out[5970];
     layer1_out[6067] <= layer0_out[11133] | layer0_out[11134];
     layer1_out[6068] <= ~layer0_out[2752];
     layer1_out[6069] <= layer0_out[8698];
     layer1_out[6070] <= layer0_out[7612] & ~layer0_out[7611];
     layer1_out[6071] <= layer0_out[794];
     layer1_out[6072] <= ~layer0_out[2044] | layer0_out[2043];
     layer1_out[6073] <= layer0_out[1751] & ~layer0_out[1752];
     layer1_out[6074] <= layer0_out[9108];
     layer1_out[6075] <= layer0_out[8156] | layer0_out[8157];
     layer1_out[6076] <= ~layer0_out[2500];
     layer1_out[6077] <= layer0_out[2065];
     layer1_out[6078] <= layer0_out[6507] & layer0_out[6508];
     layer1_out[6079] <= layer0_out[2449] & layer0_out[2450];
     layer1_out[6080] <= ~(layer0_out[4615] ^ layer0_out[4616]);
     layer1_out[6081] <= layer0_out[4634] & ~layer0_out[4635];
     layer1_out[6082] <= layer0_out[6991] & layer0_out[6992];
     layer1_out[6083] <= ~layer0_out[2025];
     layer1_out[6084] <= ~layer0_out[10248] | layer0_out[10249];
     layer1_out[6085] <= layer0_out[10722] & ~layer0_out[10721];
     layer1_out[6086] <= layer0_out[11227] & ~layer0_out[11228];
     layer1_out[6087] <= layer0_out[634] & layer0_out[635];
     layer1_out[6088] <= layer0_out[2630];
     layer1_out[6089] <= ~layer0_out[5469] | layer0_out[5470];
     layer1_out[6090] <= ~layer0_out[2432] | layer0_out[2431];
     layer1_out[6091] <= layer0_out[11650];
     layer1_out[6092] <= ~layer0_out[5586];
     layer1_out[6093] <= layer0_out[2543] & layer0_out[2544];
     layer1_out[6094] <= ~layer0_out[3795] | layer0_out[3794];
     layer1_out[6095] <= 1'b1;
     layer1_out[6096] <= ~layer0_out[8286] | layer0_out[8287];
     layer1_out[6097] <= layer0_out[1309];
     layer1_out[6098] <= layer0_out[749];
     layer1_out[6099] <= layer0_out[11770];
     layer1_out[6100] <= ~layer0_out[4698] | layer0_out[4699];
     layer1_out[6101] <= layer0_out[4658] & ~layer0_out[4657];
     layer1_out[6102] <= layer0_out[7523] & ~layer0_out[7524];
     layer1_out[6103] <= layer0_out[9802];
     layer1_out[6104] <= ~(layer0_out[4620] | layer0_out[4621]);
     layer1_out[6105] <= layer0_out[11343];
     layer1_out[6106] <= layer0_out[7424];
     layer1_out[6107] <= layer0_out[7067] & ~layer0_out[7066];
     layer1_out[6108] <= layer0_out[6466];
     layer1_out[6109] <= layer0_out[3085];
     layer1_out[6110] <= ~(layer0_out[976] & layer0_out[977]);
     layer1_out[6111] <= layer0_out[10267] & layer0_out[10268];
     layer1_out[6112] <= ~layer0_out[5726] | layer0_out[5725];
     layer1_out[6113] <= ~layer0_out[10854] | layer0_out[10855];
     layer1_out[6114] <= layer0_out[7874] & layer0_out[7875];
     layer1_out[6115] <= ~layer0_out[4962] | layer0_out[4963];
     layer1_out[6116] <= ~layer0_out[7919];
     layer1_out[6117] <= ~layer0_out[3115];
     layer1_out[6118] <= layer0_out[8753];
     layer1_out[6119] <= layer0_out[11766] & ~layer0_out[11767];
     layer1_out[6120] <= layer0_out[5946] ^ layer0_out[5947];
     layer1_out[6121] <= layer0_out[11105] & ~layer0_out[11104];
     layer1_out[6122] <= ~layer0_out[1581] | layer0_out[1580];
     layer1_out[6123] <= ~layer0_out[3324];
     layer1_out[6124] <= layer0_out[5117] & layer0_out[5118];
     layer1_out[6125] <= layer0_out[1142] & ~layer0_out[1143];
     layer1_out[6126] <= ~(layer0_out[8224] | layer0_out[8225]);
     layer1_out[6127] <= layer0_out[4921] | layer0_out[4922];
     layer1_out[6128] <= ~layer0_out[10499] | layer0_out[10500];
     layer1_out[6129] <= layer0_out[3560] & ~layer0_out[3559];
     layer1_out[6130] <= ~(layer0_out[10720] ^ layer0_out[10721]);
     layer1_out[6131] <= ~(layer0_out[3142] ^ layer0_out[3143]);
     layer1_out[6132] <= ~(layer0_out[2657] | layer0_out[2658]);
     layer1_out[6133] <= layer0_out[1549] & ~layer0_out[1548];
     layer1_out[6134] <= ~(layer0_out[9452] | layer0_out[9453]);
     layer1_out[6135] <= ~(layer0_out[3552] & layer0_out[3553]);
     layer1_out[6136] <= layer0_out[10745] & ~layer0_out[10746];
     layer1_out[6137] <= layer0_out[455];
     layer1_out[6138] <= layer0_out[3788] & ~layer0_out[3787];
     layer1_out[6139] <= layer0_out[1042] & layer0_out[1043];
     layer1_out[6140] <= layer0_out[9205] | layer0_out[9206];
     layer1_out[6141] <= layer0_out[6997] & layer0_out[6998];
     layer1_out[6142] <= layer0_out[1091] & ~layer0_out[1090];
     layer1_out[6143] <= 1'b0;
     layer1_out[6144] <= layer0_out[8525] | layer0_out[8526];
     layer1_out[6145] <= layer0_out[7215] | layer0_out[7216];
     layer1_out[6146] <= layer0_out[5780];
     layer1_out[6147] <= layer0_out[10507] & ~layer0_out[10508];
     layer1_out[6148] <= 1'b0;
     layer1_out[6149] <= ~(layer0_out[6155] | layer0_out[6156]);
     layer1_out[6150] <= layer0_out[10481] | layer0_out[10482];
     layer1_out[6151] <= layer0_out[7764];
     layer1_out[6152] <= layer0_out[8022];
     layer1_out[6153] <= layer0_out[247] & ~layer0_out[246];
     layer1_out[6154] <= layer0_out[3170] | layer0_out[3171];
     layer1_out[6155] <= layer0_out[7516] | layer0_out[7517];
     layer1_out[6156] <= layer0_out[7662];
     layer1_out[6157] <= layer0_out[8723] & ~layer0_out[8722];
     layer1_out[6158] <= layer0_out[2712] & ~layer0_out[2711];
     layer1_out[6159] <= ~layer0_out[10388];
     layer1_out[6160] <= layer0_out[7883] ^ layer0_out[7884];
     layer1_out[6161] <= layer0_out[10986];
     layer1_out[6162] <= ~layer0_out[4883] | layer0_out[4882];
     layer1_out[6163] <= ~layer0_out[6901];
     layer1_out[6164] <= ~layer0_out[4055] | layer0_out[4056];
     layer1_out[6165] <= ~layer0_out[10227];
     layer1_out[6166] <= layer0_out[5845];
     layer1_out[6167] <= layer0_out[8926] & ~layer0_out[8927];
     layer1_out[6168] <= ~(layer0_out[6703] ^ layer0_out[6704]);
     layer1_out[6169] <= layer0_out[11068] | layer0_out[11069];
     layer1_out[6170] <= layer0_out[5357] & layer0_out[5358];
     layer1_out[6171] <= 1'b0;
     layer1_out[6172] <= ~(layer0_out[8153] ^ layer0_out[8154]);
     layer1_out[6173] <= ~layer0_out[2452] | layer0_out[2451];
     layer1_out[6174] <= ~layer0_out[2988];
     layer1_out[6175] <= ~layer0_out[10754];
     layer1_out[6176] <= layer0_out[3948] | layer0_out[3949];
     layer1_out[6177] <= ~layer0_out[9958];
     layer1_out[6178] <= layer0_out[2954] ^ layer0_out[2955];
     layer1_out[6179] <= ~layer0_out[8396];
     layer1_out[6180] <= layer0_out[8696] & layer0_out[8697];
     layer1_out[6181] <= layer0_out[765];
     layer1_out[6182] <= ~(layer0_out[1582] ^ layer0_out[1583]);
     layer1_out[6183] <= ~layer0_out[11017];
     layer1_out[6184] <= layer0_out[10042];
     layer1_out[6185] <= ~layer0_out[7359];
     layer1_out[6186] <= ~(layer0_out[5811] ^ layer0_out[5812]);
     layer1_out[6187] <= layer0_out[1656] & ~layer0_out[1655];
     layer1_out[6188] <= ~layer0_out[3117] | layer0_out[3116];
     layer1_out[6189] <= ~layer0_out[3036];
     layer1_out[6190] <= layer0_out[1727] & ~layer0_out[1728];
     layer1_out[6191] <= ~layer0_out[7312];
     layer1_out[6192] <= layer0_out[10446] & layer0_out[10447];
     layer1_out[6193] <= ~(layer0_out[11753] & layer0_out[11754]);
     layer1_out[6194] <= ~layer0_out[8283] | layer0_out[8284];
     layer1_out[6195] <= ~(layer0_out[148] | layer0_out[149]);
     layer1_out[6196] <= ~layer0_out[10205];
     layer1_out[6197] <= layer0_out[5564] & layer0_out[5565];
     layer1_out[6198] <= ~(layer0_out[11669] & layer0_out[11670]);
     layer1_out[6199] <= ~(layer0_out[11811] | layer0_out[11812]);
     layer1_out[6200] <= layer0_out[10285] | layer0_out[10286];
     layer1_out[6201] <= layer0_out[8003] | layer0_out[8004];
     layer1_out[6202] <= ~(layer0_out[9517] & layer0_out[9518]);
     layer1_out[6203] <= layer0_out[6235];
     layer1_out[6204] <= ~(layer0_out[8716] ^ layer0_out[8717]);
     layer1_out[6205] <= layer0_out[11333] & ~layer0_out[11334];
     layer1_out[6206] <= layer0_out[401];
     layer1_out[6207] <= ~(layer0_out[4160] | layer0_out[4161]);
     layer1_out[6208] <= ~layer0_out[8336];
     layer1_out[6209] <= ~(layer0_out[5202] | layer0_out[5203]);
     layer1_out[6210] <= ~layer0_out[9995];
     layer1_out[6211] <= ~layer0_out[1471];
     layer1_out[6212] <= layer0_out[4976];
     layer1_out[6213] <= 1'b1;
     layer1_out[6214] <= layer0_out[7847];
     layer1_out[6215] <= layer0_out[27];
     layer1_out[6216] <= 1'b0;
     layer1_out[6217] <= ~(layer0_out[3817] & layer0_out[3818]);
     layer1_out[6218] <= layer0_out[10658] & layer0_out[10659];
     layer1_out[6219] <= layer0_out[2255] & ~layer0_out[2254];
     layer1_out[6220] <= ~layer0_out[6211];
     layer1_out[6221] <= ~layer0_out[4586] | layer0_out[4585];
     layer1_out[6222] <= layer0_out[2647] & layer0_out[2648];
     layer1_out[6223] <= ~layer0_out[2804] | layer0_out[2803];
     layer1_out[6224] <= ~(layer0_out[10888] | layer0_out[10889]);
     layer1_out[6225] <= layer0_out[6826] & layer0_out[6827];
     layer1_out[6226] <= layer0_out[8578];
     layer1_out[6227] <= ~layer0_out[1295];
     layer1_out[6228] <= layer0_out[9889];
     layer1_out[6229] <= ~layer0_out[2122] | layer0_out[2123];
     layer1_out[6230] <= ~layer0_out[836];
     layer1_out[6231] <= ~layer0_out[5538];
     layer1_out[6232] <= ~layer0_out[10581];
     layer1_out[6233] <= layer0_out[4468] & ~layer0_out[4469];
     layer1_out[6234] <= ~(layer0_out[7319] & layer0_out[7320]);
     layer1_out[6235] <= layer0_out[9821] & ~layer0_out[9820];
     layer1_out[6236] <= ~layer0_out[11308] | layer0_out[11309];
     layer1_out[6237] <= layer0_out[2869] & ~layer0_out[2870];
     layer1_out[6238] <= layer0_out[11376];
     layer1_out[6239] <= layer0_out[5148] ^ layer0_out[5149];
     layer1_out[6240] <= ~layer0_out[563] | layer0_out[564];
     layer1_out[6241] <= ~(layer0_out[5781] | layer0_out[5782]);
     layer1_out[6242] <= layer0_out[4349] & ~layer0_out[4348];
     layer1_out[6243] <= ~(layer0_out[8195] | layer0_out[8196]);
     layer1_out[6244] <= ~(layer0_out[6016] ^ layer0_out[6017]);
     layer1_out[6245] <= layer0_out[9423] & ~layer0_out[9424];
     layer1_out[6246] <= ~layer0_out[9352] | layer0_out[9353];
     layer1_out[6247] <= ~layer0_out[10710];
     layer1_out[6248] <= ~(layer0_out[11621] | layer0_out[11622]);
     layer1_out[6249] <= layer0_out[2270] & ~layer0_out[2271];
     layer1_out[6250] <= layer0_out[1075] & ~layer0_out[1074];
     layer1_out[6251] <= ~(layer0_out[4685] | layer0_out[4686]);
     layer1_out[6252] <= ~(layer0_out[11825] | layer0_out[11826]);
     layer1_out[6253] <= layer0_out[3646];
     layer1_out[6254] <= layer0_out[6241];
     layer1_out[6255] <= layer0_out[4311] | layer0_out[4312];
     layer1_out[6256] <= layer0_out[4424];
     layer1_out[6257] <= ~(layer0_out[4501] & layer0_out[4502]);
     layer1_out[6258] <= ~(layer0_out[7810] | layer0_out[7811]);
     layer1_out[6259] <= 1'b1;
     layer1_out[6260] <= ~(layer0_out[465] ^ layer0_out[466]);
     layer1_out[6261] <= layer0_out[7720];
     layer1_out[6262] <= ~(layer0_out[6239] ^ layer0_out[6240]);
     layer1_out[6263] <= layer0_out[6998];
     layer1_out[6264] <= layer0_out[2741];
     layer1_out[6265] <= ~layer0_out[10848];
     layer1_out[6266] <= layer0_out[1096];
     layer1_out[6267] <= ~(layer0_out[2359] & layer0_out[2360]);
     layer1_out[6268] <= layer0_out[671] | layer0_out[672];
     layer1_out[6269] <= layer0_out[6298] & ~layer0_out[6299];
     layer1_out[6270] <= ~(layer0_out[373] ^ layer0_out[374]);
     layer1_out[6271] <= ~layer0_out[5539];
     layer1_out[6272] <= layer0_out[11145];
     layer1_out[6273] <= layer0_out[10653] & ~layer0_out[10652];
     layer1_out[6274] <= ~(layer0_out[9137] ^ layer0_out[9138]);
     layer1_out[6275] <= ~layer0_out[7652] | layer0_out[7651];
     layer1_out[6276] <= layer0_out[4416] ^ layer0_out[4417];
     layer1_out[6277] <= layer0_out[8676];
     layer1_out[6278] <= 1'b1;
     layer1_out[6279] <= ~(layer0_out[9969] ^ layer0_out[9970]);
     layer1_out[6280] <= layer0_out[1644] & ~layer0_out[1645];
     layer1_out[6281] <= ~(layer0_out[2879] | layer0_out[2880]);
     layer1_out[6282] <= layer0_out[3795];
     layer1_out[6283] <= 1'b0;
     layer1_out[6284] <= ~layer0_out[8268] | layer0_out[8267];
     layer1_out[6285] <= ~(layer0_out[9184] & layer0_out[9185]);
     layer1_out[6286] <= layer0_out[7351] ^ layer0_out[7352];
     layer1_out[6287] <= ~(layer0_out[11680] & layer0_out[11681]);
     layer1_out[6288] <= ~layer0_out[11724];
     layer1_out[6289] <= layer0_out[4567];
     layer1_out[6290] <= layer0_out[8999] | layer0_out[9000];
     layer1_out[6291] <= layer0_out[4011];
     layer1_out[6292] <= ~layer0_out[5918];
     layer1_out[6293] <= layer0_out[7562] & layer0_out[7563];
     layer1_out[6294] <= layer0_out[3768] | layer0_out[3769];
     layer1_out[6295] <= ~layer0_out[2261];
     layer1_out[6296] <= ~layer0_out[3426];
     layer1_out[6297] <= layer0_out[3494] ^ layer0_out[3495];
     layer1_out[6298] <= layer0_out[5645];
     layer1_out[6299] <= ~layer0_out[9195];
     layer1_out[6300] <= ~layer0_out[4710] | layer0_out[4709];
     layer1_out[6301] <= layer0_out[3555];
     layer1_out[6302] <= layer0_out[11576];
     layer1_out[6303] <= layer0_out[8669] & layer0_out[8670];
     layer1_out[6304] <= layer0_out[5159] | layer0_out[5160];
     layer1_out[6305] <= ~layer0_out[9942];
     layer1_out[6306] <= ~layer0_out[9370];
     layer1_out[6307] <= layer0_out[7772] | layer0_out[7773];
     layer1_out[6308] <= ~layer0_out[3756];
     layer1_out[6309] <= layer0_out[9370] | layer0_out[9371];
     layer1_out[6310] <= layer0_out[5616];
     layer1_out[6311] <= layer0_out[6978] | layer0_out[6979];
     layer1_out[6312] <= layer0_out[196] & ~layer0_out[195];
     layer1_out[6313] <= ~layer0_out[4969];
     layer1_out[6314] <= ~layer0_out[790];
     layer1_out[6315] <= layer0_out[7796] & ~layer0_out[7795];
     layer1_out[6316] <= layer0_out[8099] | layer0_out[8100];
     layer1_out[6317] <= ~layer0_out[6048];
     layer1_out[6318] <= layer0_out[2811] & ~layer0_out[2812];
     layer1_out[6319] <= ~layer0_out[9898];
     layer1_out[6320] <= layer0_out[6960] ^ layer0_out[6961];
     layer1_out[6321] <= ~(layer0_out[3350] & layer0_out[3351]);
     layer1_out[6322] <= layer0_out[11553] & ~layer0_out[11552];
     layer1_out[6323] <= layer0_out[426] & ~layer0_out[425];
     layer1_out[6324] <= ~layer0_out[4864];
     layer1_out[6325] <= layer0_out[11862];
     layer1_out[6326] <= ~(layer0_out[316] & layer0_out[317]);
     layer1_out[6327] <= ~layer0_out[7279];
     layer1_out[6328] <= layer0_out[3535];
     layer1_out[6329] <= ~layer0_out[7667] | layer0_out[7666];
     layer1_out[6330] <= ~layer0_out[3911] | layer0_out[3910];
     layer1_out[6331] <= layer0_out[3362] & ~layer0_out[3361];
     layer1_out[6332] <= ~layer0_out[1352] | layer0_out[1353];
     layer1_out[6333] <= ~layer0_out[11147] | layer0_out[11146];
     layer1_out[6334] <= layer0_out[9279] & ~layer0_out[9280];
     layer1_out[6335] <= ~layer0_out[11641];
     layer1_out[6336] <= ~layer0_out[2825] | layer0_out[2826];
     layer1_out[6337] <= layer0_out[8070] & ~layer0_out[8071];
     layer1_out[6338] <= ~layer0_out[4044];
     layer1_out[6339] <= 1'b1;
     layer1_out[6340] <= layer0_out[1363];
     layer1_out[6341] <= ~layer0_out[5691] | layer0_out[5690];
     layer1_out[6342] <= ~layer0_out[6495];
     layer1_out[6343] <= 1'b0;
     layer1_out[6344] <= layer0_out[9364] & ~layer0_out[9365];
     layer1_out[6345] <= layer0_out[4303] & layer0_out[4304];
     layer1_out[6346] <= layer0_out[9834] & ~layer0_out[9835];
     layer1_out[6347] <= ~layer0_out[5732];
     layer1_out[6348] <= ~layer0_out[4342];
     layer1_out[6349] <= ~layer0_out[9392] | layer0_out[9391];
     layer1_out[6350] <= layer0_out[6203];
     layer1_out[6351] <= ~layer0_out[2994];
     layer1_out[6352] <= layer0_out[1995] | layer0_out[1996];
     layer1_out[6353] <= ~layer0_out[11974] | layer0_out[11973];
     layer1_out[6354] <= 1'b0;
     layer1_out[6355] <= layer0_out[6536] ^ layer0_out[6537];
     layer1_out[6356] <= layer0_out[11211] & layer0_out[11212];
     layer1_out[6357] <= ~layer0_out[3476];
     layer1_out[6358] <= ~layer0_out[7835] | layer0_out[7834];
     layer1_out[6359] <= layer0_out[5805];
     layer1_out[6360] <= ~layer0_out[4917] | layer0_out[4916];
     layer1_out[6361] <= ~layer0_out[479];
     layer1_out[6362] <= layer0_out[11939];
     layer1_out[6363] <= layer0_out[2997] ^ layer0_out[2998];
     layer1_out[6364] <= ~layer0_out[2598] | layer0_out[2599];
     layer1_out[6365] <= 1'b1;
     layer1_out[6366] <= ~layer0_out[17];
     layer1_out[6367] <= layer0_out[9095];
     layer1_out[6368] <= layer0_out[11247];
     layer1_out[6369] <= ~layer0_out[2513];
     layer1_out[6370] <= layer0_out[4274];
     layer1_out[6371] <= layer0_out[7071];
     layer1_out[6372] <= layer0_out[9437] ^ layer0_out[9438];
     layer1_out[6373] <= layer0_out[1347] | layer0_out[1348];
     layer1_out[6374] <= ~layer0_out[8144];
     layer1_out[6375] <= layer0_out[9572];
     layer1_out[6376] <= ~layer0_out[11367];
     layer1_out[6377] <= ~(layer0_out[1163] | layer0_out[1164]);
     layer1_out[6378] <= ~layer0_out[6542] | layer0_out[6541];
     layer1_out[6379] <= layer0_out[5820] | layer0_out[5821];
     layer1_out[6380] <= 1'b0;
     layer1_out[6381] <= ~layer0_out[11445];
     layer1_out[6382] <= 1'b0;
     layer1_out[6383] <= layer0_out[11483] & layer0_out[11484];
     layer1_out[6384] <= ~(layer0_out[1073] | layer0_out[1074]);
     layer1_out[6385] <= layer0_out[7157];
     layer1_out[6386] <= layer0_out[1848];
     layer1_out[6387] <= ~layer0_out[6043];
     layer1_out[6388] <= layer0_out[10947];
     layer1_out[6389] <= layer0_out[2705];
     layer1_out[6390] <= layer0_out[3397];
     layer1_out[6391] <= layer0_out[11558] & layer0_out[11559];
     layer1_out[6392] <= layer0_out[7601] & ~layer0_out[7602];
     layer1_out[6393] <= layer0_out[11779];
     layer1_out[6394] <= ~(layer0_out[1959] & layer0_out[1960]);
     layer1_out[6395] <= layer0_out[11114] & layer0_out[11115];
     layer1_out[6396] <= ~layer0_out[4393];
     layer1_out[6397] <= ~layer0_out[7130];
     layer1_out[6398] <= ~layer0_out[8550] | layer0_out[8551];
     layer1_out[6399] <= ~(layer0_out[11391] & layer0_out[11392]);
     layer1_out[6400] <= ~layer0_out[1690] | layer0_out[1689];
     layer1_out[6401] <= ~(layer0_out[4718] | layer0_out[4719]);
     layer1_out[6402] <= layer0_out[1014] & layer0_out[1015];
     layer1_out[6403] <= 1'b1;
     layer1_out[6404] <= ~layer0_out[11582];
     layer1_out[6405] <= ~layer0_out[7867];
     layer1_out[6406] <= layer0_out[1211];
     layer1_out[6407] <= ~layer0_out[5469];
     layer1_out[6408] <= layer0_out[10866] | layer0_out[10867];
     layer1_out[6409] <= layer0_out[3903];
     layer1_out[6410] <= ~layer0_out[6208] | layer0_out[6209];
     layer1_out[6411] <= ~(layer0_out[806] ^ layer0_out[807]);
     layer1_out[6412] <= layer0_out[3411];
     layer1_out[6413] <= layer0_out[1382] | layer0_out[1383];
     layer1_out[6414] <= ~layer0_out[8487];
     layer1_out[6415] <= 1'b0;
     layer1_out[6416] <= layer0_out[6258] & ~layer0_out[6257];
     layer1_out[6417] <= layer0_out[979];
     layer1_out[6418] <= layer0_out[4107] & ~layer0_out[4108];
     layer1_out[6419] <= layer0_out[10013] & layer0_out[10014];
     layer1_out[6420] <= ~(layer0_out[1474] & layer0_out[1475]);
     layer1_out[6421] <= ~layer0_out[5681];
     layer1_out[6422] <= ~(layer0_out[7188] & layer0_out[7189]);
     layer1_out[6423] <= layer0_out[8515];
     layer1_out[6424] <= ~layer0_out[10128] | layer0_out[10129];
     layer1_out[6425] <= ~layer0_out[4781] | layer0_out[4780];
     layer1_out[6426] <= ~layer0_out[3965];
     layer1_out[6427] <= ~(layer0_out[7568] | layer0_out[7569]);
     layer1_out[6428] <= layer0_out[8484] & ~layer0_out[8485];
     layer1_out[6429] <= layer0_out[11371] & layer0_out[11372];
     layer1_out[6430] <= layer0_out[4108];
     layer1_out[6431] <= layer0_out[9617];
     layer1_out[6432] <= layer0_out[6331] ^ layer0_out[6332];
     layer1_out[6433] <= 1'b1;
     layer1_out[6434] <= layer0_out[6409] | layer0_out[6410];
     layer1_out[6435] <= ~(layer0_out[7] | layer0_out[8]);
     layer1_out[6436] <= ~(layer0_out[11488] | layer0_out[11489]);
     layer1_out[6437] <= layer0_out[8241];
     layer1_out[6438] <= ~(layer0_out[8141] ^ layer0_out[8142]);
     layer1_out[6439] <= layer0_out[1844];
     layer1_out[6440] <= layer0_out[6396];
     layer1_out[6441] <= ~(layer0_out[5048] & layer0_out[5049]);
     layer1_out[6442] <= ~layer0_out[3959] | layer0_out[3958];
     layer1_out[6443] <= layer0_out[1053];
     layer1_out[6444] <= 1'b0;
     layer1_out[6445] <= layer0_out[1400];
     layer1_out[6446] <= layer0_out[6220] | layer0_out[6221];
     layer1_out[6447] <= ~layer0_out[63] | layer0_out[64];
     layer1_out[6448] <= layer0_out[3633] ^ layer0_out[3634];
     layer1_out[6449] <= layer0_out[2389];
     layer1_out[6450] <= layer0_out[9252];
     layer1_out[6451] <= ~(layer0_out[2305] | layer0_out[2306]);
     layer1_out[6452] <= layer0_out[693];
     layer1_out[6453] <= layer0_out[8637] & ~layer0_out[8636];
     layer1_out[6454] <= layer0_out[2830] & ~layer0_out[2829];
     layer1_out[6455] <= ~layer0_out[4178] | layer0_out[4177];
     layer1_out[6456] <= layer0_out[7857] & ~layer0_out[7858];
     layer1_out[6457] <= ~layer0_out[2489];
     layer1_out[6458] <= layer0_out[11088];
     layer1_out[6459] <= layer0_out[6725] ^ layer0_out[6726];
     layer1_out[6460] <= ~(layer0_out[9774] ^ layer0_out[9775]);
     layer1_out[6461] <= layer0_out[6347];
     layer1_out[6462] <= layer0_out[11954] & ~layer0_out[11953];
     layer1_out[6463] <= ~(layer0_out[5104] & layer0_out[5105]);
     layer1_out[6464] <= layer0_out[10955];
     layer1_out[6465] <= layer0_out[11849] | layer0_out[11850];
     layer1_out[6466] <= layer0_out[9379] & ~layer0_out[9380];
     layer1_out[6467] <= layer0_out[6676] & ~layer0_out[6675];
     layer1_out[6468] <= ~layer0_out[2450] | layer0_out[2451];
     layer1_out[6469] <= layer0_out[956] & layer0_out[957];
     layer1_out[6470] <= layer0_out[3972];
     layer1_out[6471] <= 1'b1;
     layer1_out[6472] <= ~(layer0_out[9860] | layer0_out[9861]);
     layer1_out[6473] <= layer0_out[11193];
     layer1_out[6474] <= ~layer0_out[6457] | layer0_out[6456];
     layer1_out[6475] <= layer0_out[3868];
     layer1_out[6476] <= layer0_out[804];
     layer1_out[6477] <= layer0_out[1775] | layer0_out[1776];
     layer1_out[6478] <= layer0_out[4660] & ~layer0_out[4661];
     layer1_out[6479] <= layer0_out[9957] ^ layer0_out[9958];
     layer1_out[6480] <= layer0_out[11383] & ~layer0_out[11382];
     layer1_out[6481] <= ~(layer0_out[7338] & layer0_out[7339]);
     layer1_out[6482] <= ~layer0_out[4523];
     layer1_out[6483] <= layer0_out[4810] & ~layer0_out[4809];
     layer1_out[6484] <= layer0_out[5327] | layer0_out[5328];
     layer1_out[6485] <= layer0_out[7520];
     layer1_out[6486] <= ~layer0_out[5969];
     layer1_out[6487] <= ~layer0_out[3066];
     layer1_out[6488] <= 1'b1;
     layer1_out[6489] <= ~layer0_out[9197];
     layer1_out[6490] <= layer0_out[3376] & layer0_out[3377];
     layer1_out[6491] <= layer0_out[413] | layer0_out[414];
     layer1_out[6492] <= ~(layer0_out[5937] ^ layer0_out[5938]);
     layer1_out[6493] <= ~layer0_out[6218] | layer0_out[6217];
     layer1_out[6494] <= ~(layer0_out[797] & layer0_out[798]);
     layer1_out[6495] <= layer0_out[2717];
     layer1_out[6496] <= ~(layer0_out[11937] ^ layer0_out[11938]);
     layer1_out[6497] <= ~(layer0_out[3710] & layer0_out[3711]);
     layer1_out[6498] <= layer0_out[10760] & ~layer0_out[10759];
     layer1_out[6499] <= ~(layer0_out[574] | layer0_out[575]);
     layer1_out[6500] <= layer0_out[11670] & layer0_out[11671];
     layer1_out[6501] <= layer0_out[4834] & ~layer0_out[4835];
     layer1_out[6502] <= ~(layer0_out[3219] | layer0_out[3220]);
     layer1_out[6503] <= ~(layer0_out[6855] | layer0_out[6856]);
     layer1_out[6504] <= ~(layer0_out[3250] & layer0_out[3251]);
     layer1_out[6505] <= layer0_out[6189] & ~layer0_out[6190];
     layer1_out[6506] <= ~layer0_out[4709];
     layer1_out[6507] <= layer0_out[11379] & ~layer0_out[11378];
     layer1_out[6508] <= layer0_out[3713] & ~layer0_out[3712];
     layer1_out[6509] <= layer0_out[3429] | layer0_out[3430];
     layer1_out[6510] <= 1'b0;
     layer1_out[6511] <= ~layer0_out[4612] | layer0_out[4611];
     layer1_out[6512] <= ~layer0_out[1268];
     layer1_out[6513] <= ~(layer0_out[594] & layer0_out[595]);
     layer1_out[6514] <= 1'b0;
     layer1_out[6515] <= layer0_out[8739] | layer0_out[8740];
     layer1_out[6516] <= layer0_out[7787] & ~layer0_out[7786];
     layer1_out[6517] <= ~layer0_out[2420] | layer0_out[2419];
     layer1_out[6518] <= ~layer0_out[9339];
     layer1_out[6519] <= layer0_out[7037] & ~layer0_out[7038];
     layer1_out[6520] <= ~(layer0_out[11606] | layer0_out[11607]);
     layer1_out[6521] <= layer0_out[8889] | layer0_out[8890];
     layer1_out[6522] <= layer0_out[3985];
     layer1_out[6523] <= ~layer0_out[6454];
     layer1_out[6524] <= ~layer0_out[3127] | layer0_out[3128];
     layer1_out[6525] <= ~(layer0_out[3729] | layer0_out[3730]);
     layer1_out[6526] <= ~(layer0_out[11440] | layer0_out[11441]);
     layer1_out[6527] <= ~layer0_out[10013];
     layer1_out[6528] <= ~layer0_out[125];
     layer1_out[6529] <= ~layer0_out[160] | layer0_out[161];
     layer1_out[6530] <= ~(layer0_out[5972] ^ layer0_out[5973]);
     layer1_out[6531] <= layer0_out[8748];
     layer1_out[6532] <= layer0_out[6065] | layer0_out[6066];
     layer1_out[6533] <= ~layer0_out[1593] | layer0_out[1594];
     layer1_out[6534] <= ~(layer0_out[4178] | layer0_out[4179]);
     layer1_out[6535] <= layer0_out[2529] & ~layer0_out[2530];
     layer1_out[6536] <= layer0_out[11732] & ~layer0_out[11731];
     layer1_out[6537] <= layer0_out[2527] & layer0_out[2528];
     layer1_out[6538] <= layer0_out[10811];
     layer1_out[6539] <= ~layer0_out[6071] | layer0_out[6072];
     layer1_out[6540] <= layer0_out[1950] & ~layer0_out[1949];
     layer1_out[6541] <= ~layer0_out[5158];
     layer1_out[6542] <= ~layer0_out[6238];
     layer1_out[6543] <= layer0_out[6194] & ~layer0_out[6193];
     layer1_out[6544] <= layer0_out[541] & layer0_out[542];
     layer1_out[6545] <= layer0_out[7519];
     layer1_out[6546] <= ~layer0_out[3217] | layer0_out[3218];
     layer1_out[6547] <= layer0_out[10333];
     layer1_out[6548] <= layer0_out[4880];
     layer1_out[6549] <= ~layer0_out[1509];
     layer1_out[6550] <= ~layer0_out[8869];
     layer1_out[6551] <= ~layer0_out[6461];
     layer1_out[6552] <= ~layer0_out[4396];
     layer1_out[6553] <= layer0_out[9725] & ~layer0_out[9724];
     layer1_out[6554] <= 1'b0;
     layer1_out[6555] <= layer0_out[7463] & ~layer0_out[7462];
     layer1_out[6556] <= ~layer0_out[8391];
     layer1_out[6557] <= ~(layer0_out[9313] ^ layer0_out[9314]);
     layer1_out[6558] <= ~layer0_out[2639] | layer0_out[2638];
     layer1_out[6559] <= layer0_out[2575] & ~layer0_out[2574];
     layer1_out[6560] <= layer0_out[6113];
     layer1_out[6561] <= layer0_out[10667] ^ layer0_out[10668];
     layer1_out[6562] <= ~layer0_out[10762] | layer0_out[10763];
     layer1_out[6563] <= ~layer0_out[6893] | layer0_out[6892];
     layer1_out[6564] <= ~(layer0_out[4572] & layer0_out[4573]);
     layer1_out[6565] <= ~layer0_out[1511] | layer0_out[1512];
     layer1_out[6566] <= layer0_out[10879];
     layer1_out[6567] <= layer0_out[7778] & ~layer0_out[7779];
     layer1_out[6568] <= layer0_out[11653] ^ layer0_out[11654];
     layer1_out[6569] <= ~layer0_out[5890];
     layer1_out[6570] <= layer0_out[10048] & ~layer0_out[10047];
     layer1_out[6571] <= ~layer0_out[3841] | layer0_out[3842];
     layer1_out[6572] <= ~(layer0_out[1913] & layer0_out[1914]);
     layer1_out[6573] <= layer0_out[5481] & layer0_out[5482];
     layer1_out[6574] <= layer0_out[6725];
     layer1_out[6575] <= layer0_out[3289];
     layer1_out[6576] <= layer0_out[1839] | layer0_out[1840];
     layer1_out[6577] <= layer0_out[10295] & ~layer0_out[10296];
     layer1_out[6578] <= layer0_out[11531];
     layer1_out[6579] <= layer0_out[7801];
     layer1_out[6580] <= ~(layer0_out[11674] ^ layer0_out[11675]);
     layer1_out[6581] <= layer0_out[4252] & ~layer0_out[4251];
     layer1_out[6582] <= layer0_out[913];
     layer1_out[6583] <= layer0_out[7977] & ~layer0_out[7978];
     layer1_out[6584] <= layer0_out[8199] & ~layer0_out[8198];
     layer1_out[6585] <= layer0_out[9784];
     layer1_out[6586] <= layer0_out[2041];
     layer1_out[6587] <= layer0_out[9359] & ~layer0_out[9358];
     layer1_out[6588] <= layer0_out[7445];
     layer1_out[6589] <= ~layer0_out[11384];
     layer1_out[6590] <= ~layer0_out[3749];
     layer1_out[6591] <= layer0_out[8298] & ~layer0_out[8297];
     layer1_out[6592] <= layer0_out[10869] ^ layer0_out[10870];
     layer1_out[6593] <= layer0_out[11386] ^ layer0_out[11387];
     layer1_out[6594] <= layer0_out[6798] ^ layer0_out[6799];
     layer1_out[6595] <= ~(layer0_out[1706] & layer0_out[1707]);
     layer1_out[6596] <= layer0_out[11724] & ~layer0_out[11725];
     layer1_out[6597] <= ~layer0_out[571];
     layer1_out[6598] <= layer0_out[10093] | layer0_out[10094];
     layer1_out[6599] <= layer0_out[2922];
     layer1_out[6600] <= ~layer0_out[7559];
     layer1_out[6601] <= ~(layer0_out[947] & layer0_out[948]);
     layer1_out[6602] <= ~(layer0_out[11920] | layer0_out[11921]);
     layer1_out[6603] <= layer0_out[6776] ^ layer0_out[6777];
     layer1_out[6604] <= ~(layer0_out[9719] | layer0_out[9720]);
     layer1_out[6605] <= ~layer0_out[396] | layer0_out[397];
     layer1_out[6606] <= layer0_out[6236] | layer0_out[6237];
     layer1_out[6607] <= layer0_out[4931] & ~layer0_out[4932];
     layer1_out[6608] <= layer0_out[7868] ^ layer0_out[7869];
     layer1_out[6609] <= ~(layer0_out[8504] ^ layer0_out[8505]);
     layer1_out[6610] <= ~layer0_out[4584];
     layer1_out[6611] <= 1'b0;
     layer1_out[6612] <= layer0_out[826] & layer0_out[827];
     layer1_out[6613] <= ~layer0_out[4380] | layer0_out[4381];
     layer1_out[6614] <= 1'b0;
     layer1_out[6615] <= layer0_out[10791] & layer0_out[10792];
     layer1_out[6616] <= layer0_out[10316];
     layer1_out[6617] <= layer0_out[8958] & ~layer0_out[8957];
     layer1_out[6618] <= layer0_out[5582];
     layer1_out[6619] <= layer0_out[7406];
     layer1_out[6620] <= ~(layer0_out[3962] | layer0_out[3963]);
     layer1_out[6621] <= ~(layer0_out[4133] | layer0_out[4134]);
     layer1_out[6622] <= layer0_out[7052];
     layer1_out[6623] <= layer0_out[7708] & layer0_out[7709];
     layer1_out[6624] <= 1'b1;
     layer1_out[6625] <= ~layer0_out[7899];
     layer1_out[6626] <= ~(layer0_out[7757] & layer0_out[7758]);
     layer1_out[6627] <= layer0_out[11237] & ~layer0_out[11236];
     layer1_out[6628] <= layer0_out[7763] & ~layer0_out[7762];
     layer1_out[6629] <= layer0_out[9879] | layer0_out[9880];
     layer1_out[6630] <= ~(layer0_out[3793] & layer0_out[3794]);
     layer1_out[6631] <= layer0_out[7399] & ~layer0_out[7400];
     layer1_out[6632] <= layer0_out[643];
     layer1_out[6633] <= ~(layer0_out[6258] & layer0_out[6259]);
     layer1_out[6634] <= ~layer0_out[8921];
     layer1_out[6635] <= ~layer0_out[818];
     layer1_out[6636] <= ~layer0_out[9619];
     layer1_out[6637] <= layer0_out[6642] & layer0_out[6643];
     layer1_out[6638] <= ~layer0_out[4458];
     layer1_out[6639] <= 1'b0;
     layer1_out[6640] <= 1'b1;
     layer1_out[6641] <= ~layer0_out[5808] | layer0_out[5809];
     layer1_out[6642] <= ~layer0_out[1220] | layer0_out[1221];
     layer1_out[6643] <= 1'b1;
     layer1_out[6644] <= ~layer0_out[5137] | layer0_out[5138];
     layer1_out[6645] <= layer0_out[6400];
     layer1_out[6646] <= layer0_out[3836] ^ layer0_out[3837];
     layer1_out[6647] <= ~(layer0_out[577] | layer0_out[578]);
     layer1_out[6648] <= layer0_out[9380] & layer0_out[9381];
     layer1_out[6649] <= ~(layer0_out[10366] | layer0_out[10367]);
     layer1_out[6650] <= ~layer0_out[1545] | layer0_out[1546];
     layer1_out[6651] <= layer0_out[4519];
     layer1_out[6652] <= ~layer0_out[1026];
     layer1_out[6653] <= ~(layer0_out[5192] ^ layer0_out[5193]);
     layer1_out[6654] <= ~layer0_out[5450];
     layer1_out[6655] <= ~(layer0_out[5426] ^ layer0_out[5427]);
     layer1_out[6656] <= layer0_out[78] | layer0_out[79];
     layer1_out[6657] <= layer0_out[11625];
     layer1_out[6658] <= layer0_out[8961];
     layer1_out[6659] <= layer0_out[4128] & ~layer0_out[4127];
     layer1_out[6660] <= ~layer0_out[991];
     layer1_out[6661] <= 1'b1;
     layer1_out[6662] <= layer0_out[4126] & ~layer0_out[4127];
     layer1_out[6663] <= layer0_out[6869];
     layer1_out[6664] <= ~(layer0_out[4144] | layer0_out[4145]);
     layer1_out[6665] <= layer0_out[7168] & ~layer0_out[7167];
     layer1_out[6666] <= ~(layer0_out[4892] | layer0_out[4893]);
     layer1_out[6667] <= ~(layer0_out[11595] & layer0_out[11596]);
     layer1_out[6668] <= layer0_out[476];
     layer1_out[6669] <= ~(layer0_out[9134] & layer0_out[9135]);
     layer1_out[6670] <= ~layer0_out[7503] | layer0_out[7502];
     layer1_out[6671] <= ~(layer0_out[8442] | layer0_out[8443]);
     layer1_out[6672] <= layer0_out[4517] & ~layer0_out[4518];
     layer1_out[6673] <= ~layer0_out[733];
     layer1_out[6674] <= layer0_out[3159];
     layer1_out[6675] <= layer0_out[7286];
     layer1_out[6676] <= layer0_out[9457];
     layer1_out[6677] <= ~(layer0_out[827] | layer0_out[828]);
     layer1_out[6678] <= ~layer0_out[9741];
     layer1_out[6679] <= ~layer0_out[5838];
     layer1_out[6680] <= ~(layer0_out[8347] ^ layer0_out[8348]);
     layer1_out[6681] <= layer0_out[7494];
     layer1_out[6682] <= layer0_out[10958] | layer0_out[10959];
     layer1_out[6683] <= ~layer0_out[9935];
     layer1_out[6684] <= ~layer0_out[10924] | layer0_out[10925];
     layer1_out[6685] <= layer0_out[11267] & ~layer0_out[11266];
     layer1_out[6686] <= layer0_out[4893] ^ layer0_out[4894];
     layer1_out[6687] <= layer0_out[6735] | layer0_out[6736];
     layer1_out[6688] <= ~(layer0_out[8690] | layer0_out[8691]);
     layer1_out[6689] <= ~layer0_out[2551];
     layer1_out[6690] <= ~(layer0_out[10556] ^ layer0_out[10557]);
     layer1_out[6691] <= ~layer0_out[2139];
     layer1_out[6692] <= layer0_out[10737];
     layer1_out[6693] <= layer0_out[4058];
     layer1_out[6694] <= ~layer0_out[5227];
     layer1_out[6695] <= layer0_out[8047];
     layer1_out[6696] <= ~layer0_out[2956] | layer0_out[2957];
     layer1_out[6697] <= layer0_out[5167];
     layer1_out[6698] <= layer0_out[11873];
     layer1_out[6699] <= layer0_out[8427] & ~layer0_out[8426];
     layer1_out[6700] <= 1'b0;
     layer1_out[6701] <= ~(layer0_out[3163] | layer0_out[3164]);
     layer1_out[6702] <= layer0_out[75] & ~layer0_out[76];
     layer1_out[6703] <= ~layer0_out[3828] | layer0_out[3829];
     layer1_out[6704] <= layer0_out[8291] & ~layer0_out[8292];
     layer1_out[6705] <= layer0_out[423] & ~layer0_out[424];
     layer1_out[6706] <= layer0_out[6205] ^ layer0_out[6206];
     layer1_out[6707] <= ~(layer0_out[2148] ^ layer0_out[2149]);
     layer1_out[6708] <= layer0_out[11560];
     layer1_out[6709] <= layer0_out[5127] & ~layer0_out[5126];
     layer1_out[6710] <= layer0_out[11985];
     layer1_out[6711] <= layer0_out[5397];
     layer1_out[6712] <= ~layer0_out[6956] | layer0_out[6955];
     layer1_out[6713] <= ~layer0_out[10131] | layer0_out[10130];
     layer1_out[6714] <= layer0_out[3406] ^ layer0_out[3407];
     layer1_out[6715] <= ~layer0_out[8287] | layer0_out[8288];
     layer1_out[6716] <= layer0_out[1372] & ~layer0_out[1371];
     layer1_out[6717] <= ~(layer0_out[3563] ^ layer0_out[3564]);
     layer1_out[6718] <= ~layer0_out[4064];
     layer1_out[6719] <= ~layer0_out[1763];
     layer1_out[6720] <= layer0_out[4608] & layer0_out[4609];
     layer1_out[6721] <= layer0_out[2066] & ~layer0_out[2067];
     layer1_out[6722] <= layer0_out[4215];
     layer1_out[6723] <= ~(layer0_out[8131] & layer0_out[8132]);
     layer1_out[6724] <= ~(layer0_out[9650] ^ layer0_out[9651]);
     layer1_out[6725] <= 1'b1;
     layer1_out[6726] <= layer0_out[11988] ^ layer0_out[11989];
     layer1_out[6727] <= ~layer0_out[10938];
     layer1_out[6728] <= ~(layer0_out[6001] | layer0_out[6002]);
     layer1_out[6729] <= ~layer0_out[2580];
     layer1_out[6730] <= layer0_out[5931] & ~layer0_out[5930];
     layer1_out[6731] <= ~layer0_out[7597];
     layer1_out[6732] <= ~layer0_out[3625];
     layer1_out[6733] <= layer0_out[3367] & ~layer0_out[3368];
     layer1_out[6734] <= layer0_out[720];
     layer1_out[6735] <= ~layer0_out[11226];
     layer1_out[6736] <= ~(layer0_out[11888] & layer0_out[11889]);
     layer1_out[6737] <= ~layer0_out[5061] | layer0_out[5060];
     layer1_out[6738] <= ~layer0_out[7641];
     layer1_out[6739] <= layer0_out[6483] & layer0_out[6484];
     layer1_out[6740] <= ~layer0_out[1597];
     layer1_out[6741] <= ~layer0_out[10932] | layer0_out[10931];
     layer1_out[6742] <= ~layer0_out[1777] | layer0_out[1778];
     layer1_out[6743] <= ~layer0_out[14];
     layer1_out[6744] <= layer0_out[5436];
     layer1_out[6745] <= layer0_out[10650] ^ layer0_out[10651];
     layer1_out[6746] <= layer0_out[9071] & layer0_out[9072];
     layer1_out[6747] <= ~layer0_out[1397] | layer0_out[1396];
     layer1_out[6748] <= ~(layer0_out[10385] ^ layer0_out[10386]);
     layer1_out[6749] <= layer0_out[6181] & layer0_out[6182];
     layer1_out[6750] <= layer0_out[6703] & ~layer0_out[6702];
     layer1_out[6751] <= ~(layer0_out[3235] ^ layer0_out[3236]);
     layer1_out[6752] <= ~layer0_out[5521];
     layer1_out[6753] <= ~layer0_out[4787];
     layer1_out[6754] <= ~layer0_out[339] | layer0_out[338];
     layer1_out[6755] <= ~layer0_out[7310] | layer0_out[7311];
     layer1_out[6756] <= layer0_out[10495] | layer0_out[10496];
     layer1_out[6757] <= ~layer0_out[4867] | layer0_out[4866];
     layer1_out[6758] <= ~layer0_out[1591];
     layer1_out[6759] <= ~(layer0_out[2629] | layer0_out[2630]);
     layer1_out[6760] <= layer0_out[4507];
     layer1_out[6761] <= 1'b0;
     layer1_out[6762] <= layer0_out[6590] & ~layer0_out[6591];
     layer1_out[6763] <= layer0_out[7811] & ~layer0_out[7812];
     layer1_out[6764] <= layer0_out[7818];
     layer1_out[6765] <= layer0_out[9675];
     layer1_out[6766] <= layer0_out[6129];
     layer1_out[6767] <= layer0_out[3700] & ~layer0_out[3699];
     layer1_out[6768] <= layer0_out[3368] & layer0_out[3369];
     layer1_out[6769] <= layer0_out[7036] & ~layer0_out[7035];
     layer1_out[6770] <= ~(layer0_out[4297] ^ layer0_out[4298]);
     layer1_out[6771] <= layer0_out[5346];
     layer1_out[6772] <= ~layer0_out[7836];
     layer1_out[6773] <= ~layer0_out[8076];
     layer1_out[6774] <= ~layer0_out[10341];
     layer1_out[6775] <= layer0_out[10035] ^ layer0_out[10036];
     layer1_out[6776] <= ~layer0_out[10394];
     layer1_out[6777] <= ~(layer0_out[6509] | layer0_out[6510]);
     layer1_out[6778] <= ~(layer0_out[10139] & layer0_out[10140]);
     layer1_out[6779] <= layer0_out[4633] ^ layer0_out[4634];
     layer1_out[6780] <= layer0_out[4022] & layer0_out[4023];
     layer1_out[6781] <= layer0_out[11338] | layer0_out[11339];
     layer1_out[6782] <= layer0_out[7236] ^ layer0_out[7237];
     layer1_out[6783] <= layer0_out[5509] ^ layer0_out[5510];
     layer1_out[6784] <= layer0_out[9744] & ~layer0_out[9743];
     layer1_out[6785] <= ~layer0_out[3336];
     layer1_out[6786] <= ~(layer0_out[7561] | layer0_out[7562]);
     layer1_out[6787] <= ~layer0_out[10789];
     layer1_out[6788] <= layer0_out[11555] & layer0_out[11556];
     layer1_out[6789] <= layer0_out[546] | layer0_out[547];
     layer1_out[6790] <= layer0_out[11033] ^ layer0_out[11034];
     layer1_out[6791] <= ~layer0_out[6346];
     layer1_out[6792] <= ~(layer0_out[3613] ^ layer0_out[3614]);
     layer1_out[6793] <= ~layer0_out[10746];
     layer1_out[6794] <= ~(layer0_out[10533] | layer0_out[10534]);
     layer1_out[6795] <= ~layer0_out[7443];
     layer1_out[6796] <= ~(layer0_out[9859] | layer0_out[9860]);
     layer1_out[6797] <= layer0_out[9560] & layer0_out[9561];
     layer1_out[6798] <= layer0_out[7286];
     layer1_out[6799] <= ~(layer0_out[6733] | layer0_out[6734]);
     layer1_out[6800] <= layer0_out[6006] & layer0_out[6007];
     layer1_out[6801] <= ~layer0_out[10349];
     layer1_out[6802] <= ~(layer0_out[5745] & layer0_out[5746]);
     layer1_out[6803] <= ~layer0_out[8944] | layer0_out[8943];
     layer1_out[6804] <= layer0_out[11861];
     layer1_out[6805] <= ~layer0_out[6692];
     layer1_out[6806] <= ~layer0_out[2709];
     layer1_out[6807] <= ~(layer0_out[1021] ^ layer0_out[1022]);
     layer1_out[6808] <= layer0_out[10839];
     layer1_out[6809] <= ~layer0_out[7729] | layer0_out[7730];
     layer1_out[6810] <= ~(layer0_out[8235] & layer0_out[8236]);
     layer1_out[6811] <= layer0_out[1196];
     layer1_out[6812] <= ~layer0_out[2213] | layer0_out[2214];
     layer1_out[6813] <= layer0_out[2168] & layer0_out[2169];
     layer1_out[6814] <= ~layer0_out[1947];
     layer1_out[6815] <= ~layer0_out[11091] | layer0_out[11092];
     layer1_out[6816] <= ~(layer0_out[6842] & layer0_out[6843]);
     layer1_out[6817] <= ~layer0_out[7494] | layer0_out[7493];
     layer1_out[6818] <= ~(layer0_out[11340] | layer0_out[11341]);
     layer1_out[6819] <= ~(layer0_out[9892] & layer0_out[9893]);
     layer1_out[6820] <= layer0_out[9973] & ~layer0_out[9972];
     layer1_out[6821] <= layer0_out[9523] & layer0_out[9524];
     layer1_out[6822] <= layer0_out[4261] & ~layer0_out[4260];
     layer1_out[6823] <= ~layer0_out[8272] | layer0_out[8271];
     layer1_out[6824] <= layer0_out[11403];
     layer1_out[6825] <= layer0_out[9324] & ~layer0_out[9323];
     layer1_out[6826] <= layer0_out[1954] & ~layer0_out[1953];
     layer1_out[6827] <= ~layer0_out[8280] | layer0_out[8281];
     layer1_out[6828] <= ~layer0_out[3016];
     layer1_out[6829] <= layer0_out[6219] | layer0_out[6220];
     layer1_out[6830] <= ~layer0_out[1420];
     layer1_out[6831] <= layer0_out[5159];
     layer1_out[6832] <= ~layer0_out[192];
     layer1_out[6833] <= layer0_out[8847] & ~layer0_out[8848];
     layer1_out[6834] <= ~layer0_out[5146] | layer0_out[5147];
     layer1_out[6835] <= ~(layer0_out[10991] ^ layer0_out[10992]);
     layer1_out[6836] <= ~(layer0_out[8715] | layer0_out[8716]);
     layer1_out[6837] <= layer0_out[4948];
     layer1_out[6838] <= 1'b0;
     layer1_out[6839] <= ~layer0_out[7934];
     layer1_out[6840] <= ~layer0_out[1513] | layer0_out[1512];
     layer1_out[6841] <= layer0_out[4172] & layer0_out[4173];
     layer1_out[6842] <= ~(layer0_out[10153] | layer0_out[10154]);
     layer1_out[6843] <= ~layer0_out[7637];
     layer1_out[6844] <= layer0_out[10682] | layer0_out[10683];
     layer1_out[6845] <= layer0_out[4166];
     layer1_out[6846] <= layer0_out[10184];
     layer1_out[6847] <= layer0_out[4378];
     layer1_out[6848] <= layer0_out[8735];
     layer1_out[6849] <= ~layer0_out[7005] | layer0_out[7004];
     layer1_out[6850] <= ~(layer0_out[1782] | layer0_out[1783]);
     layer1_out[6851] <= layer0_out[10210] | layer0_out[10211];
     layer1_out[6852] <= ~(layer0_out[10640] ^ layer0_out[10641]);
     layer1_out[6853] <= layer0_out[5057] & ~layer0_out[5058];
     layer1_out[6854] <= ~(layer0_out[5339] | layer0_out[5340]);
     layer1_out[6855] <= ~layer0_out[3970];
     layer1_out[6856] <= ~layer0_out[10282] | layer0_out[10281];
     layer1_out[6857] <= ~(layer0_out[8506] & layer0_out[8507]);
     layer1_out[6858] <= layer0_out[5081] | layer0_out[5082];
     layer1_out[6859] <= ~layer0_out[3292];
     layer1_out[6860] <= ~layer0_out[10859] | layer0_out[10860];
     layer1_out[6861] <= ~layer0_out[1204];
     layer1_out[6862] <= ~(layer0_out[10382] | layer0_out[10383]);
     layer1_out[6863] <= ~(layer0_out[7539] & layer0_out[7540]);
     layer1_out[6864] <= layer0_out[756] & layer0_out[757];
     layer1_out[6865] <= ~(layer0_out[8134] ^ layer0_out[8135]);
     layer1_out[6866] <= layer0_out[11054] & ~layer0_out[11055];
     layer1_out[6867] <= layer0_out[6111] | layer0_out[6112];
     layer1_out[6868] <= ~layer0_out[2808];
     layer1_out[6869] <= ~(layer0_out[10900] | layer0_out[10901]);
     layer1_out[6870] <= ~layer0_out[3230];
     layer1_out[6871] <= layer0_out[11048] | layer0_out[11049];
     layer1_out[6872] <= ~layer0_out[4357] | layer0_out[4358];
     layer1_out[6873] <= layer0_out[1657];
     layer1_out[6874] <= layer0_out[11589] & layer0_out[11590];
     layer1_out[6875] <= layer0_out[10416];
     layer1_out[6876] <= layer0_out[2140] ^ layer0_out[2141];
     layer1_out[6877] <= layer0_out[1378];
     layer1_out[6878] <= layer0_out[4725];
     layer1_out[6879] <= ~(layer0_out[10812] | layer0_out[10813]);
     layer1_out[6880] <= layer0_out[66];
     layer1_out[6881] <= layer0_out[10841] & ~layer0_out[10842];
     layer1_out[6882] <= layer0_out[6620] | layer0_out[6621];
     layer1_out[6883] <= ~layer0_out[10249];
     layer1_out[6884] <= ~(layer0_out[11316] ^ layer0_out[11317]);
     layer1_out[6885] <= layer0_out[816] & ~layer0_out[817];
     layer1_out[6886] <= 1'b0;
     layer1_out[6887] <= layer0_out[6341] & layer0_out[6342];
     layer1_out[6888] <= ~layer0_out[8320];
     layer1_out[6889] <= 1'b0;
     layer1_out[6890] <= layer0_out[4120];
     layer1_out[6891] <= ~layer0_out[5843];
     layer1_out[6892] <= layer0_out[11679] | layer0_out[11680];
     layer1_out[6893] <= layer0_out[5639];
     layer1_out[6894] <= ~layer0_out[712];
     layer1_out[6895] <= ~layer0_out[11471] | layer0_out[11472];
     layer1_out[6896] <= ~layer0_out[4933] | layer0_out[4932];
     layer1_out[6897] <= ~(layer0_out[6349] | layer0_out[6350]);
     layer1_out[6898] <= layer0_out[1517] & ~layer0_out[1516];
     layer1_out[6899] <= layer0_out[4658];
     layer1_out[6900] <= layer0_out[4347] & ~layer0_out[4346];
     layer1_out[6901] <= layer0_out[5664] & ~layer0_out[5665];
     layer1_out[6902] <= ~layer0_out[9152];
     layer1_out[6903] <= layer0_out[6470];
     layer1_out[6904] <= ~layer0_out[4295];
     layer1_out[6905] <= layer0_out[1712] & ~layer0_out[1713];
     layer1_out[6906] <= layer0_out[3791] & ~layer0_out[3790];
     layer1_out[6907] <= layer0_out[6996] & ~layer0_out[6995];
     layer1_out[6908] <= 1'b1;
     layer1_out[6909] <= ~layer0_out[11019] | layer0_out[11020];
     layer1_out[6910] <= layer0_out[2319] & ~layer0_out[2320];
     layer1_out[6911] <= 1'b1;
     layer1_out[6912] <= 1'b0;
     layer1_out[6913] <= layer0_out[863];
     layer1_out[6914] <= ~(layer0_out[1078] & layer0_out[1079]);
     layer1_out[6915] <= layer0_out[4389] | layer0_out[4390];
     layer1_out[6916] <= ~layer0_out[7209];
     layer1_out[6917] <= layer0_out[3157] & ~layer0_out[3158];
     layer1_out[6918] <= layer0_out[7027];
     layer1_out[6919] <= layer0_out[10112] ^ layer0_out[10113];
     layer1_out[6920] <= ~(layer0_out[8081] | layer0_out[8082]);
     layer1_out[6921] <= ~(layer0_out[7927] & layer0_out[7928]);
     layer1_out[6922] <= ~layer0_out[11243] | layer0_out[11242];
     layer1_out[6923] <= ~layer0_out[9981];
     layer1_out[6924] <= ~(layer0_out[10120] & layer0_out[10121]);
     layer1_out[6925] <= ~layer0_out[4334];
     layer1_out[6926] <= layer0_out[787] | layer0_out[788];
     layer1_out[6927] <= layer0_out[1931];
     layer1_out[6928] <= layer0_out[8734] | layer0_out[8735];
     layer1_out[6929] <= ~(layer0_out[5594] ^ layer0_out[5595]);
     layer1_out[6930] <= layer0_out[3312] | layer0_out[3313];
     layer1_out[6931] <= ~layer0_out[7266];
     layer1_out[6932] <= layer0_out[786];
     layer1_out[6933] <= layer0_out[7453] | layer0_out[7454];
     layer1_out[6934] <= ~layer0_out[5887] | layer0_out[5886];
     layer1_out[6935] <= ~layer0_out[9443];
     layer1_out[6936] <= layer0_out[1617] ^ layer0_out[1618];
     layer1_out[6937] <= ~layer0_out[1837] | layer0_out[1836];
     layer1_out[6938] <= ~layer0_out[4181];
     layer1_out[6939] <= ~layer0_out[11523];
     layer1_out[6940] <= layer0_out[6765];
     layer1_out[6941] <= layer0_out[9564];
     layer1_out[6942] <= ~layer0_out[5050];
     layer1_out[6943] <= ~(layer0_out[1066] | layer0_out[1067]);
     layer1_out[6944] <= ~(layer0_out[68] & layer0_out[69]);
     layer1_out[6945] <= layer0_out[11613];
     layer1_out[6946] <= layer0_out[10268] & layer0_out[10269];
     layer1_out[6947] <= ~layer0_out[2335] | layer0_out[2334];
     layer1_out[6948] <= ~layer0_out[5359] | layer0_out[5360];
     layer1_out[6949] <= ~layer0_out[8151];
     layer1_out[6950] <= layer0_out[9516] & ~layer0_out[9517];
     layer1_out[6951] <= ~layer0_out[5576] | layer0_out[5577];
     layer1_out[6952] <= ~(layer0_out[3407] ^ layer0_out[3408]);
     layer1_out[6953] <= layer0_out[2241] ^ layer0_out[2242];
     layer1_out[6954] <= layer0_out[10920];
     layer1_out[6955] <= layer0_out[7899];
     layer1_out[6956] <= layer0_out[11450] & ~layer0_out[11449];
     layer1_out[6957] <= layer0_out[11725];
     layer1_out[6958] <= layer0_out[8682] & ~layer0_out[8683];
     layer1_out[6959] <= layer0_out[3872];
     layer1_out[6960] <= layer0_out[9601] & layer0_out[9602];
     layer1_out[6961] <= layer0_out[50] & ~layer0_out[51];
     layer1_out[6962] <= layer0_out[8666];
     layer1_out[6963] <= ~layer0_out[5420] | layer0_out[5419];
     layer1_out[6964] <= layer0_out[10062];
     layer1_out[6965] <= ~(layer0_out[4549] & layer0_out[4550]);
     layer1_out[6966] <= ~layer0_out[8817];
     layer1_out[6967] <= ~layer0_out[2154];
     layer1_out[6968] <= layer0_out[383] & ~layer0_out[382];
     layer1_out[6969] <= ~(layer0_out[2259] ^ layer0_out[2260]);
     layer1_out[6970] <= ~layer0_out[10328];
     layer1_out[6971] <= ~layer0_out[8562];
     layer1_out[6972] <= layer0_out[3944] & layer0_out[3945];
     layer1_out[6973] <= ~layer0_out[7034];
     layer1_out[6974] <= ~(layer0_out[1518] & layer0_out[1519]);
     layer1_out[6975] <= layer0_out[6619] | layer0_out[6620];
     layer1_out[6976] <= ~(layer0_out[886] ^ layer0_out[887]);
     layer1_out[6977] <= ~layer0_out[3682] | layer0_out[3683];
     layer1_out[6978] <= layer0_out[4952];
     layer1_out[6979] <= layer0_out[9085] | layer0_out[9086];
     layer1_out[6980] <= layer0_out[3964] & layer0_out[3965];
     layer1_out[6981] <= ~layer0_out[8660] | layer0_out[8659];
     layer1_out[6982] <= ~layer0_out[6264];
     layer1_out[6983] <= layer0_out[773] | layer0_out[774];
     layer1_out[6984] <= layer0_out[7528] ^ layer0_out[7529];
     layer1_out[6985] <= ~layer0_out[2098];
     layer1_out[6986] <= layer0_out[1871];
     layer1_out[6987] <= layer0_out[3862] & layer0_out[3863];
     layer1_out[6988] <= ~layer0_out[11108];
     layer1_out[6989] <= layer0_out[3173];
     layer1_out[6990] <= ~layer0_out[4991];
     layer1_out[6991] <= layer0_out[8671] ^ layer0_out[8672];
     layer1_out[6992] <= layer0_out[3186];
     layer1_out[6993] <= ~layer0_out[4943] | layer0_out[4942];
     layer1_out[6994] <= ~layer0_out[11813];
     layer1_out[6995] <= layer0_out[4910];
     layer1_out[6996] <= ~layer0_out[10449];
     layer1_out[6997] <= layer0_out[4148] & ~layer0_out[4149];
     layer1_out[6998] <= layer0_out[10750] & layer0_out[10751];
     layer1_out[6999] <= ~(layer0_out[10673] | layer0_out[10674]);
     layer1_out[7000] <= ~layer0_out[11423];
     layer1_out[7001] <= ~layer0_out[2773];
     layer1_out[7002] <= ~layer0_out[9933];
     layer1_out[7003] <= ~layer0_out[5305];
     layer1_out[7004] <= ~layer0_out[480] | layer0_out[481];
     layer1_out[7005] <= layer0_out[7544] & layer0_out[7545];
     layer1_out[7006] <= layer0_out[10575] | layer0_out[10576];
     layer1_out[7007] <= ~layer0_out[561];
     layer1_out[7008] <= layer0_out[2034] & ~layer0_out[2033];
     layer1_out[7009] <= layer0_out[2642];
     layer1_out[7010] <= layer0_out[9231] & layer0_out[9232];
     layer1_out[7011] <= layer0_out[5941];
     layer1_out[7012] <= layer0_out[5324];
     layer1_out[7013] <= 1'b0;
     layer1_out[7014] <= ~(layer0_out[3929] & layer0_out[3930]);
     layer1_out[7015] <= 1'b1;
     layer1_out[7016] <= ~layer0_out[2201];
     layer1_out[7017] <= ~(layer0_out[11538] & layer0_out[11539]);
     layer1_out[7018] <= layer0_out[8020] & ~layer0_out[8021];
     layer1_out[7019] <= layer0_out[5850];
     layer1_out[7020] <= ~layer0_out[11468] | layer0_out[11467];
     layer1_out[7021] <= layer0_out[5223] | layer0_out[5224];
     layer1_out[7022] <= layer0_out[11193] & layer0_out[11194];
     layer1_out[7023] <= layer0_out[10368] ^ layer0_out[10369];
     layer1_out[7024] <= ~(layer0_out[1132] ^ layer0_out[1133]);
     layer1_out[7025] <= ~layer0_out[2589];
     layer1_out[7026] <= layer0_out[4001] & ~layer0_out[4002];
     layer1_out[7027] <= layer0_out[8985] & ~layer0_out[8986];
     layer1_out[7028] <= ~(layer0_out[1869] | layer0_out[1870]);
     layer1_out[7029] <= layer0_out[2069];
     layer1_out[7030] <= ~(layer0_out[5410] | layer0_out[5411]);
     layer1_out[7031] <= ~(layer0_out[3515] & layer0_out[3516]);
     layer1_out[7032] <= layer0_out[8208];
     layer1_out[7033] <= 1'b1;
     layer1_out[7034] <= ~layer0_out[3723];
     layer1_out[7035] <= 1'b0;
     layer1_out[7036] <= layer0_out[6130];
     layer1_out[7037] <= ~layer0_out[2702];
     layer1_out[7038] <= ~layer0_out[7560];
     layer1_out[7039] <= ~(layer0_out[9750] | layer0_out[9751]);
     layer1_out[7040] <= ~(layer0_out[10374] | layer0_out[10375]);
     layer1_out[7041] <= layer0_out[9945];
     layer1_out[7042] <= layer0_out[9457] & ~layer0_out[9456];
     layer1_out[7043] <= ~layer0_out[3653] | layer0_out[3654];
     layer1_out[7044] <= ~layer0_out[9764];
     layer1_out[7045] <= layer0_out[5938];
     layer1_out[7046] <= layer0_out[9887] ^ layer0_out[9888];
     layer1_out[7047] <= layer0_out[247] ^ layer0_out[248];
     layer1_out[7048] <= ~(layer0_out[10049] | layer0_out[10050]);
     layer1_out[7049] <= ~layer0_out[4098] | layer0_out[4097];
     layer1_out[7050] <= ~layer0_out[4064];
     layer1_out[7051] <= ~layer0_out[4352] | layer0_out[4351];
     layer1_out[7052] <= layer0_out[4308];
     layer1_out[7053] <= layer0_out[9341];
     layer1_out[7054] <= ~layer0_out[5077];
     layer1_out[7055] <= ~(layer0_out[8502] & layer0_out[8503]);
     layer1_out[7056] <= ~layer0_out[1387];
     layer1_out[7057] <= ~(layer0_out[7249] & layer0_out[7250]);
     layer1_out[7058] <= layer0_out[5608];
     layer1_out[7059] <= ~layer0_out[4528];
     layer1_out[7060] <= 1'b1;
     layer1_out[7061] <= ~layer0_out[10067];
     layer1_out[7062] <= layer0_out[7834];
     layer1_out[7063] <= layer0_out[5114] & ~layer0_out[5115];
     layer1_out[7064] <= layer0_out[3715] & ~layer0_out[3716];
     layer1_out[7065] <= layer0_out[9333];
     layer1_out[7066] <= ~layer0_out[504] | layer0_out[503];
     layer1_out[7067] <= layer0_out[9814] & layer0_out[9815];
     layer1_out[7068] <= layer0_out[1501] & ~layer0_out[1502];
     layer1_out[7069] <= ~(layer0_out[7058] & layer0_out[7059]);
     layer1_out[7070] <= layer0_out[11608] & ~layer0_out[11609];
     layer1_out[7071] <= 1'b1;
     layer1_out[7072] <= ~(layer0_out[8873] ^ layer0_out[8874]);
     layer1_out[7073] <= ~(layer0_out[186] & layer0_out[187]);
     layer1_out[7074] <= layer0_out[9977] & ~layer0_out[9976];
     layer1_out[7075] <= ~layer0_out[9382] | layer0_out[9381];
     layer1_out[7076] <= layer0_out[4940];
     layer1_out[7077] <= ~layer0_out[5713];
     layer1_out[7078] <= ~(layer0_out[2762] & layer0_out[2763]);
     layer1_out[7079] <= layer0_out[6363];
     layer1_out[7080] <= layer0_out[6918] & ~layer0_out[6919];
     layer1_out[7081] <= layer0_out[11358];
     layer1_out[7082] <= layer0_out[1739] & ~layer0_out[1738];
     layer1_out[7083] <= ~layer0_out[5769] | layer0_out[5768];
     layer1_out[7084] <= layer0_out[9347] & ~layer0_out[9346];
     layer1_out[7085] <= layer0_out[7152] & layer0_out[7153];
     layer1_out[7086] <= layer0_out[155];
     layer1_out[7087] <= layer0_out[968] | layer0_out[969];
     layer1_out[7088] <= ~layer0_out[3048] | layer0_out[3049];
     layer1_out[7089] <= ~(layer0_out[8422] ^ layer0_out[8423]);
     layer1_out[7090] <= layer0_out[11867] | layer0_out[11868];
     layer1_out[7091] <= layer0_out[1886] & layer0_out[1887];
     layer1_out[7092] <= ~layer0_out[10184];
     layer1_out[7093] <= layer0_out[9961];
     layer1_out[7094] <= ~layer0_out[6872];
     layer1_out[7095] <= layer0_out[4848];
     layer1_out[7096] <= ~layer0_out[10357];
     layer1_out[7097] <= layer0_out[313] ^ layer0_out[314];
     layer1_out[7098] <= ~(layer0_out[10283] | layer0_out[10284]);
     layer1_out[7099] <= ~(layer0_out[6299] & layer0_out[6300]);
     layer1_out[7100] <= ~layer0_out[7065] | layer0_out[7064];
     layer1_out[7101] <= ~(layer0_out[11989] | layer0_out[11990]);
     layer1_out[7102] <= ~layer0_out[3353];
     layer1_out[7103] <= layer0_out[856] | layer0_out[857];
     layer1_out[7104] <= ~layer0_out[2343];
     layer1_out[7105] <= layer0_out[11781];
     layer1_out[7106] <= 1'b0;
     layer1_out[7107] <= layer0_out[7932] | layer0_out[7933];
     layer1_out[7108] <= ~layer0_out[8702];
     layer1_out[7109] <= ~(layer0_out[5435] & layer0_out[5436]);
     layer1_out[7110] <= layer0_out[6115];
     layer1_out[7111] <= layer0_out[5492] | layer0_out[5493];
     layer1_out[7112] <= layer0_out[6975] & layer0_out[6976];
     layer1_out[7113] <= layer0_out[3089] & ~layer0_out[3090];
     layer1_out[7114] <= ~(layer0_out[2393] ^ layer0_out[2394]);
     layer1_out[7115] <= layer0_out[7721];
     layer1_out[7116] <= layer0_out[7505] & ~layer0_out[7504];
     layer1_out[7117] <= ~(layer0_out[10301] ^ layer0_out[10302]);
     layer1_out[7118] <= ~layer0_out[1787] | layer0_out[1786];
     layer1_out[7119] <= layer0_out[9453] | layer0_out[9454];
     layer1_out[7120] <= ~layer0_out[4167] | layer0_out[4168];
     layer1_out[7121] <= layer0_out[8808] & layer0_out[8809];
     layer1_out[7122] <= layer0_out[3961];
     layer1_out[7123] <= ~(layer0_out[11637] | layer0_out[11638]);
     layer1_out[7124] <= layer0_out[11323] | layer0_out[11324];
     layer1_out[7125] <= layer0_out[5110];
     layer1_out[7126] <= ~layer0_out[11163];
     layer1_out[7127] <= layer0_out[10511] | layer0_out[10512];
     layer1_out[7128] <= layer0_out[7483] & ~layer0_out[7484];
     layer1_out[7129] <= layer0_out[5767] | layer0_out[5768];
     layer1_out[7130] <= ~layer0_out[10729] | layer0_out[10730];
     layer1_out[7131] <= layer0_out[5145];
     layer1_out[7132] <= layer0_out[7905];
     layer1_out[7133] <= layer0_out[6412];
     layer1_out[7134] <= layer0_out[11100] & ~layer0_out[11099];
     layer1_out[7135] <= layer0_out[5240];
     layer1_out[7136] <= layer0_out[5514] | layer0_out[5515];
     layer1_out[7137] <= ~layer0_out[3193] | layer0_out[3192];
     layer1_out[7138] <= layer0_out[10293] ^ layer0_out[10294];
     layer1_out[7139] <= ~layer0_out[10398];
     layer1_out[7140] <= ~layer0_out[1975];
     layer1_out[7141] <= 1'b0;
     layer1_out[7142] <= ~(layer0_out[7275] | layer0_out[7276]);
     layer1_out[7143] <= layer0_out[5019] & ~layer0_out[5018];
     layer1_out[7144] <= ~layer0_out[8884] | layer0_out[8883];
     layer1_out[7145] <= ~(layer0_out[4293] | layer0_out[4294]);
     layer1_out[7146] <= layer0_out[3194] & ~layer0_out[3195];
     layer1_out[7147] <= layer0_out[611] ^ layer0_out[612];
     layer1_out[7148] <= ~(layer0_out[8931] ^ layer0_out[8932]);
     layer1_out[7149] <= layer0_out[2757] & ~layer0_out[2758];
     layer1_out[7150] <= ~layer0_out[6962] | layer0_out[6963];
     layer1_out[7151] <= layer0_out[8425];
     layer1_out[7152] <= layer0_out[2494] & layer0_out[2495];
     layer1_out[7153] <= layer0_out[10065] & layer0_out[10066];
     layer1_out[7154] <= layer0_out[5412] & ~layer0_out[5411];
     layer1_out[7155] <= layer0_out[3187] & ~layer0_out[3186];
     layer1_out[7156] <= layer0_out[5215] | layer0_out[5216];
     layer1_out[7157] <= layer0_out[11906];
     layer1_out[7158] <= ~(layer0_out[6621] | layer0_out[6622]);
     layer1_out[7159] <= layer0_out[8387];
     layer1_out[7160] <= layer0_out[7278] | layer0_out[7279];
     layer1_out[7161] <= layer0_out[3676] & layer0_out[3677];
     layer1_out[7162] <= 1'b1;
     layer1_out[7163] <= ~(layer0_out[282] & layer0_out[283]);
     layer1_out[7164] <= layer0_out[3305];
     layer1_out[7165] <= 1'b1;
     layer1_out[7166] <= ~layer0_out[1807];
     layer1_out[7167] <= layer0_out[9395];
     layer1_out[7168] <= layer0_out[6600] | layer0_out[6601];
     layer1_out[7169] <= ~(layer0_out[10539] & layer0_out[10540]);
     layer1_out[7170] <= layer0_out[5000] & layer0_out[5001];
     layer1_out[7171] <= 1'b1;
     layer1_out[7172] <= ~(layer0_out[4142] | layer0_out[4143]);
     layer1_out[7173] <= layer0_out[6375] | layer0_out[6376];
     layer1_out[7174] <= layer0_out[3857] & ~layer0_out[3858];
     layer1_out[7175] <= layer0_out[10214] & layer0_out[10215];
     layer1_out[7176] <= 1'b1;
     layer1_out[7177] <= layer0_out[8009] & ~layer0_out[8010];
     layer1_out[7178] <= 1'b1;
     layer1_out[7179] <= layer0_out[10502] & layer0_out[10503];
     layer1_out[7180] <= ~layer0_out[3992] | layer0_out[3991];
     layer1_out[7181] <= ~layer0_out[11610];
     layer1_out[7182] <= layer0_out[11466] & ~layer0_out[11465];
     layer1_out[7183] <= layer0_out[4674];
     layer1_out[7184] <= ~(layer0_out[10141] | layer0_out[10142]);
     layer1_out[7185] <= layer0_out[8147] & ~layer0_out[8148];
     layer1_out[7186] <= ~(layer0_out[6512] & layer0_out[6513]);
     layer1_out[7187] <= layer0_out[5464] & layer0_out[5465];
     layer1_out[7188] <= layer0_out[10680] & ~layer0_out[10681];
     layer1_out[7189] <= layer0_out[3561] & ~layer0_out[3562];
     layer1_out[7190] <= layer0_out[9591] | layer0_out[9592];
     layer1_out[7191] <= layer0_out[6218] & layer0_out[6219];
     layer1_out[7192] <= layer0_out[5317] ^ layer0_out[5318];
     layer1_out[7193] <= ~layer0_out[9420] | layer0_out[9419];
     layer1_out[7194] <= ~(layer0_out[10057] & layer0_out[10058]);
     layer1_out[7195] <= layer0_out[2819] & layer0_out[2820];
     layer1_out[7196] <= ~layer0_out[9740];
     layer1_out[7197] <= ~(layer0_out[6601] ^ layer0_out[6602]);
     layer1_out[7198] <= ~layer0_out[3038];
     layer1_out[7199] <= ~(layer0_out[9593] | layer0_out[9594]);
     layer1_out[7200] <= ~(layer0_out[1510] | layer0_out[1511]);
     layer1_out[7201] <= ~layer0_out[3457];
     layer1_out[7202] <= ~layer0_out[1464];
     layer1_out[7203] <= ~layer0_out[444];
     layer1_out[7204] <= ~layer0_out[1017];
     layer1_out[7205] <= layer0_out[5312] | layer0_out[5313];
     layer1_out[7206] <= ~(layer0_out[7003] & layer0_out[7004]);
     layer1_out[7207] <= ~layer0_out[4742];
     layer1_out[7208] <= ~layer0_out[6032] | layer0_out[6033];
     layer1_out[7209] <= layer0_out[7801];
     layer1_out[7210] <= ~layer0_out[2909] | layer0_out[2910];
     layer1_out[7211] <= ~(layer0_out[10257] | layer0_out[10258]);
     layer1_out[7212] <= layer0_out[10137] & ~layer0_out[10138];
     layer1_out[7213] <= layer0_out[2317] | layer0_out[2318];
     layer1_out[7214] <= layer0_out[3555];
     layer1_out[7215] <= ~(layer0_out[1495] | layer0_out[1496]);
     layer1_out[7216] <= ~layer0_out[6475] | layer0_out[6476];
     layer1_out[7217] <= ~layer0_out[6351];
     layer1_out[7218] <= layer0_out[524] & ~layer0_out[523];
     layer1_out[7219] <= ~layer0_out[3074] | layer0_out[3075];
     layer1_out[7220] <= layer0_out[8200];
     layer1_out[7221] <= layer0_out[5356] & ~layer0_out[5355];
     layer1_out[7222] <= ~(layer0_out[5693] & layer0_out[5694]);
     layer1_out[7223] <= layer0_out[5787] ^ layer0_out[5788];
     layer1_out[7224] <= ~(layer0_out[3019] | layer0_out[3020]);
     layer1_out[7225] <= ~(layer0_out[2818] ^ layer0_out[2819]);
     layer1_out[7226] <= layer0_out[10825];
     layer1_out[7227] <= layer0_out[4047];
     layer1_out[7228] <= ~layer0_out[473];
     layer1_out[7229] <= ~layer0_out[171];
     layer1_out[7230] <= layer0_out[6847] & ~layer0_out[6846];
     layer1_out[7231] <= layer0_out[1715];
     layer1_out[7232] <= ~layer0_out[136];
     layer1_out[7233] <= ~layer0_out[10886] | layer0_out[10887];
     layer1_out[7234] <= ~layer0_out[4742];
     layer1_out[7235] <= ~layer0_out[5110];
     layer1_out[7236] <= layer0_out[279] | layer0_out[280];
     layer1_out[7237] <= ~layer0_out[3098];
     layer1_out[7238] <= layer0_out[11643] & ~layer0_out[11642];
     layer1_out[7239] <= ~(layer0_out[10761] ^ layer0_out[10762]);
     layer1_out[7240] <= 1'b1;
     layer1_out[7241] <= 1'b1;
     layer1_out[7242] <= layer0_out[2541] & ~layer0_out[2542];
     layer1_out[7243] <= layer0_out[10510] ^ layer0_out[10511];
     layer1_out[7244] <= ~layer0_out[8264] | layer0_out[8263];
     layer1_out[7245] <= layer0_out[3290] | layer0_out[3291];
     layer1_out[7246] <= layer0_out[6399];
     layer1_out[7247] <= layer0_out[4496] & ~layer0_out[4497];
     layer1_out[7248] <= layer0_out[1478] | layer0_out[1479];
     layer1_out[7249] <= ~layer0_out[4298] | layer0_out[4299];
     layer1_out[7250] <= layer0_out[10764] | layer0_out[10765];
     layer1_out[7251] <= ~layer0_out[471];
     layer1_out[7252] <= layer0_out[11486];
     layer1_out[7253] <= layer0_out[1673] | layer0_out[1674];
     layer1_out[7254] <= layer0_out[9883] | layer0_out[9884];
     layer1_out[7255] <= layer0_out[7079] ^ layer0_out[7080];
     layer1_out[7256] <= ~layer0_out[3153] | layer0_out[3154];
     layer1_out[7257] <= layer0_out[8059] & layer0_out[8060];
     layer1_out[7258] <= layer0_out[2517];
     layer1_out[7259] <= ~layer0_out[4700] | layer0_out[4699];
     layer1_out[7260] <= ~(layer0_out[2671] ^ layer0_out[2672]);
     layer1_out[7261] <= ~(layer0_out[5331] & layer0_out[5332]);
     layer1_out[7262] <= ~(layer0_out[1934] & layer0_out[1935]);
     layer1_out[7263] <= ~layer0_out[4024];
     layer1_out[7264] <= layer0_out[11073] | layer0_out[11074];
     layer1_out[7265] <= ~layer0_out[8029] | layer0_out[8028];
     layer1_out[7266] <= ~(layer0_out[4673] ^ layer0_out[4674]);
     layer1_out[7267] <= ~layer0_out[4050];
     layer1_out[7268] <= 1'b1;
     layer1_out[7269] <= ~layer0_out[138];
     layer1_out[7270] <= layer0_out[5031] | layer0_out[5032];
     layer1_out[7271] <= ~(layer0_out[3918] & layer0_out[3919]);
     layer1_out[7272] <= ~layer0_out[6340] | layer0_out[6339];
     layer1_out[7273] <= layer0_out[1157];
     layer1_out[7274] <= ~layer0_out[11026] | layer0_out[11025];
     layer1_out[7275] <= ~layer0_out[9082];
     layer1_out[7276] <= layer0_out[3681] & layer0_out[3682];
     layer1_out[7277] <= layer0_out[6651];
     layer1_out[7278] <= ~layer0_out[1635] | layer0_out[1636];
     layer1_out[7279] <= ~layer0_out[10672] | layer0_out[10671];
     layer1_out[7280] <= layer0_out[4739] ^ layer0_out[4740];
     layer1_out[7281] <= layer0_out[4122] & ~layer0_out[4123];
     layer1_out[7282] <= ~layer0_out[4570] | layer0_out[4569];
     layer1_out[7283] <= layer0_out[686] & layer0_out[687];
     layer1_out[7284] <= layer0_out[7297];
     layer1_out[7285] <= ~layer0_out[10662] | layer0_out[10663];
     layer1_out[7286] <= layer0_out[1195];
     layer1_out[7287] <= layer0_out[5549] & ~layer0_out[5548];
     layer1_out[7288] <= ~layer0_out[1826];
     layer1_out[7289] <= layer0_out[2297];
     layer1_out[7290] <= layer0_out[3209] | layer0_out[3210];
     layer1_out[7291] <= ~layer0_out[4056];
     layer1_out[7292] <= layer0_out[8977] & layer0_out[8978];
     layer1_out[7293] <= ~layer0_out[1206] | layer0_out[1207];
     layer1_out[7294] <= ~layer0_out[2556];
     layer1_out[7295] <= ~layer0_out[519] | layer0_out[520];
     layer1_out[7296] <= layer0_out[3748] | layer0_out[3749];
     layer1_out[7297] <= layer0_out[10422] & ~layer0_out[10423];
     layer1_out[7298] <= layer0_out[8539] | layer0_out[8540];
     layer1_out[7299] <= ~layer0_out[940] | layer0_out[939];
     layer1_out[7300] <= layer0_out[5710] ^ layer0_out[5711];
     layer1_out[7301] <= layer0_out[4096] | layer0_out[4097];
     layer1_out[7302] <= layer0_out[9438];
     layer1_out[7303] <= ~(layer0_out[7210] & layer0_out[7211]);
     layer1_out[7304] <= layer0_out[5343];
     layer1_out[7305] <= ~layer0_out[5228];
     layer1_out[7306] <= layer0_out[6843];
     layer1_out[7307] <= layer0_out[8048] | layer0_out[8049];
     layer1_out[7308] <= layer0_out[3111] | layer0_out[3112];
     layer1_out[7309] <= ~(layer0_out[4289] & layer0_out[4290]);
     layer1_out[7310] <= ~(layer0_out[5505] & layer0_out[5506]);
     layer1_out[7311] <= ~layer0_out[9853] | layer0_out[9852];
     layer1_out[7312] <= layer0_out[2612];
     layer1_out[7313] <= layer0_out[4794] & ~layer0_out[4793];
     layer1_out[7314] <= layer0_out[9248] & ~layer0_out[9249];
     layer1_out[7315] <= ~layer0_out[10452];
     layer1_out[7316] <= ~layer0_out[7106];
     layer1_out[7317] <= ~layer0_out[825] | layer0_out[824];
     layer1_out[7318] <= ~layer0_out[9015];
     layer1_out[7319] <= ~layer0_out[8889];
     layer1_out[7320] <= layer0_out[3803] & layer0_out[3804];
     layer1_out[7321] <= layer0_out[7252] & ~layer0_out[7253];
     layer1_out[7322] <= layer0_out[4974] & ~layer0_out[4975];
     layer1_out[7323] <= layer0_out[1048];
     layer1_out[7324] <= layer0_out[4813];
     layer1_out[7325] <= layer0_out[11778];
     layer1_out[7326] <= layer0_out[8063] | layer0_out[8064];
     layer1_out[7327] <= ~layer0_out[11630];
     layer1_out[7328] <= ~(layer0_out[11508] ^ layer0_out[11509]);
     layer1_out[7329] <= ~(layer0_out[649] | layer0_out[650]);
     layer1_out[7330] <= layer0_out[2605] & ~layer0_out[2604];
     layer1_out[7331] <= ~(layer0_out[1685] & layer0_out[1686]);
     layer1_out[7332] <= ~layer0_out[11855] | layer0_out[11856];
     layer1_out[7333] <= ~layer0_out[2052] | layer0_out[2053];
     layer1_out[7334] <= layer0_out[8650] | layer0_out[8651];
     layer1_out[7335] <= ~(layer0_out[2941] ^ layer0_out[2942]);
     layer1_out[7336] <= layer0_out[7213] & ~layer0_out[7212];
     layer1_out[7337] <= ~(layer0_out[7224] & layer0_out[7225]);
     layer1_out[7338] <= layer0_out[8096];
     layer1_out[7339] <= ~layer0_out[3379];
     layer1_out[7340] <= 1'b0;
     layer1_out[7341] <= layer0_out[7958] & ~layer0_out[7959];
     layer1_out[7342] <= ~layer0_out[4301] | layer0_out[4302];
     layer1_out[7343] <= layer0_out[1969] & layer0_out[1970];
     layer1_out[7344] <= ~layer0_out[1543];
     layer1_out[7345] <= 1'b1;
     layer1_out[7346] <= layer0_out[8772] ^ layer0_out[8773];
     layer1_out[7347] <= ~layer0_out[2852] | layer0_out[2851];
     layer1_out[7348] <= ~layer0_out[8807];
     layer1_out[7349] <= ~(layer0_out[9510] & layer0_out[9511]);
     layer1_out[7350] <= ~(layer0_out[5354] | layer0_out[5355]);
     layer1_out[7351] <= ~layer0_out[4083] | layer0_out[4082];
     layer1_out[7352] <= layer0_out[10728] ^ layer0_out[10729];
     layer1_out[7353] <= layer0_out[6356];
     layer1_out[7354] <= ~layer0_out[10370] | layer0_out[10369];
     layer1_out[7355] <= layer0_out[2367];
     layer1_out[7356] <= ~layer0_out[2536];
     layer1_out[7357] <= layer0_out[3010];
     layer1_out[7358] <= ~layer0_out[4072];
     layer1_out[7359] <= layer0_out[10349];
     layer1_out[7360] <= layer0_out[5308] & layer0_out[5309];
     layer1_out[7361] <= ~layer0_out[3581] | layer0_out[3582];
     layer1_out[7362] <= ~layer0_out[511] | layer0_out[510];
     layer1_out[7363] <= ~layer0_out[3417] | layer0_out[3416];
     layer1_out[7364] <= layer0_out[7207] & ~layer0_out[7208];
     layer1_out[7365] <= 1'b1;
     layer1_out[7366] <= ~layer0_out[8106];
     layer1_out[7367] <= ~(layer0_out[9553] ^ layer0_out[9554]);
     layer1_out[7368] <= layer0_out[7015];
     layer1_out[7369] <= ~layer0_out[3887];
     layer1_out[7370] <= layer0_out[6381];
     layer1_out[7371] <= layer0_out[1761];
     layer1_out[7372] <= layer0_out[4876] ^ layer0_out[4877];
     layer1_out[7373] <= layer0_out[11666] | layer0_out[11667];
     layer1_out[7374] <= ~layer0_out[10162];
     layer1_out[7375] <= ~layer0_out[7872];
     layer1_out[7376] <= ~layer0_out[5303] | layer0_out[5304];
     layer1_out[7377] <= layer0_out[10548] | layer0_out[10549];
     layer1_out[7378] <= ~layer0_out[11046] | layer0_out[11047];
     layer1_out[7379] <= ~(layer0_out[3001] ^ layer0_out[3002]);
     layer1_out[7380] <= ~layer0_out[11405] | layer0_out[11406];
     layer1_out[7381] <= ~layer0_out[10890] | layer0_out[10889];
     layer1_out[7382] <= layer0_out[9577] & ~layer0_out[9576];
     layer1_out[7383] <= layer0_out[4202];
     layer1_out[7384] <= layer0_out[1823];
     layer1_out[7385] <= ~layer0_out[8954];
     layer1_out[7386] <= ~(layer0_out[6553] & layer0_out[6554]);
     layer1_out[7387] <= layer0_out[9257] & ~layer0_out[9256];
     layer1_out[7388] <= ~(layer0_out[3322] | layer0_out[3323]);
     layer1_out[7389] <= layer0_out[6035] & ~layer0_out[6036];
     layer1_out[7390] <= ~(layer0_out[5391] & layer0_out[5392]);
     layer1_out[7391] <= layer0_out[3611];
     layer1_out[7392] <= layer0_out[7780];
     layer1_out[7393] <= ~layer0_out[10402] | layer0_out[10401];
     layer1_out[7394] <= layer0_out[10750];
     layer1_out[7395] <= ~(layer0_out[628] | layer0_out[629]);
     layer1_out[7396] <= ~layer0_out[7112] | layer0_out[7111];
     layer1_out[7397] <= layer0_out[10305] & layer0_out[10306];
     layer1_out[7398] <= layer0_out[6125] & ~layer0_out[6124];
     layer1_out[7399] <= layer0_out[11010];
     layer1_out[7400] <= ~layer0_out[2845];
     layer1_out[7401] <= ~(layer0_out[4323] & layer0_out[4324]);
     layer1_out[7402] <= ~layer0_out[5452];
     layer1_out[7403] <= layer0_out[1564] & ~layer0_out[1565];
     layer1_out[7404] <= ~layer0_out[9519];
     layer1_out[7405] <= layer0_out[3216] & layer0_out[3217];
     layer1_out[7406] <= layer0_out[1972] & ~layer0_out[1973];
     layer1_out[7407] <= ~layer0_out[10989] | layer0_out[10990];
     layer1_out[7408] <= ~(layer0_out[6231] | layer0_out[6232]);
     layer1_out[7409] <= 1'b0;
     layer1_out[7410] <= ~layer0_out[1701];
     layer1_out[7411] <= ~layer0_out[1816];
     layer1_out[7412] <= ~layer0_out[10954] | layer0_out[10955];
     layer1_out[7413] <= ~(layer0_out[4918] & layer0_out[4919]);
     layer1_out[7414] <= layer0_out[9929];
     layer1_out[7415] <= layer0_out[9701] & layer0_out[9702];
     layer1_out[7416] <= layer0_out[11663] ^ layer0_out[11664];
     layer1_out[7417] <= layer0_out[6968] & layer0_out[6969];
     layer1_out[7418] <= layer0_out[9376] & ~layer0_out[9375];
     layer1_out[7419] <= layer0_out[1088];
     layer1_out[7420] <= layer0_out[4786] & layer0_out[4787];
     layer1_out[7421] <= ~layer0_out[8210] | layer0_out[8211];
     layer1_out[7422] <= ~layer0_out[8604];
     layer1_out[7423] <= ~layer0_out[339];
     layer1_out[7424] <= layer0_out[10310] & ~layer0_out[10311];
     layer1_out[7425] <= ~layer0_out[6384];
     layer1_out[7426] <= ~layer0_out[5017];
     layer1_out[7427] <= ~(layer0_out[7365] | layer0_out[7366]);
     layer1_out[7428] <= layer0_out[11314] | layer0_out[11315];
     layer1_out[7429] <= ~layer0_out[10692] | layer0_out[10693];
     layer1_out[7430] <= layer0_out[11002];
     layer1_out[7431] <= ~(layer0_out[2457] ^ layer0_out[2458]);
     layer1_out[7432] <= layer0_out[5119] & ~layer0_out[5120];
     layer1_out[7433] <= layer0_out[8011];
     layer1_out[7434] <= layer0_out[11076] | layer0_out[11077];
     layer1_out[7435] <= ~layer0_out[9565] | layer0_out[9566];
     layer1_out[7436] <= layer0_out[11441];
     layer1_out[7437] <= ~layer0_out[4110];
     layer1_out[7438] <= layer0_out[778] & layer0_out[779];
     layer1_out[7439] <= ~layer0_out[7889];
     layer1_out[7440] <= layer0_out[4010];
     layer1_out[7441] <= ~layer0_out[1792];
     layer1_out[7442] <= ~layer0_out[8383] | layer0_out[8384];
     layer1_out[7443] <= layer0_out[9080] | layer0_out[9081];
     layer1_out[7444] <= ~(layer0_out[4563] & layer0_out[4564]);
     layer1_out[7445] <= layer0_out[5963] & ~layer0_out[5964];
     layer1_out[7446] <= layer0_out[8604] & ~layer0_out[8603];
     layer1_out[7447] <= ~layer0_out[3861] | layer0_out[3862];
     layer1_out[7448] <= layer0_out[8326] & ~layer0_out[8325];
     layer1_out[7449] <= ~(layer0_out[6785] & layer0_out[6786]);
     layer1_out[7450] <= layer0_out[7585] & ~layer0_out[7586];
     layer1_out[7451] <= layer0_out[3028] & ~layer0_out[3027];
     layer1_out[7452] <= ~layer0_out[7639] | layer0_out[7638];
     layer1_out[7453] <= ~(layer0_out[10020] | layer0_out[10021]);
     layer1_out[7454] <= layer0_out[7233];
     layer1_out[7455] <= ~(layer0_out[11413] & layer0_out[11414]);
     layer1_out[7456] <= layer0_out[9144];
     layer1_out[7457] <= ~(layer0_out[6280] | layer0_out[6281]);
     layer1_out[7458] <= layer0_out[9603] & ~layer0_out[9604];
     layer1_out[7459] <= layer0_out[6493];
     layer1_out[7460] <= layer0_out[2466] & layer0_out[2467];
     layer1_out[7461] <= layer0_out[7977] & ~layer0_out[7976];
     layer1_out[7462] <= ~layer0_out[10764];
     layer1_out[7463] <= layer0_out[7815] | layer0_out[7816];
     layer1_out[7464] <= ~(layer0_out[5518] & layer0_out[5519]);
     layer1_out[7465] <= layer0_out[3990];
     layer1_out[7466] <= ~layer0_out[1076];
     layer1_out[7467] <= layer0_out[1898] ^ layer0_out[1899];
     layer1_out[7468] <= layer0_out[4357];
     layer1_out[7469] <= ~layer0_out[1520] | layer0_out[1521];
     layer1_out[7470] <= layer0_out[4355] & layer0_out[4356];
     layer1_out[7471] <= ~layer0_out[4785];
     layer1_out[7472] <= ~layer0_out[2238];
     layer1_out[7473] <= ~layer0_out[3742];
     layer1_out[7474] <= ~layer0_out[11224];
     layer1_out[7475] <= ~layer0_out[1895];
     layer1_out[7476] <= ~layer0_out[2808];
     layer1_out[7477] <= layer0_out[7384] & ~layer0_out[7385];
     layer1_out[7478] <= layer0_out[7826];
     layer1_out[7479] <= ~layer0_out[3832];
     layer1_out[7480] <= layer0_out[6102];
     layer1_out[7481] <= layer0_out[5226] | layer0_out[5227];
     layer1_out[7482] <= layer0_out[4196] ^ layer0_out[4197];
     layer1_out[7483] <= layer0_out[4286] & ~layer0_out[4287];
     layer1_out[7484] <= layer0_out[11895] ^ layer0_out[11896];
     layer1_out[7485] <= layer0_out[7891] | layer0_out[7892];
     layer1_out[7486] <= ~layer0_out[4027] | layer0_out[4026];
     layer1_out[7487] <= ~layer0_out[11130] | layer0_out[11129];
     layer1_out[7488] <= layer0_out[10254] & ~layer0_out[10255];
     layer1_out[7489] <= ~layer0_out[9224];
     layer1_out[7490] <= layer0_out[1092];
     layer1_out[7491] <= ~layer0_out[7048];
     layer1_out[7492] <= layer0_out[309];
     layer1_out[7493] <= ~layer0_out[6360];
     layer1_out[7494] <= ~layer0_out[6470];
     layer1_out[7495] <= layer0_out[7339];
     layer1_out[7496] <= 1'b0;
     layer1_out[7497] <= ~layer0_out[8456] | layer0_out[8457];
     layer1_out[7498] <= ~(layer0_out[5075] | layer0_out[5076]);
     layer1_out[7499] <= layer0_out[11896] | layer0_out[11897];
     layer1_out[7500] <= ~layer0_out[8614];
     layer1_out[7501] <= ~layer0_out[891] | layer0_out[890];
     layer1_out[7502] <= ~layer0_out[2637];
     layer1_out[7503] <= ~layer0_out[4722];
     layer1_out[7504] <= layer0_out[6994] | layer0_out[6995];
     layer1_out[7505] <= layer0_out[8072] & layer0_out[8073];
     layer1_out[7506] <= layer0_out[6033] ^ layer0_out[6034];
     layer1_out[7507] <= layer0_out[502] & ~layer0_out[501];
     layer1_out[7508] <= ~(layer0_out[188] | layer0_out[189]);
     layer1_out[7509] <= ~layer0_out[1375];
     layer1_out[7510] <= layer0_out[10048] & ~layer0_out[10049];
     layer1_out[7511] <= layer0_out[5774] & layer0_out[5775];
     layer1_out[7512] <= ~layer0_out[9678] | layer0_out[9677];
     layer1_out[7513] <= ~(layer0_out[9166] ^ layer0_out[9167]);
     layer1_out[7514] <= ~layer0_out[6251] | layer0_out[6252];
     layer1_out[7515] <= layer0_out[3960];
     layer1_out[7516] <= ~(layer0_out[4176] | layer0_out[4177]);
     layer1_out[7517] <= ~layer0_out[11969];
     layer1_out[7518] <= ~layer0_out[2177];
     layer1_out[7519] <= ~layer0_out[619];
     layer1_out[7520] <= layer0_out[7968] | layer0_out[7969];
     layer1_out[7521] <= layer0_out[2348];
     layer1_out[7522] <= layer0_out[8602] & ~layer0_out[8603];
     layer1_out[7523] <= ~layer0_out[525] | layer0_out[524];
     layer1_out[7524] <= layer0_out[9688] & ~layer0_out[9687];
     layer1_out[7525] <= ~layer0_out[5289];
     layer1_out[7526] <= layer0_out[7380] & layer0_out[7381];
     layer1_out[7527] <= layer0_out[7570] & ~layer0_out[7571];
     layer1_out[7528] <= ~(layer0_out[5211] & layer0_out[5212]);
     layer1_out[7529] <= ~(layer0_out[6580] & layer0_out[6581]);
     layer1_out[7530] <= ~layer0_out[2512];
     layer1_out[7531] <= layer0_out[5760] ^ layer0_out[5761];
     layer1_out[7532] <= layer0_out[10774] & ~layer0_out[10773];
     layer1_out[7533] <= layer0_out[8126];
     layer1_out[7534] <= layer0_out[10237] & layer0_out[10238];
     layer1_out[7535] <= layer0_out[2570] | layer0_out[2571];
     layer1_out[7536] <= ~layer0_out[865] | layer0_out[866];
     layer1_out[7537] <= layer0_out[1835];
     layer1_out[7538] <= ~layer0_out[6343] | layer0_out[6342];
     layer1_out[7539] <= layer0_out[5609] & ~layer0_out[5610];
     layer1_out[7540] <= layer0_out[6996] & layer0_out[6997];
     layer1_out[7541] <= layer0_out[11515] & ~layer0_out[11516];
     layer1_out[7542] <= layer0_out[10337];
     layer1_out[7543] <= ~layer0_out[9040];
     layer1_out[7544] <= layer0_out[6730] & layer0_out[6731];
     layer1_out[7545] <= layer0_out[3756] & ~layer0_out[3755];
     layer1_out[7546] <= ~layer0_out[9157];
     layer1_out[7547] <= ~layer0_out[9669] | layer0_out[9670];
     layer1_out[7548] <= ~layer0_out[801] | layer0_out[802];
     layer1_out[7549] <= ~(layer0_out[8433] ^ layer0_out[8434]);
     layer1_out[7550] <= ~(layer0_out[11981] | layer0_out[11982]);
     layer1_out[7551] <= ~(layer0_out[11197] & layer0_out[11198]);
     layer1_out[7552] <= layer0_out[8188];
     layer1_out[7553] <= ~(layer0_out[2533] & layer0_out[2534]);
     layer1_out[7554] <= layer0_out[1643] | layer0_out[1644];
     layer1_out[7555] <= ~layer0_out[2811] | layer0_out[2810];
     layer1_out[7556] <= ~layer0_out[11308];
     layer1_out[7557] <= layer0_out[10174];
     layer1_out[7558] <= ~layer0_out[31] | layer0_out[30];
     layer1_out[7559] <= ~(layer0_out[4438] & layer0_out[4439]);
     layer1_out[7560] <= layer0_out[10900];
     layer1_out[7561] <= ~layer0_out[7416] | layer0_out[7415];
     layer1_out[7562] <= 1'b0;
     layer1_out[7563] <= layer0_out[5616] & ~layer0_out[5615];
     layer1_out[7564] <= layer0_out[6632];
     layer1_out[7565] <= layer0_out[11686] & ~layer0_out[11687];
     layer1_out[7566] <= layer0_out[8613] & layer0_out[8614];
     layer1_out[7567] <= ~layer0_out[9534] | layer0_out[9535];
     layer1_out[7568] <= layer0_out[4539] & ~layer0_out[4540];
     layer1_out[7569] <= layer0_out[3493];
     layer1_out[7570] <= layer0_out[1983] & ~layer0_out[1982];
     layer1_out[7571] <= ~layer0_out[7362] | layer0_out[7361];
     layer1_out[7572] <= ~layer0_out[8921];
     layer1_out[7573] <= layer0_out[7061];
     layer1_out[7574] <= layer0_out[2251];
     layer1_out[7575] <= layer0_out[10391] & ~layer0_out[10392];
     layer1_out[7576] <= layer0_out[8173] & layer0_out[8174];
     layer1_out[7577] <= layer0_out[6727] ^ layer0_out[6728];
     layer1_out[7578] <= ~layer0_out[5709];
     layer1_out[7579] <= layer0_out[7989] & ~layer0_out[7990];
     layer1_out[7580] <= ~(layer0_out[11247] | layer0_out[11248]);
     layer1_out[7581] <= ~(layer0_out[1433] & layer0_out[1434]);
     layer1_out[7582] <= ~layer0_out[3404] | layer0_out[3403];
     layer1_out[7583] <= layer0_out[6371] | layer0_out[6372];
     layer1_out[7584] <= layer0_out[8174];
     layer1_out[7585] <= ~(layer0_out[10176] & layer0_out[10177]);
     layer1_out[7586] <= ~layer0_out[10088];
     layer1_out[7587] <= ~layer0_out[2259] | layer0_out[2258];
     layer1_out[7588] <= layer0_out[7713] & ~layer0_out[7714];
     layer1_out[7589] <= ~(layer0_out[9290] ^ layer0_out[9291]);
     layer1_out[7590] <= ~layer0_out[7142];
     layer1_out[7591] <= layer0_out[4072];
     layer1_out[7592] <= ~layer0_out[11519];
     layer1_out[7593] <= layer0_out[4394];
     layer1_out[7594] <= ~layer0_out[4858] | layer0_out[4859];
     layer1_out[7595] <= ~layer0_out[11926] | layer0_out[11925];
     layer1_out[7596] <= layer0_out[7725] & layer0_out[7726];
     layer1_out[7597] <= ~(layer0_out[2778] | layer0_out[2779]);
     layer1_out[7598] <= 1'b1;
     layer1_out[7599] <= ~(layer0_out[5720] & layer0_out[5721]);
     layer1_out[7600] <= layer0_out[11894];
     layer1_out[7601] <= ~(layer0_out[1679] & layer0_out[1680]);
     layer1_out[7602] <= ~layer0_out[10165] | layer0_out[10166];
     layer1_out[7603] <= layer0_out[4979] & ~layer0_out[4978];
     layer1_out[7604] <= layer0_out[11977];
     layer1_out[7605] <= layer0_out[4157] & layer0_out[4158];
     layer1_out[7606] <= ~layer0_out[11948] | layer0_out[11949];
     layer1_out[7607] <= layer0_out[366] ^ layer0_out[367];
     layer1_out[7608] <= ~layer0_out[4639];
     layer1_out[7609] <= layer0_out[9467] & ~layer0_out[9466];
     layer1_out[7610] <= layer0_out[2833] & ~layer0_out[2834];
     layer1_out[7611] <= layer0_out[5852];
     layer1_out[7612] <= layer0_out[11262] & layer0_out[11263];
     layer1_out[7613] <= ~layer0_out[7792];
     layer1_out[7614] <= ~layer0_out[9008];
     layer1_out[7615] <= layer0_out[6684] & ~layer0_out[6685];
     layer1_out[7616] <= layer0_out[4926];
     layer1_out[7617] <= layer0_out[8367];
     layer1_out[7618] <= ~layer0_out[7532];
     layer1_out[7619] <= ~layer0_out[3028] | layer0_out[3029];
     layer1_out[7620] <= layer0_out[7846] | layer0_out[7847];
     layer1_out[7621] <= ~layer0_out[1634];
     layer1_out[7622] <= layer0_out[11889] & ~layer0_out[11890];
     layer1_out[7623] <= layer0_out[7258] & ~layer0_out[7257];
     layer1_out[7624] <= layer0_out[8188] | layer0_out[8189];
     layer1_out[7625] <= ~layer0_out[1047] | layer0_out[1046];
     layer1_out[7626] <= ~layer0_out[699] | layer0_out[698];
     layer1_out[7627] <= layer0_out[10960] ^ layer0_out[10961];
     layer1_out[7628] <= ~layer0_out[10568] | layer0_out[10567];
     layer1_out[7629] <= ~layer0_out[2115] | layer0_out[2116];
     layer1_out[7630] <= ~layer0_out[6272];
     layer1_out[7631] <= layer0_out[863] & ~layer0_out[862];
     layer1_out[7632] <= layer0_out[9398] & ~layer0_out[9399];
     layer1_out[7633] <= ~(layer0_out[10851] & layer0_out[10852]);
     layer1_out[7634] <= ~(layer0_out[9646] | layer0_out[9647]);
     layer1_out[7635] <= ~layer0_out[4198] | layer0_out[4197];
     layer1_out[7636] <= layer0_out[5680];
     layer1_out[7637] <= layer0_out[4150] & layer0_out[4151];
     layer1_out[7638] <= layer0_out[8996];
     layer1_out[7639] <= layer0_out[3541];
     layer1_out[7640] <= ~layer0_out[2627];
     layer1_out[7641] <= ~layer0_out[5356] | layer0_out[5357];
     layer1_out[7642] <= ~layer0_out[5054] | layer0_out[5055];
     layer1_out[7643] <= layer0_out[5273];
     layer1_out[7644] <= layer0_out[4987] ^ layer0_out[4988];
     layer1_out[7645] <= layer0_out[6758];
     layer1_out[7646] <= ~(layer0_out[8405] & layer0_out[8406]);
     layer1_out[7647] <= ~layer0_out[842];
     layer1_out[7648] <= layer0_out[9411] | layer0_out[9412];
     layer1_out[7649] <= ~layer0_out[8062];
     layer1_out[7650] <= layer0_out[10000];
     layer1_out[7651] <= ~(layer0_out[8885] | layer0_out[8886]);
     layer1_out[7652] <= ~(layer0_out[3093] ^ layer0_out[3094]);
     layer1_out[7653] <= layer0_out[332];
     layer1_out[7654] <= layer0_out[324] & ~layer0_out[323];
     layer1_out[7655] <= ~layer0_out[3223];
     layer1_out[7656] <= ~(layer0_out[622] | layer0_out[623]);
     layer1_out[7657] <= layer0_out[4076] & ~layer0_out[4077];
     layer1_out[7658] <= ~layer0_out[6625];
     layer1_out[7659] <= layer0_out[3114];
     layer1_out[7660] <= layer0_out[2020] & ~layer0_out[2021];
     layer1_out[7661] <= layer0_out[1235] & ~layer0_out[1234];
     layer1_out[7662] <= layer0_out[3320];
     layer1_out[7663] <= layer0_out[866] ^ layer0_out[867];
     layer1_out[7664] <= ~layer0_out[6717];
     layer1_out[7665] <= ~(layer0_out[7403] & layer0_out[7404]);
     layer1_out[7666] <= layer0_out[3423] & ~layer0_out[3422];
     layer1_out[7667] <= layer0_out[3450];
     layer1_out[7668] <= layer0_out[9415];
     layer1_out[7669] <= layer0_out[5709] ^ layer0_out[5710];
     layer1_out[7670] <= 1'b0;
     layer1_out[7671] <= ~layer0_out[5038];
     layer1_out[7672] <= layer0_out[7169] ^ layer0_out[7170];
     layer1_out[7673] <= ~(layer0_out[8050] | layer0_out[8051]);
     layer1_out[7674] <= layer0_out[10782] & ~layer0_out[10781];
     layer1_out[7675] <= layer0_out[8798] & ~layer0_out[8797];
     layer1_out[7676] <= ~layer0_out[5524];
     layer1_out[7677] <= layer0_out[9489];
     layer1_out[7678] <= ~layer0_out[8466];
     layer1_out[7679] <= ~layer0_out[7718];
     layer1_out[7680] <= ~layer0_out[6248];
     layer1_out[7681] <= layer0_out[7572];
     layer1_out[7682] <= layer0_out[6319] | layer0_out[6320];
     layer1_out[7683] <= layer0_out[3374] | layer0_out[3375];
     layer1_out[7684] <= layer0_out[397];
     layer1_out[7685] <= layer0_out[7526] | layer0_out[7527];
     layer1_out[7686] <= ~layer0_out[6928] | layer0_out[6929];
     layer1_out[7687] <= ~layer0_out[6367];
     layer1_out[7688] <= ~layer0_out[6952];
     layer1_out[7689] <= layer0_out[2321];
     layer1_out[7690] <= ~layer0_out[3681];
     layer1_out[7691] <= ~layer0_out[3753] | layer0_out[3754];
     layer1_out[7692] <= layer0_out[1922];
     layer1_out[7693] <= layer0_out[6579];
     layer1_out[7694] <= layer0_out[5818];
     layer1_out[7695] <= ~(layer0_out[5556] | layer0_out[5557]);
     layer1_out[7696] <= ~layer0_out[10515] | layer0_out[10514];
     layer1_out[7697] <= layer0_out[7791];
     layer1_out[7698] <= ~(layer0_out[2163] | layer0_out[2164]);
     layer1_out[7699] <= ~(layer0_out[4228] & layer0_out[4229]);
     layer1_out[7700] <= layer0_out[7885] | layer0_out[7886];
     layer1_out[7701] <= layer0_out[5722];
     layer1_out[7702] <= layer0_out[1094] & ~layer0_out[1095];
     layer1_out[7703] <= 1'b1;
     layer1_out[7704] <= ~(layer0_out[7906] | layer0_out[7907]);
     layer1_out[7705] <= layer0_out[10829];
     layer1_out[7706] <= layer0_out[6554] ^ layer0_out[6555];
     layer1_out[7707] <= layer0_out[7481];
     layer1_out[7708] <= ~(layer0_out[8580] | layer0_out[8581]);
     layer1_out[7709] <= ~layer0_out[691];
     layer1_out[7710] <= layer0_out[11485] & ~layer0_out[11484];
     layer1_out[7711] <= layer0_out[3880] ^ layer0_out[3881];
     layer1_out[7712] <= ~layer0_out[8905] | layer0_out[8904];
     layer1_out[7713] <= layer0_out[10335];
     layer1_out[7714] <= layer0_out[8107] & ~layer0_out[8108];
     layer1_out[7715] <= layer0_out[11359];
     layer1_out[7716] <= layer0_out[4337] & layer0_out[4338];
     layer1_out[7717] <= layer0_out[9221] & ~layer0_out[9220];
     layer1_out[7718] <= layer0_out[717] | layer0_out[718];
     layer1_out[7719] <= layer0_out[10365];
     layer1_out[7720] <= ~layer0_out[7101];
     layer1_out[7721] <= ~layer0_out[10940];
     layer1_out[7722] <= ~(layer0_out[2787] & layer0_out[2788]);
     layer1_out[7723] <= ~layer0_out[11292] | layer0_out[11291];
     layer1_out[7724] <= ~(layer0_out[10925] | layer0_out[10926]);
     layer1_out[7725] <= 1'b0;
     layer1_out[7726] <= layer0_out[2795] & ~layer0_out[2794];
     layer1_out[7727] <= ~layer0_out[10225];
     layer1_out[7728] <= layer0_out[11301];
     layer1_out[7729] <= layer0_out[10107] & layer0_out[10108];
     layer1_out[7730] <= layer0_out[10515] | layer0_out[10516];
     layer1_out[7731] <= ~layer0_out[2181];
     layer1_out[7732] <= ~layer0_out[11592];
     layer1_out[7733] <= 1'b0;
     layer1_out[7734] <= layer0_out[1351] & layer0_out[1352];
     layer1_out[7735] <= ~layer0_out[2243] | layer0_out[2244];
     layer1_out[7736] <= ~layer0_out[3275];
     layer1_out[7737] <= ~layer0_out[4895];
     layer1_out[7738] <= ~(layer0_out[6884] & layer0_out[6885]);
     layer1_out[7739] <= layer0_out[3553];
     layer1_out[7740] <= ~(layer0_out[11646] & layer0_out[11647]);
     layer1_out[7741] <= ~layer0_out[1403];
     layer1_out[7742] <= ~layer0_out[5661] | layer0_out[5660];
     layer1_out[7743] <= layer0_out[433] | layer0_out[434];
     layer1_out[7744] <= layer0_out[5499] & ~layer0_out[5500];
     layer1_out[7745] <= layer0_out[2530] & layer0_out[2531];
     layer1_out[7746] <= layer0_out[2016];
     layer1_out[7747] <= layer0_out[3937] & layer0_out[3938];
     layer1_out[7748] <= ~layer0_out[511];
     layer1_out[7749] <= ~layer0_out[6623];
     layer1_out[7750] <= layer0_out[211];
     layer1_out[7751] <= ~(layer0_out[8890] & layer0_out[8891]);
     layer1_out[7752] <= ~(layer0_out[3902] | layer0_out[3903]);
     layer1_out[7753] <= layer0_out[7337] ^ layer0_out[7338];
     layer1_out[7754] <= 1'b1;
     layer1_out[7755] <= ~layer0_out[1679];
     layer1_out[7756] <= ~(layer0_out[5336] ^ layer0_out[5337]);
     layer1_out[7757] <= layer0_out[823];
     layer1_out[7758] <= layer0_out[3580] & layer0_out[3581];
     layer1_out[7759] <= ~(layer0_out[5559] | layer0_out[5560]);
     layer1_out[7760] <= ~layer0_out[3939] | layer0_out[3938];
     layer1_out[7761] <= ~layer0_out[9064];
     layer1_out[7762] <= layer0_out[615] | layer0_out[616];
     layer1_out[7763] <= ~layer0_out[3734] | layer0_out[3735];
     layer1_out[7764] <= layer0_out[1537] & ~layer0_out[1536];
     layer1_out[7765] <= layer0_out[1937] & ~layer0_out[1938];
     layer1_out[7766] <= ~layer0_out[9354] | layer0_out[9353];
     layer1_out[7767] <= ~(layer0_out[11160] | layer0_out[11161]);
     layer1_out[7768] <= layer0_out[1810];
     layer1_out[7769] <= layer0_out[6418] & ~layer0_out[6417];
     layer1_out[7770] <= layer0_out[9113];
     layer1_out[7771] <= layer0_out[1694] ^ layer0_out[1695];
     layer1_out[7772] <= layer0_out[5367];
     layer1_out[7773] <= 1'b1;
     layer1_out[7774] <= ~(layer0_out[3187] | layer0_out[3188]);
     layer1_out[7775] <= layer0_out[5828] & ~layer0_out[5829];
     layer1_out[7776] <= ~layer0_out[5358] | layer0_out[5359];
     layer1_out[7777] <= ~layer0_out[7659];
     layer1_out[7778] <= layer0_out[10233];
     layer1_out[7779] <= ~layer0_out[4903];
     layer1_out[7780] <= layer0_out[8667] | layer0_out[8668];
     layer1_out[7781] <= ~layer0_out[9687];
     layer1_out[7782] <= layer0_out[6278] & ~layer0_out[6277];
     layer1_out[7783] <= 1'b0;
     layer1_out[7784] <= layer0_out[6544] & ~layer0_out[6545];
     layer1_out[7785] <= ~(layer0_out[8374] & layer0_out[8375]);
     layer1_out[7786] <= layer0_out[4915] | layer0_out[4916];
     layer1_out[7787] <= ~layer0_out[2034] | layer0_out[2035];
     layer1_out[7788] <= ~layer0_out[3495];
     layer1_out[7789] <= ~layer0_out[5336];
     layer1_out[7790] <= layer0_out[7115] & layer0_out[7116];
     layer1_out[7791] <= layer0_out[1070] | layer0_out[1071];
     layer1_out[7792] <= ~layer0_out[1944];
     layer1_out[7793] <= ~layer0_out[653] | layer0_out[654];
     layer1_out[7794] <= layer0_out[7461] & ~layer0_out[7462];
     layer1_out[7795] <= ~(layer0_out[2134] & layer0_out[2135]);
     layer1_out[7796] <= ~(layer0_out[5142] | layer0_out[5143]);
     layer1_out[7797] <= ~layer0_out[4588];
     layer1_out[7798] <= ~layer0_out[4341] | layer0_out[4340];
     layer1_out[7799] <= layer0_out[486];
     layer1_out[7800] <= ~layer0_out[6514] | layer0_out[6513];
     layer1_out[7801] <= layer0_out[3369] & layer0_out[3370];
     layer1_out[7802] <= layer0_out[9690] ^ layer0_out[9691];
     layer1_out[7803] <= ~layer0_out[301] | layer0_out[300];
     layer1_out[7804] <= layer0_out[1426] ^ layer0_out[1427];
     layer1_out[7805] <= ~layer0_out[4628];
     layer1_out[7806] <= ~layer0_out[9897] | layer0_out[9898];
     layer1_out[7807] <= ~layer0_out[2432];
     layer1_out[7808] <= layer0_out[2252];
     layer1_out[7809] <= layer0_out[1290] & layer0_out[1291];
     layer1_out[7810] <= layer0_out[2171] | layer0_out[2172];
     layer1_out[7811] <= ~(layer0_out[9378] | layer0_out[9379]);
     layer1_out[7812] <= layer0_out[355] & ~layer0_out[356];
     layer1_out[7813] <= layer0_out[9699] | layer0_out[9700];
     layer1_out[7814] <= layer0_out[9917];
     layer1_out[7815] <= ~layer0_out[11388];
     layer1_out[7816] <= ~layer0_out[6511];
     layer1_out[7817] <= ~layer0_out[11001] | layer0_out[11002];
     layer1_out[7818] <= layer0_out[8655];
     layer1_out[7819] <= ~layer0_out[2718];
     layer1_out[7820] <= ~layer0_out[5807];
     layer1_out[7821] <= layer0_out[3571] & layer0_out[3572];
     layer1_out[7822] <= layer0_out[9101] ^ layer0_out[9102];
     layer1_out[7823] <= layer0_out[8876];
     layer1_out[7824] <= layer0_out[7446];
     layer1_out[7825] <= layer0_out[8316];
     layer1_out[7826] <= ~layer0_out[9590];
     layer1_out[7827] <= layer0_out[7387];
     layer1_out[7828] <= ~(layer0_out[7332] | layer0_out[7333]);
     layer1_out[7829] <= ~(layer0_out[8932] ^ layer0_out[8933]);
     layer1_out[7830] <= ~layer0_out[703] | layer0_out[704];
     layer1_out[7831] <= ~layer0_out[2942] | layer0_out[2943];
     layer1_out[7832] <= layer0_out[9225] & ~layer0_out[9226];
     layer1_out[7833] <= ~layer0_out[11238];
     layer1_out[7834] <= layer0_out[1625];
     layer1_out[7835] <= layer0_out[4954];
     layer1_out[7836] <= ~layer0_out[614];
     layer1_out[7837] <= ~(layer0_out[5948] ^ layer0_out[5949]);
     layer1_out[7838] <= layer0_out[57];
     layer1_out[7839] <= ~layer0_out[2801] | layer0_out[2802];
     layer1_out[7840] <= layer0_out[3007] | layer0_out[3008];
     layer1_out[7841] <= ~(layer0_out[8292] | layer0_out[8293]);
     layer1_out[7842] <= ~(layer0_out[5676] & layer0_out[5677]);
     layer1_out[7843] <= ~layer0_out[2687];
     layer1_out[7844] <= layer0_out[8061];
     layer1_out[7845] <= layer0_out[8410];
     layer1_out[7846] <= ~layer0_out[11801];
     layer1_out[7847] <= layer0_out[10082] | layer0_out[10083];
     layer1_out[7848] <= layer0_out[8505] & layer0_out[8506];
     layer1_out[7849] <= layer0_out[6983];
     layer1_out[7850] <= layer0_out[3433] & ~layer0_out[3434];
     layer1_out[7851] <= layer0_out[11567];
     layer1_out[7852] <= layer0_out[4029];
     layer1_out[7853] <= layer0_out[1256] | layer0_out[1257];
     layer1_out[7854] <= ~layer0_out[1951];
     layer1_out[7855] <= ~layer0_out[3800];
     layer1_out[7856] <= layer0_out[5444] & ~layer0_out[5445];
     layer1_out[7857] <= 1'b1;
     layer1_out[7858] <= ~layer0_out[9418] | layer0_out[9417];
     layer1_out[7859] <= ~layer0_out[1784] | layer0_out[1785];
     layer1_out[7860] <= ~(layer0_out[18] | layer0_out[19]);
     layer1_out[7861] <= layer0_out[8064] & ~layer0_out[8065];
     layer1_out[7862] <= ~layer0_out[9692];
     layer1_out[7863] <= ~layer0_out[10270] | layer0_out[10269];
     layer1_out[7864] <= ~layer0_out[10827];
     layer1_out[7865] <= ~(layer0_out[8978] | layer0_out[8979]);
     layer1_out[7866] <= layer0_out[10684] & ~layer0_out[10685];
     layer1_out[7867] <= ~layer0_out[821];
     layer1_out[7868] <= layer0_out[7514];
     layer1_out[7869] <= 1'b1;
     layer1_out[7870] <= layer0_out[9641];
     layer1_out[7871] <= layer0_out[4304] | layer0_out[4305];
     layer1_out[7872] <= ~(layer0_out[11313] & layer0_out[11314]);
     layer1_out[7873] <= layer0_out[7118] & ~layer0_out[7117];
     layer1_out[7874] <= layer0_out[9258] & ~layer0_out[9259];
     layer1_out[7875] <= layer0_out[3483] & layer0_out[3484];
     layer1_out[7876] <= ~(layer0_out[11929] & layer0_out[11930]);
     layer1_out[7877] <= layer0_out[593] & layer0_out[594];
     layer1_out[7878] <= 1'b0;
     layer1_out[7879] <= ~(layer0_out[1112] ^ layer0_out[1113]);
     layer1_out[7880] <= layer0_out[11474] | layer0_out[11475];
     layer1_out[7881] <= ~(layer0_out[8301] | layer0_out[8302]);
     layer1_out[7882] <= ~(layer0_out[3041] ^ layer0_out[3042]);
     layer1_out[7883] <= ~(layer0_out[10984] ^ layer0_out[10985]);
     layer1_out[7884] <= layer0_out[6661];
     layer1_out[7885] <= ~(layer0_out[1734] & layer0_out[1735]);
     layer1_out[7886] <= layer0_out[3487] & ~layer0_out[3488];
     layer1_out[7887] <= layer0_out[1238] ^ layer0_out[1239];
     layer1_out[7888] <= layer0_out[30];
     layer1_out[7889] <= ~layer0_out[8031] | layer0_out[8030];
     layer1_out[7890] <= ~(layer0_out[2423] ^ layer0_out[2424]);
     layer1_out[7891] <= layer0_out[8609] & ~layer0_out[8610];
     layer1_out[7892] <= layer0_out[7302] & layer0_out[7303];
     layer1_out[7893] <= ~layer0_out[7924];
     layer1_out[7894] <= layer0_out[4370];
     layer1_out[7895] <= ~(layer0_out[11838] & layer0_out[11839]);
     layer1_out[7896] <= ~layer0_out[6385];
     layer1_out[7897] <= ~layer0_out[4379] | layer0_out[4378];
     layer1_out[7898] <= layer0_out[2332];
     layer1_out[7899] <= layer0_out[11142];
     layer1_out[7900] <= ~layer0_out[309];
     layer1_out[7901] <= ~(layer0_out[2046] | layer0_out[2047]);
     layer1_out[7902] <= layer0_out[4641] & layer0_out[4642];
     layer1_out[7903] <= layer0_out[3329] & ~layer0_out[3330];
     layer1_out[7904] <= ~(layer0_out[624] & layer0_out[625]);
     layer1_out[7905] <= layer0_out[11191];
     layer1_out[7906] <= ~(layer0_out[5076] | layer0_out[5077]);
     layer1_out[7907] <= layer0_out[5992] | layer0_out[5993];
     layer1_out[7908] <= layer0_out[165];
     layer1_out[7909] <= layer0_out[3919] ^ layer0_out[3920];
     layer1_out[7910] <= ~(layer0_out[6275] & layer0_out[6276]);
     layer1_out[7911] <= layer0_out[292] | layer0_out[293];
     layer1_out[7912] <= ~layer0_out[4824] | layer0_out[4823];
     layer1_out[7913] <= 1'b1;
     layer1_out[7914] <= ~layer0_out[9088];
     layer1_out[7915] <= 1'b0;
     layer1_out[7916] <= 1'b0;
     layer1_out[7917] <= layer0_out[6146];
     layer1_out[7918] <= layer0_out[1147];
     layer1_out[7919] <= layer0_out[10364] | layer0_out[10365];
     layer1_out[7920] <= ~layer0_out[7911] | layer0_out[7912];
     layer1_out[7921] <= 1'b0;
     layer1_out[7922] <= ~(layer0_out[894] & layer0_out[895]);
     layer1_out[7923] <= layer0_out[9735] ^ layer0_out[9736];
     layer1_out[7924] <= layer0_out[11764] & ~layer0_out[11765];
     layer1_out[7925] <= ~layer0_out[3175];
     layer1_out[7926] <= 1'b1;
     layer1_out[7927] <= layer0_out[1781];
     layer1_out[7928] <= layer0_out[2158];
     layer1_out[7929] <= layer0_out[3997] | layer0_out[3998];
     layer1_out[7930] <= ~layer0_out[10855];
     layer1_out[7931] <= ~layer0_out[11869];
     layer1_out[7932] <= layer0_out[6243] & ~layer0_out[6244];
     layer1_out[7933] <= ~layer0_out[4726] | layer0_out[4727];
     layer1_out[7934] <= layer0_out[2008] & ~layer0_out[2007];
     layer1_out[7935] <= 1'b0;
     layer1_out[7936] <= 1'b0;
     layer1_out[7937] <= layer0_out[3000];
     layer1_out[7938] <= layer0_out[9822];
     layer1_out[7939] <= layer0_out[11636];
     layer1_out[7940] <= ~layer0_out[4236];
     layer1_out[7941] <= 1'b1;
     layer1_out[7942] <= layer0_out[10545];
     layer1_out[7943] <= ~layer0_out[8617];
     layer1_out[7944] <= layer0_out[5065];
     layer1_out[7945] <= layer0_out[7226] & ~layer0_out[7227];
     layer1_out[7946] <= layer0_out[361];
     layer1_out[7947] <= ~(layer0_out[2727] ^ layer0_out[2728]);
     layer1_out[7948] <= ~layer0_out[2281];
     layer1_out[7949] <= ~(layer0_out[4629] | layer0_out[4630]);
     layer1_out[7950] <= layer0_out[4679];
     layer1_out[7951] <= ~(layer0_out[11157] & layer0_out[11158]);
     layer1_out[7952] <= layer0_out[6229] | layer0_out[6230];
     layer1_out[7953] <= layer0_out[7745] & ~layer0_out[7746];
     layer1_out[7954] <= layer0_out[8002] & layer0_out[8003];
     layer1_out[7955] <= layer0_out[3676] & ~layer0_out[3675];
     layer1_out[7956] <= ~layer0_out[1484] | layer0_out[1483];
     layer1_out[7957] <= layer0_out[9047] & ~layer0_out[9048];
     layer1_out[7958] <= layer0_out[7077] | layer0_out[7078];
     layer1_out[7959] <= layer0_out[2394] & layer0_out[2395];
     layer1_out[7960] <= layer0_out[538] & ~layer0_out[537];
     layer1_out[7961] <= layer0_out[2917] & layer0_out[2918];
     layer1_out[7962] <= ~(layer0_out[10239] | layer0_out[10240]);
     layer1_out[7963] <= layer0_out[11694];
     layer1_out[7964] <= ~layer0_out[3469];
     layer1_out[7965] <= ~layer0_out[10904];
     layer1_out[7966] <= ~layer0_out[8395];
     layer1_out[7967] <= layer0_out[10032];
     layer1_out[7968] <= ~layer0_out[4409];
     layer1_out[7969] <= layer0_out[8364] | layer0_out[8365];
     layer1_out[7970] <= ~(layer0_out[7897] & layer0_out[7898]);
     layer1_out[7971] <= ~(layer0_out[5590] & layer0_out[5591]);
     layer1_out[7972] <= ~layer0_out[918] | layer0_out[917];
     layer1_out[7973] <= ~layer0_out[335] | layer0_out[336];
     layer1_out[7974] <= layer0_out[2073];
     layer1_out[7975] <= layer0_out[185];
     layer1_out[7976] <= layer0_out[3128];
     layer1_out[7977] <= layer0_out[11349];
     layer1_out[7978] <= layer0_out[1626] & layer0_out[1627];
     layer1_out[7979] <= ~(layer0_out[2728] & layer0_out[2729]);
     layer1_out[7980] <= ~(layer0_out[10414] | layer0_out[10415]);
     layer1_out[7981] <= ~layer0_out[8109];
     layer1_out[7982] <= layer0_out[7342] | layer0_out[7343];
     layer1_out[7983] <= layer0_out[6226] & layer0_out[6227];
     layer1_out[7984] <= ~(layer0_out[746] ^ layer0_out[747]);
     layer1_out[7985] <= ~(layer0_out[4027] ^ layer0_out[4028]);
     layer1_out[7986] <= layer0_out[11182];
     layer1_out[7987] <= ~layer0_out[1241];
     layer1_out[7988] <= 1'b1;
     layer1_out[7989] <= layer0_out[8481];
     layer1_out[7990] <= ~(layer0_out[10229] & layer0_out[10230]);
     layer1_out[7991] <= layer0_out[2878] & ~layer0_out[2879];
     layer1_out[7992] <= layer0_out[3439] & layer0_out[3440];
     layer1_out[7993] <= ~layer0_out[10947];
     layer1_out[7994] <= ~(layer0_out[737] ^ layer0_out[738]);
     layer1_out[7995] <= ~layer0_out[3349] | layer0_out[3350];
     layer1_out[7996] <= layer0_out[11950];
     layer1_out[7997] <= layer0_out[7545];
     layer1_out[7998] <= 1'b0;
     layer1_out[7999] <= layer0_out[788];
     layer1_out[8000] <= ~layer0_out[7131] | layer0_out[7132];
     layer1_out[8001] <= ~(layer0_out[2612] & layer0_out[2613]);
     layer1_out[8002] <= layer0_out[4639] | layer0_out[4640];
     layer1_out[8003] <= ~(layer0_out[734] & layer0_out[735]);
     layer1_out[8004] <= ~layer0_out[6087] | layer0_out[6088];
     layer1_out[8005] <= layer0_out[9482];
     layer1_out[8006] <= layer0_out[1416] & ~layer0_out[1415];
     layer1_out[8007] <= ~(layer0_out[9729] | layer0_out[9730]);
     layer1_out[8008] <= ~layer0_out[11282] | layer0_out[11283];
     layer1_out[8009] <= ~layer0_out[1563];
     layer1_out[8010] <= ~layer0_out[6503];
     layer1_out[8011] <= ~(layer0_out[3684] & layer0_out[3685]);
     layer1_out[8012] <= layer0_out[6916];
     layer1_out[8013] <= layer0_out[4649];
     layer1_out[8014] <= layer0_out[6532] & layer0_out[6533];
     layer1_out[8015] <= layer0_out[7068] & ~layer0_out[7069];
     layer1_out[8016] <= layer0_out[7581];
     layer1_out[8017] <= ~layer0_out[11965];
     layer1_out[8018] <= ~(layer0_out[5691] & layer0_out[5692]);
     layer1_out[8019] <= layer0_out[402] & layer0_out[403];
     layer1_out[8020] <= ~layer0_out[8386] | layer0_out[8387];
     layer1_out[8021] <= ~(layer0_out[2538] ^ layer0_out[2539]);
     layer1_out[8022] <= ~layer0_out[4908];
     layer1_out[8023] <= layer0_out[980] | layer0_out[981];
     layer1_out[8024] <= ~(layer0_out[745] & layer0_out[746]);
     layer1_out[8025] <= ~(layer0_out[202] ^ layer0_out[203]);
     layer1_out[8026] <= ~(layer0_out[10352] | layer0_out[10353]);
     layer1_out[8027] <= layer0_out[11622] & ~layer0_out[11623];
     layer1_out[8028] <= ~(layer0_out[8054] & layer0_out[8055]);
     layer1_out[8029] <= ~(layer0_out[8363] & layer0_out[8364]);
     layer1_out[8030] <= ~layer0_out[2476] | layer0_out[2477];
     layer1_out[8031] <= layer0_out[5339] & ~layer0_out[5338];
     layer1_out[8032] <= layer0_out[9844] & ~layer0_out[9845];
     layer1_out[8033] <= layer0_out[9148] & ~layer0_out[9147];
     layer1_out[8034] <= layer0_out[6611];
     layer1_out[8035] <= layer0_out[10853];
     layer1_out[8036] <= layer0_out[7153] ^ layer0_out[7154];
     layer1_out[8037] <= ~layer0_out[5667];
     layer1_out[8038] <= layer0_out[7732];
     layer1_out[8039] <= layer0_out[5891];
     layer1_out[8040] <= ~(layer0_out[1353] ^ layer0_out[1354]);
     layer1_out[8041] <= layer0_out[4865] ^ layer0_out[4866];
     layer1_out[8042] <= layer0_out[7861] & layer0_out[7862];
     layer1_out[8043] <= ~layer0_out[10585];
     layer1_out[8044] <= layer0_out[8870] & layer0_out[8871];
     layer1_out[8045] <= layer0_out[11750] & layer0_out[11751];
     layer1_out[8046] <= layer0_out[10035];
     layer1_out[8047] <= layer0_out[6246] & layer0_out[6247];
     layer1_out[8048] <= ~(layer0_out[5824] ^ layer0_out[5825]);
     layer1_out[8049] <= layer0_out[2841] ^ layer0_out[2842];
     layer1_out[8050] <= ~(layer0_out[1383] & layer0_out[1384]);
     layer1_out[8051] <= layer0_out[4766] & ~layer0_out[4767];
     layer1_out[8052] <= ~layer0_out[11840] | layer0_out[11841];
     layer1_out[8053] <= layer0_out[7392];
     layer1_out[8054] <= layer0_out[3072] & layer0_out[3073];
     layer1_out[8055] <= layer0_out[3755] & ~layer0_out[3754];
     layer1_out[8056] <= layer0_out[5080] & ~layer0_out[5081];
     layer1_out[8057] <= ~(layer0_out[7490] | layer0_out[7491]);
     layer1_out[8058] <= ~layer0_out[9536] | layer0_out[9535];
     layer1_out[8059] <= layer0_out[1955] ^ layer0_out[1956];
     layer1_out[8060] <= ~(layer0_out[2889] | layer0_out[2890]);
     layer1_out[8061] <= layer0_out[5598] & layer0_out[5599];
     layer1_out[8062] <= layer0_out[4457] & ~layer0_out[4456];
     layer1_out[8063] <= layer0_out[2781] & ~layer0_out[2782];
     layer1_out[8064] <= layer0_out[10547] & ~layer0_out[10546];
     layer1_out[8065] <= layer0_out[6478] & ~layer0_out[6479];
     layer1_out[8066] <= layer0_out[1508];
     layer1_out[8067] <= layer0_out[10456] | layer0_out[10457];
     layer1_out[8068] <= layer0_out[5996];
     layer1_out[8069] <= ~(layer0_out[6637] & layer0_out[6638]);
     layer1_out[8070] <= ~(layer0_out[7870] & layer0_out[7871]);
     layer1_out[8071] <= 1'b0;
     layer1_out[8072] <= layer0_out[10620] & ~layer0_out[10619];
     layer1_out[8073] <= layer0_out[8255];
     layer1_out[8074] <= layer0_out[11262];
     layer1_out[8075] <= ~layer0_out[874];
     layer1_out[8076] <= layer0_out[5923] | layer0_out[5924];
     layer1_out[8077] <= ~(layer0_out[10983] ^ layer0_out[10984]);
     layer1_out[8078] <= layer0_out[3649];
     layer1_out[8079] <= ~layer0_out[3654] | layer0_out[3655];
     layer1_out[8080] <= ~(layer0_out[7155] | layer0_out[7156]);
     layer1_out[8081] <= layer0_out[8945] & layer0_out[8946];
     layer1_out[8082] <= ~(layer0_out[444] & layer0_out[445]);
     layer1_out[8083] <= layer0_out[6839] ^ layer0_out[6840];
     layer1_out[8084] <= layer0_out[10743];
     layer1_out[8085] <= ~layer0_out[2453];
     layer1_out[8086] <= layer0_out[1252] & ~layer0_out[1253];
     layer1_out[8087] <= layer0_out[7888] | layer0_out[7889];
     layer1_out[8088] <= ~layer0_out[853];
     layer1_out[8089] <= layer0_out[3970];
     layer1_out[8090] <= layer0_out[11199] ^ layer0_out[11200];
     layer1_out[8091] <= ~layer0_out[10019] | layer0_out[10020];
     layer1_out[8092] <= layer0_out[11327];
     layer1_out[8093] <= layer0_out[10069] | layer0_out[10070];
     layer1_out[8094] <= ~layer0_out[2396] | layer0_out[2395];
     layer1_out[8095] <= layer0_out[1125];
     layer1_out[8096] <= ~layer0_out[6851] | layer0_out[6852];
     layer1_out[8097] <= ~layer0_out[8662];
     layer1_out[8098] <= ~layer0_out[8935];
     layer1_out[8099] <= layer0_out[11389];
     layer1_out[8100] <= 1'b0;
     layer1_out[8101] <= ~(layer0_out[3892] ^ layer0_out[3893]);
     layer1_out[8102] <= ~(layer0_out[1930] & layer0_out[1931]);
     layer1_out[8103] <= layer0_out[11448] | layer0_out[11449];
     layer1_out[8104] <= ~(layer0_out[11858] & layer0_out[11859]);
     layer1_out[8105] <= ~layer0_out[11784];
     layer1_out[8106] <= ~(layer0_out[4790] | layer0_out[4791]);
     layer1_out[8107] <= ~(layer0_out[5108] ^ layer0_out[5109]);
     layer1_out[8108] <= ~layer0_out[9804] | layer0_out[9805];
     layer1_out[8109] <= ~(layer0_out[7812] ^ layer0_out[7813]);
     layer1_out[8110] <= ~layer0_out[6275] | layer0_out[6274];
     layer1_out[8111] <= layer0_out[11679];
     layer1_out[8112] <= layer0_out[11971] & ~layer0_out[11970];
     layer1_out[8113] <= layer0_out[8302];
     layer1_out[8114] <= ~layer0_out[10009];
     layer1_out[8115] <= layer0_out[118];
     layer1_out[8116] <= ~layer0_out[1130] | layer0_out[1129];
     layer1_out[8117] <= layer0_out[11093] & ~layer0_out[11092];
     layer1_out[8118] <= layer0_out[303] & layer0_out[304];
     layer1_out[8119] <= layer0_out[5617] | layer0_out[5618];
     layer1_out[8120] <= 1'b0;
     layer1_out[8121] <= ~layer0_out[11097];
     layer1_out[8122] <= ~(layer0_out[8508] & layer0_out[8509]);
     layer1_out[8123] <= layer0_out[2901] & layer0_out[2902];
     layer1_out[8124] <= ~layer0_out[10625];
     layer1_out[8125] <= layer0_out[4153] ^ layer0_out[4154];
     layer1_out[8126] <= layer0_out[3834] | layer0_out[3835];
     layer1_out[8127] <= layer0_out[4458];
     layer1_out[8128] <= ~layer0_out[6729] | layer0_out[6728];
     layer1_out[8129] <= layer0_out[755];
     layer1_out[8130] <= layer0_out[8376];
     layer1_out[8131] <= layer0_out[3422];
     layer1_out[8132] <= layer0_out[2338] | layer0_out[2339];
     layer1_out[8133] <= ~layer0_out[3385] | layer0_out[3384];
     layer1_out[8134] <= ~(layer0_out[7590] ^ layer0_out[7591]);
     layer1_out[8135] <= ~layer0_out[5676] | layer0_out[5675];
     layer1_out[8136] <= layer0_out[11919] & ~layer0_out[11918];
     layer1_out[8137] <= ~(layer0_out[4405] & layer0_out[4406]);
     layer1_out[8138] <= ~layer0_out[1551] | layer0_out[1550];
     layer1_out[8139] <= ~layer0_out[8168];
     layer1_out[8140] <= layer0_out[9862];
     layer1_out[8141] <= layer0_out[7524];
     layer1_out[8142] <= ~(layer0_out[8170] | layer0_out[8171]);
     layer1_out[8143] <= ~(layer0_out[5101] | layer0_out[5102]);
     layer1_out[8144] <= layer0_out[8368];
     layer1_out[8145] <= ~layer0_out[4566];
     layer1_out[8146] <= 1'b1;
     layer1_out[8147] <= layer0_out[2146] & ~layer0_out[2147];
     layer1_out[8148] <= layer0_out[11602] | layer0_out[11603];
     layer1_out[8149] <= ~layer0_out[11564];
     layer1_out[8150] <= layer0_out[1030];
     layer1_out[8151] <= ~layer0_out[11082];
     layer1_out[8152] <= 1'b0;
     layer1_out[8153] <= ~layer0_out[11536];
     layer1_out[8154] <= ~layer0_out[11997];
     layer1_out[8155] <= layer0_out[8518];
     layer1_out[8156] <= ~(layer0_out[8746] | layer0_out[8747]);
     layer1_out[8157] <= layer0_out[11303] & ~layer0_out[11302];
     layer1_out[8158] <= layer0_out[11841];
     layer1_out[8159] <= ~layer0_out[1449];
     layer1_out[8160] <= ~layer0_out[7783];
     layer1_out[8161] <= layer0_out[8443];
     layer1_out[8162] <= 1'b0;
     layer1_out[8163] <= layer0_out[4583] & ~layer0_out[4584];
     layer1_out[8164] <= layer0_out[10090];
     layer1_out[8165] <= layer0_out[596];
     layer1_out[8166] <= layer0_out[9306];
     layer1_out[8167] <= ~layer0_out[11296];
     layer1_out[8168] <= ~layer0_out[4227] | layer0_out[4226];
     layer1_out[8169] <= layer0_out[6535];
     layer1_out[8170] <= ~(layer0_out[7414] & layer0_out[7415]);
     layer1_out[8171] <= ~layer0_out[507] | layer0_out[506];
     layer1_out[8172] <= ~layer0_out[4754] | layer0_out[4755];
     layer1_out[8173] <= layer0_out[2131];
     layer1_out[8174] <= layer0_out[11697];
     layer1_out[8175] <= layer0_out[4795] & ~layer0_out[4796];
     layer1_out[8176] <= layer0_out[5160] | layer0_out[5161];
     layer1_out[8177] <= layer0_out[6111];
     layer1_out[8178] <= layer0_out[8521] ^ layer0_out[8522];
     layer1_out[8179] <= 1'b0;
     layer1_out[8180] <= layer0_out[5805];
     layer1_out[8181] <= layer0_out[7257];
     layer1_out[8182] <= ~layer0_out[11747];
     layer1_out[8183] <= layer0_out[6993];
     layer1_out[8184] <= layer0_out[1338] & ~layer0_out[1337];
     layer1_out[8185] <= layer0_out[6468];
     layer1_out[8186] <= ~layer0_out[7342];
     layer1_out[8187] <= ~layer0_out[5117] | layer0_out[5116];
     layer1_out[8188] <= layer0_out[7874];
     layer1_out[8189] <= ~layer0_out[2416] | layer0_out[2415];
     layer1_out[8190] <= ~(layer0_out[2474] | layer0_out[2475]);
     layer1_out[8191] <= ~layer0_out[1119] | layer0_out[1118];
     layer1_out[8192] <= layer0_out[2905];
     layer1_out[8193] <= layer0_out[10536] & layer0_out[10537];
     layer1_out[8194] <= layer0_out[10019];
     layer1_out[8195] <= layer0_out[5578] | layer0_out[5579];
     layer1_out[8196] <= layer0_out[107] | layer0_out[108];
     layer1_out[8197] <= layer0_out[6410] | layer0_out[6411];
     layer1_out[8198] <= ~layer0_out[5407] | layer0_out[5406];
     layer1_out[8199] <= layer0_out[9513];
     layer1_out[8200] <= ~(layer0_out[1566] & layer0_out[1567]);
     layer1_out[8201] <= layer0_out[8918] & ~layer0_out[8917];
     layer1_out[8202] <= ~(layer0_out[6312] ^ layer0_out[6313]);
     layer1_out[8203] <= ~layer0_out[3303];
     layer1_out[8204] <= layer0_out[9005] & layer0_out[9006];
     layer1_out[8205] <= ~layer0_out[4515];
     layer1_out[8206] <= ~(layer0_out[10935] ^ layer0_out[10936]);
     layer1_out[8207] <= layer0_out[8695] | layer0_out[8696];
     layer1_out[8208] <= ~layer0_out[7121] | layer0_out[7120];
     layer1_out[8209] <= layer0_out[9833];
     layer1_out[8210] <= ~layer0_out[190] | layer0_out[189];
     layer1_out[8211] <= layer0_out[2846] & layer0_out[2847];
     layer1_out[8212] <= layer0_out[5028];
     layer1_out[8213] <= layer0_out[2609] & layer0_out[2610];
     layer1_out[8214] <= layer0_out[10430] & layer0_out[10431];
     layer1_out[8215] <= layer0_out[11071] & layer0_out[11072];
     layer1_out[8216] <= ~layer0_out[1662];
     layer1_out[8217] <= layer0_out[8008] & layer0_out[8009];
     layer1_out[8218] <= ~(layer0_out[5795] ^ layer0_out[5796]);
     layer1_out[8219] <= ~layer0_out[9428] | layer0_out[9429];
     layer1_out[8220] <= layer0_out[8560];
     layer1_out[8221] <= ~layer0_out[1423] | layer0_out[1422];
     layer1_out[8222] <= layer0_out[1170] & layer0_out[1171];
     layer1_out[8223] <= layer0_out[851] | layer0_out[852];
     layer1_out[8224] <= ~layer0_out[9029];
     layer1_out[8225] <= layer0_out[9569] & ~layer0_out[9568];
     layer1_out[8226] <= ~layer0_out[10161];
     layer1_out[8227] <= ~layer0_out[8635] | layer0_out[8634];
     layer1_out[8228] <= ~(layer0_out[5014] & layer0_out[5015]);
     layer1_out[8229] <= layer0_out[6090] & layer0_out[6091];
     layer1_out[8230] <= ~(layer0_out[1394] & layer0_out[1395]);
     layer1_out[8231] <= layer0_out[992] | layer0_out[993];
     layer1_out[8232] <= ~layer0_out[2832];
     layer1_out[8233] <= ~layer0_out[9426];
     layer1_out[8234] <= ~layer0_out[7456];
     layer1_out[8235] <= layer0_out[5383];
     layer1_out[8236] <= ~layer0_out[440];
     layer1_out[8237] <= layer0_out[2497] ^ layer0_out[2498];
     layer1_out[8238] <= layer0_out[6078] & ~layer0_out[6077];
     layer1_out[8239] <= layer0_out[7528] & ~layer0_out[7527];
     layer1_out[8240] <= layer0_out[1485] & ~layer0_out[1486];
     layer1_out[8241] <= layer0_out[2894] & ~layer0_out[2895];
     layer1_out[8242] <= layer0_out[4691] & ~layer0_out[4692];
     layer1_out[8243] <= ~layer0_out[1909] | layer0_out[1910];
     layer1_out[8244] <= layer0_out[8223];
     layer1_out[8245] <= layer0_out[4766];
     layer1_out[8246] <= ~layer0_out[6166] | layer0_out[6167];
     layer1_out[8247] <= layer0_out[522];
     layer1_out[8248] <= ~(layer0_out[6348] | layer0_out[6349]);
     layer1_out[8249] <= ~layer0_out[127];
     layer1_out[8250] <= ~layer0_out[11416] | layer0_out[11415];
     layer1_out[8251] <= layer0_out[9476] | layer0_out[9477];
     layer1_out[8252] <= ~layer0_out[7022];
     layer1_out[8253] <= ~layer0_out[9452];
     layer1_out[8254] <= ~(layer0_out[4619] | layer0_out[4620]);
     layer1_out[8255] <= ~(layer0_out[3009] ^ layer0_out[3010]);
     layer1_out[8256] <= ~(layer0_out[6935] & layer0_out[6936]);
     layer1_out[8257] <= layer0_out[5918];
     layer1_out[8258] <= layer0_out[5865] | layer0_out[5866];
     layer1_out[8259] <= ~layer0_out[2895];
     layer1_out[8260] <= layer0_out[4814] ^ layer0_out[4815];
     layer1_out[8261] <= layer0_out[3423] & layer0_out[3424];
     layer1_out[8262] <= ~(layer0_out[7567] & layer0_out[7568]);
     layer1_out[8263] <= layer0_out[7649] & layer0_out[7650];
     layer1_out[8264] <= layer0_out[10154];
     layer1_out[8265] <= layer0_out[2374];
     layer1_out[8266] <= ~(layer0_out[9886] ^ layer0_out[9887]);
     layer1_out[8267] <= layer0_out[10702] ^ layer0_out[10703];
     layer1_out[8268] <= ~layer0_out[8417] | layer0_out[8416];
     layer1_out[8269] <= layer0_out[9320] & ~layer0_out[9321];
     layer1_out[8270] <= layer0_out[6190] & layer0_out[6191];
     layer1_out[8271] <= ~(layer0_out[7656] | layer0_out[7657]);
     layer1_out[8272] <= ~layer0_out[368];
     layer1_out[8273] <= layer0_out[11919];
     layer1_out[8274] <= ~layer0_out[8852];
     layer1_out[8275] <= ~layer0_out[3764] | layer0_out[3763];
     layer1_out[8276] <= ~layer0_out[7482];
     layer1_out[8277] <= ~layer0_out[4906];
     layer1_out[8278] <= ~layer0_out[179] | layer0_out[178];
     layer1_out[8279] <= layer0_out[9784] & ~layer0_out[9783];
     layer1_out[8280] <= ~layer0_out[8676];
     layer1_out[8281] <= layer0_out[1066] & ~layer0_out[1065];
     layer1_out[8282] <= layer0_out[1271];
     layer1_out[8283] <= layer0_out[6058] ^ layer0_out[6059];
     layer1_out[8284] <= ~layer0_out[10180];
     layer1_out[8285] <= layer0_out[3819] & ~layer0_out[3818];
     layer1_out[8286] <= layer0_out[1286];
     layer1_out[8287] <= layer0_out[550] & layer0_out[551];
     layer1_out[8288] <= ~(layer0_out[2292] ^ layer0_out[2293]);
     layer1_out[8289] <= ~(layer0_out[6386] | layer0_out[6387]);
     layer1_out[8290] <= layer0_out[1925] & ~layer0_out[1924];
     layer1_out[8291] <= ~(layer0_out[9680] & layer0_out[9681]);
     layer1_out[8292] <= layer0_out[9174] & layer0_out[9175];
     layer1_out[8293] <= ~(layer0_out[10554] & layer0_out[10555]);
     layer1_out[8294] <= 1'b1;
     layer1_out[8295] <= ~layer0_out[772];
     layer1_out[8296] <= ~(layer0_out[1705] | layer0_out[1706]);
     layer1_out[8297] <= ~layer0_out[3932];
     layer1_out[8298] <= ~(layer0_out[3980] & layer0_out[3981]);
     layer1_out[8299] <= ~layer0_out[6396] | layer0_out[6397];
     layer1_out[8300] <= ~layer0_out[7060] | layer0_out[7059];
     layer1_out[8301] <= ~layer0_out[3807];
     layer1_out[8302] <= layer0_out[5544] & layer0_out[5545];
     layer1_out[8303] <= ~(layer0_out[5191] | layer0_out[5192]);
     layer1_out[8304] <= ~(layer0_out[1748] | layer0_out[1749]);
     layer1_out[8305] <= layer0_out[2189] & layer0_out[2190];
     layer1_out[8306] <= layer0_out[10583] & ~layer0_out[10582];
     layer1_out[8307] <= layer0_out[930] | layer0_out[931];
     layer1_out[8308] <= ~(layer0_out[3215] & layer0_out[3216]);
     layer1_out[8309] <= ~layer0_out[4507] | layer0_out[4506];
     layer1_out[8310] <= layer0_out[8830] & ~layer0_out[8829];
     layer1_out[8311] <= ~layer0_out[7268];
     layer1_out[8312] <= layer0_out[9945] & ~layer0_out[9944];
     layer1_out[8313] <= ~layer0_out[5205];
     layer1_out[8314] <= ~(layer0_out[3946] & layer0_out[3947]);
     layer1_out[8315] <= layer0_out[4105];
     layer1_out[8316] <= ~layer0_out[10479];
     layer1_out[8317] <= ~(layer0_out[9760] | layer0_out[9761]);
     layer1_out[8318] <= ~layer0_out[6325] | layer0_out[6326];
     layer1_out[8319] <= ~layer0_out[10180];
     layer1_out[8320] <= layer0_out[546];
     layer1_out[8321] <= layer0_out[1774] & ~layer0_out[1773];
     layer1_out[8322] <= layer0_out[1963] & layer0_out[1964];
     layer1_out[8323] <= 1'b1;
     layer1_out[8324] <= 1'b0;
     layer1_out[8325] <= ~(layer0_out[926] | layer0_out[927]);
     layer1_out[8326] <= layer0_out[4975] | layer0_out[4976];
     layer1_out[8327] <= layer0_out[8193];
     layer1_out[8328] <= layer0_out[9395] & ~layer0_out[9394];
     layer1_out[8329] <= 1'b0;
     layer1_out[8330] <= layer0_out[10225];
     layer1_out[8331] <= ~layer0_out[3703] | layer0_out[3702];
     layer1_out[8332] <= layer0_out[10043];
     layer1_out[8333] <= layer0_out[2103] & ~layer0_out[2102];
     layer1_out[8334] <= ~(layer0_out[3674] ^ layer0_out[3675]);
     layer1_out[8335] <= ~layer0_out[8952] | layer0_out[8953];
     layer1_out[8336] <= layer0_out[8455];
     layer1_out[8337] <= layer0_out[9509];
     layer1_out[8338] <= layer0_out[11547] & ~layer0_out[11548];
     layer1_out[8339] <= layer0_out[4919] & ~layer0_out[4920];
     layer1_out[8340] <= layer0_out[6305];
     layer1_out[8341] <= layer0_out[2211];
     layer1_out[8342] <= ~layer0_out[9234] | layer0_out[9235];
     layer1_out[8343] <= layer0_out[7824] & ~layer0_out[7823];
     layer1_out[8344] <= layer0_out[9138] & layer0_out[9139];
     layer1_out[8345] <= layer0_out[2308] & ~layer0_out[2309];
     layer1_out[8346] <= ~(layer0_out[2220] | layer0_out[2221]);
     layer1_out[8347] <= layer0_out[2071] | layer0_out[2072];
     layer1_out[8348] <= layer0_out[11537] & layer0_out[11538];
     layer1_out[8349] <= ~layer0_out[2921];
     layer1_out[8350] <= ~layer0_out[380] | layer0_out[379];
     layer1_out[8351] <= ~(layer0_out[6633] ^ layer0_out[6634]);
     layer1_out[8352] <= layer0_out[1157] | layer0_out[1158];
     layer1_out[8353] <= layer0_out[5869] | layer0_out[5870];
     layer1_out[8354] <= ~(layer0_out[11749] ^ layer0_out[11750]);
     layer1_out[8355] <= ~layer0_out[1868];
     layer1_out[8356] <= layer0_out[1022] & ~layer0_out[1023];
     layer1_out[8357] <= ~layer0_out[6157] | layer0_out[6156];
     layer1_out[8358] <= ~layer0_out[10484];
     layer1_out[8359] <= layer0_out[2257];
     layer1_out[8360] <= layer0_out[796] | layer0_out[797];
     layer1_out[8361] <= ~layer0_out[6697];
     layer1_out[8362] <= ~layer0_out[10551];
     layer1_out[8363] <= ~layer0_out[4521] | layer0_out[4520];
     layer1_out[8364] <= layer0_out[4480] ^ layer0_out[4481];
     layer1_out[8365] <= ~layer0_out[7986] | layer0_out[7987];
     layer1_out[8366] <= layer0_out[6913];
     layer1_out[8367] <= layer0_out[137] | layer0_out[138];
     layer1_out[8368] <= layer0_out[11798];
     layer1_out[8369] <= ~layer0_out[11464] | layer0_out[11463];
     layer1_out[8370] <= 1'b1;
     layer1_out[8371] <= layer0_out[10424] | layer0_out[10425];
     layer1_out[8372] <= layer0_out[82] & layer0_out[83];
     layer1_out[8373] <= layer0_out[1893] & layer0_out[1894];
     layer1_out[8374] <= ~layer0_out[5259];
     layer1_out[8375] <= layer0_out[2282] ^ layer0_out[2283];
     layer1_out[8376] <= layer0_out[238] & ~layer0_out[237];
     layer1_out[8377] <= layer0_out[4116];
     layer1_out[8378] <= layer0_out[8441] & ~layer0_out[8442];
     layer1_out[8379] <= ~(layer0_out[3442] ^ layer0_out[3443]);
     layer1_out[8380] <= ~(layer0_out[10115] ^ layer0_out[10116]);
     layer1_out[8381] <= layer0_out[7580];
     layer1_out[8382] <= layer0_out[6956] ^ layer0_out[6957];
     layer1_out[8383] <= ~(layer0_out[6165] ^ layer0_out[6166]);
     layer1_out[8384] <= layer0_out[3596] & ~layer0_out[3595];
     layer1_out[8385] <= layer0_out[7510];
     layer1_out[8386] <= layer0_out[6222];
     layer1_out[8387] <= layer0_out[1219];
     layer1_out[8388] <= ~(layer0_out[3281] ^ layer0_out[3282]);
     layer1_out[8389] <= layer0_out[6641];
     layer1_out[8390] <= layer0_out[2622];
     layer1_out[8391] <= ~layer0_out[4900];
     layer1_out[8392] <= layer0_out[11803] & ~layer0_out[11804];
     layer1_out[8393] <= ~layer0_out[10028] | layer0_out[10029];
     layer1_out[8394] <= layer0_out[8433];
     layer1_out[8395] <= ~layer0_out[10798];
     layer1_out[8396] <= layer0_out[11753];
     layer1_out[8397] <= layer0_out[3310] & ~layer0_out[3309];
     layer1_out[8398] <= layer0_out[4387] & ~layer0_out[4388];
     layer1_out[8399] <= layer0_out[10435];
     layer1_out[8400] <= ~layer0_out[9554];
     layer1_out[8401] <= layer0_out[9824] & ~layer0_out[9823];
     layer1_out[8402] <= ~layer0_out[8528];
     layer1_out[8403] <= 1'b1;
     layer1_out[8404] <= layer0_out[9297];
     layer1_out[8405] <= ~layer0_out[34] | layer0_out[35];
     layer1_out[8406] <= layer0_out[2267] & layer0_out[2268];
     layer1_out[8407] <= ~layer0_out[7177] | layer0_out[7176];
     layer1_out[8408] <= layer0_out[4421];
     layer1_out[8409] <= layer0_out[10787];
     layer1_out[8410] <= layer0_out[4544];
     layer1_out[8411] <= layer0_out[6599];
     layer1_out[8412] <= layer0_out[7979] & ~layer0_out[7980];
     layer1_out[8413] <= layer0_out[4205];
     layer1_out[8414] <= ~layer0_out[7202];
     layer1_out[8415] <= ~layer0_out[5541] | layer0_out[5542];
     layer1_out[8416] <= layer0_out[10341];
     layer1_out[8417] <= layer0_out[5419] & ~layer0_out[5418];
     layer1_out[8418] <= ~layer0_out[4089] | layer0_out[4088];
     layer1_out[8419] <= ~layer0_out[11411];
     layer1_out[8420] <= layer0_out[98];
     layer1_out[8421] <= ~(layer0_out[6913] ^ layer0_out[6914]);
     layer1_out[8422] <= layer0_out[741] ^ layer0_out[742];
     layer1_out[8423] <= ~(layer0_out[10716] | layer0_out[10717]);
     layer1_out[8424] <= layer0_out[1686] | layer0_out[1687];
     layer1_out[8425] <= layer0_out[6284];
     layer1_out[8426] <= layer0_out[1764] | layer0_out[1765];
     layer1_out[8427] <= ~layer0_out[252] | layer0_out[253];
     layer1_out[8428] <= layer0_out[7747] & ~layer0_out[7746];
     layer1_out[8429] <= layer0_out[146] & ~layer0_out[145];
     layer1_out[8430] <= layer0_out[11500];
     layer1_out[8431] <= ~layer0_out[9978] | layer0_out[9977];
     layer1_out[8432] <= 1'b1;
     layer1_out[8433] <= layer0_out[7595] & ~layer0_out[7594];
     layer1_out[8434] <= layer0_out[9386];
     layer1_out[8435] <= ~(layer0_out[3558] | layer0_out[3559]);
     layer1_out[8436] <= 1'b0;
     layer1_out[8437] <= layer0_out[6173] ^ layer0_out[6174];
     layer1_out[8438] <= ~(layer0_out[1192] | layer0_out[1193]);
     layer1_out[8439] <= ~layer0_out[245] | layer0_out[246];
     layer1_out[8440] <= ~layer0_out[11079];
     layer1_out[8441] <= 1'b1;
     layer1_out[8442] <= layer0_out[11715] ^ layer0_out[11716];
     layer1_out[8443] <= layer0_out[7875] & layer0_out[7876];
     layer1_out[8444] <= ~(layer0_out[3789] ^ layer0_out[3790]);
     layer1_out[8445] <= layer0_out[4358] ^ layer0_out[4359];
     layer1_out[8446] <= layer0_out[8586];
     layer1_out[8447] <= layer0_out[3735];
     layer1_out[8448] <= layer0_out[1264] & ~layer0_out[1265];
     layer1_out[8449] <= layer0_out[6693];
     layer1_out[8450] <= ~layer0_out[7464];
     layer1_out[8451] <= ~layer0_out[3295] | layer0_out[3294];
     layer1_out[8452] <= layer0_out[4238] & ~layer0_out[4239];
     layer1_out[8453] <= ~layer0_out[5789];
     layer1_out[8454] <= ~layer0_out[9462] | layer0_out[9463];
     layer1_out[8455] <= ~layer0_out[4644] | layer0_out[4643];
     layer1_out[8456] <= ~layer0_out[3594];
     layer1_out[8457] <= layer0_out[2774];
     layer1_out[8458] <= ~layer0_out[10121];
     layer1_out[8459] <= layer0_out[7045] & ~layer0_out[7046];
     layer1_out[8460] <= ~(layer0_out[9769] & layer0_out[9770]);
     layer1_out[8461] <= layer0_out[2600];
     layer1_out[8462] <= ~(layer0_out[3015] & layer0_out[3016]);
     layer1_out[8463] <= layer0_out[8911] & ~layer0_out[8912];
     layer1_out[8464] <= layer0_out[1978] | layer0_out[1979];
     layer1_out[8465] <= layer0_out[8015] ^ layer0_out[8016];
     layer1_out[8466] <= ~layer0_out[11633];
     layer1_out[8467] <= layer0_out[9803];
     layer1_out[8468] <= ~layer0_out[11842];
     layer1_out[8469] <= ~layer0_out[9401] | layer0_out[9402];
     layer1_out[8470] <= layer0_out[1561] | layer0_out[1562];
     layer1_out[8471] <= ~layer0_out[9002] | layer0_out[9001];
     layer1_out[8472] <= ~layer0_out[5365] | layer0_out[5364];
     layer1_out[8473] <= ~layer0_out[10118] | layer0_out[10119];
     layer1_out[8474] <= layer0_out[7704] & ~layer0_out[7703];
     layer1_out[8475] <= ~layer0_out[11028];
     layer1_out[8476] <= layer0_out[2827] | layer0_out[2828];
     layer1_out[8477] <= layer0_out[10934];
     layer1_out[8478] <= ~layer0_out[7150];
     layer1_out[8479] <= ~layer0_out[2547];
     layer1_out[8480] <= ~(layer0_out[1513] & layer0_out[1514]);
     layer1_out[8481] <= layer0_out[4407];
     layer1_out[8482] <= layer0_out[6731] | layer0_out[6732];
     layer1_out[8483] <= ~layer0_out[4684];
     layer1_out[8484] <= ~layer0_out[1929];
     layer1_out[8485] <= ~layer0_out[11189];
     layer1_out[8486] <= ~layer0_out[8869];
     layer1_out[8487] <= layer0_out[3632] & ~layer0_out[3633];
     layer1_out[8488] <= 1'b0;
     layer1_out[8489] <= layer0_out[370] & ~layer0_out[369];
     layer1_out[8490] <= layer0_out[6636] ^ layer0_out[6637];
     layer1_out[8491] <= 1'b0;
     layer1_out[8492] <= layer0_out[10928] | layer0_out[10929];
     layer1_out[8493] <= ~layer0_out[10527];
     layer1_out[8494] <= layer0_out[3526];
     layer1_out[8495] <= ~(layer0_out[3049] | layer0_out[3050]);
     layer1_out[8496] <= layer0_out[8841] & ~layer0_out[8842];
     layer1_out[8497] <= layer0_out[11647] | layer0_out[11648];
     layer1_out[8498] <= layer0_out[5953];
     layer1_out[8499] <= layer0_out[6566] & ~layer0_out[6567];
     layer1_out[8500] <= ~(layer0_out[5059] | layer0_out[5060]);
     layer1_out[8501] <= layer0_out[3713];
     layer1_out[8502] <= layer0_out[8198] & ~layer0_out[8197];
     layer1_out[8503] <= ~layer0_out[6841];
     layer1_out[8504] <= layer0_out[2967] | layer0_out[2968];
     layer1_out[8505] <= ~layer0_out[9843] | layer0_out[9842];
     layer1_out[8506] <= layer0_out[464] & ~layer0_out[463];
     layer1_out[8507] <= layer0_out[5352] & layer0_out[5353];
     layer1_out[8508] <= ~layer0_out[7716] | layer0_out[7715];
     layer1_out[8509] <= layer0_out[2366] & layer0_out[2367];
     layer1_out[8510] <= layer0_out[4619];
     layer1_out[8511] <= ~layer0_out[9307];
     layer1_out[8512] <= 1'b0;
     layer1_out[8513] <= 1'b0;
     layer1_out[8514] <= ~layer0_out[1917];
     layer1_out[8515] <= ~layer0_out[10657];
     layer1_out[8516] <= ~layer0_out[2872] | layer0_out[2871];
     layer1_out[8517] <= ~layer0_out[7001];
     layer1_out[8518] <= ~layer0_out[8411] | layer0_out[8412];
     layer1_out[8519] <= layer0_out[2362] | layer0_out[2363];
     layer1_out[8520] <= ~(layer0_out[3459] | layer0_out[3460]);
     layer1_out[8521] <= ~layer0_out[5659];
     layer1_out[8522] <= layer0_out[4690] & ~layer0_out[4691];
     layer1_out[8523] <= layer0_out[11126];
     layer1_out[8524] <= layer0_out[7126];
     layer1_out[8525] <= layer0_out[3112] & ~layer0_out[3113];
     layer1_out[8526] <= ~(layer0_out[8588] ^ layer0_out[8589]);
     layer1_out[8527] <= layer0_out[163] & ~layer0_out[162];
     layer1_out[8528] <= layer0_out[10096];
     layer1_out[8529] <= ~layer0_out[6627];
     layer1_out[8530] <= ~layer0_out[10723];
     layer1_out[8531] <= layer0_out[2653] & ~layer0_out[2654];
     layer1_out[8532] <= layer0_out[46] & ~layer0_out[47];
     layer1_out[8533] <= ~layer0_out[889] | layer0_out[890];
     layer1_out[8534] <= layer0_out[9608] | layer0_out[9609];
     layer1_out[8535] <= layer0_out[9560] & ~layer0_out[9559];
     layer1_out[8536] <= layer0_out[2861] ^ layer0_out[2862];
     layer1_out[8537] <= ~layer0_out[3458];
     layer1_out[8538] <= ~(layer0_out[8205] & layer0_out[8206]);
     layer1_out[8539] <= ~layer0_out[3203] | layer0_out[3204];
     layer1_out[8540] <= 1'b1;
     layer1_out[8541] <= layer0_out[3120];
     layer1_out[8542] <= layer0_out[662];
     layer1_out[8543] <= layer0_out[11268] ^ layer0_out[11269];
     layer1_out[8544] <= layer0_out[5088];
     layer1_out[8545] <= ~layer0_out[4720];
     layer1_out[8546] <= ~layer0_out[95];
     layer1_out[8547] <= ~layer0_out[10951];
     layer1_out[8548] <= layer0_out[8270];
     layer1_out[8549] <= ~layer0_out[3517];
     layer1_out[8550] <= layer0_out[11520] & layer0_out[11521];
     layer1_out[8551] <= layer0_out[7841] & layer0_out[7842];
     layer1_out[8552] <= ~layer0_out[620];
     layer1_out[8553] <= ~(layer0_out[7830] & layer0_out[7831]);
     layer1_out[8554] <= ~(layer0_out[2840] | layer0_out[2841]);
     layer1_out[8555] <= layer0_out[877] | layer0_out[878];
     layer1_out[8556] <= ~layer0_out[2299];
     layer1_out[8557] <= layer0_out[1051] | layer0_out[1052];
     layer1_out[8558] <= layer0_out[11727] & layer0_out[11728];
     layer1_out[8559] <= layer0_out[1612] & ~layer0_out[1611];
     layer1_out[8560] <= layer0_out[8389] & ~layer0_out[8390];
     layer1_out[8561] <= ~(layer0_out[1598] ^ layer0_out[1599]);
     layer1_out[8562] <= layer0_out[6933] & layer0_out[6934];
     layer1_out[8563] <= ~(layer0_out[8395] & layer0_out[8396]);
     layer1_out[8564] <= ~(layer0_out[324] & layer0_out[325]);
     layer1_out[8565] <= ~layer0_out[10303];
     layer1_out[8566] <= layer0_out[8358] & ~layer0_out[8359];
     layer1_out[8567] <= layer0_out[10776];
     layer1_out[8568] <= ~layer0_out[2899] | layer0_out[2898];
     layer1_out[8569] <= ~layer0_out[4521] | layer0_out[4522];
     layer1_out[8570] <= 1'b0;
     layer1_out[8571] <= 1'b1;
     layer1_out[8572] <= ~layer0_out[4808] | layer0_out[4807];
     layer1_out[8573] <= ~layer0_out[2134] | layer0_out[2133];
     layer1_out[8574] <= ~(layer0_out[2927] & layer0_out[2928]);
     layer1_out[8575] <= layer0_out[5483] | layer0_out[5484];
     layer1_out[8576] <= ~layer0_out[11771];
     layer1_out[8577] <= ~layer0_out[4871];
     layer1_out[8578] <= ~layer0_out[3855] | layer0_out[3856];
     layer1_out[8579] <= layer0_out[5304];
     layer1_out[8580] <= ~(layer0_out[6168] & layer0_out[6169]);
     layer1_out[8581] <= ~(layer0_out[10943] | layer0_out[10944]);
     layer1_out[8582] <= ~layer0_out[8251];
     layer1_out[8583] <= ~layer0_out[11959];
     layer1_out[8584] <= layer0_out[6803];
     layer1_out[8585] <= 1'b0;
     layer1_out[8586] <= layer0_out[10727] | layer0_out[10728];
     layer1_out[8587] <= layer0_out[6597] | layer0_out[6598];
     layer1_out[8588] <= ~layer0_out[7600] | layer0_out[7599];
     layer1_out[8589] <= ~layer0_out[8963];
     layer1_out[8590] <= ~layer0_out[8240] | layer0_out[8239];
     layer1_out[8591] <= layer0_out[4748];
     layer1_out[8592] <= 1'b0;
     layer1_out[8593] <= ~layer0_out[8145];
     layer1_out[8594] <= layer0_out[6326] | layer0_out[6327];
     layer1_out[8595] <= 1'b0;
     layer1_out[8596] <= layer0_out[110] & ~layer0_out[111];
     layer1_out[8597] <= layer0_out[6520] & layer0_out[6521];
     layer1_out[8598] <= layer0_out[2005];
     layer1_out[8599] <= ~(layer0_out[10606] | layer0_out[10607]);
     layer1_out[8600] <= ~(layer0_out[2302] | layer0_out[2303]);
     layer1_out[8601] <= layer0_out[2650] & ~layer0_out[2649];
     layer1_out[8602] <= ~(layer0_out[307] ^ layer0_out[308]);
     layer1_out[8603] <= ~(layer0_out[6800] ^ layer0_out[6801]);
     layer1_out[8604] <= layer0_out[11162] & ~layer0_out[11161];
     layer1_out[8605] <= layer0_out[3678] | layer0_out[3679];
     layer1_out[8606] <= layer0_out[9136] & layer0_out[9137];
     layer1_out[8607] <= layer0_out[6526];
     layer1_out[8608] <= ~layer0_out[915] | layer0_out[914];
     layer1_out[8609] <= layer0_out[5210] & layer0_out[5211];
     layer1_out[8610] <= ~layer0_out[5752];
     layer1_out[8611] <= layer0_out[2730] | layer0_out[2731];
     layer1_out[8612] <= ~(layer0_out[701] & layer0_out[702]);
     layer1_out[8613] <= layer0_out[5509];
     layer1_out[8614] <= ~(layer0_out[2360] ^ layer0_out[2361]);
     layer1_out[8615] <= layer0_out[5593] ^ layer0_out[5594];
     layer1_out[8616] <= layer0_out[2969] & layer0_out[2970];
     layer1_out[8617] <= layer0_out[104];
     layer1_out[8618] <= layer0_out[295];
     layer1_out[8619] <= layer0_out[4981] & ~layer0_out[4982];
     layer1_out[8620] <= ~(layer0_out[11395] ^ layer0_out[11396]);
     layer1_out[8621] <= ~(layer0_out[11435] ^ layer0_out[11436]);
     layer1_out[8622] <= ~layer0_out[5600];
     layer1_out[8623] <= ~layer0_out[4538];
     layer1_out[8624] <= layer0_out[2239] | layer0_out[2240];
     layer1_out[8625] <= layer0_out[8779] ^ layer0_out[8780];
     layer1_out[8626] <= layer0_out[527] & layer0_out[528];
     layer1_out[8627] <= ~(layer0_out[4382] ^ layer0_out[4383]);
     layer1_out[8628] <= ~(layer0_out[11427] | layer0_out[11428]);
     layer1_out[8629] <= layer0_out[8455];
     layer1_out[8630] <= ~layer0_out[7760] | layer0_out[7759];
     layer1_out[8631] <= ~layer0_out[3275];
     layer1_out[8632] <= ~layer0_out[2024];
     layer1_out[8633] <= ~layer0_out[6425];
     layer1_out[8634] <= ~layer0_out[929];
     layer1_out[8635] <= ~layer0_out[7374];
     layer1_out[8636] <= layer0_out[10466] & ~layer0_out[10467];
     layer1_out[8637] <= layer0_out[6105];
     layer1_out[8638] <= ~layer0_out[2267] | layer0_out[2266];
     layer1_out[8639] <= layer0_out[3231];
     layer1_out[8640] <= layer0_out[10657] & ~layer0_out[10656];
     layer1_out[8641] <= ~layer0_out[1670] | layer0_out[1671];
     layer1_out[8642] <= layer0_out[2673];
     layer1_out[8643] <= ~layer0_out[5479];
     layer1_out[8644] <= layer0_out[2143] & layer0_out[2144];
     layer1_out[8645] <= ~(layer0_out[4195] & layer0_out[4196]);
     layer1_out[8646] <= ~layer0_out[4188];
     layer1_out[8647] <= layer0_out[2881] & layer0_out[2882];
     layer1_out[8648] <= layer0_out[7308] & ~layer0_out[7307];
     layer1_out[8649] <= layer0_out[3271] & ~layer0_out[3272];
     layer1_out[8650] <= layer0_out[1775];
     layer1_out[8651] <= ~layer0_out[8345];
     layer1_out[8652] <= layer0_out[1024];
     layer1_out[8653] <= layer0_out[11668];
     layer1_out[8654] <= layer0_out[5467];
     layer1_out[8655] <= ~(layer0_out[10119] ^ layer0_out[10120]);
     layer1_out[8656] <= layer0_out[6999] & layer0_out[7000];
     layer1_out[8657] <= ~layer0_out[10307];
     layer1_out[8658] <= layer0_out[4605] & ~layer0_out[4604];
     layer1_out[8659] <= layer0_out[2595] & ~layer0_out[2594];
     layer1_out[8660] <= layer0_out[1820] & ~layer0_out[1821];
     layer1_out[8661] <= layer0_out[1897] ^ layer0_out[1898];
     layer1_out[8662] <= layer0_out[4526];
     layer1_out[8663] <= layer0_out[11095];
     layer1_out[8664] <= layer0_out[7465];
     layer1_out[8665] <= layer0_out[8646] | layer0_out[8647];
     layer1_out[8666] <= ~layer0_out[10610];
     layer1_out[8667] <= ~(layer0_out[4324] & layer0_out[4325]);
     layer1_out[8668] <= ~(layer0_out[2569] & layer0_out[2570]);
     layer1_out[8669] <= 1'b0;
     layer1_out[8670] <= ~layer0_out[11586];
     layer1_out[8671] <= ~layer0_out[6775];
     layer1_out[8672] <= ~layer0_out[4553];
     layer1_out[8673] <= ~(layer0_out[6308] & layer0_out[6309]);
     layer1_out[8674] <= ~(layer0_out[454] ^ layer0_out[455]);
     layer1_out[8675] <= layer0_out[1855];
     layer1_out[8676] <= layer0_out[3282] | layer0_out[3283];
     layer1_out[8677] <= layer0_out[8976];
     layer1_out[8678] <= layer0_out[3334] | layer0_out[3335];
     layer1_out[8679] <= layer0_out[3573];
     layer1_out[8680] <= layer0_out[115] & ~layer0_out[114];
     layer1_out[8681] <= ~layer0_out[2729] | layer0_out[2730];
     layer1_out[8682] <= ~layer0_out[5867];
     layer1_out[8683] <= ~layer0_out[6488];
     layer1_out[8684] <= layer0_out[7013] & ~layer0_out[7012];
     layer1_out[8685] <= layer0_out[2985] & layer0_out[2986];
     layer1_out[8686] <= layer0_out[6679] & ~layer0_out[6680];
     layer1_out[8687] <= ~layer0_out[879];
     layer1_out[8688] <= layer0_out[495] & layer0_out[496];
     layer1_out[8689] <= layer0_out[4181];
     layer1_out[8690] <= 1'b0;
     layer1_out[8691] <= ~(layer0_out[8463] & layer0_out[8464]);
     layer1_out[8692] <= ~layer0_out[5549] | layer0_out[5550];
     layer1_out[8693] <= layer0_out[2050];
     layer1_out[8694] <= layer0_out[3285];
     layer1_out[8695] <= ~layer0_out[11573];
     layer1_out[8696] <= ~layer0_out[9343] | layer0_out[9342];
     layer1_out[8697] <= layer0_out[2749] ^ layer0_out[2750];
     layer1_out[8698] <= ~layer0_out[11215];
     layer1_out[8699] <= ~layer0_out[11505] | layer0_out[11504];
     layer1_out[8700] <= ~layer0_out[3499];
     layer1_out[8701] <= ~(layer0_out[11978] ^ layer0_out[11979]);
     layer1_out[8702] <= layer0_out[10790] & ~layer0_out[10791];
     layer1_out[8703] <= layer0_out[2156] & layer0_out[2157];
     layer1_out[8704] <= 1'b0;
     layer1_out[8705] <= 1'b1;
     layer1_out[8706] <= layer0_out[7866] ^ layer0_out[7867];
     layer1_out[8707] <= layer0_out[8523] | layer0_out[8524];
     layer1_out[8708] <= ~layer0_out[10525];
     layer1_out[8709] <= ~layer0_out[2979];
     layer1_out[8710] <= layer0_out[8300] & ~layer0_out[8301];
     layer1_out[8711] <= ~(layer0_out[11174] ^ layer0_out[11175]);
     layer1_out[8712] <= layer0_out[4312] & layer0_out[4313];
     layer1_out[8713] <= layer0_out[9532];
     layer1_out[8714] <= layer0_out[5835];
     layer1_out[8715] <= layer0_out[9814] & ~layer0_out[9813];
     layer1_out[8716] <= layer0_out[6429];
     layer1_out[8717] <= ~layer0_out[2903] | layer0_out[2902];
     layer1_out[8718] <= layer0_out[10189] & ~layer0_out[10188];
     layer1_out[8719] <= ~layer0_out[9348];
     layer1_out[8720] <= ~layer0_out[7980];
     layer1_out[8721] <= layer0_out[2992];
     layer1_out[8722] <= ~layer0_out[2160];
     layer1_out[8723] <= layer0_out[7988];
     layer1_out[8724] <= ~layer0_out[9912] | layer0_out[9911];
     layer1_out[8725] <= layer0_out[5273];
     layer1_out[8726] <= ~layer0_out[7322] | layer0_out[7323];
     layer1_out[8727] <= layer0_out[7566] & ~layer0_out[7567];
     layer1_out[8728] <= ~(layer0_out[2857] & layer0_out[2858]);
     layer1_out[8729] <= layer0_out[5174] & ~layer0_out[5175];
     layer1_out[8730] <= ~layer0_out[6300] | layer0_out[6301];
     layer1_out[8731] <= ~layer0_out[7382];
     layer1_out[8732] <= ~(layer0_out[374] & layer0_out[375]);
     layer1_out[8733] <= ~(layer0_out[6004] ^ layer0_out[6005]);
     layer1_out[8734] <= layer0_out[1181];
     layer1_out[8735] <= layer0_out[5997];
     layer1_out[8736] <= layer0_out[2298] & ~layer0_out[2297];
     layer1_out[8737] <= layer0_out[101] & ~layer0_out[100];
     layer1_out[8738] <= ~layer0_out[2991] | layer0_out[2990];
     layer1_out[8739] <= 1'b0;
     layer1_out[8740] <= layer0_out[1855] | layer0_out[1856];
     layer1_out[8741] <= layer0_out[919];
     layer1_out[8742] <= ~(layer0_out[571] ^ layer0_out[572]);
     layer1_out[8743] <= ~layer0_out[8655];
     layer1_out[8744] <= ~(layer0_out[5129] | layer0_out[5130]);
     layer1_out[8745] <= layer0_out[5915] | layer0_out[5916];
     layer1_out[8746] <= layer0_out[6199] ^ layer0_out[6200];
     layer1_out[8747] <= layer0_out[11275];
     layer1_out[8748] <= ~(layer0_out[9545] | layer0_out[9546]);
     layer1_out[8749] <= layer0_out[1444];
     layer1_out[8750] <= layer0_out[7593] & ~layer0_out[7594];
     layer1_out[8751] <= layer0_out[2480];
     layer1_out[8752] <= layer0_out[9780];
     layer1_out[8753] <= ~(layer0_out[1333] | layer0_out[1334]);
     layer1_out[8754] <= ~(layer0_out[7737] & layer0_out[7738]);
     layer1_out[8755] <= layer0_out[8804];
     layer1_out[8756] <= ~(layer0_out[2844] | layer0_out[2845]);
     layer1_out[8757] <= ~layer0_out[16];
     layer1_out[8758] <= layer0_out[10846];
     layer1_out[8759] <= ~layer0_out[11000];
     layer1_out[8760] <= ~(layer0_out[10102] & layer0_out[10103]);
     layer1_out[8761] <= ~(layer0_out[10648] & layer0_out[10649]);
     layer1_out[8762] <= ~(layer0_out[10073] | layer0_out[10074]);
     layer1_out[8763] <= layer0_out[11524] & ~layer0_out[11525];
     layer1_out[8764] <= layer0_out[697] | layer0_out[698];
     layer1_out[8765] <= ~layer0_out[4747] | layer0_out[4746];
     layer1_out[8766] <= ~layer0_out[3615] | layer0_out[3614];
     layer1_out[8767] <= ~layer0_out[7331];
     layer1_out[8768] <= ~layer0_out[3366];
     layer1_out[8769] <= ~layer0_out[9265];
     layer1_out[8770] <= layer0_out[5311] & ~layer0_out[5310];
     layer1_out[8771] <= ~(layer0_out[8319] & layer0_out[8320]);
     layer1_out[8772] <= ~layer0_out[3464] | layer0_out[3465];
     layer1_out[8773] <= layer0_out[9295] & ~layer0_out[9294];
     layer1_out[8774] <= layer0_out[8249] ^ layer0_out[8250];
     layer1_out[8775] <= layer0_out[3860] & ~layer0_out[3861];
     layer1_out[8776] <= layer0_out[6584] & layer0_out[6585];
     layer1_out[8777] <= ~(layer0_out[223] & layer0_out[224]);
     layer1_out[8778] <= layer0_out[162];
     layer1_out[8779] <= layer0_out[10171];
     layer1_out[8780] <= ~layer0_out[2384] | layer0_out[2385];
     layer1_out[8781] <= layer0_out[10513] | layer0_out[10514];
     layer1_out[8782] <= layer0_out[5829];
     layer1_out[8783] <= layer0_out[973] & layer0_out[974];
     layer1_out[8784] <= ~(layer0_out[9685] & layer0_out[9686]);
     layer1_out[8785] <= layer0_out[4471];
     layer1_out[8786] <= layer0_out[5450] & layer0_out[5451];
     layer1_out[8787] <= ~layer0_out[7686];
     layer1_out[8788] <= ~(layer0_out[387] & layer0_out[388]);
     layer1_out[8789] <= ~layer0_out[11879];
     layer1_out[8790] <= layer0_out[8105];
     layer1_out[8791] <= ~layer0_out[6559] | layer0_out[6558];
     layer1_out[8792] <= ~layer0_out[1466] | layer0_out[1467];
     layer1_out[8793] <= layer0_out[6132] & layer0_out[6133];
     layer1_out[8794] <= layer0_out[2930];
     layer1_out[8795] <= ~(layer0_out[9574] ^ layer0_out[9575]);
     layer1_out[8796] <= layer0_out[2067];
     layer1_out[8797] <= layer0_out[9962] | layer0_out[9963];
     layer1_out[8798] <= ~layer0_out[9062] | layer0_out[9061];
     layer1_out[8799] <= layer0_out[5582];
     layer1_out[8800] <= ~(layer0_out[4320] | layer0_out[4321]);
     layer1_out[8801] <= ~(layer0_out[11759] & layer0_out[11760]);
     layer1_out[8802] <= layer0_out[8810];
     layer1_out[8803] <= layer0_out[8730] & ~layer0_out[8731];
     layer1_out[8804] <= ~layer0_out[3744];
     layer1_out[8805] <= ~(layer0_out[9267] & layer0_out[9268]);
     layer1_out[8806] <= ~(layer0_out[1904] ^ layer0_out[1905]);
     layer1_out[8807] <= layer0_out[1226] & ~layer0_out[1225];
     layer1_out[8808] <= ~layer0_out[11066];
     layer1_out[8809] <= ~layer0_out[6805];
     layer1_out[8810] <= layer0_out[10664] | layer0_out[10665];
     layer1_out[8811] <= ~(layer0_out[1845] ^ layer0_out[1846]);
     layer1_out[8812] <= layer0_out[5687] & ~layer0_out[5688];
     layer1_out[8813] <= layer0_out[11902] & layer0_out[11903];
     layer1_out[8814] <= layer0_out[5380];
     layer1_out[8815] <= ~(layer0_out[799] & layer0_out[800]);
     layer1_out[8816] <= layer0_out[5428];
     layer1_out[8817] <= ~layer0_out[373] | layer0_out[372];
     layer1_out[8818] <= layer0_out[7336];
     layer1_out[8819] <= layer0_out[11579] & layer0_out[11580];
     layer1_out[8820] <= ~layer0_out[4874];
     layer1_out[8821] <= ~(layer0_out[11736] & layer0_out[11737]);
     layer1_out[8822] <= ~layer0_out[235] | layer0_out[234];
     layer1_out[8823] <= ~layer0_out[1086];
     layer1_out[8824] <= 1'b0;
     layer1_out[8825] <= ~layer0_out[10769];
     layer1_out[8826] <= layer0_out[4189] ^ layer0_out[4190];
     layer1_out[8827] <= layer0_out[1432] & ~layer0_out[1431];
     layer1_out[8828] <= layer0_out[5052] & ~layer0_out[5053];
     layer1_out[8829] <= ~layer0_out[4770] | layer0_out[4771];
     layer1_out[8830] <= layer0_out[10804] & ~layer0_out[10805];
     layer1_out[8831] <= ~layer0_out[7604] | layer0_out[7605];
     layer1_out[8832] <= layer0_out[5217];
     layer1_out[8833] <= layer0_out[3750] | layer0_out[3751];
     layer1_out[8834] <= layer0_out[10607] & layer0_out[10608];
     layer1_out[8835] <= ~(layer0_out[9984] & layer0_out[9985]);
     layer1_out[8836] <= layer0_out[4904] & ~layer0_out[4903];
     layer1_out[8837] <= 1'b1;
     layer1_out[8838] <= layer0_out[3362] ^ layer0_out[3363];
     layer1_out[8839] <= ~layer0_out[3569];
     layer1_out[8840] <= ~layer0_out[8963];
     layer1_out[8841] <= ~layer0_out[3252];
     layer1_out[8842] <= ~layer0_out[1471] | layer0_out[1472];
     layer1_out[8843] <= layer0_out[2396] & ~layer0_out[2397];
     layer1_out[8844] <= layer0_out[8022];
     layer1_out[8845] <= layer0_out[11741];
     layer1_out[8846] <= layer0_out[9653];
     layer1_out[8847] <= ~layer0_out[2602];
     layer1_out[8848] <= ~layer0_out[11930];
     layer1_out[8849] <= layer0_out[2182] & layer0_out[2183];
     layer1_out[8850] <= layer0_out[6121] & ~layer0_out[6120];
     layer1_out[8851] <= ~layer0_out[256];
     layer1_out[8852] <= layer0_out[9505];
     layer1_out[8853] <= layer0_out[4081];
     layer1_out[8854] <= 1'b0;
     layer1_out[8855] <= ~layer0_out[8760];
     layer1_out[8856] <= layer0_out[1730];
     layer1_out[8857] <= ~layer0_out[3890] | layer0_out[3891];
     layer1_out[8858] <= layer0_out[3846] | layer0_out[3847];
     layer1_out[8859] <= ~layer0_out[8214] | layer0_out[8213];
     layer1_out[8860] <= layer0_out[9526] & ~layer0_out[9525];
     layer1_out[8861] <= ~layer0_out[2480] | layer0_out[2481];
     layer1_out[8862] <= layer0_out[4406] | layer0_out[4407];
     layer1_out[8863] <= ~(layer0_out[5477] & layer0_out[5478]);
     layer1_out[8864] <= layer0_out[2578];
     layer1_out[8865] <= layer0_out[10770] | layer0_out[10771];
     layer1_out[8866] <= ~(layer0_out[1273] | layer0_out[1274]);
     layer1_out[8867] <= ~layer0_out[9471] | layer0_out[9472];
     layer1_out[8868] <= layer0_out[11082];
     layer1_out[8869] <= ~layer0_out[5906];
     layer1_out[8870] <= layer0_out[4682] | layer0_out[4683];
     layer1_out[8871] <= ~layer0_out[3118] | layer0_out[3117];
     layer1_out[8872] <= layer0_out[9857];
     layer1_out[8873] <= ~layer0_out[5486];
     layer1_out[8874] <= ~layer0_out[1231];
     layer1_out[8875] <= layer0_out[8019];
     layer1_out[8876] <= ~layer0_out[2634] | layer0_out[2633];
     layer1_out[8877] <= layer0_out[9223];
     layer1_out[8878] <= layer0_out[9037];
     layer1_out[8879] <= layer0_out[9975] & layer0_out[9976];
     layer1_out[8880] <= layer0_out[11439] | layer0_out[11440];
     layer1_out[8881] <= ~layer0_out[305];
     layer1_out[8882] <= layer0_out[6870] & ~layer0_out[6871];
     layer1_out[8883] <= ~(layer0_out[6606] & layer0_out[6607]);
     layer1_out[8884] <= layer0_out[1027] ^ layer0_out[1028];
     layer1_out[8885] <= ~layer0_out[2541] | layer0_out[2540];
     layer1_out[8886] <= layer0_out[10501] | layer0_out[10502];
     layer1_out[8887] <= ~(layer0_out[9495] | layer0_out[9496]);
     layer1_out[8888] <= layer0_out[7818] | layer0_out[7819];
     layer1_out[8889] <= ~(layer0_out[310] | layer0_out[311]);
     layer1_out[8890] <= ~(layer0_out[6546] ^ layer0_out[6547]);
     layer1_out[8891] <= ~(layer0_out[4446] & layer0_out[4447]);
     layer1_out[8892] <= ~layer0_out[3063];
     layer1_out[8893] <= ~(layer0_out[10411] | layer0_out[10412]);
     layer1_out[8894] <= layer0_out[131] & layer0_out[132];
     layer1_out[8895] <= ~layer0_out[8534];
     layer1_out[8896] <= layer0_out[11461] & ~layer0_out[11462];
     layer1_out[8897] <= layer0_out[11995];
     layer1_out[8898] <= layer0_out[1669] ^ layer0_out[1670];
     layer1_out[8899] <= ~(layer0_out[9625] & layer0_out[9626]);
     layer1_out[8900] <= ~layer0_out[8826];
     layer1_out[8901] <= layer0_out[11941];
     layer1_out[8902] <= ~layer0_out[4016];
     layer1_out[8903] <= layer0_out[6547] | layer0_out[6548];
     layer1_out[8904] <= ~layer0_out[10523] | layer0_out[10522];
     layer1_out[8905] <= ~(layer0_out[7928] | layer0_out[7929]);
     layer1_out[8906] <= ~layer0_out[4433];
     layer1_out[8907] <= layer0_out[11166];
     layer1_out[8908] <= ~(layer0_out[11139] ^ layer0_out[11140]);
     layer1_out[8909] <= ~layer0_out[10857];
     layer1_out[8910] <= ~(layer0_out[6054] & layer0_out[6055]);
     layer1_out[8911] <= ~layer0_out[10085] | layer0_out[10084];
     layer1_out[8912] <= layer0_out[1938] & ~layer0_out[1939];
     layer1_out[8913] <= layer0_out[9228];
     layer1_out[8914] <= layer0_out[10605] & ~layer0_out[10606];
     layer1_out[8915] <= ~layer0_out[997] | layer0_out[998];
     layer1_out[8916] <= ~(layer0_out[6761] ^ layer0_out[6762]);
     layer1_out[8917] <= layer0_out[1932] ^ layer0_out[1933];
     layer1_out[8918] <= ~(layer0_out[774] | layer0_out[775]);
     layer1_out[8919] <= layer0_out[2408];
     layer1_out[8920] <= ~(layer0_out[8434] & layer0_out[8435]);
     layer1_out[8921] <= ~layer0_out[860] | layer0_out[861];
     layer1_out[8922] <= ~layer0_out[5401] | layer0_out[5400];
     layer1_out[8923] <= layer0_out[2593] & layer0_out[2594];
     layer1_out[8924] <= layer0_out[1888];
     layer1_out[8925] <= ~layer0_out[10324];
     layer1_out[8926] <= layer0_out[11017] & ~layer0_out[11016];
     layer1_out[8927] <= layer0_out[560];
     layer1_out[8928] <= layer0_out[3560] | layer0_out[3561];
     layer1_out[8929] <= layer0_out[834];
     layer1_out[8930] <= ~layer0_out[4459];
     layer1_out[8931] <= layer0_out[10877] & ~layer0_out[10876];
     layer1_out[8932] <= ~layer0_out[9222] | layer0_out[9221];
     layer1_out[8933] <= ~layer0_out[2893];
     layer1_out[8934] <= ~layer0_out[10033];
     layer1_out[8935] <= layer0_out[11993] & ~layer0_out[11992];
     layer1_out[8936] <= 1'b0;
     layer1_out[8937] <= 1'b0;
     layer1_out[8938] <= layer0_out[11353];
     layer1_out[8939] <= ~(layer0_out[8849] | layer0_out[8850]);
     layer1_out[8940] <= ~layer0_out[3398] | layer0_out[3399];
     layer1_out[8941] <= ~layer0_out[11881];
     layer1_out[8942] <= layer0_out[8366] ^ layer0_out[8367];
     layer1_out[8943] <= ~layer0_out[9683];
     layer1_out[8944] <= ~(layer0_out[4452] | layer0_out[4453]);
     layer1_out[8945] <= ~layer0_out[3391];
     layer1_out[8946] <= layer0_out[5776] | layer0_out[5777];
     layer1_out[8947] <= layer0_out[10316] | layer0_out[10317];
     layer1_out[8948] <= layer0_out[6903] & ~layer0_out[6904];
     layer1_out[8949] <= layer0_out[11205] & ~layer0_out[11204];
     layer1_out[8950] <= layer0_out[6202] & ~layer0_out[6201];
     layer1_out[8951] <= ~(layer0_out[5739] | layer0_out[5740]);
     layer1_out[8952] <= ~layer0_out[4798];
     layer1_out[8953] <= ~layer0_out[10105] | layer0_out[10106];
     layer1_out[8954] <= 1'b1;
     layer1_out[8955] <= ~layer0_out[8557];
     layer1_out[8956] <= ~layer0_out[8186];
     layer1_out[8957] <= layer0_out[11293] & ~layer0_out[11294];
     layer1_out[8958] <= layer0_out[11217];
     layer1_out[8959] <= layer0_out[7591] & layer0_out[7592];
     layer1_out[8960] <= layer0_out[7607] | layer0_out[7608];
     layer1_out[8961] <= layer0_out[8475] & layer0_out[8476];
     layer1_out[8962] <= ~layer0_out[598];
     layer1_out[8963] <= layer0_out[1003] & ~layer0_out[1002];
     layer1_out[8964] <= layer0_out[10198] & layer0_out[10199];
     layer1_out[8965] <= ~layer0_out[4821];
     layer1_out[8966] <= layer0_out[1890];
     layer1_out[8967] <= layer0_out[5841] & layer0_out[5842];
     layer1_out[8968] <= layer0_out[5417];
     layer1_out[8969] <= ~(layer0_out[2227] ^ layer0_out[2228]);
     layer1_out[8970] <= layer0_out[7764];
     layer1_out[8971] <= ~layer0_out[6672] | layer0_out[6673];
     layer1_out[8972] <= ~(layer0_out[11167] | layer0_out[11168]);
     layer1_out[8973] <= layer0_out[10754] & layer0_out[10755];
     layer1_out[8974] <= ~(layer0_out[1035] & layer0_out[1036]);
     layer1_out[8975] <= ~layer0_out[5611];
     layer1_out[8976] <= layer0_out[1402];
     layer1_out[8977] <= layer0_out[3146];
     layer1_out[8978] <= ~(layer0_out[7340] & layer0_out[7341]);
     layer1_out[8979] <= 1'b1;
     layer1_out[8980] <= layer0_out[1537] & ~layer0_out[1538];
     layer1_out[8981] <= ~(layer0_out[11061] | layer0_out[11062]);
     layer1_out[8982] <= layer0_out[9033];
     layer1_out[8983] <= ~layer0_out[10380];
     layer1_out[8984] <= layer0_out[1588];
     layer1_out[8985] <= ~layer0_out[4454] | layer0_out[4453];
     layer1_out[8986] <= layer0_out[5632] ^ layer0_out[5633];
     layer1_out[8987] <= ~(layer0_out[4007] | layer0_out[4008]);
     layer1_out[8988] <= ~(layer0_out[11594] & layer0_out[11595]);
     layer1_out[8989] <= ~(layer0_out[238] & layer0_out[239]);
     layer1_out[8990] <= ~layer0_out[11407];
     layer1_out[8991] <= layer0_out[10197] | layer0_out[10198];
     layer1_out[8992] <= ~layer0_out[5727];
     layer1_out[8993] <= layer0_out[4702];
     layer1_out[8994] <= 1'b1;
     layer1_out[8995] <= ~(layer0_out[2930] & layer0_out[2931]);
     layer1_out[8996] <= ~layer0_out[5753];
     layer1_out[8997] <= ~layer0_out[5065];
     layer1_out[8998] <= layer0_out[8135];
     layer1_out[8999] <= ~(layer0_out[9041] ^ layer0_out[9042]);
     layer1_out[9000] <= layer0_out[9714] & ~layer0_out[9715];
     layer1_out[9001] <= layer0_out[8184] & ~layer0_out[8183];
     layer1_out[9002] <= ~(layer0_out[9492] & layer0_out[9493]);
     layer1_out[9003] <= layer0_out[8398] & layer0_out[8399];
     layer1_out[9004] <= layer0_out[936] & layer0_out[937];
     layer1_out[9005] <= layer0_out[7698] ^ layer0_out[7699];
     layer1_out[9006] <= layer0_out[10967];
     layer1_out[9007] <= ~layer0_out[10572];
     layer1_out[9008] <= ~(layer0_out[2743] ^ layer0_out[2744]);
     layer1_out[9009] <= layer0_out[8751] | layer0_out[8752];
     layer1_out[9010] <= ~(layer0_out[5669] | layer0_out[5670]);
     layer1_out[9011] <= layer0_out[6889] ^ layer0_out[6890];
     layer1_out[9012] <= ~layer0_out[6521];
     layer1_out[9013] <= layer0_out[7146] & ~layer0_out[7147];
     layer1_out[9014] <= layer0_out[7831] ^ layer0_out[7832];
     layer1_out[9015] <= layer0_out[3231];
     layer1_out[9016] <= layer0_out[11661] ^ layer0_out[11662];
     layer1_out[9017] <= ~layer0_out[7433] | layer0_out[7432];
     layer1_out[9018] <= ~layer0_out[1057];
     layer1_out[9019] <= ~layer0_out[11996];
     layer1_out[9020] <= ~(layer0_out[10231] & layer0_out[10232]);
     layer1_out[9021] <= ~layer0_out[2156];
     layer1_out[9022] <= ~layer0_out[11297];
     layer1_out[9023] <= layer0_out[6572] & ~layer0_out[6571];
     layer1_out[9024] <= ~layer0_out[11709];
     layer1_out[9025] <= layer0_out[8796];
     layer1_out[9026] <= ~(layer0_out[7600] ^ layer0_out[7601]);
     layer1_out[9027] <= 1'b1;
     layer1_out[9028] <= ~layer0_out[2566];
     layer1_out[9029] <= layer0_out[1453] & ~layer0_out[1454];
     layer1_out[9030] <= 1'b1;
     layer1_out[9031] <= layer0_out[9299] | layer0_out[9300];
     layer1_out[9032] <= ~(layer0_out[3099] & layer0_out[3100]);
     layer1_out[9033] <= ~layer0_out[7469];
     layer1_out[9034] <= ~(layer0_out[9159] | layer0_out[9160]);
     layer1_out[9035] <= layer0_out[2224];
     layer1_out[9036] <= layer0_out[10915] & ~layer0_out[10914];
     layer1_out[9037] <= layer0_out[810];
     layer1_out[9038] <= layer0_out[7744] & ~layer0_out[7743];
     layer1_out[9039] <= layer0_out[9181] & layer0_out[9182];
     layer1_out[9040] <= ~(layer0_out[10472] ^ layer0_out[10473]);
     layer1_out[9041] <= layer0_out[3905] & layer0_out[3906];
     layer1_out[9042] <= ~layer0_out[1863];
     layer1_out[9043] <= ~(layer0_out[6831] & layer0_out[6832]);
     layer1_out[9044] <= ~(layer0_out[5975] | layer0_out[5976]);
     layer1_out[9045] <= layer0_out[5898];
     layer1_out[9046] <= ~layer0_out[7196];
     layer1_out[9047] <= layer0_out[498];
     layer1_out[9048] <= ~layer0_out[147] | layer0_out[148];
     layer1_out[9049] <= layer0_out[5091];
     layer1_out[9050] <= layer0_out[10883] | layer0_out[10884];
     layer1_out[9051] <= layer0_out[8040] | layer0_out[8041];
     layer1_out[9052] <= ~layer0_out[10961] | layer0_out[10962];
     layer1_out[9053] <= layer0_out[8645];
     layer1_out[9054] <= ~layer0_out[1895];
     layer1_out[9055] <= ~layer0_out[5483] | layer0_out[5482];
     layer1_out[9056] <= layer0_out[4400] | layer0_out[4401];
     layer1_out[9057] <= layer0_out[115] | layer0_out[116];
     layer1_out[9058] <= ~(layer0_out[10588] & layer0_out[10589]);
     layer1_out[9059] <= ~(layer0_out[2584] & layer0_out[2585]);
     layer1_out[9060] <= ~layer0_out[10428];
     layer1_out[9061] <= layer0_out[11969] & ~layer0_out[11968];
     layer1_out[9062] <= ~(layer0_out[1421] ^ layer0_out[1422]);
     layer1_out[9063] <= ~layer0_out[684];
     layer1_out[9064] <= ~layer0_out[11287];
     layer1_out[9065] <= layer0_out[2000];
     layer1_out[9066] <= ~(layer0_out[6631] | layer0_out[6632]);
     layer1_out[9067] <= ~layer0_out[5218];
     layer1_out[9068] <= layer0_out[5250] & ~layer0_out[5251];
     layer1_out[9069] <= layer0_out[11875] ^ layer0_out[11876];
     layer1_out[9070] <= ~layer0_out[11209];
     layer1_out[9071] <= ~layer0_out[6737];
     layer1_out[9072] <= ~layer0_out[6851];
     layer1_out[9073] <= layer0_out[10335];
     layer1_out[9074] <= ~layer0_out[11023] | layer0_out[11022];
     layer1_out[9075] <= layer0_out[8470] & ~layer0_out[8469];
     layer1_out[9076] <= layer0_out[3951];
     layer1_out[9077] <= layer0_out[512] ^ layer0_out[513];
     layer1_out[9078] <= ~layer0_out[10297];
     layer1_out[9079] <= layer0_out[8132] ^ layer0_out[8133];
     layer1_out[9080] <= layer0_out[147] & ~layer0_out[146];
     layer1_out[9081] <= layer0_out[3279];
     layer1_out[9082] <= 1'b1;
     layer1_out[9083] <= ~layer0_out[3619];
     layer1_out[9084] <= ~layer0_out[7983];
     layer1_out[9085] <= layer0_out[5927];
     layer1_out[9086] <= layer0_out[5458] | layer0_out[5459];
     layer1_out[9087] <= ~layer0_out[10157] | layer0_out[10156];
     layer1_out[9088] <= layer0_out[5184];
     layer1_out[9089] <= ~(layer0_out[4362] & layer0_out[4363]);
     layer1_out[9090] <= ~layer0_out[11189];
     layer1_out[9091] <= layer0_out[3435] & ~layer0_out[3436];
     layer1_out[9092] <= layer0_out[9250] ^ layer0_out[9251];
     layer1_out[9093] <= ~layer0_out[4416] | layer0_out[4415];
     layer1_out[9094] <= layer0_out[9546];
     layer1_out[9095] <= ~layer0_out[4774];
     layer1_out[9096] <= layer0_out[6060] & ~layer0_out[6061];
     layer1_out[9097] <= layer0_out[9] & layer0_out[10];
     layer1_out[9098] <= layer0_out[10172] & ~layer0_out[10173];
     layer1_out[9099] <= layer0_out[7681] & layer0_out[7682];
     layer1_out[9100] <= ~(layer0_out[9927] & layer0_out[9928]);
     layer1_out[9101] <= layer0_out[9450] & ~layer0_out[9451];
     layer1_out[9102] <= layer0_out[5839];
     layer1_out[9103] <= layer0_out[399];
     layer1_out[9104] <= layer0_out[10843];
     layer1_out[9105] <= layer0_out[3091] & layer0_out[3092];
     layer1_out[9106] <= layer0_out[8764];
     layer1_out[9107] <= ~layer0_out[4240];
     layer1_out[9108] <= ~layer0_out[7557] | layer0_out[7556];
     layer1_out[9109] <= ~layer0_out[10636];
     layer1_out[9110] <= layer0_out[6899] & layer0_out[6900];
     layer1_out[9111] <= ~(layer0_out[3415] & layer0_out[3416]);
     layer1_out[9112] <= ~layer0_out[8837];
     layer1_out[9113] <= layer0_out[3782] & ~layer0_out[3781];
     layer1_out[9114] <= layer0_out[4902];
     layer1_out[9115] <= layer0_out[2617];
     layer1_out[9116] <= layer0_out[3833] | layer0_out[3834];
     layer1_out[9117] <= ~layer0_out[7005] | layer0_out[7006];
     layer1_out[9118] <= layer0_out[9890] & ~layer0_out[9891];
     layer1_out[9119] <= ~(layer0_out[8599] & layer0_out[8600]);
     layer1_out[9120] <= layer0_out[7674] | layer0_out[7675];
     layer1_out[9121] <= layer0_out[950];
     layer1_out[9122] <= layer0_out[11437] & layer0_out[11438];
     layer1_out[9123] <= ~layer0_out[6226];
     layer1_out[9124] <= layer0_out[10849];
     layer1_out[9125] <= ~(layer0_out[3982] & layer0_out[3983]);
     layer1_out[9126] <= layer0_out[4232] | layer0_out[4233];
     layer1_out[9127] <= 1'b1;
     layer1_out[9128] <= ~layer0_out[5399] | layer0_out[5398];
     layer1_out[9129] <= layer0_out[3156] & ~layer0_out[3157];
     layer1_out[9130] <= ~layer0_out[4764];
     layer1_out[9131] <= layer0_out[3669] & ~layer0_out[3670];
     layer1_out[9132] <= ~layer0_out[6713];
     layer1_out[9133] <= layer0_out[587] & ~layer0_out[586];
     layer1_out[9134] <= layer0_out[2209];
     layer1_out[9135] <= layer0_out[11738];
     layer1_out[9136] <= layer0_out[6695] | layer0_out[6696];
     layer1_out[9137] <= ~layer0_out[5045] | layer0_out[5046];
     layer1_out[9138] <= layer0_out[6629] | layer0_out[6630];
     layer1_out[9139] <= layer0_out[10747] & ~layer0_out[10748];
     layer1_out[9140] <= layer0_out[3510] & layer0_out[3511];
     layer1_out[9141] <= layer0_out[8691] & ~layer0_out[8692];
     layer1_out[9142] <= layer0_out[5023];
     layer1_out[9143] <= layer0_out[219] & ~layer0_out[220];
     layer1_out[9144] <= ~(layer0_out[4535] | layer0_out[4536]);
     layer1_out[9145] <= ~(layer0_out[1589] ^ layer0_out[1590]);
     layer1_out[9146] <= layer0_out[3109] & layer0_out[3110];
     layer1_out[9147] <= layer0_out[7176];
     layer1_out[9148] <= 1'b0;
     layer1_out[9149] <= layer0_out[7277] & layer0_out[7278];
     layer1_out[9150] <= ~(layer0_out[1205] & layer0_out[1206]);
     layer1_out[9151] <= ~layer0_out[11650];
     layer1_out[9152] <= layer0_out[5832];
     layer1_out[9153] <= ~layer0_out[4632] | layer0_out[4633];
     layer1_out[9154] <= ~(layer0_out[5701] | layer0_out[5702]);
     layer1_out[9155] <= ~layer0_out[205];
     layer1_out[9156] <= ~layer0_out[3674] | layer0_out[3673];
     layer1_out[9157] <= layer0_out[4379] & layer0_out[4380];
     layer1_out[9158] <= layer0_out[9845] | layer0_out[9846];
     layer1_out[9159] <= ~layer0_out[2150];
     layer1_out[9160] <= ~layer0_out[580] | layer0_out[581];
     layer1_out[9161] <= layer0_out[8576] & ~layer0_out[8575];
     layer1_out[9162] <= ~(layer0_out[2804] & layer0_out[2805]);
     layer1_out[9163] <= ~(layer0_out[450] | layer0_out[451]);
     layer1_out[9164] <= layer0_out[5800];
     layer1_out[9165] <= ~layer0_out[4360];
     layer1_out[9166] <= ~layer0_out[10001];
     layer1_out[9167] <= ~layer0_out[8639];
     layer1_out[9168] <= layer0_out[11890] & ~layer0_out[11891];
     layer1_out[9169] <= ~(layer0_out[9695] & layer0_out[9696]);
     layer1_out[9170] <= layer0_out[11996];
     layer1_out[9171] <= ~layer0_out[7033];
     layer1_out[9172] <= layer0_out[6183] & ~layer0_out[6182];
     layer1_out[9173] <= ~layer0_out[5677] | layer0_out[5678];
     layer1_out[9174] <= layer0_out[3821];
     layer1_out[9175] <= layer0_out[6963] ^ layer0_out[6964];
     layer1_out[9176] <= ~(layer0_out[8778] & layer0_out[8779]);
     layer1_out[9177] <= ~layer0_out[7351] | layer0_out[7350];
     layer1_out[9178] <= layer0_out[9610];
     layer1_out[9179] <= layer0_out[449] & ~layer0_out[450];
     layer1_out[9180] <= layer0_out[3765] & ~layer0_out[3764];
     layer1_out[9181] <= layer0_out[5712] & ~layer0_out[5711];
     layer1_out[9182] <= ~layer0_out[9798];
     layer1_out[9183] <= layer0_out[3499] ^ layer0_out[3500];
     layer1_out[9184] <= ~(layer0_out[2417] ^ layer0_out[2418]);
     layer1_out[9185] <= ~layer0_out[5009] | layer0_out[5010];
     layer1_out[9186] <= ~layer0_out[2059];
     layer1_out[9187] <= ~(layer0_out[10347] & layer0_out[10348]);
     layer1_out[9188] <= layer0_out[1128];
     layer1_out[9189] <= ~layer0_out[5647];
     layer1_out[9190] <= ~layer0_out[9794];
     layer1_out[9191] <= layer0_out[3175] & ~layer0_out[3174];
     layer1_out[9192] <= layer0_out[5098];
     layer1_out[9193] <= ~(layer0_out[3651] | layer0_out[3652]);
     layer1_out[9194] <= ~layer0_out[3949];
     layer1_out[9195] <= layer0_out[8833] | layer0_out[8834];
     layer1_out[9196] <= layer0_out[9240];
     layer1_out[9197] <= layer0_out[5425] & layer0_out[5426];
     layer1_out[9198] <= layer0_out[44] & ~layer0_out[43];
     layer1_out[9199] <= ~layer0_out[7705];
     layer1_out[9200] <= ~layer0_out[1919];
     layer1_out[9201] <= ~layer0_out[3486] | layer0_out[3485];
     layer1_out[9202] <= layer0_out[2593];
     layer1_out[9203] <= 1'b1;
     layer1_out[9204] <= layer0_out[84] & ~layer0_out[85];
     layer1_out[9205] <= ~(layer0_out[1603] | layer0_out[1604]);
     layer1_out[9206] <= ~layer0_out[6624];
     layer1_out[9207] <= layer0_out[6373] | layer0_out[6374];
     layer1_out[9208] <= ~layer0_out[10124];
     layer1_out[9209] <= ~layer0_out[7174];
     layer1_out[9210] <= layer0_out[9339];
     layer1_out[9211] <= 1'b0;
     layer1_out[9212] <= ~(layer0_out[3639] & layer0_out[3640]);
     layer1_out[9213] <= layer0_out[8408];
     layer1_out[9214] <= 1'b0;
     layer1_out[9215] <= ~layer0_out[11408] | layer0_out[11409];
     layer1_out[9216] <= layer0_out[4599] ^ layer0_out[4600];
     layer1_out[9217] <= layer0_out[8134];
     layer1_out[9218] <= layer0_out[2910] & ~layer0_out[2911];
     layer1_out[9219] <= ~layer0_out[1859];
     layer1_out[9220] <= ~layer0_out[4430];
     layer1_out[9221] <= ~layer0_out[2346];
     layer1_out[9222] <= 1'b1;
     layer1_out[9223] <= ~layer0_out[6683];
     layer1_out[9224] <= ~(layer0_out[8818] ^ layer0_out[8819]);
     layer1_out[9225] <= ~layer0_out[7727];
     layer1_out[9226] <= layer0_out[1004];
     layer1_out[9227] <= layer0_out[1527] & layer0_out[1528];
     layer1_out[9228] <= layer0_out[2205] ^ layer0_out[2206];
     layer1_out[9229] <= layer0_out[5987] & ~layer0_out[5986];
     layer1_out[9230] <= layer0_out[9387] & layer0_out[9388];
     layer1_out[9231] <= layer0_out[4509] & ~layer0_out[4510];
     layer1_out[9232] <= ~(layer0_out[708] ^ layer0_out[709]);
     layer1_out[9233] <= ~layer0_out[870];
     layer1_out[9234] <= ~layer0_out[9758] | layer0_out[9759];
     layer1_out[9235] <= layer0_out[7526];
     layer1_out[9236] <= layer0_out[3694];
     layer1_out[9237] <= layer0_out[7325] | layer0_out[7326];
     layer1_out[9238] <= layer0_out[2055];
     layer1_out[9239] <= layer0_out[9210] ^ layer0_out[9211];
     layer1_out[9240] <= layer0_out[6164];
     layer1_out[9241] <= layer0_out[11635] & ~layer0_out[11634];
     layer1_out[9242] <= layer0_out[3031];
     layer1_out[9243] <= ~(layer0_out[10541] & layer0_out[10542]);
     layer1_out[9244] <= layer0_out[7489];
     layer1_out[9245] <= layer0_out[10538] | layer0_out[10539];
     layer1_out[9246] <= layer0_out[518] & ~layer0_out[517];
     layer1_out[9247] <= layer0_out[11123];
     layer1_out[9248] <= layer0_out[6588];
     layer1_out[9249] <= layer0_out[1228] ^ layer0_out[1229];
     layer1_out[9250] <= layer0_out[11677];
     layer1_out[9251] <= layer0_out[8273] & ~layer0_out[8274];
     layer1_out[9252] <= ~layer0_out[6799];
     layer1_out[9253] <= ~(layer0_out[660] ^ layer0_out[661]);
     layer1_out[9254] <= ~layer0_out[458];
     layer1_out[9255] <= layer0_out[10206];
     layer1_out[9256] <= ~layer0_out[8499];
     layer1_out[9257] <= layer0_out[5452] | layer0_out[5453];
     layer1_out[9258] <= ~layer0_out[7268];
     layer1_out[9259] <= layer0_out[5932] & ~layer0_out[5933];
     layer1_out[9260] <= ~layer0_out[1183] | layer0_out[1182];
     layer1_out[9261] <= layer0_out[5754] & layer0_out[5755];
     layer1_out[9262] <= layer0_out[9397] | layer0_out[9398];
     layer1_out[9263] <= layer0_out[4541] & layer0_out[4542];
     layer1_out[9264] <= ~layer0_out[9297];
     layer1_out[9265] <= layer0_out[11967];
     layer1_out[9266] <= ~(layer0_out[8462] & layer0_out[8463]);
     layer1_out[9267] <= ~layer0_out[781];
     layer1_out[9268] <= layer0_out[7974] & ~layer0_out[7975];
     layer1_out[9269] <= layer0_out[4838] & ~layer0_out[4837];
     layer1_out[9270] <= layer0_out[4062] | layer0_out[4063];
     layer1_out[9271] <= ~(layer0_out[2063] | layer0_out[2064]);
     layer1_out[9272] <= ~(layer0_out[9703] | layer0_out[9704]);
     layer1_out[9273] <= ~layer0_out[7411];
     layer1_out[9274] <= ~layer0_out[7803];
     layer1_out[9275] <= ~layer0_out[3097];
     layer1_out[9276] <= layer0_out[4024] & layer0_out[4025];
     layer1_out[9277] <= layer0_out[8042] ^ layer0_out[8043];
     layer1_out[9278] <= layer0_out[5456] | layer0_out[5457];
     layer1_out[9279] <= layer0_out[1084] & ~layer0_out[1085];
     layer1_out[9280] <= layer0_out[5869] & ~layer0_out[5868];
     layer1_out[9281] <= layer0_out[2166] & ~layer0_out[2167];
     layer1_out[9282] <= ~(layer0_out[1341] & layer0_out[1342]);
     layer1_out[9283] <= layer0_out[32];
     layer1_out[9284] <= layer0_out[10695];
     layer1_out[9285] <= ~layer0_out[1232] | layer0_out[1233];
     layer1_out[9286] <= ~layer0_out[7459];
     layer1_out[9287] <= ~layer0_out[5] | layer0_out[4];
     layer1_out[9288] <= ~layer0_out[7450] | layer0_out[7449];
     layer1_out[9289] <= ~layer0_out[6254];
     layer1_out[9290] <= layer0_out[10761];
     layer1_out[9291] <= layer0_out[6133];
     layer1_out[9292] <= layer0_out[3062] & ~layer0_out[3061];
     layer1_out[9293] <= ~layer0_out[8681];
     layer1_out[9294] <= layer0_out[4764];
     layer1_out[9295] <= ~layer0_out[351] | layer0_out[352];
     layer1_out[9296] <= layer0_out[5290];
     layer1_out[9297] <= ~layer0_out[1318] | layer0_out[1317];
     layer1_out[9298] <= layer0_out[2281] & ~layer0_out[2280];
     layer1_out[9299] <= ~layer0_out[4209];
     layer1_out[9300] <= ~(layer0_out[1427] ^ layer0_out[1428]);
     layer1_out[9301] <= layer0_out[10079] & layer0_out[10080];
     layer1_out[9302] <= layer0_out[9455];
     layer1_out[9303] <= 1'b1;
     layer1_out[9304] <= 1'b1;
     layer1_out[9305] <= layer0_out[3738] & ~layer0_out[3737];
     layer1_out[9306] <= ~layer0_out[7401] | layer0_out[7400];
     layer1_out[9307] <= layer0_out[7606] | layer0_out[7607];
     layer1_out[9308] <= layer0_out[9799] | layer0_out[9800];
     layer1_out[9309] <= ~(layer0_out[11854] & layer0_out[11855]);
     layer1_out[9310] <= ~(layer0_out[11900] | layer0_out[11901]);
     layer1_out[9311] <= layer0_out[3064] & ~layer0_out[3065];
     layer1_out[9312] <= ~layer0_out[7548];
     layer1_out[9313] <= ~layer0_out[3779] | layer0_out[3780];
     layer1_out[9314] <= layer0_out[8119];
     layer1_out[9315] <= ~layer0_out[2539] | layer0_out[2540];
     layer1_out[9316] <= ~layer0_out[11241];
     layer1_out[9317] <= ~(layer0_out[7965] | layer0_out[7966]);
     layer1_out[9318] <= 1'b0;
     layer1_out[9319] <= layer0_out[6529] & layer0_out[6530];
     layer1_out[9320] <= ~(layer0_out[2173] ^ layer0_out[2174]);
     layer1_out[9321] <= layer0_out[1919] & layer0_out[1920];
     layer1_out[9322] <= layer0_out[1455];
     layer1_out[9323] <= layer0_out[5989] & layer0_out[5990];
     layer1_out[9324] <= layer0_out[2865];
     layer1_out[9325] <= ~(layer0_out[4229] & layer0_out[4230]);
     layer1_out[9326] <= layer0_out[108] | layer0_out[109];
     layer1_out[9327] <= layer0_out[6135] & ~layer0_out[6136];
     layer1_out[9328] <= ~layer0_out[9115] | layer0_out[9116];
     layer1_out[9329] <= layer0_out[6259] & ~layer0_out[6260];
     layer1_out[9330] <= ~layer0_out[11834];
     layer1_out[9331] <= 1'b0;
     layer1_out[9332] <= 1'b1;
     layer1_out[9333] <= layer0_out[3413] | layer0_out[3414];
     layer1_out[9334] <= layer0_out[3911] | layer0_out[3912];
     layer1_out[9335] <= layer0_out[8861];
     layer1_out[9336] <= ~(layer0_out[7473] & layer0_out[7474]);
     layer1_out[9337] <= layer0_out[7509] & ~layer0_out[7508];
     layer1_out[9338] <= layer0_out[4712] | layer0_out[4713];
     layer1_out[9339] <= layer0_out[6149];
     layer1_out[9340] <= ~layer0_out[3344];
     layer1_out[9341] <= layer0_out[3612] & ~layer0_out[3613];
     layer1_out[9342] <= layer0_out[9597];
     layer1_out[9343] <= ~layer0_out[7542];
     layer1_out[9344] <= ~layer0_out[2645];
     layer1_out[9345] <= ~(layer0_out[5558] | layer0_out[5559]);
     layer1_out[9346] <= layer0_out[3311];
     layer1_out[9347] <= ~(layer0_out[8512] | layer0_out[8513]);
     layer1_out[9348] <= layer0_out[9521] & layer0_out[9522];
     layer1_out[9349] <= ~(layer0_out[5935] & layer0_out[5936]);
     layer1_out[9350] <= layer0_out[9185] & ~layer0_out[9186];
     layer1_out[9351] <= ~layer0_out[7471];
     layer1_out[9352] <= layer0_out[1330];
     layer1_out[9353] <= ~layer0_out[4888];
     layer1_out[9354] <= layer0_out[8722] & ~layer0_out[8721];
     layer1_out[9355] <= 1'b0;
     layer1_out[9356] <= ~(layer0_out[6490] | layer0_out[6491]);
     layer1_out[9357] <= layer0_out[958] & layer0_out[959];
     layer1_out[9358] <= ~(layer0_out[8495] | layer0_out[8496]);
     layer1_out[9359] <= layer0_out[9921] & ~layer0_out[9922];
     layer1_out[9360] <= ~(layer0_out[2273] & layer0_out[2274]);
     layer1_out[9361] <= layer0_out[11689] & ~layer0_out[11688];
     layer1_out[9362] <= ~layer0_out[10813];
     layer1_out[9363] <= layer0_out[9512];
     layer1_out[9364] <= ~(layer0_out[2057] & layer0_out[2058]);
     layer1_out[9365] <= layer0_out[8429] | layer0_out[8430];
     layer1_out[9366] <= ~layer0_out[3771] | layer0_out[3772];
     layer1_out[9367] <= ~layer0_out[1614] | layer0_out[1615];
     layer1_out[9368] <= ~(layer0_out[9526] & layer0_out[9527]);
     layer1_out[9369] <= layer0_out[6699];
     layer1_out[9370] <= layer0_out[5046] | layer0_out[5047];
     layer1_out[9371] <= ~(layer0_out[11554] | layer0_out[11555]);
     layer1_out[9372] <= layer0_out[10815] ^ layer0_out[10816];
     layer1_out[9373] <= layer0_out[7984] & layer0_out[7985];
     layer1_out[9374] <= ~layer0_out[128];
     layer1_out[9375] <= layer0_out[8644];
     layer1_out[9376] <= layer0_out[1856] & layer0_out[1857];
     layer1_out[9377] <= ~layer0_out[5877];
     layer1_out[9378] <= ~layer0_out[7456];
     layer1_out[9379] <= layer0_out[8628];
     layer1_out[9380] <= ~layer0_out[882] | layer0_out[883];
     layer1_out[9381] <= layer0_out[7362] | layer0_out[7363];
     layer1_out[9382] <= ~layer0_out[10571];
     layer1_out[9383] <= layer0_out[11318] & layer0_out[11319];
     layer1_out[9384] <= layer0_out[1469] & ~layer0_out[1470];
     layer1_out[9385] <= ~layer0_out[1299] | layer0_out[1298];
     layer1_out[9386] <= ~layer0_out[7950];
     layer1_out[9387] <= ~layer0_out[10804] | layer0_out[10803];
     layer1_out[9388] <= ~layer0_out[8674];
     layer1_out[9389] <= ~(layer0_out[8598] & layer0_out[8599]);
     layer1_out[9390] <= ~layer0_out[3600] | layer0_out[3601];
     layer1_out[9391] <= ~layer0_out[11906] | layer0_out[11907];
     layer1_out[9392] <= ~layer0_out[1680];
     layer1_out[9393] <= layer0_out[11129];
     layer1_out[9394] <= layer0_out[5954];
     layer1_out[9395] <= layer0_out[452];
     layer1_out[9396] <= ~layer0_out[2261] | layer0_out[2260];
     layer1_out[9397] <= layer0_out[9079];
     layer1_out[9398] <= ~layer0_out[5043] | layer0_out[5042];
     layer1_out[9399] <= layer0_out[7988];
     layer1_out[9400] <= layer0_out[3045] | layer0_out[3046];
     layer1_out[9401] <= layer0_out[3344] & ~layer0_out[3345];
     layer1_out[9402] <= layer0_out[4774] & ~layer0_out[4773];
     layer1_out[9403] <= ~(layer0_out[8624] & layer0_out[8625]);
     layer1_out[9404] <= ~(layer0_out[11879] | layer0_out[11880]);
     layer1_out[9405] <= ~layer0_out[2454];
     layer1_out[9406] <= layer0_out[7683];
     layer1_out[9407] <= ~(layer0_out[2185] | layer0_out[2186]);
     layer1_out[9408] <= layer0_out[8038];
     layer1_out[9409] <= ~layer0_out[5902] | layer0_out[5903];
     layer1_out[9410] <= layer0_out[1344];
     layer1_out[9411] <= ~(layer0_out[10808] ^ layer0_out[10809]);
     layer1_out[9412] <= ~(layer0_out[1235] ^ layer0_out[1236]);
     layer1_out[9413] <= ~(layer0_out[5128] & layer0_out[5129]);
     layer1_out[9414] <= ~(layer0_out[2700] | layer0_out[2701]);
     layer1_out[9415] <= layer0_out[8476] ^ layer0_out[8477];
     layer1_out[9416] <= ~layer0_out[6740];
     layer1_out[9417] <= layer0_out[8555];
     layer1_out[9418] <= layer0_out[5209];
     layer1_out[9419] <= ~layer0_out[2361];
     layer1_out[9420] <= ~layer0_out[3347];
     layer1_out[9421] <= 1'b1;
     layer1_out[9422] <= ~layer0_out[3466];
     layer1_out[9423] <= ~layer0_out[9676] | layer0_out[9677];
     layer1_out[9424] <= layer0_out[7465] ^ layer0_out[7466];
     layer1_out[9425] <= ~(layer0_out[10418] | layer0_out[10419]);
     layer1_out[9426] <= ~layer0_out[1041] | layer0_out[1040];
     layer1_out[9427] <= layer0_out[6223] ^ layer0_out[6224];
     layer1_out[9428] <= layer0_out[9242] & layer0_out[9243];
     layer1_out[9429] <= layer0_out[1456];
     layer1_out[9430] <= ~layer0_out[7894];
     layer1_out[9431] <= layer0_out[5502] & ~layer0_out[5501];
     layer1_out[9432] <= layer0_out[113] & ~layer0_out[114];
     layer1_out[9433] <= layer0_out[7112] | layer0_out[7113];
     layer1_out[9434] <= ~(layer0_out[8740] ^ layer0_out[8741]);
     layer1_out[9435] <= ~layer0_out[1030];
     layer1_out[9436] <= layer0_out[6823];
     layer1_out[9437] <= ~(layer0_out[4720] & layer0_out[4721]);
     layer1_out[9438] <= ~layer0_out[11512] | layer0_out[11511];
     layer1_out[9439] <= layer0_out[2325] & layer0_out[2326];
     layer1_out[9440] <= ~layer0_out[9143] | layer0_out[9144];
     layer1_out[9441] <= layer0_out[10677] ^ layer0_out[10678];
     layer1_out[9442] <= layer0_out[460] & ~layer0_out[459];
     layer1_out[9443] <= layer0_out[9605] ^ layer0_out[9606];
     layer1_out[9444] <= 1'b0;
     layer1_out[9445] <= layer0_out[2470];
     layer1_out[9446] <= layer0_out[464];
     layer1_out[9447] <= layer0_out[6015] | layer0_out[6016];
     layer1_out[9448] <= ~(layer0_out[9749] ^ layer0_out[9750]);
     layer1_out[9449] <= layer0_out[6041] & layer0_out[6042];
     layer1_out[9450] <= ~(layer0_out[1063] | layer0_out[1064]);
     layer1_out[9451] <= layer0_out[9119];
     layer1_out[9452] <= ~layer0_out[4804];
     layer1_out[9453] <= ~layer0_out[8950];
     layer1_out[9454] <= ~(layer0_out[632] | layer0_out[633]);
     layer1_out[9455] <= layer0_out[9656] ^ layer0_out[9657];
     layer1_out[9456] <= layer0_out[8982];
     layer1_out[9457] <= layer0_out[5320] | layer0_out[5321];
     layer1_out[9458] <= ~layer0_out[7147];
     layer1_out[9459] <= layer0_out[4950];
     layer1_out[9460] <= layer0_out[8707] & layer0_out[8708];
     layer1_out[9461] <= layer0_out[7135];
     layer1_out[9462] <= ~layer0_out[3776] | layer0_out[3777];
     layer1_out[9463] <= ~layer0_out[31];
     layer1_out[9464] <= ~(layer0_out[10573] & layer0_out[10574]);
     layer1_out[9465] <= ~layer0_out[2262];
     layer1_out[9466] <= ~layer0_out[6031];
     layer1_out[9467] <= ~layer0_out[245];
     layer1_out[9468] <= layer0_out[3051];
     layer1_out[9469] <= layer0_out[3147] & layer0_out[3148];
     layer1_out[9470] <= layer0_out[6442];
     layer1_out[9471] <= ~(layer0_out[1244] & layer0_out[1245]);
     layer1_out[9472] <= layer0_out[4156] | layer0_out[4157];
     layer1_out[9473] <= ~layer0_out[4790];
     layer1_out[9474] <= layer0_out[3761];
     layer1_out[9475] <= layer0_out[8069] & layer0_out[8070];
     layer1_out[9476] <= layer0_out[3626];
     layer1_out[9477] <= ~layer0_out[5144] | layer0_out[5143];
     layer1_out[9478] <= layer0_out[1795];
     layer1_out[9479] <= 1'b1;
     layer1_out[9480] <= layer0_out[5378];
     layer1_out[9481] <= ~layer0_out[3693] | layer0_out[3694];
     layer1_out[9482] <= 1'b1;
     layer1_out[9483] <= layer0_out[11346] ^ layer0_out[11347];
     layer1_out[9484] <= layer0_out[9140] & ~layer0_out[9141];
     layer1_out[9485] <= ~layer0_out[4640] | layer0_out[4641];
     layer1_out[9486] <= ~(layer0_out[6256] & layer0_out[6257]);
     layer1_out[9487] <= layer0_out[472] & ~layer0_out[473];
     layer1_out[9488] <= 1'b0;
     layer1_out[9489] <= ~layer0_out[8954] | layer0_out[8953];
     layer1_out[9490] <= ~layer0_out[6716];
     layer1_out[9491] <= 1'b1;
     layer1_out[9492] <= 1'b0;
     layer1_out[9493] <= layer0_out[6535];
     layer1_out[9494] <= layer0_out[2989] & ~layer0_out[2990];
     layer1_out[9495] <= layer0_out[2640] ^ layer0_out[2641];
     layer1_out[9496] <= layer0_out[3486] & layer0_out[3487];
     layer1_out[9497] <= layer0_out[2247] & ~layer0_out[2248];
     layer1_out[9498] <= ~layer0_out[8501];
     layer1_out[9499] <= ~layer0_out[5794] | layer0_out[5795];
     layer1_out[9500] <= layer0_out[1765] | layer0_out[1766];
     layer1_out[9501] <= 1'b1;
     layer1_out[9502] <= layer0_out[8994] & ~layer0_out[8995];
     layer1_out[9503] <= ~(layer0_out[4617] & layer0_out[4618]);
     layer1_out[9504] <= layer0_out[8997] & layer0_out[8998];
     layer1_out[9505] <= ~layer0_out[11651] | layer0_out[11652];
     layer1_out[9506] <= layer0_out[1253] & ~layer0_out[1254];
     layer1_out[9507] <= ~(layer0_out[5430] & layer0_out[5431]);
     layer1_out[9508] <= ~(layer0_out[4225] & layer0_out[4226]);
     layer1_out[9509] <= ~(layer0_out[5122] & layer0_out[5123]);
     layer1_out[9510] <= ~(layer0_out[5182] ^ layer0_out[5183]);
     layer1_out[9511] <= ~layer0_out[11169];
     layer1_out[9512] <= layer0_out[5810];
     layer1_out[9513] <= layer0_out[4777] & ~layer0_out[4778];
     layer1_out[9514] <= ~(layer0_out[10384] & layer0_out[10385]);
     layer1_out[9515] <= ~layer0_out[5404] | layer0_out[5405];
     layer1_out[9516] <= layer0_out[5100];
     layer1_out[9517] <= ~layer0_out[7053];
     layer1_out[9518] <= ~layer0_out[6705];
     layer1_out[9519] <= ~layer0_out[9192] | layer0_out[9193];
     layer1_out[9520] <= layer0_out[7615] | layer0_out[7616];
     layer1_out[9521] <= layer0_out[7229];
     layer1_out[9522] <= layer0_out[8005];
     layer1_out[9523] <= ~layer0_out[6092];
     layer1_out[9524] <= ~layer0_out[8143] | layer0_out[8142];
     layer1_out[9525] <= layer0_out[469];
     layer1_out[9526] <= layer0_out[599] & layer0_out[600];
     layer1_out[9527] <= layer0_out[6076] ^ layer0_out[6077];
     layer1_out[9528] <= ~(layer0_out[9529] & layer0_out[9530]);
     layer1_out[9529] <= ~layer0_out[6651] | layer0_out[6650];
     layer1_out[9530] <= layer0_out[5373];
     layer1_out[9531] <= ~(layer0_out[3103] | layer0_out[3104]);
     layer1_out[9532] <= ~layer0_out[8218];
     layer1_out[9533] <= ~layer0_out[5638] | layer0_out[5637];
     layer1_out[9534] <= layer0_out[9831];
     layer1_out[9535] <= layer0_out[4276];
     layer1_out[9536] <= layer0_out[4831] & ~layer0_out[4832];
     layer1_out[9537] <= ~layer0_out[8079];
     layer1_out[9538] <= layer0_out[1293];
     layer1_out[9539] <= ~layer0_out[388];
     layer1_out[9540] <= layer0_out[8386] & ~layer0_out[8385];
     layer1_out[9541] <= ~layer0_out[7994] | layer0_out[7993];
     layer1_out[9542] <= layer0_out[2916] | layer0_out[2917];
     layer1_out[9543] <= ~(layer0_out[10923] & layer0_out[10924]);
     layer1_out[9544] <= layer0_out[11253] & ~layer0_out[11252];
     layer1_out[9545] <= layer0_out[2095] ^ layer0_out[2096];
     layer1_out[9546] <= layer0_out[1409] & ~layer0_out[1408];
     layer1_out[9547] <= ~(layer0_out[3338] & layer0_out[3339]);
     layer1_out[9548] <= ~(layer0_out[3728] & layer0_out[3729]);
     layer1_out[9549] <= layer0_out[4308];
     layer1_out[9550] <= layer0_out[7296] & layer0_out[7297];
     layer1_out[9551] <= layer0_out[3056] & ~layer0_out[3057];
     layer1_out[9552] <= 1'b1;
     layer1_out[9553] <= layer0_out[6029];
     layer1_out[9554] <= ~layer0_out[7498] | layer0_out[7499];
     layer1_out[9555] <= ~layer0_out[5115];
     layer1_out[9556] <= layer0_out[685];
     layer1_out[9557] <= ~layer0_out[1882];
     layer1_out[9558] <= ~(layer0_out[4068] & layer0_out[4069]);
     layer1_out[9559] <= 1'b1;
     layer1_out[9560] <= ~layer0_out[9131] | layer0_out[9130];
     layer1_out[9561] <= layer0_out[5592];
     layer1_out[9562] <= layer0_out[7920];
     layer1_out[9563] <= layer0_out[5957] | layer0_out[5958];
     layer1_out[9564] <= layer0_out[4676];
     layer1_out[9565] <= layer0_out[5345] & ~layer0_out[5346];
     layer1_out[9566] <= ~layer0_out[2914] | layer0_out[2915];
     layer1_out[9567] <= layer0_out[5070] & layer0_out[5071];
     layer1_out[9568] <= layer0_out[7915];
     layer1_out[9569] <= ~(layer0_out[7010] ^ layer0_out[7011]);
     layer1_out[9570] <= ~layer0_out[11256];
     layer1_out[9571] <= layer0_out[7408] | layer0_out[7409];
     layer1_out[9572] <= ~layer0_out[4935];
     layer1_out[9573] <= 1'b1;
     layer1_out[9574] <= 1'b0;
     layer1_out[9575] <= ~layer0_out[4759];
     layer1_out[9576] <= ~layer0_out[3331];
     layer1_out[9577] <= ~(layer0_out[5648] & layer0_out[5649]);
     layer1_out[9578] <= layer0_out[4839] & ~layer0_out[4838];
     layer1_out[9579] <= ~(layer0_out[1434] ^ layer0_out[1435]);
     layer1_out[9580] <= ~(layer0_out[4435] & layer0_out[4436]);
     layer1_out[9581] <= layer0_out[5465] & layer0_out[5466];
     layer1_out[9582] <= layer0_out[3101] ^ layer0_out[3102];
     layer1_out[9583] <= layer0_out[6286];
     layer1_out[9584] <= layer0_out[4436] & layer0_out[4437];
     layer1_out[9585] <= ~(layer0_out[8279] | layer0_out[8280]);
     layer1_out[9586] <= layer0_out[10116];
     layer1_out[9587] <= layer0_out[9106] & ~layer0_out[9105];
     layer1_out[9588] <= layer0_out[4801];
     layer1_out[9589] <= layer0_out[8016] | layer0_out[8017];
     layer1_out[9590] <= ~layer0_out[909];
     layer1_out[9591] <= layer0_out[10785];
     layer1_out[9592] <= ~layer0_out[1759];
     layer1_out[9593] <= layer0_out[6307] & ~layer0_out[6306];
     layer1_out[9594] <= ~layer0_out[1144];
     layer1_out[9595] <= ~layer0_out[2796] | layer0_out[2797];
     layer1_out[9596] <= layer0_out[896] & layer0_out[897];
     layer1_out[9597] <= ~layer0_out[10699];
     layer1_out[9598] <= layer0_out[3665];
     layer1_out[9599] <= ~layer0_out[5793] | layer0_out[5794];
     layer1_out[9600] <= layer0_out[3330] | layer0_out[3331];
     layer1_out[9601] <= layer0_out[7357] & layer0_out[7358];
     layer1_out[9602] <= ~layer0_out[640];
     layer1_out[9603] <= ~layer0_out[11934] | layer0_out[11935];
     layer1_out[9604] <= ~layer0_out[6516];
     layer1_out[9605] <= ~layer0_out[9890] | layer0_out[9889];
     layer1_out[9606] <= layer0_out[6188];
     layer1_out[9607] <= layer0_out[7816] & layer0_out[7817];
     layer1_out[9608] <= layer0_out[9403];
     layer1_out[9609] <= ~layer0_out[10875];
     layer1_out[9610] <= layer0_out[5248];
     layer1_out[9611] <= ~layer0_out[11910];
     layer1_out[9612] <= layer0_out[8532];
     layer1_out[9613] <= layer0_out[4994] & layer0_out[4995];
     layer1_out[9614] <= layer0_out[11110] | layer0_out[11111];
     layer1_out[9615] <= layer0_out[7246];
     layer1_out[9616] <= layer0_out[8785] | layer0_out[8786];
     layer1_out[9617] <= layer0_out[3850] & ~layer0_out[3849];
     layer1_out[9618] <= layer0_out[8323] & layer0_out[8324];
     layer1_out[9619] <= ~layer0_out[6126];
     layer1_out[9620] <= layer0_out[1942] & ~layer0_out[1941];
     layer1_out[9621] <= layer0_out[3107] & layer0_out[3108];
     layer1_out[9622] <= layer0_out[7663];
     layer1_out[9623] <= layer0_out[8032];
     layer1_out[9624] <= ~layer0_out[11000] | layer0_out[11001];
     layer1_out[9625] <= ~layer0_out[783];
     layer1_out[9626] <= layer0_out[4208] | layer0_out[4209];
     layer1_out[9627] <= layer0_out[3724] & ~layer0_out[3725];
     layer1_out[9628] <= ~layer0_out[7879];
     layer1_out[9629] <= ~layer0_out[7044] | layer0_out[7043];
     layer1_out[9630] <= layer0_out[5960];
     layer1_out[9631] <= layer0_out[768];
     layer1_out[9632] <= layer0_out[500];
     layer1_out[9633] <= ~(layer0_out[3396] & layer0_out[3397]);
     layer1_out[9634] <= layer0_out[3802];
     layer1_out[9635] <= ~layer0_out[9439];
     layer1_out[9636] <= layer0_out[9876] & ~layer0_out[9877];
     layer1_out[9637] <= layer0_out[7517] & layer0_out[7518];
     layer1_out[9638] <= 1'b0;
     layer1_out[9639] <= ~layer0_out[10780] | layer0_out[10781];
     layer1_out[9640] <= layer0_out[6762];
     layer1_out[9641] <= layer0_out[3845] | layer0_out[3846];
     layer1_out[9642] <= ~layer0_out[11156];
     layer1_out[9643] <= layer0_out[11903] & ~layer0_out[11904];
     layer1_out[9644] <= ~layer0_out[5098];
     layer1_out[9645] <= ~(layer0_out[1761] & layer0_out[1762]);
     layer1_out[9646] <= layer0_out[1700] & ~layer0_out[1699];
     layer1_out[9647] <= layer0_out[11585];
     layer1_out[9648] <= layer0_out[325] & ~layer0_out[326];
     layer1_out[9649] <= ~layer0_out[3917] | layer0_out[3916];
     layer1_out[9650] <= ~layer0_out[10996];
     layer1_out[9651] <= layer0_out[3165];
     layer1_out[9652] <= layer0_out[7487] | layer0_out[7488];
     layer1_out[9653] <= ~(layer0_out[1077] | layer0_out[1078]);
     layer1_out[9654] <= ~(layer0_out[5421] & layer0_out[5422]);
     layer1_out[9655] <= ~(layer0_out[9694] & layer0_out[9695]);
     layer1_out[9656] <= ~(layer0_out[6098] | layer0_out[6099]);
     layer1_out[9657] <= ~layer0_out[4301] | layer0_out[4300];
     layer1_out[9658] <= ~(layer0_out[2685] ^ layer0_out[2686]);
     layer1_out[9659] <= layer0_out[2061] | layer0_out[2062];
     layer1_out[9660] <= ~layer0_out[4959];
     layer1_out[9661] <= ~layer0_out[9093];
     layer1_out[9662] <= layer0_out[1123] | layer0_out[1124];
     layer1_out[9663] <= ~layer0_out[2525] | layer0_out[2526];
     layer1_out[9664] <= ~layer0_out[6815];
     layer1_out[9665] <= ~layer0_out[380];
     layer1_out[9666] <= layer0_out[3299] & ~layer0_out[3300];
     layer1_out[9667] <= ~(layer0_out[10379] | layer0_out[10380]);
     layer1_out[9668] <= layer0_out[3386] & layer0_out[3387];
     layer1_out[9669] <= ~(layer0_out[1345] | layer0_out[1346]);
     layer1_out[9670] <= ~(layer0_out[4769] | layer0_out[4770]);
     layer1_out[9671] <= layer0_out[9123] & ~layer0_out[9124];
     layer1_out[9672] <= layer0_out[10709] | layer0_out[10710];
     layer1_out[9673] <= ~layer0_out[9705];
     layer1_out[9674] <= layer0_out[10028];
     layer1_out[9675] <= layer0_out[11048];
     layer1_out[9676] <= layer0_out[2688] & ~layer0_out[2687];
     layer1_out[9677] <= ~layer0_out[11469];
     layer1_out[9678] <= layer0_out[5362];
     layer1_out[9679] <= ~layer0_out[5293];
     layer1_out[9680] <= ~layer0_out[10613];
     layer1_out[9681] <= layer0_out[11748];
     layer1_out[9682] <= ~layer0_out[11986];
     layer1_out[9683] <= ~layer0_out[1734];
     layer1_out[9684] <= layer0_out[664] & ~layer0_out[663];
     layer1_out[9685] <= layer0_out[8053] & ~layer0_out[8052];
     layer1_out[9686] <= layer0_out[334] & layer0_out[335];
     layer1_out[9687] <= ~layer0_out[6145] | layer0_out[6144];
     layer1_out[9688] <= layer0_out[11528];
     layer1_out[9689] <= layer0_out[6209] ^ layer0_out[6210];
     layer1_out[9690] <= ~layer0_out[4040] | layer0_out[4041];
     layer1_out[9691] <= ~(layer0_out[4693] ^ layer0_out[4694]);
     layer1_out[9692] <= 1'b0;
     layer1_out[9693] <= layer0_out[10155];
     layer1_out[9694] <= layer0_out[9440] | layer0_out[9441];
     layer1_out[9695] <= ~layer0_out[4762];
     layer1_out[9696] <= layer0_out[8503];
     layer1_out[9697] <= layer0_out[4203];
     layer1_out[9698] <= ~layer0_out[8710];
     layer1_out[9699] <= layer0_out[7826];
     layer1_out[9700] <= layer0_out[2560] & ~layer0_out[2559];
     layer1_out[9701] <= ~(layer0_out[1964] & layer0_out[1965]);
     layer1_out[9702] <= layer0_out[2933] | layer0_out[2934];
     layer1_out[9703] <= ~layer0_out[10118] | layer0_out[10117];
     layer1_out[9704] <= ~layer0_out[7183];
     layer1_out[9705] <= ~(layer0_out[2720] & layer0_out[2721]);
     layer1_out[9706] <= ~layer0_out[2995];
     layer1_out[9707] <= layer0_out[3672];
     layer1_out[9708] <= ~layer0_out[8643];
     layer1_out[9709] <= ~(layer0_out[6648] & layer0_out[6649]);
     layer1_out[9710] <= layer0_out[963] & ~layer0_out[964];
     layer1_out[9711] <= layer0_out[4409];
     layer1_out[9712] <= ~layer0_out[2494];
     layer1_out[9713] <= 1'b1;
     layer1_out[9714] <= layer0_out[3197] & ~layer0_out[3198];
     layer1_out[9715] <= layer0_out[4700] & ~layer0_out[4701];
     layer1_out[9716] <= ~layer0_out[9201];
     layer1_out[9717] <= layer0_out[10687] & ~layer0_out[10688];
     layer1_out[9718] <= layer0_out[7506];
     layer1_out[9719] <= layer0_out[9263] & ~layer0_out[9262];
     layer1_out[9720] <= ~(layer0_out[579] & layer0_out[580]);
     layer1_out[9721] <= ~layer0_out[3586];
     layer1_out[9722] <= layer0_out[6495] & ~layer0_out[6494];
     layer1_out[9723] <= ~layer0_out[8253];
     layer1_out[9724] <= ~layer0_out[4701];
     layer1_out[9725] <= 1'b0;
     layer1_out[9726] <= layer0_out[555] | layer0_out[556];
     layer1_out[9727] <= layer0_out[6855] & ~layer0_out[6854];
     layer1_out[9728] <= ~(layer0_out[6882] ^ layer0_out[6883]);
     layer1_out[9729] <= ~layer0_out[7327];
     layer1_out[9730] <= layer0_out[10099] & ~layer0_out[10100];
     layer1_out[9731] <= ~layer0_out[9466];
     layer1_out[9732] <= layer0_out[531] | layer0_out[532];
     layer1_out[9733] <= ~(layer0_out[9027] | layer0_out[9028]);
     layer1_out[9734] <= ~layer0_out[1350] | layer0_out[1349];
     layer1_out[9735] <= layer0_out[8340] & ~layer0_out[8341];
     layer1_out[9736] <= ~layer0_out[6771];
     layer1_out[9737] <= layer0_out[7642] & layer0_out[7643];
     layer1_out[9738] <= ~(layer0_out[3002] ^ layer0_out[3003]);
     layer1_out[9739] <= ~(layer0_out[5964] ^ layer0_out[5965]);
     layer1_out[9740] <= layer0_out[9543] & ~layer0_out[9544];
     layer1_out[9741] <= layer0_out[5351];
     layer1_out[9742] <= layer0_out[7495] | layer0_out[7496];
     layer1_out[9743] <= layer0_out[8378] | layer0_out[8379];
     layer1_out[9744] <= ~(layer0_out[4017] & layer0_out[4018]);
     layer1_out[9745] <= layer0_out[3866] | layer0_out[3867];
     layer1_out[9746] <= layer0_out[8861] ^ layer0_out[8862];
     layer1_out[9747] <= ~layer0_out[6080];
     layer1_out[9748] <= layer0_out[1848] & ~layer0_out[1847];
     layer1_out[9749] <= layer0_out[3617];
     layer1_out[9750] <= ~layer0_out[1177];
     layer1_out[9751] <= layer0_out[4373];
     layer1_out[9752] <= layer0_out[4500] & ~layer0_out[4499];
     layer1_out[9753] <= ~layer0_out[2849] | layer0_out[2850];
     layer1_out[9754] <= layer0_out[995];
     layer1_out[9755] <= ~layer0_out[9205];
     layer1_out[9756] <= ~layer0_out[1073] | layer0_out[1072];
     layer1_out[9757] <= layer0_out[5629];
     layer1_out[9758] <= layer0_out[8742] & ~layer0_out[8743];
     layer1_out[9759] <= layer0_out[6678] & ~layer0_out[6677];
     layer1_out[9760] <= ~layer0_out[5690];
     layer1_out[9761] <= ~(layer0_out[666] | layer0_out[667]);
     layer1_out[9762] <= ~(layer0_out[5131] & layer0_out[5132]);
     layer1_out[9763] <= ~layer0_out[577] | layer0_out[576];
     layer1_out[9764] <= layer0_out[7250] | layer0_out[7251];
     layer1_out[9765] <= ~(layer0_out[6474] & layer0_out[6475]);
     layer1_out[9766] <= layer0_out[7895];
     layer1_out[9767] <= layer0_out[6893];
     layer1_out[9768] <= layer0_out[5992];
     layer1_out[9769] <= layer0_out[9900];
     layer1_out[9770] <= ~layer0_out[840] | layer0_out[841];
     layer1_out[9771] <= ~(layer0_out[7505] & layer0_out[7506]);
     layer1_out[9772] <= layer0_out[9504] | layer0_out[9505];
     layer1_out[9773] <= ~layer0_out[2120] | layer0_out[2121];
     layer1_out[9774] <= layer0_out[8522];
     layer1_out[9775] <= layer0_out[6332] | layer0_out[6333];
     layer1_out[9776] <= layer0_out[3047];
     layer1_out[9777] <= layer0_out[10497] | layer0_out[10498];
     layer1_out[9778] <= ~layer0_out[4542] | layer0_out[4543];
     layer1_out[9779] <= layer0_out[2150];
     layer1_out[9780] <= ~layer0_out[2704];
     layer1_out[9781] <= layer0_out[6666];
     layer1_out[9782] <= layer0_out[1787] & layer0_out[1788];
     layer1_out[9783] <= ~layer0_out[9207];
     layer1_out[9784] <= layer0_out[6715];
     layer1_out[9785] <= layer0_out[10535] | layer0_out[10536];
     layer1_out[9786] <= layer0_out[1252] & ~layer0_out[1251];
     layer1_out[9787] <= ~layer0_out[6452] | layer0_out[6453];
     layer1_out[9788] <= layer0_out[7858] | layer0_out[7859];
     layer1_out[9789] <= layer0_out[5621];
     layer1_out[9790] <= layer0_out[7069];
     layer1_out[9791] <= ~(layer0_out[4414] | layer0_out[4415]);
     layer1_out[9792] <= layer0_out[488] & ~layer0_out[487];
     layer1_out[9793] <= ~(layer0_out[5282] & layer0_out[5283]);
     layer1_out[9794] <= ~(layer0_out[10562] ^ layer0_out[10563]);
     layer1_out[9795] <= layer0_out[2323] & ~layer0_out[2324];
     layer1_out[9796] <= ~(layer0_out[10005] & layer0_out[10006]);
     layer1_out[9797] <= ~(layer0_out[10300] | layer0_out[10301]);
     layer1_out[9798] <= ~layer0_out[11563] | layer0_out[11562];
     layer1_out[9799] <= ~layer0_out[1772];
     layer1_out[9800] <= ~layer0_out[6155];
     layer1_out[9801] <= layer0_out[9026];
     layer1_out[9802] <= layer0_out[10905];
     layer1_out[9803] <= layer0_out[8726] & ~layer0_out[8725];
     layer1_out[9804] <= ~(layer0_out[10719] & layer0_out[10720]);
     layer1_out[9805] <= layer0_out[3409] & ~layer0_out[3408];
     layer1_out[9806] <= layer0_out[2349] | layer0_out[2350];
     layer1_out[9807] <= ~(layer0_out[6056] ^ layer0_out[6057]);
     layer1_out[9808] <= layer0_out[5487] & layer0_out[5488];
     layer1_out[9809] <= ~(layer0_out[1405] ^ layer0_out[1406]);
     layer1_out[9810] <= ~(layer0_out[6659] | layer0_out[6660]);
     layer1_out[9811] <= 1'b1;
     layer1_out[9812] <= layer0_out[11479];
     layer1_out[9813] <= layer0_out[10387] & ~layer0_out[10388];
     layer1_out[9814] <= layer0_out[8155];
     layer1_out[9815] <= layer0_out[11060] & ~layer0_out[11061];
     layer1_out[9816] <= ~layer0_out[6246];
     layer1_out[9817] <= layer0_out[11831] | layer0_out[11832];
     layer1_out[9818] <= ~(layer0_out[8143] ^ layer0_out[8144]);
     layer1_out[9819] <= layer0_out[2814];
     layer1_out[9820] <= ~(layer0_out[3709] & layer0_out[3710]);
     layer1_out[9821] <= layer0_out[2130];
     layer1_out[9822] <= ~(layer0_out[6934] ^ layer0_out[6935]);
     layer1_out[9823] <= ~(layer0_out[9936] | layer0_out[9937]);
     layer1_out[9824] <= layer0_out[9410] & layer0_out[9411];
     layer1_out[9825] <= layer0_out[3322] & ~layer0_out[3321];
     layer1_out[9826] <= ~(layer0_out[6574] & layer0_out[6575]);
     layer1_out[9827] <= layer0_out[8182] & ~layer0_out[8181];
     layer1_out[9828] <= ~(layer0_out[4694] & layer0_out[4695]);
     layer1_out[9829] <= ~(layer0_out[10978] | layer0_out[10979]);
     layer1_out[9830] <= layer0_out[1896];
     layer1_out[9831] <= layer0_out[876];
     layer1_out[9832] <= layer0_out[8874];
     layer1_out[9833] <= ~layer0_out[7384];
     layer1_out[9834] <= 1'b0;
     layer1_out[9835] <= layer0_out[5179] & ~layer0_out[5180];
     layer1_out[9836] <= ~layer0_out[8259];
     layer1_out[9837] <= ~(layer0_out[1323] & layer0_out[1324]);
     layer1_out[9838] <= ~(layer0_out[5422] & layer0_out[5423]);
     layer1_out[9839] <= ~(layer0_out[7880] | layer0_out[7881]);
     layer1_out[9840] <= 1'b1;
     layer1_out[9841] <= layer0_out[4799] & ~layer0_out[4800];
     layer1_out[9842] <= layer0_out[1057];
     layer1_out[9843] <= 1'b0;
     layer1_out[9844] <= layer0_out[3169];
     layer1_out[9845] <= ~layer0_out[998];
     layer1_out[9846] <= ~layer0_out[5796];
     layer1_out[9847] <= layer0_out[11028] | layer0_out[11029];
     layer1_out[9848] <= ~layer0_out[10376];
     layer1_out[9849] <= layer0_out[1785] ^ layer0_out[1786];
     layer1_out[9850] <= 1'b1;
     layer1_out[9851] <= layer0_out[8810];
     layer1_out[9852] <= ~layer0_out[11401];
     layer1_out[9853] <= layer0_out[5930];
     layer1_out[9854] <= ~(layer0_out[1973] | layer0_out[1974]);
     layer1_out[9855] <= ~layer0_out[3292] | layer0_out[3293];
     layer1_out[9856] <= layer0_out[8899] & ~layer0_out[8900];
     layer1_out[9857] <= layer0_out[4200] & ~layer0_out[4201];
     layer1_out[9858] <= layer0_out[8791] & ~layer0_out[8792];
     layer1_out[9859] <= ~(layer0_out[305] | layer0_out[306]);
     layer1_out[9860] <= layer0_out[3132] & ~layer0_out[3133];
     layer1_out[9861] <= layer0_out[8472] | layer0_out[8473];
     layer1_out[9862] <= layer0_out[1772];
     layer1_out[9863] <= ~(layer0_out[5534] | layer0_out[5535]);
     layer1_out[9864] <= layer0_out[5527] & ~layer0_out[5528];
     layer1_out[9865] <= layer0_out[2075] & ~layer0_out[2076];
     layer1_out[9866] <= layer0_out[3269] & ~layer0_out[3270];
     layer1_out[9867] <= layer0_out[1992] & ~layer0_out[1993];
     layer1_out[9868] <= layer0_out[10655] & ~layer0_out[10654];
     layer1_out[9869] <= 1'b1;
     layer1_out[9870] <= ~layer0_out[10222];
     layer1_out[9871] <= layer0_out[10069];
     layer1_out[9872] <= layer0_out[9669] & ~layer0_out[9668];
     layer1_out[9873] <= layer0_out[9344];
     layer1_out[9874] <= layer0_out[11086];
     layer1_out[9875] <= 1'b1;
     layer1_out[9876] <= ~layer0_out[3603];
     layer1_out[9877] <= ~(layer0_out[4913] ^ layer0_out[4914]);
     layer1_out[9878] <= ~layer0_out[6830] | layer0_out[6831];
     layer1_out[9879] <= ~layer0_out[10734] | layer0_out[10735];
     layer1_out[9880] <= ~(layer0_out[8621] & layer0_out[8622]);
     layer1_out[9881] <= ~(layer0_out[8474] & layer0_out[8475]);
     layer1_out[9882] <= layer0_out[5813] | layer0_out[5814];
     layer1_out[9883] <= ~(layer0_out[11003] | layer0_out[11004]);
     layer1_out[9884] <= layer0_out[2117] ^ layer0_out[2118];
     layer1_out[9885] <= ~layer0_out[2504] | layer0_out[2505];
     layer1_out[9886] <= ~layer0_out[10212];
     layer1_out[9887] <= ~(layer0_out[7828] | layer0_out[7829]);
     layer1_out[9888] <= ~(layer0_out[6586] & layer0_out[6587]);
     layer1_out[9889] <= ~layer0_out[299];
     layer1_out[9890] <= ~layer0_out[2659];
     layer1_out[9891] <= ~layer0_out[11312] | layer0_out[11311];
     layer1_out[9892] <= layer0_out[6361] & layer0_out[6362];
     layer1_out[9893] <= ~layer0_out[9053] | layer0_out[9054];
     layer1_out[9894] <= ~layer0_out[3767];
     layer1_out[9895] <= ~layer0_out[5446] | layer0_out[5445];
     layer1_out[9896] <= layer0_out[11829] & ~layer0_out[11828];
     layer1_out[9897] <= ~layer0_out[8795];
     layer1_out[9898] <= ~layer0_out[2053] | layer0_out[2054];
     layer1_out[9899] <= layer0_out[70];
     layer1_out[9900] <= layer0_out[11125];
     layer1_out[9901] <= layer0_out[1768];
     layer1_out[9902] <= layer0_out[5137];
     layer1_out[9903] <= layer0_out[4578] ^ layer0_out[4579];
     layer1_out[9904] <= ~layer0_out[2113];
     layer1_out[9905] <= layer0_out[6068] & ~layer0_out[6069];
     layer1_out[9906] <= layer0_out[9869] | layer0_out[9870];
     layer1_out[9907] <= layer0_out[390] | layer0_out[391];
     layer1_out[9908] <= layer0_out[4601] & layer0_out[4602];
     layer1_out[9909] <= layer0_out[7703];
     layer1_out[9910] <= ~(layer0_out[2693] & layer0_out[2694]);
     layer1_out[9911] <= layer0_out[10187];
     layer1_out[9912] <= layer0_out[2041] | layer0_out[2042];
     layer1_out[9913] <= layer0_out[11120];
     layer1_out[9914] <= ~layer0_out[7785];
     layer1_out[9915] <= layer0_out[9638] | layer0_out[9639];
     layer1_out[9916] <= ~(layer0_out[3454] ^ layer0_out[3455]);
     layer1_out[9917] <= ~layer0_out[1120] | layer0_out[1121];
     layer1_out[9918] <= ~(layer0_out[6773] | layer0_out[6774]);
     layer1_out[9919] <= ~layer0_out[10441] | layer0_out[10442];
     layer1_out[9920] <= ~(layer0_out[4460] | layer0_out[4461]);
     layer1_out[9921] <= ~layer0_out[2848];
     layer1_out[9922] <= layer0_out[8067] & ~layer0_out[8066];
     layer1_out[9923] <= layer0_out[7564] ^ layer0_out[7565];
     layer1_out[9924] <= ~(layer0_out[7690] & layer0_out[7691]);
     layer1_out[9925] <= layer0_out[6890] & ~layer0_out[6891];
     layer1_out[9926] <= layer0_out[2245];
     layer1_out[9927] <= ~(layer0_out[6180] ^ layer0_out[6181]);
     layer1_out[9928] <= ~layer0_out[2790];
     layer1_out[9929] <= layer0_out[7712] ^ layer0_out[7713];
     layer1_out[9930] <= layer0_out[1216] | layer0_out[1217];
     layer1_out[9931] <= ~(layer0_out[4792] | layer0_out[4793]);
     layer1_out[9932] <= layer0_out[7239] ^ layer0_out[7240];
     layer1_out[9933] <= ~layer0_out[11763] | layer0_out[11764];
     layer1_out[9934] <= ~layer0_out[11075];
     layer1_out[9935] <= ~layer0_out[6594];
     layer1_out[9936] <= layer0_out[5747];
     layer1_out[9937] <= ~(layer0_out[6069] ^ layer0_out[6070]);
     layer1_out[9938] <= ~layer0_out[5496] | layer0_out[5497];
     layer1_out[9939] <= ~layer0_out[2241];
     layer1_out[9940] <= ~layer0_out[7730] | layer0_out[7731];
     layer1_out[9941] <= ~layer0_out[2624];
     layer1_out[9942] <= layer0_out[420];
     layer1_out[9943] <= layer0_out[294] & ~layer0_out[293];
     layer1_out[9944] <= ~layer0_out[3428];
     layer1_out[9945] <= ~layer0_out[716];
     layer1_out[9946] <= layer0_out[4859] | layer0_out[4860];
     layer1_out[9947] <= layer0_out[8671];
     layer1_out[9948] <= layer0_out[2666] & ~layer0_out[2667];
     layer1_out[9949] <= ~layer0_out[8665];
     layer1_out[9950] <= layer0_out[11053] & ~layer0_out[11052];
     layer1_out[9951] <= ~layer0_out[3431];
     layer1_out[9952] <= ~layer0_out[7555] | layer0_out[7556];
     layer1_out[9953] <= layer0_out[10674];
     layer1_out[9954] <= layer0_out[11557] & ~layer0_out[11558];
     layer1_out[9955] <= layer0_out[11925] & ~layer0_out[11924];
     layer1_out[9956] <= layer0_out[5986] & ~layer0_out[5985];
     layer1_out[9957] <= ~layer0_out[11103];
     layer1_out[9958] <= ~layer0_out[4048] | layer0_out[4049];
     layer1_out[9959] <= ~layer0_out[551];
     layer1_out[9960] <= ~layer0_out[6640] | layer0_out[6639];
     layer1_out[9961] <= layer0_out[1114];
     layer1_out[9962] <= ~layer0_out[5862];
     layer1_out[9963] <= layer0_out[8693];
     layer1_out[9964] <= layer0_out[7346] & ~layer0_out[7345];
     layer1_out[9965] <= ~layer0_out[3982];
     layer1_out[9966] <= layer0_out[952] | layer0_out[953];
     layer1_out[9967] <= ~layer0_out[4636];
     layer1_out[9968] <= layer0_out[9133] & ~layer0_out[9134];
     layer1_out[9969] <= ~layer0_out[1843] | layer0_out[1842];
     layer1_out[9970] <= ~layer0_out[9327];
     layer1_out[9971] <= layer0_out[7876] & ~layer0_out[7877];
     layer1_out[9972] <= ~layer0_out[6644];
     layer1_out[9973] <= ~layer0_out[11117];
     layer1_out[9974] <= layer0_out[6936] & ~layer0_out[6937];
     layer1_out[9975] <= layer0_out[6369] & ~layer0_out[6368];
     layer1_out[9976] <= layer0_out[11714] ^ layer0_out[11715];
     layer1_out[9977] <= 1'b1;
     layer1_out[9978] <= ~(layer0_out[8648] & layer0_out[8649]);
     layer1_out[9979] <= ~layer0_out[7577];
     layer1_out[9980] <= ~layer0_out[112];
     layer1_out[9981] <= ~layer0_out[4085] | layer0_out[4084];
     layer1_out[9982] <= layer0_out[11566] & ~layer0_out[11565];
     layer1_out[9983] <= layer0_out[3902] & ~layer0_out[3901];
     layer1_out[9984] <= layer0_out[2333];
     layer1_out[9985] <= layer0_out[7758] | layer0_out[7759];
     layer1_out[9986] <= ~layer0_out[2122] | layer0_out[2121];
     layer1_out[9987] <= layer0_out[3336];
     layer1_out[9988] <= layer0_out[9874] & ~layer0_out[9875];
     layer1_out[9989] <= ~(layer0_out[11762] | layer0_out[11763]);
     layer1_out[9990] <= ~layer0_out[5667];
     layer1_out[9991] <= layer0_out[4851];
     layer1_out[9992] <= ~layer0_out[7714] | layer0_out[7715];
     layer1_out[9993] <= ~(layer0_out[11829] ^ layer0_out[11830]);
     layer1_out[9994] <= ~layer0_out[8518] | layer0_out[8517];
     layer1_out[9995] <= layer0_out[595] & layer0_out[596];
     layer1_out[9996] <= layer0_out[1538] | layer0_out[1539];
     layer1_out[9997] <= ~layer0_out[5000];
     layer1_out[9998] <= ~layer0_out[9659] | layer0_out[9660];
     layer1_out[9999] <= ~layer0_out[1873] | layer0_out[1872];
     layer1_out[10000] <= layer0_out[11145] & ~layer0_out[11146];
     layer1_out[10001] <= layer0_out[9753] & ~layer0_out[9754];
     layer1_out[10002] <= layer0_out[8596] & layer0_out[8597];
     layer1_out[10003] <= ~layer0_out[6884];
     layer1_out[10004] <= layer0_out[2468] & layer0_out[2469];
     layer1_out[10005] <= ~layer0_out[5287] | layer0_out[5288];
     layer1_out[10006] <= layer0_out[5002];
     layer1_out[10007] <= 1'b1;
     layer1_out[10008] <= ~(layer0_out[7802] ^ layer0_out[7803]);
     layer1_out[10009] <= ~layer0_out[3179] | layer0_out[3180];
     layer1_out[10010] <= layer0_out[4044] & layer0_out[4045];
     layer1_out[10011] <= ~layer0_out[7140];
     layer1_out[10012] <= ~layer0_out[6573];
     layer1_out[10013] <= layer0_out[4107] & ~layer0_out[4106];
     layer1_out[10014] <= ~(layer0_out[9771] & layer0_out[9772]);
     layer1_out[10015] <= layer0_out[9790] & ~layer0_out[9791];
     layer1_out[10016] <= ~layer0_out[3039] | layer0_out[3038];
     layer1_out[10017] <= ~(layer0_out[7293] | layer0_out[7294]);
     layer1_out[10018] <= layer0_out[11458] & layer0_out[11459];
     layer1_out[10019] <= layer0_out[6425];
     layer1_out[10020] <= ~(layer0_out[1553] ^ layer0_out[1554]);
     layer1_out[10021] <= ~layer0_out[10298];
     layer1_out[10022] <= layer0_out[4753];
     layer1_out[10023] <= layer0_out[5944] & layer0_out[5945];
     layer1_out[10024] <= layer0_out[7995] & ~layer0_out[7996];
     layer1_out[10025] <= layer0_out[6841] | layer0_out[6842];
     layer1_out[10026] <= ~(layer0_out[7474] & layer0_out[7475]);
     layer1_out[10027] <= ~layer0_out[11057];
     layer1_out[10028] <= layer0_out[341];
     layer1_out[10029] <= ~(layer0_out[6011] ^ layer0_out[6012]);
     layer1_out[10030] <= ~layer0_out[10542] | layer0_out[10543];
     layer1_out[10031] <= layer0_out[10195];
     layer1_out[10032] <= layer0_out[8773];
     layer1_out[10033] <= layer0_out[11354] | layer0_out[11355];
     layer1_out[10034] <= ~(layer0_out[681] ^ layer0_out[682]);
     layer1_out[10035] <= layer0_out[10018] & ~layer0_out[10017];
     layer1_out[10036] <= ~(layer0_out[3878] ^ layer0_out[3879]);
     layer1_out[10037] <= ~layer0_out[10309] | layer0_out[10308];
     layer1_out[10038] <= layer0_out[5385] ^ layer0_out[5386];
     layer1_out[10039] <= layer0_out[8277] & ~layer0_out[8276];
     layer1_out[10040] <= 1'b1;
     layer1_out[10041] <= layer0_out[11499];
     layer1_out[10042] <= layer0_out[7098] | layer0_out[7099];
     layer1_out[10043] <= layer0_out[674];
     layer1_out[10044] <= ~layer0_out[3900] | layer0_out[3899];
     layer1_out[10045] <= layer0_out[1262] & layer0_out[1263];
     layer1_out[10046] <= layer0_out[9501] & layer0_out[9502];
     layer1_out[10047] <= ~(layer0_out[5074] | layer0_out[5075]);
     layer1_out[10048] <= ~(layer0_out[11935] & layer0_out[11936]);
     layer1_out[10049] <= layer0_out[1070];
     layer1_out[10050] <= ~layer0_out[4502];
     layer1_out[10051] <= ~layer0_out[10974];
     layer1_out[10052] <= ~layer0_out[11133] | layer0_out[11132];
     layer1_out[10053] <= ~layer0_out[2805] | layer0_out[2806];
     layer1_out[10054] <= ~layer0_out[7047] | layer0_out[7048];
     layer1_out[10055] <= ~layer0_out[2617];
     layer1_out[10056] <= layer0_out[11673];
     layer1_out[10057] <= ~(layer0_out[619] & layer0_out[620]);
     layer1_out[10058] <= layer0_out[9614];
     layer1_out[10059] <= ~layer0_out[4937];
     layer1_out[10060] <= ~layer0_out[346];
     layer1_out[10061] <= ~layer0_out[3297];
     layer1_out[10062] <= layer0_out[2761];
     layer1_out[10063] <= layer0_out[6937] | layer0_out[6938];
     layer1_out[10064] <= ~(layer0_out[11038] & layer0_out[11039]);
     layer1_out[10065] <= ~(layer0_out[1310] & layer0_out[1311]);
     layer1_out[10066] <= layer0_out[6212] ^ layer0_out[6213];
     layer1_out[10067] <= ~layer0_out[11497];
     layer1_out[10068] <= ~(layer0_out[3873] | layer0_out[3874]);
     layer1_out[10069] <= ~layer0_out[6370];
     layer1_out[10070] <= ~(layer0_out[11601] & layer0_out[11602]);
     layer1_out[10071] <= layer0_out[6150] & layer0_out[6151];
     layer1_out[10072] <= ~layer0_out[5602];
     layer1_out[10073] <= ~layer0_out[9765] | layer0_out[9764];
     layer1_out[10074] <= 1'b0;
     layer1_out[10075] <= ~(layer0_out[2002] & layer0_out[2003]);
     layer1_out[10076] <= ~layer0_out[7629] | layer0_out[7628];
     layer1_out[10077] <= layer0_out[5486];
     layer1_out[10078] <= ~layer0_out[6476];
     layer1_out[10079] <= ~(layer0_out[5274] & layer0_out[5275]);
     layer1_out[10080] <= layer0_out[9675] & layer0_out[9676];
     layer1_out[10081] <= ~layer0_out[7319] | layer0_out[7318];
     layer1_out[10082] <= ~layer0_out[7572];
     layer1_out[10083] <= ~layer0_out[9483];
     layer1_out[10084] <= layer0_out[4519];
     layer1_out[10085] <= layer0_out[6605] & layer0_out[6606];
     layer1_out[10086] <= ~layer0_out[1981] | layer0_out[1980];
     layer1_out[10087] <= ~layer0_out[3054] | layer0_out[3055];
     layer1_out[10088] <= ~layer0_out[8613] | layer0_out[8612];
     layer1_out[10089] <= ~layer0_out[3789];
     layer1_out[10090] <= ~layer0_out[10585];
     layer1_out[10091] <= layer0_out[7170];
     layer1_out[10092] <= layer0_out[11031] & layer0_out[11032];
     layer1_out[10093] <= layer0_out[1824] | layer0_out[1825];
     layer1_out[10094] <= 1'b0;
     layer1_out[10095] <= ~(layer0_out[11115] & layer0_out[11116]);
     layer1_out[10096] <= layer0_out[6720] & layer0_out[6721];
     layer1_out[10097] <= 1'b1;
     layer1_out[10098] <= layer0_out[4311];
     layer1_out[10099] <= layer0_out[10744] & ~layer0_out[10743];
     layer1_out[10100] <= ~layer0_out[3118];
     layer1_out[10101] <= layer0_out[10454] & ~layer0_out[10455];
     layer1_out[10102] <= layer0_out[1525] ^ layer0_out[1526];
     layer1_out[10103] <= ~(layer0_out[7202] & layer0_out[7203]);
     layer1_out[10104] <= layer0_out[10641] & ~layer0_out[10642];
     layer1_out[10105] <= ~(layer0_out[3839] ^ layer0_out[3840]);
     layer1_out[10106] <= ~(layer0_out[7678] & layer0_out[7679]);
     layer1_out[10107] <= layer0_out[5036];
     layer1_out[10108] <= layer0_out[7735] & ~layer0_out[7736];
     layer1_out[10109] <= ~layer0_out[8347];
     layer1_out[10110] <= ~layer0_out[7130];
     layer1_out[10111] <= ~(layer0_out[11745] & layer0_out[11746]);
     layer1_out[10112] <= ~layer0_out[4114] | layer0_out[4115];
     layer1_out[10113] <= ~(layer0_out[6777] | layer0_out[6778]);
     layer1_out[10114] <= layer0_out[3003] | layer0_out[3004];
     layer1_out[10115] <= layer0_out[7401] ^ layer0_out[7402];
     layer1_out[10116] <= ~layer0_out[8004] | layer0_out[8005];
     layer1_out[10117] <= layer0_out[8494] ^ layer0_out[8495];
     layer1_out[10118] <= ~(layer0_out[515] | layer0_out[516]);
     layer1_out[10119] <= ~layer0_out[11050] | layer0_out[11051];
     layer1_out[10120] <= ~(layer0_out[6152] & layer0_out[6153]);
     layer1_out[10121] <= layer0_out[420] & ~layer0_out[419];
     layer1_out[10122] <= layer0_out[5381] | layer0_out[5382];
     layer1_out[10123] <= ~(layer0_out[2852] & layer0_out[2853]);
     layer1_out[10124] <= ~(layer0_out[10751] & layer0_out[10752]);
     layer1_out[10125] <= ~layer0_out[6085] | layer0_out[6084];
     layer1_out[10126] <= ~(layer0_out[2939] | layer0_out[2940]);
     layer1_out[10127] <= ~(layer0_out[6685] | layer0_out[6686]);
     layer1_out[10128] <= ~layer0_out[7947] | layer0_out[7946];
     layer1_out[10129] <= layer0_out[427] ^ layer0_out[428];
     layer1_out[10130] <= ~layer0_out[1370];
     layer1_out[10131] <= layer0_out[6140];
     layer1_out[10132] <= layer0_out[5822] & ~layer0_out[5821];
     layer1_out[10133] <= ~layer0_out[2101];
     layer1_out[10134] <= layer0_out[222] & ~layer0_out[223];
     layer1_out[10135] <= layer0_out[613] & ~layer0_out[612];
     layer1_out[10136] <= layer0_out[4990] | layer0_out[4991];
     layer1_out[10137] <= ~(layer0_out[8332] | layer0_out[8333]);
     layer1_out[10138] <= layer0_out[12] ^ layer0_out[13];
     layer1_out[10139] <= ~layer0_out[8031];
     layer1_out[10140] <= layer0_out[10505];
     layer1_out[10141] <= ~layer0_out[10885] | layer0_out[10884];
     layer1_out[10142] <= layer0_out[10990] | layer0_out[10991];
     layer1_out[10143] <= layer0_out[9233];
     layer1_out[10144] <= ~layer0_out[10634] | layer0_out[10633];
     layer1_out[10145] <= 1'b0;
     layer1_out[10146] <= ~layer0_out[7751] | layer0_out[7750];
     layer1_out[10147] <= ~(layer0_out[1147] | layer0_out[1148]);
     layer1_out[10148] <= layer0_out[4505] & ~layer0_out[4506];
     layer1_out[10149] <= layer0_out[10339] & layer0_out[10340];
     layer1_out[10150] <= layer0_out[9661];
     layer1_out[10151] <= layer0_out[6171] | layer0_out[6172];
     layer1_out[10152] <= ~layer0_out[218];
     layer1_out[10153] <= ~layer0_out[129] | layer0_out[130];
     layer1_out[10154] <= layer0_out[1191];
     layer1_out[10155] <= layer0_out[6390] & ~layer0_out[6391];
     layer1_out[10156] <= layer0_out[11796] & ~layer0_out[11797];
     layer1_out[10157] <= ~layer0_out[8632] | layer0_out[8633];
     layer1_out[10158] <= ~layer0_out[2750] | layer0_out[2751];
     layer1_out[10159] <= layer0_out[6497];
     layer1_out[10160] <= ~(layer0_out[6266] & layer0_out[6267]);
     layer1_out[10161] <= ~(layer0_out[11549] & layer0_out[11550]);
     layer1_out[10162] <= layer0_out[6817] & layer0_out[6818];
     layer1_out[10163] <= ~(layer0_out[8941] ^ layer0_out[8942]);
     layer1_out[10164] <= 1'b0;
     layer1_out[10165] <= ~layer0_out[3356] | layer0_out[3355];
     layer1_out[10166] <= layer0_out[9189] | layer0_out[9190];
     layer1_out[10167] <= ~layer0_out[4271] | layer0_out[4270];
     layer1_out[10168] <= layer0_out[780] & ~layer0_out[779];
     layer1_out[10169] <= layer0_out[10353] & ~layer0_out[10354];
     layer1_out[10170] <= layer0_out[10836] & ~layer0_out[10837];
     layer1_out[10171] <= ~(layer0_out[4998] & layer0_out[4999]);
     layer1_out[10172] <= ~(layer0_out[8092] | layer0_out[8093]);
     layer1_out[10173] <= layer0_out[8790] & ~layer0_out[8791];
     layer1_out[10174] <= ~layer0_out[1743] | layer0_out[1742];
     layer1_out[10175] <= ~layer0_out[11580];
     layer1_out[10176] <= ~layer0_out[11799] | layer0_out[11798];
     layer1_out[10177] <= layer0_out[409] & ~layer0_out[410];
     layer1_out[10178] <= layer0_out[9732];
     layer1_out[10179] <= ~layer0_out[4111] | layer0_out[4112];
     layer1_out[10180] <= 1'b1;
     layer1_out[10181] <= layer0_out[5652] & layer0_out[5653];
     layer1_out[10182] <= layer0_out[7935] | layer0_out[7936];
     layer1_out[10183] <= ~layer0_out[7781];
     layer1_out[10184] <= ~layer0_out[11245] | layer0_out[11244];
     layer1_out[10185] <= ~(layer0_out[11045] | layer0_out[11046]);
     layer1_out[10186] <= layer0_out[8629] & layer0_out[8630];
     layer1_out[10187] <= layer0_out[7623] & ~layer0_out[7624];
     layer1_out[10188] <= ~layer0_out[1659];
     layer1_out[10189] <= layer0_out[6643];
     layer1_out[10190] <= ~layer0_out[6556];
     layer1_out[10191] <= ~(layer0_out[5939] & layer0_out[5940]);
     layer1_out[10192] <= layer0_out[337] | layer0_out[338];
     layer1_out[10193] <= 1'b1;
     layer1_out[10194] <= ~(layer0_out[7407] ^ layer0_out[7408]);
     layer1_out[10195] <= ~layer0_out[3747];
     layer1_out[10196] <= ~layer0_out[1463];
     layer1_out[10197] <= ~layer0_out[4708];
     layer1_out[10198] <= ~(layer0_out[3224] | layer0_out[3225]);
     layer1_out[10199] <= ~(layer0_out[4493] | layer0_out[4494]);
     layer1_out[10200] <= layer0_out[11215] | layer0_out[11216];
     layer1_out[10201] <= ~layer0_out[3202];
     layer1_out[10202] <= layer0_out[6946];
     layer1_out[10203] <= ~(layer0_out[3301] | layer0_out[3302]);
     layer1_out[10204] <= 1'b0;
     layer1_out[10205] <= ~(layer0_out[7765] & layer0_out[7766]);
     layer1_out[10206] <= layer0_out[5755] | layer0_out[5756];
     layer1_out[10207] <= layer0_out[2957] & ~layer0_out[2958];
     layer1_out[10208] <= ~layer0_out[6667];
     layer1_out[10209] <= layer0_out[2133];
     layer1_out[10210] <= ~(layer0_out[601] | layer0_out[602]);
     layer1_out[10211] <= layer0_out[9405] & layer0_out[9406];
     layer1_out[10212] <= layer0_out[2042];
     layer1_out[10213] <= layer0_out[9525] & ~layer0_out[9524];
     layer1_out[10214] <= layer0_out[3637] | layer0_out[3638];
     layer1_out[10215] <= layer0_out[4169] & layer0_out[4170];
     layer1_out[10216] <= ~(layer0_out[5825] & layer0_out[5826]);
     layer1_out[10217] <= ~layer0_out[1777];
     layer1_out[10218] <= ~layer0_out[6824] | layer0_out[6825];
     layer1_out[10219] <= ~layer0_out[9929] | layer0_out[9930];
     layer1_out[10220] <= layer0_out[4651] & ~layer0_out[4652];
     layer1_out[10221] <= ~layer0_out[9430];
     layer1_out[10222] <= ~(layer0_out[8127] & layer0_out[8128]);
     layer1_out[10223] <= layer0_out[3894];
     layer1_out[10224] <= ~layer0_out[7031];
     layer1_out[10225] <= ~(layer0_out[8415] | layer0_out[8416]);
     layer1_out[10226] <= ~layer0_out[793];
     layer1_out[10227] <= ~layer0_out[7552] | layer0_out[7553];
     layer1_out[10228] <= layer0_out[9847] & ~layer0_out[9846];
     layer1_out[10229] <= ~(layer0_out[9678] & layer0_out[9679]);
     layer1_out[10230] <= layer0_out[9679] & layer0_out[9680];
     layer1_out[10231] <= ~layer0_out[2198];
     layer1_out[10232] <= ~layer0_out[11683] | layer0_out[11682];
     layer1_out[10233] <= ~(layer0_out[311] | layer0_out[312]);
     layer1_out[10234] <= ~(layer0_out[4806] ^ layer0_out[4807]);
     layer1_out[10235] <= layer0_out[7436] & ~layer0_out[7437];
     layer1_out[10236] <= ~(layer0_out[6330] & layer0_out[6331]);
     layer1_out[10237] <= layer0_out[3248] & layer0_out[3249];
     layer1_out[10238] <= layer0_out[3034] & ~layer0_out[3033];
     layer1_out[10239] <= ~(layer0_out[10145] & layer0_out[10146]);
     layer1_out[10240] <= layer0_out[611];
     layer1_out[10241] <= ~(layer0_out[7652] ^ layer0_out[7653]);
     layer1_out[10242] <= layer0_out[1831] ^ layer0_out[1832];
     layer1_out[10243] <= layer0_out[8226] ^ layer0_out[8227];
     layer1_out[10244] <= ~layer0_out[7630] | layer0_out[7629];
     layer1_out[10245] <= ~(layer0_out[9121] | layer0_out[9122]);
     layer1_out[10246] <= ~layer0_out[6932] | layer0_out[6933];
     layer1_out[10247] <= layer0_out[8023] ^ layer0_out[8024];
     layer1_out[10248] <= ~(layer0_out[7733] ^ layer0_out[7734]);
     layer1_out[10249] <= layer0_out[10733] | layer0_out[10734];
     layer1_out[10250] <= layer0_out[6022];
     layer1_out[10251] <= 1'b1;
     layer1_out[10252] <= layer0_out[11165] & ~layer0_out[11164];
     layer1_out[10253] <= layer0_out[3667] & ~layer0_out[3668];
     layer1_out[10254] <= layer0_out[3880];
     layer1_out[10255] <= ~layer0_out[941];
     layer1_out[10256] <= layer0_out[3854] & ~layer0_out[3853];
     layer1_out[10257] <= ~layer0_out[4320];
     layer1_out[10258] <= ~layer0_out[11649] | layer0_out[11648];
     layer1_out[10259] <= layer0_out[2184] | layer0_out[2185];
     layer1_out[10260] <= ~(layer0_out[10367] | layer0_out[10368]);
     layer1_out[10261] <= layer0_out[1207];
     layer1_out[10262] <= ~layer0_out[11273] | layer0_out[11274];
     layer1_out[10263] <= ~(layer0_out[493] ^ layer0_out[494]);
     layer1_out[10264] <= ~layer0_out[11786];
     layer1_out[10265] <= ~layer0_out[5663];
     layer1_out[10266] <= ~layer0_out[9394];
     layer1_out[10267] <= layer0_out[1882] & ~layer0_out[1881];
     layer1_out[10268] <= ~layer0_out[404] | layer0_out[405];
     layer1_out[10269] <= layer0_out[4476] & ~layer0_out[4477];
     layer1_out[10270] <= layer0_out[6543] & ~layer0_out[6544];
     layer1_out[10271] <= ~layer0_out[11392] | layer0_out[11393];
     layer1_out[10272] <= layer0_out[7118] & layer0_out[7119];
     layer1_out[10273] <= ~layer0_out[1806];
     layer1_out[10274] <= 1'b0;
     layer1_out[10275] <= ~(layer0_out[9408] | layer0_out[9409]);
     layer1_out[10276] <= layer0_out[10630] | layer0_out[10631];
     layer1_out[10277] <= ~(layer0_out[2597] ^ layer0_out[2598]);
     layer1_out[10278] <= ~(layer0_out[815] | layer0_out[816]);
     layer1_out[10279] <= layer0_out[3570] & ~layer0_out[3571];
     layer1_out[10280] <= ~layer0_out[1457];
     layer1_out[10281] <= ~(layer0_out[7957] | layer0_out[7958]);
     layer1_out[10282] <= ~(layer0_out[9903] | layer0_out[9904]);
     layer1_out[10283] <= ~layer0_out[10665] | layer0_out[10666];
     layer1_out[10284] <= ~layer0_out[10128] | layer0_out[10127];
     layer1_out[10285] <= ~layer0_out[5234];
     layer1_out[10286] <= ~(layer0_out[9491] & layer0_out[9492]);
     layer1_out[10287] <= ~(layer0_out[10644] | layer0_out[10645]);
     layer1_out[10288] <= ~(layer0_out[3460] & layer0_out[3461]);
     layer1_out[10289] <= layer0_out[4412] & layer0_out[4413];
     layer1_out[10290] <= ~layer0_out[3784];
     layer1_out[10291] <= layer0_out[6743];
     layer1_out[10292] <= ~(layer0_out[6335] | layer0_out[6336]);
     layer1_out[10293] <= layer0_out[1186] & layer0_out[1187];
     layer1_out[10294] <= layer0_out[1509] & ~layer0_out[1508];
     layer1_out[10295] <= layer0_out[10820] ^ layer0_out[10821];
     layer1_out[10296] <= layer0_out[9569] & ~layer0_out[9570];
     layer1_out[10297] <= layer0_out[835] & layer0_out[836];
     layer1_out[10298] <= 1'b1;
     layer1_out[10299] <= layer0_out[2607];
     layer1_out[10300] <= ~(layer0_out[9124] | layer0_out[9125]);
     layer1_out[10301] <= layer0_out[1687] & layer0_out[1688];
     layer1_out[10302] <= ~layer0_out[2817] | layer0_out[2816];
     layer1_out[10303] <= ~(layer0_out[8244] ^ layer0_out[8245]);
     layer1_out[10304] <= ~layer0_out[3809] | layer0_out[3810];
     layer1_out[10305] <= ~(layer0_out[5686] ^ layer0_out[5687]);
     layer1_out[10306] <= ~(layer0_out[5685] & layer0_out[5686]);
     layer1_out[10307] <= layer0_out[3434] ^ layer0_out[3435];
     layer1_out[10308] <= ~layer0_out[10971] | layer0_out[10972];
     layer1_out[10309] <= layer0_out[10181] & ~layer0_out[10182];
     layer1_out[10310] <= ~layer0_out[8371];
     layer1_out[10311] <= layer0_out[10592];
     layer1_out[10312] <= ~(layer0_out[5103] | layer0_out[5104]);
     layer1_out[10313] <= layer0_out[7716];
     layer1_out[10314] <= ~layer0_out[1102];
     layer1_out[10315] <= ~layer0_out[6602] | layer0_out[6603];
     layer1_out[10316] <= ~(layer0_out[25] ^ layer0_out[26]);
     layer1_out[10317] <= ~(layer0_out[11008] | layer0_out[11009]);
     layer1_out[10318] <= ~layer0_out[9544];
     layer1_out[10319] <= layer0_out[5443] ^ layer0_out[5444];
     layer1_out[10320] <= layer0_out[11762];
     layer1_out[10321] <= layer0_out[7588] & layer0_out[7589];
     layer1_out[10322] <= ~(layer0_out[8123] & layer0_out[8124]);
     layer1_out[10323] <= ~(layer0_out[6825] | layer0_out[6826]);
     layer1_out[10324] <= 1'b1;
     layer1_out[10325] <= layer0_out[11973] & ~layer0_out[11972];
     layer1_out[10326] <= layer0_out[5696];
     layer1_out[10327] <= layer0_out[2277];
     layer1_out[10328] <= layer0_out[1660] ^ layer0_out[1661];
     layer1_out[10329] <= ~layer0_out[11830];
     layer1_out[10330] <= ~(layer0_out[9727] & layer0_out[9728]);
     layer1_out[10331] <= ~layer0_out[7047] | layer0_out[7046];
     layer1_out[10332] <= ~layer0_out[2430];
     layer1_out[10333] <= ~layer0_out[9116];
     layer1_out[10334] <= 1'b1;
     layer1_out[10335] <= ~layer0_out[2428];
     layer1_out[10336] <= layer0_out[7190];
     layer1_out[10337] <= ~(layer0_out[9302] | layer0_out[9303]);
     layer1_out[10338] <= layer0_out[5322] & ~layer0_out[5323];
     layer1_out[10339] <= ~(layer0_out[7364] ^ layer0_out[7365]);
     layer1_out[10340] <= ~layer0_out[5817];
     layer1_out[10341] <= layer0_out[2544] & ~layer0_out[2545];
     layer1_out[10342] <= ~(layer0_out[4419] ^ layer0_out[4420]);
     layer1_out[10343] <= layer0_out[4282] & ~layer0_out[4283];
     layer1_out[10344] <= ~layer0_out[5955];
     layer1_out[10345] <= layer0_out[2110] | layer0_out[2111];
     layer1_out[10346] <= layer0_out[3469] | layer0_out[3470];
     layer1_out[10347] <= layer0_out[6117] & layer0_out[6118];
     layer1_out[10348] <= layer0_out[3318] & layer0_out[3319];
     layer1_out[10349] <= ~layer0_out[2370];
     layer1_out[10350] <= ~layer0_out[8840] | layer0_out[8839];
     layer1_out[10351] <= ~(layer0_out[6002] | layer0_out[6003]);
     layer1_out[10352] <= ~(layer0_out[4074] & layer0_out[4075]);
     layer1_out[10353] <= ~layer0_out[11356] | layer0_out[11357];
     layer1_out[10354] <= ~layer0_out[6711] | layer0_out[6712];
     layer1_out[10355] <= ~layer0_out[6807] | layer0_out[6808];
     layer1_out[10356] <= layer0_out[3622] | layer0_out[3623];
     layer1_out[10357] <= ~layer0_out[2713] | layer0_out[2714];
     layer1_out[10358] <= layer0_out[2436] & layer0_out[2437];
     layer1_out[10359] <= ~(layer0_out[11884] ^ layer0_out[11885]);
     layer1_out[10360] <= ~layer0_out[2399];
     layer1_out[10361] <= layer0_out[1369];
     layer1_out[10362] <= ~layer0_out[1647];
     layer1_out[10363] <= ~(layer0_out[7509] | layer0_out[7510]);
     layer1_out[10364] <= ~layer0_out[9811];
     layer1_out[10365] <= ~(layer0_out[2495] | layer0_out[2496]);
     layer1_out[10366] <= layer0_out[7436] & ~layer0_out[7435];
     layer1_out[10367] <= ~(layer0_out[2752] & layer0_out[2753]);
     layer1_out[10368] <= ~(layer0_out[5399] & layer0_out[5400]);
     layer1_out[10369] <= layer0_out[7218] & ~layer0_out[7217];
     layer1_out[10370] <= ~layer0_out[0] | layer0_out[2];
     layer1_out[10371] <= 1'b1;
     layer1_out[10372] <= ~(layer0_out[1703] & layer0_out[1704]);
     layer1_out[10373] <= ~layer0_out[5041];
     layer1_out[10374] <= layer0_out[7596];
     layer1_out[10375] <= ~layer0_out[5653];
     layer1_out[10376] <= ~(layer0_out[6856] & layer0_out[6857]);
     layer1_out[10377] <= layer0_out[10551];
     layer1_out[10378] <= ~layer0_out[8128] | layer0_out[8129];
     layer1_out[10379] <= ~layer0_out[2774];
     layer1_out[10380] <= ~(layer0_out[11426] ^ layer0_out[11427]);
     layer1_out[10381] <= ~layer0_out[1985] | layer0_out[1986];
     layer1_out[10382] <= 1'b1;
     layer1_out[10383] <= ~(layer0_out[9666] ^ layer0_out[9667]);
     layer1_out[10384] <= layer0_out[2307] ^ layer0_out[2308];
     layer1_out[10385] <= ~(layer0_out[11844] & layer0_out[11845]);
     layer1_out[10386] <= ~(layer0_out[2858] | layer0_out[2859]);
     layer1_out[10387] <= layer0_out[4146] ^ layer0_out[4147];
     layer1_out[10388] <= layer0_out[10681] | layer0_out[10682];
     layer1_out[10389] <= ~(layer0_out[2306] & layer0_out[2307]);
     layer1_out[10390] <= ~layer0_out[5783];
     layer1_out[10391] <= layer0_out[435] & ~layer0_out[434];
     layer1_out[10392] <= layer0_out[4762] & ~layer0_out[4761];
     layer1_out[10393] <= layer0_out[2652];
     layer1_out[10394] <= ~layer0_out[1104] | layer0_out[1103];
     layer1_out[10395] <= ~layer0_out[10748];
     layer1_out[10396] <= 1'b0;
     layer1_out[10397] <= ~layer0_out[8697];
     layer1_out[10398] <= layer0_out[10243];
     layer1_out[10399] <= ~(layer0_out[5229] & layer0_out[5230]);
     layer1_out[10400] <= layer0_out[1379] & layer0_out[1380];
     layer1_out[10401] <= ~layer0_out[9410];
     layer1_out[10402] <= layer0_out[9620] | layer0_out[9621];
     layer1_out[10403] <= layer0_out[5182] & ~layer0_out[5181];
     layer1_out[10404] <= layer0_out[263];
     layer1_out[10405] <= layer0_out[10983];
     layer1_out[10406] <= ~layer0_out[8162];
     layer1_out[10407] <= layer0_out[9258];
     layer1_out[10408] <= ~(layer0_out[4606] | layer0_out[4607]);
     layer1_out[10409] <= ~(layer0_out[9480] | layer0_out[9481]);
     layer1_out[10410] <= layer0_out[11414] & ~layer0_out[11415];
     layer1_out[10411] <= ~layer0_out[2780] | layer0_out[2781];
     layer1_out[10412] <= ~(layer0_out[6487] | layer0_out[6488]);
     layer1_out[10413] <= ~layer0_out[5871] | layer0_out[5870];
     layer1_out[10414] <= layer0_out[5353] & ~layer0_out[5354];
     layer1_out[10415] <= ~layer0_out[10697];
     layer1_out[10416] <= layer0_out[11384] ^ layer0_out[11385];
     layer1_out[10417] <= layer0_out[2291];
     layer1_out[10418] <= layer0_out[5028];
     layer1_out[10419] <= layer0_out[41] & ~layer0_out[42];
     layer1_out[10420] <= layer0_out[2048] | layer0_out[2049];
     layer1_out[10421] <= layer0_out[11434];
     layer1_out[10422] <= layer0_out[7878] | layer0_out[7879];
     layer1_out[10423] <= ~(layer0_out[10490] & layer0_out[10491]);
     layer1_out[10424] <= 1'b1;
     layer1_out[10425] <= layer0_out[11672] & ~layer0_out[11671];
     layer1_out[10426] <= ~(layer0_out[4947] & layer0_out[4948]);
     layer1_out[10427] <= layer0_out[9681] | layer0_out[9682];
     layer1_out[10428] <= layer0_out[943];
     layer1_out[10429] <= layer0_out[7979];
     layer1_out[10430] <= ~layer0_out[1204] | layer0_out[1203];
     layer1_out[10431] <= layer0_out[11185];
     layer1_out[10432] <= layer0_out[1684] & ~layer0_out[1683];
     layer1_out[10433] <= ~layer0_out[5446];
     layer1_out[10434] <= ~(layer0_out[6430] | layer0_out[6431]);
     layer1_out[10435] <= 1'b1;
     layer1_out[10436] <= layer0_out[5855] & ~layer0_out[5854];
     layer1_out[10437] <= ~(layer0_out[3496] & layer0_out[3497]);
     layer1_out[10438] <= ~layer0_out[5652];
     layer1_out[10439] <= layer0_out[10965] & ~layer0_out[10964];
     layer1_out[10440] <= layer0_out[6051];
     layer1_out[10441] <= layer0_out[2951];
     layer1_out[10442] <= layer0_out[9244] & ~layer0_out[9243];
     layer1_out[10443] <= ~layer0_out[8737];
     layer1_out[10444] <= ~(layer0_out[7248] & layer0_out[7249]);
     layer1_out[10445] <= ~(layer0_out[4397] | layer0_out[4398]);
     layer1_out[10446] <= ~(layer0_out[8351] & layer0_out[8352]);
     layer1_out[10447] <= ~(layer0_out[10125] & layer0_out[10126]);
     layer1_out[10448] <= 1'b0;
     layer1_out[10449] <= layer0_out[359];
     layer1_out[10450] <= ~(layer0_out[3524] ^ layer0_out[3525]);
     layer1_out[10451] <= layer0_out[11977] | layer0_out[11978];
     layer1_out[10452] <= ~layer0_out[7711] | layer0_out[7712];
     layer1_out[10453] <= 1'b1;
     layer1_out[10454] <= ~layer0_out[334] | layer0_out[333];
     layer1_out[10455] <= ~layer0_out[2295] | layer0_out[2294];
     layer1_out[10456] <= layer0_out[2776] & ~layer0_out[2777];
     layer1_out[10457] <= layer0_out[5816] ^ layer0_out[5817];
     layer1_out[10458] <= layer0_out[6408] | layer0_out[6409];
     layer1_out[10459] <= layer0_out[10460] & ~layer0_out[10459];
     layer1_out[10460] <= ~layer0_out[5247];
     layer1_out[10461] <= layer0_out[11150] ^ layer0_out[11151];
     layer1_out[10462] <= layer0_out[839];
     layer1_out[10463] <= layer0_out[6261];
     layer1_out[10464] <= ~layer0_out[8956];
     layer1_out[10465] <= layer0_out[3980];
     layer1_out[10466] <= layer0_out[9628] & layer0_out[9629];
     layer1_out[10467] <= ~layer0_out[4233];
     layer1_out[10468] <= layer0_out[2976];
     layer1_out[10469] <= layer0_out[11872] & ~layer0_out[11871];
     layer1_out[10470] <= ~(layer0_out[8214] ^ layer0_out[8215]);
     layer1_out[10471] <= ~layer0_out[4899];
     layer1_out[10472] <= 1'b0;
     layer1_out[10473] <= ~layer0_out[9208] | layer0_out[9209];
     layer1_out[10474] <= layer0_out[10450] & ~layer0_out[10449];
     layer1_out[10475] <= ~(layer0_out[935] & layer0_out[936]);
     layer1_out[10476] <= ~layer0_out[3413];
     layer1_out[10477] <= layer0_out[10230] & ~layer0_out[10231];
     layer1_out[10478] <= layer0_out[8452] & layer0_out[8453];
     layer1_out[10479] <= ~layer0_out[330] | layer0_out[329];
     layer1_out[10480] <= layer0_out[4675] & ~layer0_out[4676];
     layer1_out[10481] <= ~(layer0_out[2850] | layer0_out[2851]);
     layer1_out[10482] <= layer0_out[11922] & ~layer0_out[11923];
     layer1_out[10483] <= ~layer0_out[2144];
     layer1_out[10484] <= ~layer0_out[11684] | layer0_out[11685];
     layer1_out[10485] <= layer0_out[5991];
     layer1_out[10486] <= layer0_out[5130];
     layer1_out[10487] <= layer0_out[8306];
     layer1_out[10488] <= layer0_out[7398];
     layer1_out[10489] <= 1'b1;
     layer1_out[10490] <= layer0_out[4575];
     layer1_out[10491] <= ~layer0_out[821];
     layer1_out[10492] <= ~(layer0_out[6252] & layer0_out[6253]);
     layer1_out[10493] <= ~layer0_out[5510];
     layer1_out[10494] <= layer0_out[9502];
     layer1_out[10495] <= ~layer0_out[709] | layer0_out[710];
     layer1_out[10496] <= layer0_out[1025] ^ layer0_out[1026];
     layer1_out[10497] <= ~layer0_out[8873];
     layer1_out[10498] <= ~(layer0_out[5947] ^ layer0_out[5948]);
     layer1_out[10499] <= layer0_out[8824];
     layer1_out[10500] <= 1'b0;
     layer1_out[10501] <= ~layer0_out[4706];
     layer1_out[10502] <= ~(layer0_out[10956] & layer0_out[10957]);
     layer1_out[10503] <= layer0_out[7490] & ~layer0_out[7489];
     layer1_out[10504] <= 1'b0;
     layer1_out[10505] <= ~(layer0_out[8172] & layer0_out[8173]);
     layer1_out[10506] <= layer0_out[4486] & ~layer0_out[4487];
     layer1_out[10507] <= layer0_out[4086] | layer0_out[4087];
     layer1_out[10508] <= ~(layer0_out[10026] ^ layer0_out[10027]);
     layer1_out[10509] <= ~layer0_out[1307];
     layer1_out[10510] <= layer0_out[4262];
     layer1_out[10511] <= ~(layer0_out[3228] & layer0_out[3229]);
     layer1_out[10512] <= ~(layer0_out[7756] & layer0_out[7757]);
     layer1_out[10513] <= ~(layer0_out[4136] & layer0_out[4137]);
     layer1_out[10514] <= ~layer0_out[11693];
     layer1_out[10515] <= layer0_out[4025] & layer0_out[4026];
     layer1_out[10516] <= layer0_out[6353];
     layer1_out[10517] <= layer0_out[668];
     layer1_out[10518] <= ~layer0_out[1728];
     layer1_out[10519] <= ~(layer0_out[3698] | layer0_out[3699]);
     layer1_out[10520] <= layer0_out[9566] | layer0_out[9567];
     layer1_out[10521] <= ~(layer0_out[6263] | layer0_out[6264]);
     layer1_out[10522] <= layer0_out[2556] ^ layer0_out[2557];
     layer1_out[10523] <= ~layer0_out[5067];
     layer1_out[10524] <= ~(layer0_out[22] ^ layer0_out[23]);
     layer1_out[10525] <= layer0_out[10628] & ~layer0_out[10627];
     layer1_out[10526] <= layer0_out[144];
     layer1_out[10527] <= layer0_out[4071] & ~layer0_out[4070];
     layer1_out[10528] <= layer0_out[4627] | layer0_out[4628];
     layer1_out[10529] <= layer0_out[7617];
     layer1_out[10530] <= layer0_out[4653];
     layer1_out[10531] <= layer0_out[2284] | layer0_out[2285];
     layer1_out[10532] <= ~(layer0_out[6942] | layer0_out[6943]);
     layer1_out[10533] <= layer0_out[5619] & ~layer0_out[5618];
     layer1_out[10534] <= ~(layer0_out[6433] & layer0_out[6434]);
     layer1_out[10535] <= layer0_out[9317] & ~layer0_out[9318];
     layer1_out[10536] <= layer0_out[2112] & ~layer0_out[2111];
     layer1_out[10537] <= ~layer0_out[6447];
     layer1_out[10538] <= layer0_out[1122] & ~layer0_out[1121];
     layer1_out[10539] <= layer0_out[11787] & ~layer0_out[11788];
     layer1_out[10540] <= ~layer0_out[560];
     layer1_out[10541] <= ~(layer0_out[3257] | layer0_out[3258]);
     layer1_out[10542] <= ~layer0_out[10778];
     layer1_out[10543] <= ~layer0_out[11965];
     layer1_out[10544] <= layer0_out[10565] & ~layer0_out[10564];
     layer1_out[10545] <= layer0_out[10423] ^ layer0_out[10424];
     layer1_out[10546] <= layer0_out[96] ^ layer0_out[97];
     layer1_out[10547] <= ~layer0_out[9528];
     layer1_out[10548] <= layer0_out[1542] & ~layer0_out[1543];
     layer1_out[10549] <= layer0_out[174] & ~layer0_out[173];
     layer1_out[10550] <= ~layer0_out[11722] | layer0_out[11721];
     layer1_out[10551] <= layer0_out[5563];
     layer1_out[10552] <= 1'b0;
     layer1_out[10553] <= ~(layer0_out[3604] & layer0_out[3605]);
     layer1_out[10554] <= layer0_out[5294];
     layer1_out[10555] <= layer0_out[5459] ^ layer0_out[5460];
     layer1_out[10556] <= layer0_out[4306];
     layer1_out[10557] <= ~layer0_out[9021];
     layer1_out[10558] <= layer0_out[1661] | layer0_out[1662];
     layer1_out[10559] <= layer0_out[408] & ~layer0_out[409];
     layer1_out[10560] <= layer0_out[493];
     layer1_out[10561] <= layer0_out[9264] & layer0_out[9265];
     layer1_out[10562] <= ~(layer0_out[9902] ^ layer0_out[9903]);
     layer1_out[10563] <= layer0_out[4360];
     layer1_out[10564] <= ~layer0_out[2833] | layer0_out[2832];
     layer1_out[10565] <= ~(layer0_out[1169] | layer0_out[1170]);
     layer1_out[10566] <= ~layer0_out[7179] | layer0_out[7180];
     layer1_out[10567] <= layer0_out[973];
     layer1_out[10568] <= layer0_out[117];
     layer1_out[10569] <= layer0_out[11870];
     layer1_out[10570] <= layer0_out[4965] ^ layer0_out[4966];
     layer1_out[10571] <= ~layer0_out[5280];
     layer1_out[10572] <= layer0_out[5716] & layer0_out[5717];
     layer1_out[10573] <= ~layer0_out[2578] | layer0_out[2579];
     layer1_out[10574] <= ~(layer0_out[11271] & layer0_out[11272]);
     layer1_out[10575] <= layer0_out[1098] & layer0_out[1099];
     layer1_out[10576] <= ~layer0_out[1436] | layer0_out[1437];
     layer1_out[10577] <= layer0_out[3101];
     layer1_out[10578] <= layer0_out[8631];
     layer1_out[10579] <= layer0_out[6834] & layer0_out[6835];
     layer1_out[10580] <= layer0_out[6730] & ~layer0_out[6729];
     layer1_out[10581] <= ~(layer0_out[299] | layer0_out[300]);
     layer1_out[10582] <= ~layer0_out[7998] | layer0_out[7997];
     layer1_out[10583] <= layer0_out[9621] & layer0_out[9622];
     layer1_out[10584] <= ~layer0_out[8479] | layer0_out[8480];
     layer1_out[10585] <= ~(layer0_out[11500] ^ layer0_out[11501]);
     layer1_out[10586] <= 1'b0;
     layer1_out[10587] <= ~(layer0_out[3110] | layer0_out[3111]);
     layer1_out[10588] <= ~layer0_out[5282];
     layer1_out[10589] <= layer0_out[3080];
     layer1_out[10590] <= layer0_out[3557];
     layer1_out[10591] <= ~layer0_out[2419];
     layer1_out[10592] <= layer0_out[3261] & ~layer0_out[3262];
     layer1_out[10593] <= ~layer0_out[887];
     layer1_out[10594] <= ~layer0_out[8372];
     layer1_out[10595] <= ~(layer0_out[8822] ^ layer0_out[8823]);
     layer1_out[10596] <= ~(layer0_out[5792] | layer0_out[5793]);
     layer1_out[10597] <= layer0_out[11237] & layer0_out[11238];
     layer1_out[10598] <= ~(layer0_out[9232] | layer0_out[9233]);
     layer1_out[10599] <= ~layer0_out[1552];
     layer1_out[10600] <= ~layer0_out[3055] | layer0_out[3056];
     layer1_out[10601] <= ~layer0_out[5390];
     layer1_out[10602] <= layer0_out[6582] | layer0_out[6583];
     layer1_out[10603] <= ~layer0_out[11275];
     layer1_out[10604] <= layer0_out[8642];
     layer1_out[10605] <= ~layer0_out[7468];
     layer1_out[10606] <= layer0_out[10280] & layer0_out[10281];
     layer1_out[10607] <= layer0_out[10374] & ~layer0_out[10373];
     layer1_out[10608] <= ~layer0_out[1174];
     layer1_out[10609] <= ~layer0_out[3308];
     layer1_out[10610] <= ~(layer0_out[7073] & layer0_out[7074]);
     layer1_out[10611] <= ~layer0_out[11606];
     layer1_out[10612] <= layer0_out[5111];
     layer1_out[10613] <= ~layer0_out[7051];
     layer1_out[10614] <= layer0_out[7891] & ~layer0_out[7890];
     layer1_out[10615] <= ~layer0_out[7808];
     layer1_out[10616] <= ~layer0_out[4090] | layer0_out[4091];
     layer1_out[10617] <= ~layer0_out[5004];
     layer1_out[10618] <= ~layer0_out[2820];
     layer1_out[10619] <= ~layer0_out[4746] | layer0_out[4745];
     layer1_out[10620] <= ~(layer0_out[3522] | layer0_out[3523]);
     layer1_out[10621] <= layer0_out[4686] | layer0_out[4687];
     layer1_out[10622] <= layer0_out[3102] | layer0_out[3103];
     layer1_out[10623] <= ~(layer0_out[7848] | layer0_out[7849]);
     layer1_out[10624] <= layer0_out[7425];
     layer1_out[10625] <= ~layer0_out[9577] | layer0_out[9578];
     layer1_out[10626] <= ~(layer0_out[8445] | layer0_out[8446]);
     layer1_out[10627] <= ~layer0_out[1701];
     layer1_out[10628] <= ~layer0_out[3154] | layer0_out[3155];
     layer1_out[10629] <= layer0_out[7856] & ~layer0_out[7857];
     layer1_out[10630] <= ~(layer0_out[724] & layer0_out[725]);
     layer1_out[10631] <= ~layer0_out[4855];
     layer1_out[10632] <= layer0_out[243] & layer0_out[244];
     layer1_out[10633] <= layer0_out[8243] & ~layer0_out[8244];
     layer1_out[10634] <= ~layer0_out[6177] | layer0_out[6178];
     layer1_out[10635] <= ~layer0_out[11064] | layer0_out[11063];
     layer1_out[10636] <= layer0_out[4945] & layer0_out[4946];
     layer1_out[10637] <= ~(layer0_out[10519] & layer0_out[10520]);
     layer1_out[10638] <= layer0_out[11459] & layer0_out[11460];
     layer1_out[10639] <= layer0_out[5845];
     layer1_out[10640] <= layer0_out[8836] & ~layer0_out[8835];
     layer1_out[10641] <= layer0_out[3343] & ~layer0_out[3342];
     layer1_out[10642] <= layer0_out[9913] & ~layer0_out[9912];
     layer1_out[10643] <= layer0_out[4571];
     layer1_out[10644] <= 1'b0;
     layer1_out[10645] <= 1'b0;
     layer1_out[10646] <= ~layer0_out[2377];
     layer1_out[10647] <= ~layer0_out[3544] | layer0_out[3545];
     layer1_out[10648] <= layer0_out[7309];
     layer1_out[10649] <= layer0_out[8259] | layer0_out[8260];
     layer1_out[10650] <= ~layer0_out[3242];
     layer1_out[10651] <= ~layer0_out[3077];
     layer1_out[10652] <= 1'b1;
     layer1_out[10653] <= layer0_out[11342] ^ layer0_out[11343];
     layer1_out[10654] <= ~layer0_out[6328] | layer0_out[6329];
     layer1_out[10655] <= ~(layer0_out[10217] | layer0_out[10218]);
     layer1_out[10656] <= ~layer0_out[3162];
     layer1_out[10657] <= layer0_out[232];
     layer1_out[10658] <= layer0_out[1602] & ~layer0_out[1601];
     layer1_out[10659] <= ~(layer0_out[6712] & layer0_out[6713]);
     layer1_out[10660] <= 1'b0;
     layer1_out[10661] <= layer0_out[2233] & ~layer0_out[2232];
     layer1_out[10662] <= ~layer0_out[9988];
     layer1_out[10663] <= ~layer0_out[1310] | layer0_out[1309];
     layer1_out[10664] <= ~(layer0_out[11786] ^ layer0_out[11787]);
     layer1_out[10665] <= layer0_out[3984];
     layer1_out[10666] <= layer0_out[3896];
     layer1_out[10667] <= layer0_out[1890] & ~layer0_out[1891];
     layer1_out[10668] <= layer0_out[10372] & layer0_out[10373];
     layer1_out[10669] <= layer0_out[2554];
     layer1_out[10670] <= layer0_out[1263] ^ layer0_out[1264];
     layer1_out[10671] <= layer0_out[11187];
     layer1_out[10672] <= layer0_out[5032] & ~layer0_out[5033];
     layer1_out[10673] <= ~layer0_out[3234];
     layer1_out[10674] <= layer0_out[10789];
     layer1_out[10675] <= 1'b1;
     layer1_out[10676] <= layer0_out[5320] & ~layer0_out[5319];
     layer1_out[10677] <= ~layer0_out[5204];
     layer1_out[10678] <= ~(layer0_out[3450] ^ layer0_out[3451]);
     layer1_out[10679] <= ~layer0_out[5943];
     layer1_out[10680] <= layer0_out[4132];
     layer1_out[10681] <= layer0_out[1755] | layer0_out[1756];
     layer1_out[10682] <= ~layer0_out[2614];
     layer1_out[10683] <= layer0_out[11045];
     layer1_out[10684] <= layer0_out[7196] | layer0_out[7197];
     layer1_out[10685] <= layer0_out[7451] & layer0_out[7452];
     layer1_out[10686] <= 1'b1;
     layer1_out[10687] <= layer0_out[9556] ^ layer0_out[9557];
     layer1_out[10688] <= ~layer0_out[6098];
     layer1_out[10689] <= layer0_out[4391] & ~layer0_out[4390];
     layer1_out[10690] <= ~(layer0_out[8122] & layer0_out[8123]);
     layer1_out[10691] <= ~layer0_out[4688];
     layer1_out[10692] <= 1'b1;
     layer1_out[10693] <= ~(layer0_out[647] ^ layer0_out[648]);
     layer1_out[10694] <= layer0_out[10631] ^ layer0_out[10632];
     layer1_out[10695] <= ~(layer0_out[5155] | layer0_out[5156]);
     layer1_out[10696] <= layer0_out[6354] & ~layer0_out[6355];
     layer1_out[10697] <= ~layer0_out[443] | layer0_out[442];
     layer1_out[10698] <= layer0_out[39] | layer0_out[40];
     layer1_out[10699] <= layer0_out[1326];
     layer1_out[10700] <= 1'b0;
     layer1_out[10701] <= ~layer0_out[8078];
     layer1_out[10702] <= layer0_out[4352];
     layer1_out[10703] <= ~layer0_out[372];
     layer1_out[10704] <= layer0_out[10034];
     layer1_out[10705] <= ~layer0_out[3734];
     layer1_out[10706] <= layer0_out[11429] | layer0_out[11430];
     layer1_out[10707] <= layer0_out[10471];
     layer1_out[10708] <= 1'b0;
     layer1_out[10709] <= ~layer0_out[3382] | layer0_out[3383];
     layer1_out[10710] <= ~layer0_out[8166];
     layer1_out[10711] <= layer0_out[7371] & ~layer0_out[7370];
     layer1_out[10712] <= layer0_out[3214];
     layer1_out[10713] <= layer0_out[5936];
     layer1_out[10714] <= layer0_out[7844] & ~layer0_out[7843];
     layer1_out[10715] <= layer0_out[10175] & layer0_out[10176];
     layer1_out[10716] <= ~(layer0_out[4130] | layer0_out[4131]);
     layer1_out[10717] <= ~layer0_out[5030] | layer0_out[5029];
     layer1_out[10718] <= ~layer0_out[5875] | layer0_out[5876];
     layer1_out[10719] <= ~layer0_out[8112] | layer0_out[8111];
     layer1_out[10720] <= layer0_out[4474];
     layer1_out[10721] <= layer0_out[8744] ^ layer0_out[8745];
     layer1_out[10722] <= ~layer0_out[8483];
     layer1_out[10723] <= ~(layer0_out[8966] & layer0_out[8967]);
     layer1_out[10724] <= layer0_out[900];
     layer1_out[10725] <= layer0_out[8404];
     layer1_out[10726] <= ~layer0_out[4523];
     layer1_out[10727] <= ~(layer0_out[4391] & layer0_out[4392]);
     layer1_out[10728] <= layer0_out[2081];
     layer1_out[10729] <= layer0_out[9014] & ~layer0_out[9013];
     layer1_out[10730] <= ~(layer0_out[5773] ^ layer0_out[5774]);
     layer1_out[10731] <= layer0_out[3418] & ~layer0_out[3419];
     layer1_out[10732] <= layer0_out[925] & ~layer0_out[924];
     layer1_out[10733] <= ~(layer0_out[10722] & layer0_out[10723]);
     layer1_out[10734] <= ~layer0_out[1580] | layer0_out[1579];
     layer1_out[10735] <= layer0_out[6083] & ~layer0_out[6082];
     layer1_out[10736] <= ~(layer0_out[1459] | layer0_out[1460]);
     layer1_out[10737] <= layer0_out[6751];
     layer1_out[10738] <= layer0_out[7627];
     layer1_out[10739] <= ~layer0_out[7838] | layer0_out[7837];
     layer1_out[10740] <= layer0_out[7303] | layer0_out[7304];
     layer1_out[10741] <= ~(layer0_out[1272] & layer0_out[1273]);
     layer1_out[10742] <= ~(layer0_out[3719] ^ layer0_out[3720]);
     layer1_out[10743] <= layer0_out[5194] & ~layer0_out[5195];
     layer1_out[10744] <= ~(layer0_out[3588] & layer0_out[3589]);
     layer1_out[10745] <= layer0_out[330] & ~layer0_out[331];
     layer1_out[10746] <= layer0_out[9776];
     layer1_out[10747] <= layer0_out[10114] & layer0_out[10115];
     layer1_out[10748] <= ~layer0_out[2364] | layer0_out[2365];
     layer1_out[10749] <= layer0_out[10255];
     layer1_out[10750] <= ~layer0_out[5982] | layer0_out[5983];
     layer1_out[10751] <= layer0_out[4890];
     layer1_out[10752] <= ~layer0_out[7017];
     layer1_out[10753] <= ~(layer0_out[6723] & layer0_out[6724]);
     layer1_out[10754] <= layer0_out[8247] | layer0_out[8248];
     layer1_out[10755] <= layer0_out[7534] & ~layer0_out[7533];
     layer1_out[10756] <= ~(layer0_out[4184] | layer0_out[4185]);
     layer1_out[10757] <= ~layer0_out[2372] | layer0_out[2371];
     layer1_out[10758] <= layer0_out[284] | layer0_out[285];
     layer1_out[10759] <= ~(layer0_out[6064] | layer0_out[6065]);
     layer1_out[10760] <= ~layer0_out[11620];
     layer1_out[10761] <= ~layer0_out[1438] | layer0_out[1439];
     layer1_out[10762] <= ~layer0_out[11956] | layer0_out[11955];
     layer1_out[10763] <= layer0_out[5494] ^ layer0_out[5495];
     layer1_out[10764] <= ~(layer0_out[7247] | layer0_out[7248]);
     layer1_out[10765] <= layer0_out[3708] ^ layer0_out[3709];
     layer1_out[10766] <= ~layer0_out[9950] | layer0_out[9949];
     layer1_out[10767] <= layer0_out[9809] & ~layer0_out[9808];
     layer1_out[10768] <= ~layer0_out[499] | layer0_out[500];
     layer1_out[10769] <= layer0_out[11062] | layer0_out[11063];
     layer1_out[10770] <= layer0_out[2742] & layer0_out[2743];
     layer1_out[10771] <= ~layer0_out[2091] | layer0_out[2090];
     layer1_out[10772] <= ~layer0_out[6600];
     layer1_out[10773] <= layer0_out[5896];
     layer1_out[10774] <= layer0_out[7911] & ~layer0_out[7910];
     layer1_out[10775] <= layer0_out[6964] | layer0_out[6965];
     layer1_out[10776] <= layer0_out[7026];
     layer1_out[10777] <= layer0_out[7273] & ~layer0_out[7272];
     layer1_out[10778] <= ~layer0_out[4758] | layer0_out[4757];
     layer1_out[10779] <= ~layer0_out[4444];
     layer1_out[10780] <= layer0_out[1506] | layer0_out[1507];
     layer1_out[10781] <= layer0_out[227] & layer0_out[228];
     layer1_out[10782] <= layer0_out[1291];
     layer1_out[10783] <= ~(layer0_out[8161] & layer0_out[8162]);
     layer1_out[10784] <= ~(layer0_out[4365] | layer0_out[4366]);
     layer1_out[10785] <= ~(layer0_out[807] & layer0_out[808]);
     layer1_out[10786] <= ~layer0_out[2745] | layer0_out[2746];
     layer1_out[10787] <= 1'b0;
     layer1_out[10788] <= layer0_out[11289] & layer0_out[11290];
     layer1_out[10789] <= layer0_out[3816];
     layer1_out[10790] <= layer0_out[2109] | layer0_out[2110];
     layer1_out[10791] <= layer0_out[7767];
     layer1_out[10792] <= layer0_out[4266] ^ layer0_out[4267];
     layer1_out[10793] <= layer0_out[8179];
     layer1_out[10794] <= ~layer0_out[9334];
     layer1_out[10795] <= ~layer0_out[2436] | layer0_out[2435];
     layer1_out[10796] <= layer0_out[8363] & ~layer0_out[8362];
     layer1_out[10797] <= ~(layer0_out[4128] | layer0_out[4129]);
     layer1_out[10798] <= layer0_out[9595] & ~layer0_out[9596];
     layer1_out[10799] <= layer0_out[10902] & ~layer0_out[10903];
     layer1_out[10800] <= ~layer0_out[5661];
     layer1_out[10801] <= ~(layer0_out[475] & layer0_out[476]);
     layer1_out[10802] <= layer0_out[6003] ^ layer0_out[6004];
     layer1_out[10803] <= layer0_out[3022] & layer0_out[3023];
     layer1_out[10804] <= layer0_out[8987];
     layer1_out[10805] <= ~layer0_out[2596] | layer0_out[2597];
     layer1_out[10806] <= layer0_out[7939] & ~layer0_out[7940];
     layer1_out[10807] <= layer0_out[240] & layer0_out[241];
     layer1_out[10808] <= ~layer0_out[10588] | layer0_out[10587];
     layer1_out[10809] <= 1'b1;
     layer1_out[10810] <= ~layer0_out[6444] | layer0_out[6445];
     layer1_out[10811] <= ~layer0_out[350] | layer0_out[349];
     layer1_out[10812] <= ~layer0_out[11703];
     layer1_out[10813] <= layer0_out[10971];
     layer1_out[10814] <= ~layer0_out[5270];
     layer1_out[10815] <= layer0_out[6109];
     layer1_out[10816] <= ~(layer0_out[11765] & layer0_out[11766]);
     layer1_out[10817] <= ~layer0_out[7926] | layer0_out[7925];
     layer1_out[10818] <= ~(layer0_out[10402] & layer0_out[10403]);
     layer1_out[10819] <= ~layer0_out[6925] | layer0_out[6924];
     layer1_out[10820] <= ~(layer0_out[2275] ^ layer0_out[2276]);
     layer1_out[10821] <= layer0_out[4175];
     layer1_out[10822] <= 1'b1;
     layer1_out[10823] <= 1'b0;
     layer1_out[10824] <= layer0_out[9522] & ~layer0_out[9523];
     layer1_out[10825] <= layer0_out[1853] & layer0_out[1854];
     layer1_out[10826] <= ~layer0_out[6092] | layer0_out[6091];
     layer1_out[10827] <= ~layer0_out[5526];
     layer1_out[10828] <= ~layer0_out[8541] | layer0_out[8542];
     layer1_out[10829] <= layer0_out[3529] | layer0_out[3530];
     layer1_out[10830] <= 1'b1;
     layer1_out[10831] <= layer0_out[10628];
     layer1_out[10832] <= layer0_out[11065];
     layer1_out[10833] <= layer0_out[11488];
     layer1_out[10834] <= ~(layer0_out[4536] | layer0_out[4537]);
     layer1_out[10835] <= layer0_out[6035];
     layer1_out[10836] <= ~layer0_out[9738] | layer0_out[9739];
     layer1_out[10837] <= ~layer0_out[10464] | layer0_out[10465];
     layer1_out[10838] <= layer0_out[9180];
     layer1_out[10839] <= layer0_out[6629] & ~layer0_out[6628];
     layer1_out[10840] <= ~layer0_out[1766];
     layer1_out[10841] <= layer0_out[11175] & ~layer0_out[11176];
     layer1_out[10842] <= layer0_out[1965] & ~layer0_out[1966];
     layer1_out[10843] <= ~layer0_out[22];
     layer1_out[10844] <= ~layer0_out[4805];
     layer1_out[10845] <= ~layer0_out[7728];
     layer1_out[10846] <= ~(layer0_out[4551] & layer0_out[4552]);
     layer1_out[10847] <= ~(layer0_out[1429] & layer0_out[1430]);
     layer1_out[10848] <= ~layer0_out[1083] | layer0_out[1082];
     layer1_out[10849] <= ~layer0_out[2407] | layer0_out[2406];
     layer1_out[10850] <= layer0_out[7];
     layer1_out[10851] <= layer0_out[2622] | layer0_out[2623];
     layer1_out[10852] <= layer0_out[4030];
     layer1_out[10853] <= ~(layer0_out[1684] & layer0_out[1685]);
     layer1_out[10854] <= layer0_out[2162] & ~layer0_out[2163];
     layer1_out[10855] <= ~(layer0_out[1392] & layer0_out[1393]);
     layer1_out[10856] <= ~layer0_out[3000] | layer0_out[3001];
     layer1_out[10857] <= layer0_out[5694] & layer0_out[5695];
     layer1_out[10858] <= layer0_out[7770];
     layer1_out[10859] <= layer0_out[8239] & ~layer0_out[8238];
     layer1_out[10860] <= layer0_out[4510];
     layer1_out[10861] <= layer0_out[5370];
     layer1_out[10862] <= layer0_out[9321];
     layer1_out[10863] <= layer0_out[7514] & layer0_out[7515];
     layer1_out[10864] <= layer0_out[8468] & ~layer0_out[8469];
     layer1_out[10865] <= ~(layer0_out[7080] ^ layer0_out[7081]);
     layer1_out[10866] <= layer0_out[7613] ^ layer0_out[7614];
     layer1_out[10867] <= layer0_out[4227];
     layer1_out[10868] <= layer0_out[2230] & ~layer0_out[2229];
     layer1_out[10869] <= ~layer0_out[5683];
     layer1_out[10870] <= layer0_out[9726] & layer0_out[9727];
     layer1_out[10871] <= ~(layer0_out[3984] | layer0_out[3985]);
     layer1_out[10872] <= ~layer0_out[53];
     layer1_out[10873] <= ~layer0_out[1244];
     layer1_out[10874] <= layer0_out[5249] & layer0_out[5250];
     layer1_out[10875] <= ~(layer0_out[2391] & layer0_out[2392]);
     layer1_out[10876] <= layer0_out[1314] & layer0_out[1315];
     layer1_out[10877] <= ~layer0_out[4143];
     layer1_out[10878] <= layer0_out[10319] & layer0_out[10320];
     layer1_out[10879] <= 1'b1;
     layer1_out[10880] <= layer0_out[1445] & ~layer0_out[1446];
     layer1_out[10881] <= layer0_out[4165] | layer0_out[4166];
     layer1_out[10882] <= 1'b1;
     layer1_out[10883] <= ~(layer0_out[7222] & layer0_out[7223]);
     layer1_out[10884] <= ~(layer0_out[6828] & layer0_out[6829]);
     layer1_out[10885] <= layer0_out[4344] & ~layer0_out[4343];
     layer1_out[10886] <= ~layer0_out[10503] | layer0_out[10504];
     layer1_out[10887] <= ~(layer0_out[1741] & layer0_out[1742]);
     layer1_out[10888] <= layer0_out[9880] & layer0_out[9881];
     layer1_out[10889] <= ~(layer0_out[10270] | layer0_out[10271]);
     layer1_out[10890] <= ~layer0_out[9357] | layer0_out[9356];
     layer1_out[10891] <= layer0_out[7598];
     layer1_out[10892] <= layer0_out[9293] ^ layer0_out[9294];
     layer1_out[10893] <= layer0_out[523];
     layer1_out[10894] <= layer0_out[2411] & ~layer0_out[2412];
     layer1_out[10895] <= ~layer0_out[1542] | layer0_out[1541];
     layer1_out[10896] <= ~layer0_out[6407] | layer0_out[6408];
     layer1_out[10897] <= ~layer0_out[5232];
     layer1_out[10898] <= ~layer0_out[6769];
     layer1_out[10899] <= ~layer0_out[3352] | layer0_out[3351];
     layer1_out[10900] <= layer0_out[5152];
     layer1_out[10901] <= layer0_out[4085] & ~layer0_out[4086];
     layer1_out[10902] <= ~layer0_out[1713] | layer0_out[1714];
     layer1_out[10903] <= ~(layer0_out[4735] | layer0_out[4736]);
     layer1_out[10904] <= ~(layer0_out[2866] & layer0_out[2867]);
     layer1_out[10905] <= ~(layer0_out[4061] & layer0_out[4062]);
     layer1_out[10906] <= ~layer0_out[6659];
     layer1_out[10907] <= layer0_out[547] | layer0_out[548];
     layer1_out[10908] <= ~layer0_out[9540];
     layer1_out[10909] <= layer0_out[10986] & layer0_out[10987];
     layer1_out[10910] <= ~(layer0_out[6392] | layer0_out[6393]);
     layer1_out[10911] <= layer0_out[202];
     layer1_out[10912] <= ~layer0_out[5403];
     layer1_out[10913] <= ~(layer0_out[10052] | layer0_out[10053]);
     layer1_out[10914] <= layer0_out[11566] | layer0_out[11567];
     layer1_out[10915] <= ~layer0_out[505];
     layer1_out[10916] <= ~layer0_out[3742];
     layer1_out[10917] <= layer0_out[2925] & layer0_out[2926];
     layer1_out[10918] <= ~layer0_out[5889];
     layer1_out[10919] <= layer0_out[10910] | layer0_out[10911];
     layer1_out[10920] <= ~(layer0_out[10390] & layer0_out[10391]);
     layer1_out[10921] <= layer0_out[11135] & ~layer0_out[11134];
     layer1_out[10922] <= layer0_out[11882] & layer0_out[11883];
     layer1_out[10923] <= ~(layer0_out[1011] & layer0_out[1012]);
     layer1_out[10924] <= layer0_out[11540];
     layer1_out[10925] <= 1'b1;
     layer1_out[10926] <= layer0_out[10793] & ~layer0_out[10792];
     layer1_out[10927] <= ~layer0_out[2304] | layer0_out[2305];
     layer1_out[10928] <= layer0_out[9199] & ~layer0_out[9200];
     layer1_out[10929] <= ~layer0_out[7975] | layer0_out[7976];
     layer1_out[10930] <= layer0_out[9986] & layer0_out[9987];
     layer1_out[10931] <= ~layer0_out[4010] | layer0_out[4011];
     layer1_out[10932] <= ~layer0_out[10516] | layer0_out[10517];
     layer1_out[10933] <= layer0_out[6562] ^ layer0_out[6563];
     layer1_out[10934] <= layer0_out[2835] | layer0_out[2836];
     layer1_out[10935] <= ~layer0_out[7610];
     layer1_out[10936] <= layer0_out[11395];
     layer1_out[10937] <= ~layer0_out[9299];
     layer1_out[10938] <= layer0_out[11109];
     layer1_out[10939] <= ~layer0_out[5011] | layer0_out[5012];
     layer1_out[10940] <= ~(layer0_out[11604] | layer0_out[11605]);
     layer1_out[10941] <= layer0_out[8651] & ~layer0_out[8652];
     layer1_out[10942] <= layer0_out[4855] & layer0_out[4856];
     layer1_out[10943] <= ~(layer0_out[8760] ^ layer0_out[8761]);
     layer1_out[10944] <= layer0_out[9190] & layer0_out[9191];
     layer1_out[10945] <= ~layer0_out[10740];
     layer1_out[10946] <= ~layer0_out[10885];
     layer1_out[10947] <= ~(layer0_out[4467] & layer0_out[4468]);
     layer1_out[10948] <= ~layer0_out[6523] | layer0_out[6524];
     layer1_out[10949] <= ~layer0_out[4809] | layer0_out[4808];
     layer1_out[10950] <= layer0_out[8552] & layer0_out[8553];
     layer1_out[10951] <= ~(layer0_out[5953] | layer0_out[5954]);
     layer1_out[10952] <= layer0_out[6281] & layer0_out[6282];
     layer1_out[10953] <= ~layer0_out[9630];
     layer1_out[10954] <= layer0_out[1979] & ~layer0_out[1980];
     layer1_out[10955] <= ~layer0_out[4373];
     layer1_out[10956] <= 1'b0;
     layer1_out[10957] <= ~(layer0_out[1499] & layer0_out[1500]);
     layer1_out[10958] <= ~layer0_out[5472] | layer0_out[5473];
     layer1_out[10959] <= ~layer0_out[7079];
     layer1_out[10960] <= layer0_out[5541];
     layer1_out[10961] <= ~layer0_out[3632];
     layer1_out[10962] <= layer0_out[3451];
     layer1_out[10963] <= layer0_out[2485];
     layer1_out[10964] <= ~(layer0_out[10425] | layer0_out[10426]);
     layer1_out[10965] <= ~layer0_out[5919] | layer0_out[5920];
     layer1_out[10966] <= ~layer0_out[9862];
     layer1_out[10967] <= layer0_out[8789] & ~layer0_out[8790];
     layer1_out[10968] <= ~layer0_out[274];
     layer1_out[10969] <= layer0_out[94];
     layer1_out[10970] <= layer0_out[10811];
     layer1_out[10971] <= ~(layer0_out[11067] | layer0_out[11068]);
     layer1_out[10972] <= ~(layer0_out[1152] | layer0_out[1153]);
     layer1_out[10973] <= layer0_out[4054] | layer0_out[4055];
     layer1_out[10974] <= ~layer0_out[6287] | layer0_out[6286];
     layer1_out[10975] <= layer0_out[1068];
     layer1_out[10976] <= layer0_out[1020] & ~layer0_out[1019];
     layer1_out[10977] <= ~layer0_out[467] | layer0_out[468];
     layer1_out[10978] <= ~layer0_out[8238];
     layer1_out[10979] <= layer0_out[11479] & ~layer0_out[11478];
     layer1_out[10980] <= ~layer0_out[3183];
     layer1_out[10981] <= layer0_out[3023] & layer0_out[3024];
     layer1_out[10982] <= ~(layer0_out[1148] | layer0_out[1149]);
     layer1_out[10983] <= ~layer0_out[9594] | layer0_out[9595];
     layer1_out[10984] <= layer0_out[8628] & ~layer0_out[8629];
     layer1_out[10985] <= ~layer0_out[11898];
     layer1_out[10986] <= layer0_out[4369] | layer0_out[4370];
     layer1_out[10987] <= layer0_out[3265] & ~layer0_out[3264];
     layer1_out[10988] <= layer0_out[8601] ^ layer0_out[8602];
     layer1_out[10989] <= layer0_out[4885] ^ layer0_out[4886];
     layer1_out[10990] <= layer0_out[9811] | layer0_out[9812];
     layer1_out[10991] <= layer0_out[9364] & ~layer0_out[9363];
     layer1_out[10992] <= ~(layer0_out[10568] | layer0_out[10569]);
     layer1_out[10993] <= layer0_out[9488];
     layer1_out[10994] <= 1'b0;
     layer1_out[10995] <= 1'b0;
     layer1_out[10996] <= layer0_out[6074];
     layer1_out[10997] <= layer0_out[11035] | layer0_out[11036];
     layer1_out[10998] <= ~(layer0_out[485] | layer0_out[486]);
     layer1_out[10999] <= layer0_out[3778] & layer0_out[3779];
     layer1_out[11000] <= layer0_out[4095];
     layer1_out[11001] <= 1'b0;
     layer1_out[11002] <= ~layer0_out[7625];
     layer1_out[11003] <= layer0_out[8012];
     layer1_out[11004] <= layer0_out[10] & layer0_out[11];
     layer1_out[11005] <= ~(layer0_out[11569] & layer0_out[11570]);
     layer1_out[11006] <= layer0_out[19] | layer0_out[20];
     layer1_out[11007] <= ~(layer0_out[10279] & layer0_out[10280]);
     layer1_out[11008] <= ~layer0_out[11037];
     layer1_out[11009] <= layer0_out[9479];
     layer1_out[11010] <= layer0_out[5539] | layer0_out[5540];
     layer1_out[11011] <= layer0_out[2800];
     layer1_out[11012] <= layer0_out[9274] & ~layer0_out[9273];
     layer1_out[11013] <= layer0_out[1911] & layer0_out[1912];
     layer1_out[11014] <= ~(layer0_out[1575] & layer0_out[1576]);
     layer1_out[11015] <= ~layer0_out[6266];
     layer1_out[11016] <= layer0_out[5573] & ~layer0_out[5572];
     layer1_out[11017] <= layer0_out[1583] & layer0_out[1584];
     layer1_out[11018] <= layer0_out[7877] & ~layer0_out[7878];
     layer1_out[11019] <= ~layer0_out[11809] | layer0_out[11810];
     layer1_out[11020] <= layer0_out[5781];
     layer1_out[11021] <= layer0_out[5699];
     layer1_out[11022] <= ~(layer0_out[2353] | layer0_out[2354]);
     layer1_out[11023] <= layer0_out[4874];
     layer1_out[11024] <= ~layer0_out[4649] | layer0_out[4650];
     layer1_out[11025] <= layer0_out[2427];
     layer1_out[11026] <= layer0_out[10416] ^ layer0_out[10417];
     layer1_out[11027] <= layer0_out[9623] & layer0_out[9624];
     layer1_out[11028] <= ~layer0_out[9580] | layer0_out[9581];
     layer1_out[11029] <= ~layer0_out[7912];
     layer1_out[11030] <= layer0_out[1289] & ~layer0_out[1288];
     layer1_out[11031] <= ~(layer0_out[3942] & layer0_out[3943]);
     layer1_out[11032] <= layer0_out[7693];
     layer1_out[11033] <= layer0_out[7998] & layer0_out[7999];
     layer1_out[11034] <= ~(layer0_out[11225] & layer0_out[11226]);
     layer1_out[11035] <= ~(layer0_out[3327] & layer0_out[3328]);
     layer1_out[11036] <= layer0_out[4776];
     layer1_out[11037] <= ~layer0_out[9787];
     layer1_out[11038] <= ~(layer0_out[3266] ^ layer0_out[3267]);
     layer1_out[11039] <= layer0_out[9603] & ~layer0_out[9602];
     layer1_out[11040] <= layer0_out[6674] | layer0_out[6675];
     layer1_out[11041] <= 1'b0;
     layer1_out[11042] <= layer0_out[393];
     layer1_out[11043] <= layer0_out[7627] & ~layer0_out[7628];
     layer1_out[11044] <= layer0_out[8493] & ~layer0_out[8492];
     layer1_out[11045] <= ~layer0_out[9813];
     layer1_out[11046] <= layer0_out[2175] | layer0_out[2176];
     layer1_out[11047] <= ~layer0_out[3511] | layer0_out[3512];
     layer1_out[11048] <= layer0_out[11277] & ~layer0_out[11278];
     layer1_out[11049] <= layer0_out[9070] ^ layer0_out[9071];
     layer1_out[11050] <= layer0_out[9643];
     layer1_out[11051] <= layer0_out[1622] & ~layer0_out[1623];
     layer1_out[11052] <= ~(layer0_out[9429] ^ layer0_out[9430]);
     layer1_out[11053] <= ~(layer0_out[6421] ^ layer0_out[6422]);
     layer1_out[11054] <= layer0_out[1374] & ~layer0_out[1375];
     layer1_out[11055] <= layer0_out[11691] & ~layer0_out[11690];
     layer1_out[11056] <= layer0_out[602] | layer0_out[603];
     layer1_out[11057] <= layer0_out[9329];
     layer1_out[11058] <= layer0_out[3566] & layer0_out[3567];
     layer1_out[11059] <= ~(layer0_out[6528] ^ layer0_out[6529]);
     layer1_out[11060] <= ~layer0_out[8414];
     layer1_out[11061] <= ~layer0_out[6604];
     layer1_out[11062] <= ~layer0_out[1114];
     layer1_out[11063] <= ~layer0_out[5087] | layer0_out[5086];
     layer1_out[11064] <= ~layer0_out[10623];
     layer1_out[11065] <= ~layer0_out[11857];
     layer1_out[11066] <= ~layer0_out[5997];
     layer1_out[11067] <= ~(layer0_out[5455] | layer0_out[5456]);
     layer1_out[11068] <= layer0_out[3930] | layer0_out[3931];
     layer1_out[11069] <= ~layer0_out[11686];
     layer1_out[11070] <= ~(layer0_out[1835] & layer0_out[1836]);
     layer1_out[11071] <= ~layer0_out[8278];
     layer1_out[11072] <= layer0_out[34];
     layer1_out[11073] <= ~layer0_out[4001];
     layer1_out[11074] <= layer0_out[10052];
     layer1_out[11075] <= ~layer0_out[8236];
     layer1_out[11076] <= ~(layer0_out[10881] & layer0_out[10882]);
     layer1_out[11077] <= layer0_out[1193] ^ layer0_out[1194];
     layer1_out[11078] <= ~(layer0_out[10386] | layer0_out[10387]);
     layer1_out[11079] <= ~layer0_out[2212];
     layer1_out[11080] <= ~layer0_out[4315] | layer0_out[4314];
     layer1_out[11081] <= ~layer0_out[292];
     layer1_out[11082] <= ~layer0_out[4383];
     layer1_out[11083] <= layer0_out[3719] & ~layer0_out[3718];
     layer1_out[11084] <= layer0_out[7678] & ~layer0_out[7677];
     layer1_out[11085] <= layer0_out[6169] & ~layer0_out[6170];
     layer1_out[11086] <= layer0_out[3521] & layer0_out[3522];
     layer1_out[11087] <= layer0_out[2586] & ~layer0_out[2585];
     layer1_out[11088] <= ~layer0_out[4419];
     layer1_out[11089] <= layer0_out[8470] | layer0_out[8471];
     layer1_out[11090] <= layer0_out[6039] | layer0_out[6040];
     layer1_out[11091] <= ~(layer0_out[8113] & layer0_out[8114]);
     layer1_out[11092] <= ~(layer0_out[726] | layer0_out[727]);
     layer1_out[11093] <= ~layer0_out[1150] | layer0_out[1151];
     layer1_out[11094] <= layer0_out[5787];
     layer1_out[11095] <= ~(layer0_out[1227] & layer0_out[1228]);
     layer1_out[11096] <= layer0_out[10993] | layer0_out[10994];
     layer1_out[11097] <= ~layer0_out[3426];
     layer1_out[11098] <= ~layer0_out[4756] | layer0_out[4755];
     layer1_out[11099] <= layer0_out[7767];
     layer1_out[11100] <= ~layer0_out[4617] | layer0_out[4616];
     layer1_out[11101] <= ~layer0_out[4158] | layer0_out[4159];
     layer1_out[11102] <= ~layer0_out[11916] | layer0_out[11917];
     layer1_out[11103] <= ~layer0_out[6787];
     layer1_out[11104] <= layer0_out[4665];
     layer1_out[11105] <= ~layer0_out[4431];
     layer1_out[11106] <= layer0_out[4220] & ~layer0_out[4219];
     layer1_out[11107] <= ~(layer0_out[8083] & layer0_out[8084]);
     layer1_out[11108] <= layer0_out[498];
     layer1_out[11109] <= layer0_out[11391];
     layer1_out[11110] <= layer0_out[10901] | layer0_out[10902];
     layer1_out[11111] <= 1'b0;
     layer1_out[11112] <= layer0_out[5025];
     layer1_out[11113] <= layer0_out[423] & ~layer0_out[422];
     layer1_out[11114] <= layer0_out[11704] & ~layer0_out[11705];
     layer1_out[11115] <= layer0_out[296] & layer0_out[297];
     layer1_out[11116] <= ~layer0_out[9874] | layer0_out[9873];
     layer1_out[11117] <= ~(layer0_out[2620] & layer0_out[2621]);
     layer1_out[11118] <= layer0_out[3848];
     layer1_out[11119] <= layer0_out[1185];
     layer1_out[11120] <= ~(layer0_out[6818] | layer0_out[6819]);
     layer1_out[11121] <= layer0_out[5007];
     layer1_out[11122] <= ~layer0_out[2076];
     layer1_out[11123] <= ~(layer0_out[9583] | layer0_out[9584]);
     layer1_out[11124] <= ~(layer0_out[11080] & layer0_out[11081]);
     layer1_out[11125] <= ~layer0_out[4512];
     layer1_out[11126] <= layer0_out[11279] | layer0_out[11280];
     layer1_out[11127] <= ~layer0_out[6196];
     layer1_out[11128] <= ~(layer0_out[2329] | layer0_out[2330]);
     layer1_out[11129] <= ~layer0_out[9725];
     layer1_out[11130] <= layer0_out[2855] & ~layer0_out[2856];
     layer1_out[11131] <= layer0_out[11349];
     layer1_out[11132] <= layer0_out[6350] & layer0_out[6351];
     layer1_out[11133] <= layer0_out[4194] & ~layer0_out[4195];
     layer1_out[11134] <= layer0_out[8864] & ~layer0_out[8865];
     layer1_out[11135] <= ~layer0_out[5933];
     layer1_out[11136] <= layer0_out[4224] ^ layer0_out[4225];
     layer1_out[11137] <= layer0_out[7427];
     layer1_out[11138] <= ~(layer0_out[4336] | layer0_out[4337]);
     layer1_out[11139] <= ~layer0_out[3467] | layer0_out[3468];
     layer1_out[11140] <= layer0_out[7596] & layer0_out[7597];
     layer1_out[11141] <= ~layer0_out[873] | layer0_out[874];
     layer1_out[11142] <= ~(layer0_out[9938] ^ layer0_out[9939]);
     layer1_out[11143] <= ~layer0_out[10655];
     layer1_out[11144] <= ~layer0_out[8066];
     layer1_out[11145] <= layer0_out[9734] & layer0_out[9735];
     layer1_out[11146] <= layer0_out[4846] & layer0_out[4847];
     layer1_out[11147] <= layer0_out[2502];
     layer1_out[11148] <= layer0_out[124];
     layer1_out[11149] <= layer0_out[10457];
     layer1_out[11150] <= 1'b1;
     layer1_out[11151] <= layer0_out[8893];
     layer1_out[11152] <= ~layer0_out[2456] | layer0_out[2455];
     layer1_out[11153] <= layer0_out[6857] & layer0_out[6858];
     layer1_out[11154] <= layer0_out[8321];
     layer1_out[11155] <= ~layer0_out[7833] | layer0_out[7832];
     layer1_out[11156] <= layer0_out[3297] | layer0_out[3298];
     layer1_out[11157] <= layer0_out[1588];
     layer1_out[11158] <= ~layer0_out[4734];
     layer1_out[11159] <= ~(layer0_out[771] | layer0_out[772]);
     layer1_out[11160] <= ~layer0_out[8242];
     layer1_out[11161] <= layer0_out[7741] | layer0_out[7742];
     layer1_out[11162] <= ~layer0_out[6506];
     layer1_out[11163] <= layer0_out[970] & ~layer0_out[971];
     layer1_out[11164] <= ~layer0_out[1550] | layer0_out[1549];
     layer1_out[11165] <= layer0_out[9458] ^ layer0_out[9459];
     layer1_out[11166] <= 1'b0;
     layer1_out[11167] <= layer0_out[10558] ^ layer0_out[10559];
     layer1_out[11168] <= layer0_out[4467] & ~layer0_out[4466];
     layer1_out[11169] <= layer0_out[3508];
     layer1_out[11170] <= layer0_out[6566];
     layer1_out[11171] <= layer0_out[10010];
     layer1_out[11172] <= ~layer0_out[2696];
     layer1_out[11173] <= ~layer0_out[1441];
     layer1_out[11174] <= ~layer0_out[2118];
     layer1_out[11175] <= ~layer0_out[10566];
     layer1_out[11176] <= layer0_out[10132] & layer0_out[10133];
     layer1_out[11177] <= ~(layer0_out[4775] & layer0_out[4776]);
     layer1_out[11178] <= ~(layer0_out[6654] ^ layer0_out[6655]);
     layer1_out[11179] <= ~layer0_out[7006];
     layer1_out[11180] <= ~layer0_out[7105] | layer0_out[7104];
     layer1_out[11181] <= layer0_out[340] | layer0_out[341];
     layer1_out[11182] <= ~(layer0_out[49] | layer0_out[50]);
     layer1_out[11183] <= layer0_out[5512];
     layer1_out[11184] <= layer0_out[4318] & layer0_out[4319];
     layer1_out[11185] <= 1'b1;
     layer1_out[11186] <= layer0_out[3327];
     layer1_out[11187] <= layer0_out[1846];
     layer1_out[11188] <= ~(layer0_out[10962] | layer0_out[10963]);
     layer1_out[11189] <= layer0_out[997];
     layer1_out[11190] <= ~(layer0_out[3954] & layer0_out[3955]);
     layer1_out[11191] <= ~(layer0_out[5480] | layer0_out[5481]);
     layer1_out[11192] <= ~layer0_out[1320];
     layer1_out[11193] <= layer0_out[10287] | layer0_out[10288];
     layer1_out[11194] <= 1'b1;
     layer1_out[11195] <= layer0_out[133] ^ layer0_out[134];
     layer1_out[11196] <= layer0_out[8257] & ~layer0_out[8256];
     layer1_out[11197] <= layer0_out[3644];
     layer1_out[11198] <= ~layer0_out[921] | layer0_out[922];
     layer1_out[11199] <= ~layer0_out[9132];
     layer1_out[11200] <= layer0_out[8575] & ~layer0_out[8574];
     layer1_out[11201] <= layer0_out[10495];
     layer1_out[11202] <= ~layer0_out[10598];
     layer1_out[11203] <= ~layer0_out[7583] | layer0_out[7582];
     layer1_out[11204] <= ~(layer0_out[6560] & layer0_out[6561]);
     layer1_out[11205] <= ~layer0_out[8030];
     layer1_out[11206] <= layer0_out[554];
     layer1_out[11207] <= ~(layer0_out[10927] | layer0_out[10928]);
     layer1_out[11208] <= ~layer0_out[7220];
     layer1_out[11209] <= ~layer0_out[4564] | layer0_out[4565];
     layer1_out[11210] <= ~(layer0_out[4743] & layer0_out[4744]);
     layer1_out[11211] <= layer0_out[11546] & ~layer0_out[11545];
     layer1_out[11212] <= ~layer0_out[7129];
     layer1_out[11213] <= ~layer0_out[4844];
     layer1_out[11214] <= layer0_out[6646];
     layer1_out[11215] <= ~layer0_out[636];
     layer1_out[11216] <= layer0_out[7416] ^ layer0_out[7417];
     layer1_out[11217] <= ~layer0_out[1001];
     layer1_out[11218] <= layer0_out[646] & layer0_out[647];
     layer1_out[11219] <= ~(layer0_out[7243] | layer0_out[7244]);
     layer1_out[11220] <= ~(layer0_out[10936] | layer0_out[10937]);
     layer1_out[11221] <= ~layer0_out[4993];
     layer1_out[11222] <= layer0_out[8337];
     layer1_out[11223] <= ~layer0_out[2345];
     layer1_out[11224] <= layer0_out[7280] | layer0_out[7281];
     layer1_out[11225] <= layer0_out[6213];
     layer1_out[11226] <= layer0_out[2487];
     layer1_out[11227] <= layer0_out[8991] & layer0_out[8992];
     layer1_out[11228] <= layer0_out[4212] ^ layer0_out[4213];
     layer1_out[11229] <= layer0_out[271] & ~layer0_out[270];
     layer1_out[11230] <= ~(layer0_out[4977] & layer0_out[4978]);
     layer1_out[11231] <= ~layer0_out[9671];
     layer1_out[11232] <= ~(layer0_out[7261] | layer0_out[7262]);
     layer1_out[11233] <= ~(layer0_out[7670] | layer0_out[7671]);
     layer1_out[11234] <= layer0_out[6358];
     layer1_out[11235] <= ~layer0_out[10002];
     layer1_out[11236] <= layer0_out[2444] & ~layer0_out[2445];
     layer1_out[11237] <= layer0_out[1874];
     layer1_out[11238] <= ~layer0_out[7530] | layer0_out[7531];
     layer1_out[11239] <= 1'b1;
     layer1_out[11240] <= layer0_out[11180];
     layer1_out[11241] <= ~layer0_out[9732] | layer0_out[9731];
     layer1_out[11242] <= ~(layer0_out[1560] | layer0_out[1561]);
     layer1_out[11243] <= 1'b0;
     layer1_out[11244] <= layer0_out[3955] ^ layer0_out[3956];
     layer1_out[11245] <= ~layer0_out[9366] | layer0_out[9367];
     layer1_out[11246] <= ~layer0_out[4375];
     layer1_out[11247] <= ~(layer0_out[8171] & layer0_out[8172]);
     layer1_out[11248] <= layer0_out[10712] & ~layer0_out[10711];
     layer1_out[11249] <= ~(layer0_out[4422] | layer0_out[4423]);
     layer1_out[11250] <= layer0_out[9598] ^ layer0_out[9599];
     layer1_out[11251] <= ~layer0_out[503];
     layer1_out[11252] <= layer0_out[8755];
     layer1_out[11253] <= ~(layer0_out[11492] | layer0_out[11493]);
     layer1_out[11254] <= ~layer0_out[1125] | layer0_out[1126];
     layer1_out[11255] <= ~layer0_out[5045];
     layer1_out[11256] <= layer0_out[180];
     layer1_out[11257] <= ~(layer0_out[10106] ^ layer0_out[10107]);
     layer1_out[11258] <= 1'b0;
     layer1_out[11259] <= ~layer0_out[9699] | layer0_out[9698];
     layer1_out[11260] <= layer0_out[4450] ^ layer0_out[4451];
     layer1_out[11261] <= layer0_out[220];
     layer1_out[11262] <= ~(layer0_out[1808] | layer0_out[1809]);
     layer1_out[11263] <= ~(layer0_out[4972] ^ layer0_out[4973]);
     layer1_out[11264] <= layer0_out[5238] & layer0_out[5239];
     layer1_out[11265] <= ~layer0_out[5852];
     layer1_out[11266] <= layer0_out[11210] & ~layer0_out[11211];
     layer1_out[11267] <= layer0_out[6638] & ~layer0_out[6639];
     layer1_out[11268] <= ~layer0_out[7323];
     layer1_out[11269] <= layer0_out[4823];
     layer1_out[11270] <= layer0_out[3706] | layer0_out[3707];
     layer1_out[11271] <= ~layer0_out[417] | layer0_out[416];
     layer1_out[11272] <= ~(layer0_out[177] | layer0_out[178]);
     layer1_out[11273] <= ~layer0_out[753];
     layer1_out[11274] <= layer0_out[1411];
     layer1_out[11275] <= layer0_out[7475];
     layer1_out[11276] <= layer0_out[327] | layer0_out[328];
     layer1_out[11277] <= layer0_out[5016];
     layer1_out[11278] <= layer0_out[3474] & layer0_out[3475];
     layer1_out[11279] <= layer0_out[1988] & layer0_out[1989];
     layer1_out[11280] <= layer0_out[710] & layer0_out[711];
     layer1_out[11281] <= ~layer0_out[10113];
     layer1_out[11282] <= ~layer0_out[11837];
     layer1_out[11283] <= layer0_out[6232];
     layer1_out[11284] <= ~layer0_out[4751];
     layer1_out[11285] <= layer0_out[435];
     layer1_out[11286] <= layer0_out[3432] ^ layer0_out[3433];
     layer1_out[11287] <= ~layer0_out[8329] | layer0_out[8330];
     layer1_out[11288] <= layer0_out[7908];
     layer1_out[11289] <= ~layer0_out[3925];
     layer1_out[11290] <= layer0_out[7203] | layer0_out[7204];
     layer1_out[11291] <= 1'b1;
     layer1_out[11292] <= ~layer0_out[4879] | layer0_out[4880];
     layer1_out[11293] <= ~(layer0_out[9076] & layer0_out[9077]);
     layer1_out[11294] <= ~layer0_out[1639];
     layer1_out[11295] <= layer0_out[4488] & layer0_out[4489];
     layer1_out[11296] <= layer0_out[3137] & ~layer0_out[3138];
     layer1_out[11297] <= layer0_out[2698] | layer0_out[2699];
     layer1_out[11298] <= ~(layer0_out[8322] & layer0_out[8323]);
     layer1_out[11299] <= ~layer0_out[678];
     layer1_out[11300] <= ~layer0_out[1698] | layer0_out[1697];
     layer1_out[11301] <= layer0_out[7181] & layer0_out[7182];
     layer1_out[11302] <= layer0_out[9825];
     layer1_out[11303] <= ~(layer0_out[2715] & layer0_out[2716]);
     layer1_out[11304] <= ~layer0_out[7532];
     layer1_out[11305] <= layer0_out[1570] ^ layer0_out[1571];
     layer1_out[11306] <= layer0_out[11590] & ~layer0_out[11591];
     layer1_out[11307] <= 1'b0;
     layer1_out[11308] <= layer0_out[1226] & layer0_out[1227];
     layer1_out[11309] <= ~layer0_out[2464] | layer0_out[2463];
     layer1_out[11310] <= ~layer0_out[11654];
     layer1_out[11311] <= layer0_out[2568] & ~layer0_out[2567];
     layer1_out[11312] <= ~layer0_out[1442];
     layer1_out[11313] <= ~layer0_out[2789];
     layer1_out[11314] <= layer0_out[6404] & layer0_out[6405];
     layer1_out[11315] <= layer0_out[4917];
     layer1_out[11316] <= layer0_out[1884];
     layer1_out[11317] <= ~layer0_out[6508];
     layer1_out[11318] <= layer0_out[7368] | layer0_out[7369];
     layer1_out[11319] <= ~layer0_out[7603];
     layer1_out[11320] <= ~(layer0_out[11149] ^ layer0_out[11150]);
     layer1_out[11321] <= layer0_out[2332] & ~layer0_out[2331];
     layer1_out[11322] <= ~layer0_out[7709] | layer0_out[7710];
     layer1_out[11323] <= layer0_out[11707] | layer0_out[11708];
     layer1_out[11324] <= ~(layer0_out[7668] & layer0_out[7669]);
     layer1_out[11325] <= ~(layer0_out[5328] & layer0_out[5329]);
     layer1_out[11326] <= ~(layer0_out[3606] | layer0_out[3607]);
     layer1_out[11327] <= ~layer0_out[6449];
     layer1_out[11328] <= layer0_out[4042];
     layer1_out[11329] <= layer0_out[79] & layer0_out[80];
     layer1_out[11330] <= ~layer0_out[2414];
     layer1_out[11331] <= ~(layer0_out[9287] | layer0_out[9288]);
     layer1_out[11332] <= ~layer0_out[8449] | layer0_out[8448];
     layer1_out[11333] <= layer0_out[7398] & ~layer0_out[7397];
     layer1_out[11334] <= ~layer0_out[2509];
     layer1_out[11335] <= layer0_out[2962] & ~layer0_out[2963];
     layer1_out[11336] <= layer0_out[5623] & ~layer0_out[5622];
     layer1_out[11337] <= ~(layer0_out[7301] ^ layer0_out[7302]);
     layer1_out[11338] <= ~layer0_out[3489];
     layer1_out[11339] <= ~(layer0_out[4498] | layer0_out[4499]);
     layer1_out[11340] <= ~(layer0_out[11628] | layer0_out[11629]);
     layer1_out[11341] <= ~layer0_out[2761];
     layer1_out[11342] <= ~layer0_out[10164];
     layer1_out[11343] <= layer0_out[7040];
     layer1_out[11344] <= ~layer0_out[3548] | layer0_out[3547];
     layer1_out[11345] <= layer0_out[4245] & ~layer0_out[4246];
     layer1_out[11346] <= layer0_out[7733];
     layer1_out[11347] <= layer0_out[1990];
     layer1_out[11348] <= layer0_out[1248] & layer0_out[1249];
     layer1_out[11349] <= ~layer0_out[2074] | layer0_out[2073];
     layer1_out[11350] <= layer0_out[10597] & layer0_out[10598];
     layer1_out[11351] <= ~layer0_out[3629] | layer0_out[3630];
     layer1_out[11352] <= layer0_out[5134];
     layer1_out[11353] <= layer0_out[1486] | layer0_out[1487];
     layer1_out[11354] <= layer0_out[854] & ~layer0_out[855];
     layer1_out[11355] <= ~(layer0_out[7055] ^ layer0_out[7056]);
     layer1_out[11356] <= layer0_out[8857] ^ layer0_out[8858];
     layer1_out[11357] <= ~(layer0_out[10136] & layer0_out[10137]);
     layer1_out[11358] <= layer0_out[2810];
     layer1_out[11359] <= layer0_out[10654];
     layer1_out[11360] <= 1'b1;
     layer1_out[11361] <= 1'b1;
     layer1_out[11362] <= ~(layer0_out[3743] & layer0_out[3744]);
     layer1_out[11363] <= ~layer0_out[6539];
     layer1_out[11364] <= layer0_out[11471];
     layer1_out[11365] <= ~layer0_out[5671] | layer0_out[5672];
     layer1_out[11366] <= 1'b0;
     layer1_out[11367] <= layer0_out[5791];
     layer1_out[11368] <= layer0_out[4292];
     layer1_out[11369] <= ~layer0_out[5416];
     layer1_out[11370] <= layer0_out[10801] & layer0_out[10802];
     layer1_out[11371] <= layer0_out[7569];
     layer1_out[11372] <= layer0_out[2167];
     layer1_out[11373] <= layer0_out[3543];
     layer1_out[11374] <= layer0_out[8046] | layer0_out[8047];
     layer1_out[11375] <= layer0_out[7086] & layer0_out[7087];
     layer1_out[11376] <= ~layer0_out[6669];
     layer1_out[11377] <= ~layer0_out[6038];
     layer1_out[11378] <= layer0_out[10918] | layer0_out[10919];
     layer1_out[11379] <= 1'b1;
     layer1_out[11380] <= layer0_out[10594];
     layer1_out[11381] <= layer0_out[5168];
     layer1_out[11382] <= 1'b0;
     layer1_out[11383] <= layer0_out[5556] & ~layer0_out[5555];
     layer1_out[11384] <= ~layer0_out[8842];
     layer1_out[11385] <= layer0_out[1723] ^ layer0_out[1724];
     layer1_out[11386] <= ~layer0_out[10839];
     layer1_out[11387] <= layer0_out[1829];
     layer1_out[11388] <= ~layer0_out[4291];
     layer1_out[11389] <= layer0_out[4110] & ~layer0_out[4109];
     layer1_out[11390] <= layer0_out[6492];
     layer1_out[11391] <= layer0_out[1900];
     layer1_out[11392] <= layer0_out[6191];
     layer1_out[11393] <= layer0_out[9606] | layer0_out[9607];
     layer1_out[11394] <= layer0_out[2909];
     layer1_out[11395] <= layer0_out[9319];
     layer1_out[11396] <= ~layer0_out[5971];
     layer1_out[11397] <= ~(layer0_out[944] ^ layer0_out[945]);
     layer1_out[11398] <= layer0_out[2829];
     layer1_out[11399] <= ~layer0_out[10098] | layer0_out[10099];
     layer1_out[11400] <= ~(layer0_out[7238] | layer0_out[7239]);
     layer1_out[11401] <= ~layer0_out[7648] | layer0_out[7649];
     layer1_out[11402] <= layer0_out[11222];
     layer1_out[11403] <= layer0_out[7020];
     layer1_out[11404] <= layer0_out[1177];
     layer1_out[11405] <= layer0_out[3059] & ~layer0_out[3058];
     layer1_out[11406] <= layer0_out[3831];
     layer1_out[11407] <= ~(layer0_out[174] & layer0_out[175]);
     layer1_out[11408] <= ~(layer0_out[7684] & layer0_out[7685]);
     layer1_out[11409] <= ~(layer0_out[4443] ^ layer0_out[4444]);
     layer1_out[11410] <= layer0_out[11944] & ~layer0_out[11945];
     layer1_out[11411] <= ~layer0_out[3828];
     layer1_out[11412] <= ~layer0_out[8117];
     layer1_out[11413] <= layer0_out[11138] ^ layer0_out[11139];
     layer1_out[11414] <= layer0_out[6852] & layer0_out[6853];
     layer1_out[11415] <= layer0_out[5388];
     layer1_out[11416] <= 1'b1;
     layer1_out[11417] <= ~(layer0_out[8285] & layer0_out[8286]);
     layer1_out[11418] <= ~layer0_out[5096];
     layer1_out[11419] <= layer0_out[4582] & ~layer0_out[4581];
     layer1_out[11420] <= ~layer0_out[1203];
     layer1_out[11421] <= ~(layer0_out[682] ^ layer0_out[683]);
     layer1_out[11422] <= 1'b0;
     layer1_out[11423] <= ~(layer0_out[9274] | layer0_out[9275]);
     layer1_out[11424] <= layer0_out[5535];
     layer1_out[11425] <= layer0_out[8757] & layer0_out[8758];
     layer1_out[11426] <= ~layer0_out[732];
     layer1_out[11427] <= ~layer0_out[7097];
     layer1_out[11428] <= layer0_out[9684] ^ layer0_out[9685];
     layer1_out[11429] <= ~(layer0_out[9736] & layer0_out[9737]);
     layer1_out[11430] <= ~layer0_out[8894] | layer0_out[8893];
     layer1_out[11431] <= ~layer0_out[2669] | layer0_out[2670];
     layer1_out[11432] <= layer0_out[10685] & ~layer0_out[10686];
     layer1_out[11433] <= ~(layer0_out[5374] | layer0_out[5375]);
     layer1_out[11434] <= layer0_out[2603] & ~layer0_out[2604];
     layer1_out[11435] <= ~layer0_out[184] | layer0_out[183];
     layer1_out[11436] <= ~layer0_out[6439] | layer0_out[6440];
     layer1_out[11437] <= ~layer0_out[11355];
     layer1_out[11438] <= 1'b0;
     layer1_out[11439] <= ~(layer0_out[6159] | layer0_out[6160]);
     layer1_out[11440] <= ~layer0_out[6749];
     layer1_out[11441] <= layer0_out[3180] | layer0_out[3181];
     layer1_out[11442] <= layer0_out[6683] & layer0_out[6684];
     layer1_out[11443] <= ~layer0_out[9414];
     layer1_out[11444] <= layer0_out[2606] & ~layer0_out[2605];
     layer1_out[11445] <= layer0_out[192] ^ layer0_out[193];
     layer1_out[11446] <= ~layer0_out[3823];
     layer1_out[11447] <= layer0_out[6944] & ~layer0_out[6945];
     layer1_out[11448] <= layer0_out[3815];
     layer1_out[11449] <= 1'b0;
     layer1_out[11450] <= layer0_out[10888];
     layer1_out[11451] <= layer0_out[3904] & layer0_out[3905];
     layer1_out[11452] <= layer0_out[7630] | layer0_out[7631];
     layer1_out[11453] <= ~layer0_out[1250] | layer0_out[1251];
     layer1_out[11454] <= layer0_out[7373];
     layer1_out[11455] <= layer0_out[7688];
     layer1_out[11456] <= ~(layer0_out[2708] & layer0_out[2709]);
     layer1_out[11457] <= ~layer0_out[5135];
     layer1_out[11458] <= layer0_out[6468] & layer0_out[6469];
     layer1_out[11459] <= layer0_out[6018];
     layer1_out[11460] <= 1'b0;
     layer1_out[11461] <= layer0_out[9044] ^ layer0_out[9045];
     layer1_out[11462] <= layer0_out[5900] | layer0_out[5901];
     layer1_out[11463] <= layer0_out[5800];
     layer1_out[11464] <= ~(layer0_out[7515] ^ layer0_out[7516]);
     layer1_out[11465] <= layer0_out[1967] & ~layer0_out[1968];
     layer1_out[11466] <= layer0_out[5657];
     layer1_out[11467] <= 1'b1;
     layer1_out[11468] <= ~layer0_out[2309];
     layer1_out[11469] <= ~layer0_out[4989];
     layer1_out[11470] <= layer0_out[11644] & ~layer0_out[11645];
     layer1_out[11471] <= ~layer0_out[6041] | layer0_out[6040];
     layer1_out[11472] <= layer0_out[2425];
     layer1_out[11473] <= ~layer0_out[1223];
     layer1_out[11474] <= ~layer0_out[255];
     layer1_out[11475] <= ~(layer0_out[3133] | layer0_out[3134]);
     layer1_out[11476] <= layer0_out[2358] & layer0_out[2359];
     layer1_out[11477] <= layer0_out[911] & layer0_out[912];
     layer1_out[11478] <= ~(layer0_out[5761] | layer0_out[5762]);
     layer1_out[11479] <= layer0_out[10439];
     layer1_out[11480] <= ~layer0_out[1382];
     layer1_out[11481] <= 1'b0;
     layer1_out[11482] <= ~layer0_out[8393] | layer0_out[8392];
     layer1_out[11483] <= ~layer0_out[763];
     layer1_out[11484] <= layer0_out[11730] & ~layer0_out[11729];
     layer1_out[11485] <= ~layer0_out[11041];
     layer1_out[11486] <= layer0_out[8291] & ~layer0_out[8290];
     layer1_out[11487] <= layer0_out[3639] & ~layer0_out[3638];
     layer1_out[11488] <= ~(layer0_out[6269] | layer0_out[6270]);
     layer1_out[11489] <= layer0_out[834] ^ layer0_out[835];
     layer1_out[11490] <= ~layer0_out[5253] | layer0_out[5252];
     layer1_out[11491] <= layer0_out[5561] & ~layer0_out[5560];
     layer1_out[11492] <= ~layer0_out[2383];
     layer1_out[11493] <= layer0_out[4050] ^ layer0_out[4051];
     layer1_out[11494] <= layer0_out[6474] & ~layer0_out[6473];
     layer1_out[11495] <= ~layer0_out[10894] | layer0_out[10893];
     layer1_out[11496] <= 1'b1;
     layer1_out[11497] <= ~layer0_out[1287] | layer0_out[1288];
     layer1_out[11498] <= ~layer0_out[8299] | layer0_out[8298];
     layer1_out[11499] <= layer0_out[1212];
     layer1_out[11500] <= layer0_out[3538] & layer0_out[3539];
     layer1_out[11501] <= ~(layer0_out[8084] & layer0_out[8085]);
     layer1_out[11502] <= 1'b0;
     layer1_out[11503] <= 1'b1;
     layer1_out[11504] <= ~(layer0_out[946] | layer0_out[947]);
     layer1_out[11505] <= layer0_out[9214];
     layer1_out[11506] <= layer0_out[8678] & layer0_out[8679];
     layer1_out[11507] <= layer0_out[3605] | layer0_out[3606];
     layer1_out[11508] <= layer0_out[4402] | layer0_out[4403];
     layer1_out[11509] <= layer0_out[11065] ^ layer0_out[11066];
     layer1_out[11510] <= layer0_out[6698];
     layer1_out[11511] <= ~layer0_out[11315];
     layer1_out[11512] <= ~(layer0_out[4971] | layer0_out[4972]);
     layer1_out[11513] <= layer0_out[11795] & ~layer0_out[11796];
     layer1_out[11514] <= layer0_out[10547] & layer0_out[10548];
     layer1_out[11515] <= layer0_out[9548] & ~layer0_out[9549];
     layer1_out[11516] <= ~(layer0_out[9028] | layer0_out[9029]);
     layer1_out[11517] <= layer0_out[5068];
     layer1_out[11518] <= layer0_out[844];
     layer1_out[11519] <= 1'b1;
     layer1_out[11520] <= ~layer0_out[105];
     layer1_out[11521] <= layer0_out[187];
     layer1_out[11522] <= layer0_out[4132];
     layer1_out[11523] <= layer0_out[4368];
     layer1_out[11524] <= ~layer0_out[6908];
     layer1_out[11525] <= ~layer0_out[5177];
     layer1_out[11526] <= layer0_out[10603] | layer0_out[10604];
     layer1_out[11527] <= ~(layer0_out[10320] & layer0_out[10321]);
     layer1_out[11528] <= ~layer0_out[4245];
     layer1_out[11529] <= ~layer0_out[9585] | layer0_out[9586];
     layer1_out[11530] <= layer0_out[6564] | layer0_out[6565];
     layer1_out[11531] <= ~(layer0_out[272] ^ layer0_out[273]);
     layer1_out[11532] <= layer0_out[4596] & ~layer0_out[4597];
     layer1_out[11533] <= layer0_out[9897];
     layer1_out[11534] <= ~layer0_out[590];
     layer1_out[11535] <= ~layer0_out[3800];
     layer1_out[11536] <= ~layer0_out[11251];
     layer1_out[11537] <= layer0_out[733] | layer0_out[734];
     layer1_out[11538] <= ~layer0_out[10290] | layer0_out[10291];
     layer1_out[11539] <= ~layer0_out[4171] | layer0_out[4170];
     layer1_out[11540] <= layer0_out[11662] & layer0_out[11663];
     layer1_out[11541] <= ~layer0_out[3171];
     layer1_out[11542] <= layer0_out[8289] ^ layer0_out[8290];
     layer1_out[11543] <= layer0_out[10242] & layer0_out[10243];
     layer1_out[11544] <= ~layer0_out[9276];
     layer1_out[11545] <= layer0_out[1850] ^ layer0_out[1851];
     layer1_out[11546] <= ~layer0_out[10775] | layer0_out[10774];
     layer1_out[11547] <= ~layer0_out[10726] | layer0_out[10727];
     layer1_out[11548] <= 1'b0;
     layer1_out[11549] <= ~layer0_out[2461] | layer0_out[2462];
     layer1_out[11550] <= layer0_out[540] & ~layer0_out[539];
     layer1_out[11551] <= layer0_out[8807];
     layer1_out[11552] <= ~layer0_out[6578] | layer0_out[6577];
     layer1_out[11553] <= layer0_out[1132];
     layer1_out[11554] <= layer0_out[9336] & ~layer0_out[9335];
     layer1_out[11555] <= ~layer0_out[5135] | layer0_out[5134];
     layer1_out[11556] <= layer0_out[8925];
     layer1_out[11557] <= layer0_out[7981];
     layer1_out[11558] <= 1'b1;
     layer1_out[11559] <= layer0_out[11911] & ~layer0_out[11912];
     layer1_out[11560] <= ~layer0_out[10716] | layer0_out[10715];
     layer1_out[11561] <= layer0_out[3973];
     layer1_out[11562] <= layer0_out[215] & ~layer0_out[214];
     layer1_out[11563] <= ~layer0_out[1481] | layer0_out[1482];
     layer1_out[11564] <= layer0_out[9414] & ~layer0_out[9413];
     layer1_out[11565] <= ~layer0_out[5003];
     layer1_out[11566] <= layer0_out[6573] & ~layer0_out[6574];
     layer1_out[11567] <= layer0_out[10528];
     layer1_out[11568] <= ~layer0_out[673];
     layer1_out[11569] <= ~layer0_out[8024];
     layer1_out[11570] <= layer0_out[8093] | layer0_out[8094];
     layer1_out[11571] <= ~(layer0_out[11417] ^ layer0_out[11418]);
     layer1_out[11572] <= layer0_out[4954];
     layer1_out[11573] <= layer0_out[11881] & ~layer0_out[11880];
     layer1_out[11574] <= ~layer0_out[10213];
     layer1_out[11575] <= layer0_out[4500];
     layer1_out[11576] <= layer0_out[1220];
     layer1_out[11577] <= ~layer0_out[7789];
     layer1_out[11578] <= layer0_out[4427] & layer0_out[4428];
     layer1_out[11579] <= layer0_out[921];
     layer1_out[11580] <= ~(layer0_out[1277] | layer0_out[1278]);
     layer1_out[11581] <= layer0_out[8908];
     layer1_out[11582] <= layer0_out[8702] | layer0_out[8703];
     layer1_out[11583] <= ~(layer0_out[9626] ^ layer0_out[9627]);
     layer1_out[11584] <= layer0_out[1246] | layer0_out[1247];
     layer1_out[11585] <= ~(layer0_out[5757] & layer0_out[5758]);
     layer1_out[11586] <= layer0_out[11776];
     layer1_out[11587] <= layer0_out[10929];
     layer1_out[11588] <= ~(layer0_out[362] & layer0_out[363]);
     layer1_out[11589] <= ~layer0_out[6100];
     layer1_out[11590] <= layer0_out[2164];
     layer1_out[11591] <= layer0_out[8421] & ~layer0_out[8420];
     layer1_out[11592] <= ~layer0_out[8085];
     layer1_out[11593] <= ~layer0_out[11495];
     layer1_out[11594] <= 1'b1;
     layer1_out[11595] <= layer0_out[7804] ^ layer0_out[7805];
     layer1_out[11596] <= layer0_out[4890];
     layer1_out[11597] <= 1'b1;
     layer1_out[11598] <= ~(layer0_out[9867] & layer0_out[9868]);
     layer1_out[11599] <= ~layer0_out[8923];
     layer1_out[11600] <= layer0_out[5095] & ~layer0_out[5096];
     layer1_out[11601] <= 1'b0;
     layer1_out[11602] <= layer0_out[1788];
     layer1_out[11603] <= ~(layer0_out[3583] | layer0_out[3584]);
     layer1_out[11604] <= ~layer0_out[782];
     layer1_out[11605] <= layer0_out[1472] & ~layer0_out[1473];
     layer1_out[11606] <= ~(layer0_out[11974] | layer0_out[11975]);
     layer1_out[11607] <= layer0_out[9407] & layer0_out[9408];
     layer1_out[11608] <= layer0_out[4508] | layer0_out[4509];
     layer1_out[11609] <= layer0_out[1526] & ~layer0_out[1527];
     layer1_out[11610] <= ~layer0_out[418];
     layer1_out[11611] <= layer0_out[7288] ^ layer0_out[7289];
     layer1_out[11612] <= ~layer0_out[3421];
     layer1_out[11613] <= ~(layer0_out[8745] | layer0_out[8746]);
     layer1_out[11614] <= ~layer0_out[4255];
     layer1_out[11615] <= layer0_out[9017] & ~layer0_out[9016];
     layer1_out[11616] <= layer0_out[6522];
     layer1_out[11617] <= layer0_out[1393] & ~layer0_out[1394];
     layer1_out[11618] <= ~(layer0_out[9308] & layer0_out[9309]);
     layer1_out[11619] <= layer0_out[7438] & layer0_out[7439];
     layer1_out[11620] <= ~(layer0_out[9575] | layer0_out[9576]);
     layer1_out[11621] <= ~layer0_out[10481] | layer0_out[10480];
     layer1_out[11622] <= ~(layer0_out[1229] | layer0_out[1230]);
     layer1_out[11623] <= layer0_out[6103];
     layer1_out[11624] <= ~(layer0_out[9549] & layer0_out[9550]);
     layer1_out[11625] <= layer0_out[8661] & ~layer0_out[8660];
     layer1_out[11626] <= layer0_out[2966] & layer0_out[2967];
     layer1_out[11627] <= ~layer0_out[8119] | layer0_out[8120];
     layer1_out[11628] <= layer0_out[10878];
     layer1_out[11629] <= ~layer0_out[7941];
     layer1_out[11630] <= layer0_out[8845];
     layer1_out[11631] <= layer0_out[4715] & ~layer0_out[4714];
     layer1_out[11632] <= layer0_out[1217] ^ layer0_out[1218];
     layer1_out[11633] <= ~(layer0_out[11502] & layer0_out[11503]);
     layer1_out[11634] <= layer0_out[11326];
     layer1_out[11635] <= layer0_out[8927] | layer0_out[8928];
     layer1_out[11636] <= ~layer0_out[8816];
     layer1_out[11637] <= ~layer0_out[11445];
     layer1_out[11638] <= layer0_out[8617] & ~layer0_out[8616];
     layer1_out[11639] <= ~layer0_out[5788];
     layer1_out[11640] <= ~layer0_out[1215];
     layer1_out[11641] <= layer0_out[9403];
     layer1_out[11642] <= layer0_out[8010] | layer0_out[8011];
     layer1_out[11643] <= ~layer0_out[10736];
     layer1_out[11644] <= layer0_out[2171];
     layer1_out[11645] <= ~layer0_out[3871] | layer0_out[3872];
     layer1_out[11646] <= layer0_out[7855];
     layer1_out[11647] <= layer0_out[2524] | layer0_out[2525];
     layer1_out[11648] <= layer0_out[4366];
     layer1_out[11649] <= layer0_out[9165] & layer0_out[9166];
     layer1_out[11650] <= ~layer0_out[3508];
     layer1_out[11651] <= layer0_out[3558];
     layer1_out[11652] <= ~(layer0_out[7578] ^ layer0_out[7579]);
     layer1_out[11653] <= ~(layer0_out[6238] ^ layer0_out[6239]);
     layer1_out[11654] <= ~layer0_out[7672] | layer0_out[7671];
     layer1_out[11655] <= ~layer0_out[7503] | layer0_out[7504];
     layer1_out[11656] <= 1'b1;
     layer1_out[11657] <= layer0_out[4271];
     layer1_out[11658] <= ~layer0_out[1802];
     layer1_out[11659] <= ~(layer0_out[7520] | layer0_out[7521]);
     layer1_out[11660] <= ~layer0_out[941] | layer0_out[942];
     layer1_out[11661] <= layer0_out[10289];
     layer1_out[11662] <= 1'b0;
     layer1_out[11663] <= ~layer0_out[9368];
     layer1_out[11664] <= layer0_out[4668];
     layer1_out[11665] <= ~layer0_out[6911];
     layer1_out[11666] <= layer0_out[8359] & layer0_out[8360];
     layer1_out[11667] <= layer0_out[6592];
     layer1_out[11668] <= ~(layer0_out[8592] ^ layer0_out[8593]);
     layer1_out[11669] <= layer0_out[1261];
     layer1_out[11670] <= ~(layer0_out[5736] & layer0_out[5737]);
     layer1_out[11671] <= layer0_out[102] & layer0_out[103];
     layer1_out[11672] <= layer0_out[2037] ^ layer0_out[2038];
     layer1_out[11673] <= layer0_out[11975] & layer0_out[11976];
     layer1_out[11674] <= ~(layer0_out[9926] & layer0_out[9927]);
     layer1_out[11675] <= ~(layer0_out[9592] | layer0_out[9593]);
     layer1_out[11676] <= ~layer0_out[7680] | layer0_out[7681];
     layer1_out[11677] <= layer0_out[9597];
     layer1_out[11678] <= ~(layer0_out[9757] & layer0_out[9758]);
     layer1_out[11679] <= ~(layer0_out[11137] ^ layer0_out[11138]);
     layer1_out[11680] <= ~layer0_out[2416];
     layer1_out[11681] <= layer0_out[10071];
     layer1_out[11682] <= ~layer0_out[688] | layer0_out[689];
     layer1_out[11683] <= ~(layer0_out[7328] | layer0_out[7329]);
     layer1_out[11684] <= layer0_out[3908] & ~layer0_out[3907];
     layer1_out[11685] <= layer0_out[4258] ^ layer0_out[4259];
     layer1_out[11686] <= ~layer0_out[9260];
     layer1_out[11687] <= ~layer0_out[8920] | layer0_out[8919];
     layer1_out[11688] <= ~layer0_out[229];
     layer1_out[11689] <= layer0_out[2141] & ~layer0_out[2142];
     layer1_out[11690] <= layer0_out[9280] ^ layer0_out[9281];
     layer1_out[11691] <= ~(layer0_out[2203] & layer0_out[2204]);
     layer1_out[11692] <= ~(layer0_out[6595] | layer0_out[6596]);
     layer1_out[11693] <= layer0_out[5092];
     layer1_out[11694] <= ~layer0_out[9247];
     layer1_out[11695] <= ~layer0_out[5600];
     layer1_out[11696] <= layer0_out[6047] & layer0_out[6048];
     layer1_out[11697] <= 1'b0;
     layer1_out[11698] <= ~(layer0_out[2812] & layer0_out[2813]);
     layer1_out[11699] <= ~layer0_out[10421] | layer0_out[10422];
     layer1_out[11700] <= layer0_out[8552];
     layer1_out[11701] <= ~(layer0_out[5005] ^ layer0_out[5006]);
     layer1_out[11702] <= ~(layer0_out[4104] & layer0_out[4105]);
     layer1_out[11703] <= ~layer0_out[6096];
     layer1_out[11704] <= ~layer0_out[3630];
     layer1_out[11705] <= layer0_out[5683] & layer0_out[5684];
     layer1_out[11706] <= layer0_out[5236] & ~layer0_out[5235];
     layer1_out[11707] <= layer0_out[10288] | layer0_out[10289];
     layer1_out[11708] <= layer0_out[10554];
     layer1_out[11709] <= ~(layer0_out[10897] ^ layer0_out[10898]);
     layer1_out[11710] <= ~layer0_out[5763];
     layer1_out[11711] <= layer0_out[3340] ^ layer0_out[3341];
     layer1_out[11712] <= ~(layer0_out[3314] & layer0_out[3315]);
     layer1_out[11713] <= ~(layer0_out[6477] & layer0_out[6478]);
     layer1_out[11714] <= ~layer0_out[3724];
     layer1_out[11715] <= layer0_out[642];
     layer1_out[11716] <= ~layer0_out[9160] | layer0_out[9161];
     layer1_out[11717] <= ~(layer0_out[9418] & layer0_out[9419]);
     layer1_out[11718] <= ~layer0_out[6036] | layer0_out[6037];
     layer1_out[11719] <= ~(layer0_out[7116] ^ layer0_out[7117]);
     layer1_out[11720] <= ~(layer0_out[3812] & layer0_out[3813]);
     layer1_out[11721] <= layer0_out[5350];
     layer1_out[11722] <= ~layer0_out[5858] | layer0_out[5857];
     layer1_out[11723] <= layer0_out[4815] & layer0_out[4816];
     layer1_out[11724] <= ~(layer0_out[5654] | layer0_out[5655]);
     layer1_out[11725] <= layer0_out[8898] & ~layer0_out[8897];
     layer1_out[11726] <= layer0_out[2078] & layer0_out[2079];
     layer1_out[11727] <= layer0_out[5154];
     layer1_out[11728] <= ~(layer0_out[3044] & layer0_out[3045]);
     layer1_out[11729] <= ~layer0_out[10089] | layer0_out[10088];
     layer1_out[11730] <= 1'b0;
     layer1_out[11731] <= ~layer0_out[815];
     layer1_out[11732] <= ~layer0_out[25] | layer0_out[24];
     layer1_out[11733] <= layer0_out[11404] | layer0_out[11405];
     layer1_out[11734] <= layer0_out[1137] | layer0_out[1138];
     layer1_out[11735] <= layer0_out[1643] & ~layer0_out[1642];
     layer1_out[11736] <= ~layer0_out[4180];
     layer1_out[11737] <= ~layer0_out[7044] | layer0_out[7045];
     layer1_out[11738] <= ~(layer0_out[5022] | layer0_out[5023]);
     layer1_out[11739] <= layer0_out[2815];
     layer1_out[11740] <= layer0_out[3026] & ~layer0_out[3027];
     layer1_out[11741] <= ~(layer0_out[10714] & layer0_out[10715]);
     layer1_out[11742] <= ~(layer0_out[2856] | layer0_out[2857]);
     layer1_out[11743] <= ~layer0_out[2783] | layer0_out[2782];
     layer1_out[11744] <= layer0_out[4985] ^ layer0_out[4986];
     layer1_out[11745] <= layer0_out[2569];
     layer1_out[11746] <= layer0_out[10911] | layer0_out[10912];
     layer1_out[11747] <= ~layer0_out[2737] | layer0_out[2738];
     layer1_out[11748] <= ~layer0_out[8230] | layer0_out[8231];
     layer1_out[11749] <= ~layer0_out[6551] | layer0_out[6552];
     layer1_out[11750] <= layer0_out[3762];
     layer1_out[11751] <= layer0_out[7414];
     layer1_out[11752] <= ~layer0_out[1305];
     layer1_out[11753] <= layer0_out[10833] | layer0_out[10834];
     layer1_out[11754] <= layer0_out[4214] & ~layer0_out[4213];
     layer1_out[11755] <= ~layer0_out[9432] | layer0_out[9431];
     layer1_out[11756] <= ~(layer0_out[5497] | layer0_out[5498]);
     layer1_out[11757] <= layer0_out[933] & ~layer0_out[934];
     layer1_out[11758] <= layer0_out[2814];
     layer1_out[11759] <= ~(layer0_out[5566] | layer0_out[5567]);
     layer1_out[11760] <= ~layer0_out[6208] | layer0_out[6207];
     layer1_out[11761] <= ~layer0_out[1007] | layer0_out[1006];
     layer1_out[11762] <= ~(layer0_out[8666] ^ layer0_out[8667]);
     layer1_out[11763] <= layer0_out[4693];
     layer1_out[11764] <= ~layer0_out[8606];
     layer1_out[11765] <= ~layer0_out[5517];
     layer1_out[11766] <= ~(layer0_out[1950] & layer0_out[1951]);
     layer1_out[11767] <= ~layer0_out[3588] | layer0_out[3587];
     layer1_out[11768] <= layer0_out[5854];
     layer1_out[11769] <= layer0_out[11659];
     layer1_out[11770] <= layer0_out[185] | layer0_out[186];
     layer1_out[11771] <= ~layer0_out[5534];
     layer1_out[11772] <= ~layer0_out[4947];
     layer1_out[11773] <= layer0_out[2215] & layer0_out[2216];
     layer1_out[11774] <= ~layer0_out[1850] | layer0_out[1849];
     layer1_out[11775] <= layer0_out[510] & ~layer0_out[509];
     layer1_out[11776] <= ~layer0_out[6611];
     layer1_out[11777] <= layer0_out[11570] & ~layer0_out[11571];
     layer1_out[11778] <= ~(layer0_out[6585] & layer0_out[6586]);
     layer1_out[11779] <= layer0_out[9446];
     layer1_out[11780] <= layer0_out[6970];
     layer1_out[11781] <= layer0_out[2101];
     layer1_out[11782] <= ~(layer0_out[4230] & layer0_out[4231]);
     layer1_out[11783] <= layer0_out[9643] & ~layer0_out[9642];
     layer1_out[11784] <= ~layer0_out[6940] | layer0_out[6941];
     layer1_out[11785] <= layer0_out[4140] & ~layer0_out[4139];
     layer1_out[11786] <= ~layer0_out[6309] | layer0_out[6310];
     layer1_out[11787] <= layer0_out[0];
     layer1_out[11788] <= ~layer0_out[10070] | layer0_out[10071];
     layer1_out[11789] <= ~layer0_out[2351];
     layer1_out[11790] <= layer0_out[10355] & ~layer0_out[10356];
     layer1_out[11791] <= layer0_out[11587];
     layer1_out[11792] <= layer0_out[798] & layer0_out[799];
     layer1_out[11793] <= ~layer0_out[10627] | layer0_out[10626];
     layer1_out[11794] <= layer0_out[1304] ^ layer0_out[1305];
     layer1_out[11795] <= layer0_out[10151] ^ layer0_out[10152];
     layer1_out[11796] <= layer0_out[11219] & ~layer0_out[11220];
     layer1_out[11797] <= layer0_out[4317];
     layer1_out[11798] <= layer0_out[4280];
     layer1_out[11799] <= layer0_out[2019] ^ layer0_out[2020];
     layer1_out[11800] <= ~layer0_out[4751] | layer0_out[4752];
     layer1_out[11801] <= layer0_out[11638];
     layer1_out[11802] <= layer0_out[2414] & ~layer0_out[2413];
     layer1_out[11803] <= layer0_out[4053] | layer0_out[4054];
     layer1_out[11804] <= ~layer0_out[10868] | layer0_out[10869];
     layer1_out[11805] <= layer0_out[983] & layer0_out[984];
     layer1_out[11806] <= ~layer0_out[9865];
     layer1_out[11807] <= ~layer0_out[11078];
     layer1_out[11808] <= layer0_out[11328];
     layer1_out[11809] <= layer0_out[4315] & ~layer0_out[4316];
     layer1_out[11810] <= ~layer0_out[10459];
     layer1_out[11811] <= ~layer0_out[3181];
     layer1_out[11812] <= layer0_out[3008] & ~layer0_out[3009];
     layer1_out[11813] <= layer0_out[8959];
     layer1_out[11814] <= ~layer0_out[4112] | layer0_out[4113];
     layer1_out[11815] <= layer0_out[9065];
     layer1_out[11816] <= layer0_out[3122];
     layer1_out[11817] <= ~(layer0_out[257] | layer0_out[258]);
     layer1_out[11818] <= ~(layer0_out[9640] & layer0_out[9641]);
     layer1_out[11819] <= ~layer0_out[5267];
     layer1_out[11820] <= ~layer0_out[10029];
     layer1_out[11821] <= ~layer0_out[3738] | layer0_out[3739];
     layer1_out[11822] <= ~layer0_out[11007];
     layer1_out[11823] <= layer0_out[10144] | layer0_out[10145];
     layer1_out[11824] <= layer0_out[6740] | layer0_out[6741];
     layer1_out[11825] <= layer0_out[8251];
     layer1_out[11826] <= layer0_out[2212] | layer0_out[2213];
     layer1_out[11827] <= ~layer0_out[2725];
     layer1_out[11828] <= ~layer0_out[1696] | layer0_out[1697];
     layer1_out[11829] <= layer0_out[7583] & layer0_out[7584];
     layer1_out[11830] <= layer0_out[6014] | layer0_out[6015];
     layer1_out[11831] <= ~layer0_out[7127];
     layer1_out[11832] <= ~(layer0_out[8388] ^ layer0_out[8389]);
     layer1_out[11833] <= ~layer0_out[7019];
     layer1_out[11834] <= layer0_out[460] & ~layer0_out[461];
     layer1_out[11835] <= 1'b0;
     layer1_out[11836] <= ~layer0_out[9970];
     layer1_out[11837] <= layer0_out[11531];
     layer1_out[11838] <= ~(layer0_out[11894] ^ layer0_out[11895]);
     layer1_out[11839] <= layer0_out[8761];
     layer1_out[11840] <= ~(layer0_out[8813] | layer0_out[8814]);
     layer1_out[11841] <= layer0_out[680] | layer0_out[681];
     layer1_out[11842] <= ~layer0_out[8096];
     layer1_out[11843] <= 1'b0;
     layer1_out[11844] <= ~layer0_out[2908];
     layer1_out[11845] <= layer0_out[11077] | layer0_out[11078];
     layer1_out[11846] <= ~layer0_out[1610] | layer0_out[1611];
     layer1_out[11847] <= layer0_out[6178];
     layer1_out[11848] <= layer0_out[3011] & layer0_out[3012];
     layer1_out[11849] <= ~layer0_out[4155];
     layer1_out[11850] <= ~(layer0_out[7691] ^ layer0_out[7692]);
     layer1_out[11851] <= layer0_out[9486];
     layer1_out[11852] <= layer0_out[9292] | layer0_out[9293];
     layer1_out[11853] <= layer0_out[7807] | layer0_out[7808];
     layer1_out[11854] <= ~(layer0_out[11917] ^ layer0_out[11918]);
     layer1_out[11855] <= ~layer0_out[10399] | layer0_out[10400];
     layer1_out[11856] <= layer0_out[9106] & ~layer0_out[9107];
     layer1_out[11857] <= ~(layer0_out[229] | layer0_out[230]);
     layer1_out[11858] <= layer0_out[1424] | layer0_out[1425];
     layer1_out[11859] <= layer0_out[7305] & layer0_out[7306];
     layer1_out[11860] <= ~layer0_out[7813];
     layer1_out[11861] <= ~layer0_out[268];
     layer1_out[11862] <= ~layer0_out[2227];
     layer1_out[11863] <= ~layer0_out[10977];
     layer1_out[11864] <= ~layer0_out[47] | layer0_out[48];
     layer1_out[11865] <= layer0_out[9605] & ~layer0_out[9604];
     layer1_out[11866] <= layer0_out[8991];
     layer1_out[11867] <= layer0_out[2662] & ~layer0_out[2661];
     layer1_out[11868] <= layer0_out[7134];
     layer1_out[11869] <= layer0_out[3777] & layer0_out[3778];
     layer1_out[11870] <= ~layer0_out[4817];
     layer1_out[11871] <= layer0_out[10622] ^ layer0_out[10623];
     layer1_out[11872] <= layer0_out[5093] & layer0_out[5094];
     layer1_out[11873] <= 1'b1;
     layer1_out[11874] <= ~layer0_out[5172];
     layer1_out[11875] <= layer0_out[7397] & ~layer0_out[7396];
     layer1_out[11876] <= ~(layer0_out[5297] & layer0_out[5298]);
     layer1_out[11877] <= layer0_out[6549];
     layer1_out[11878] <= layer0_out[3437] & ~layer0_out[3436];
     layer1_out[11879] <= ~(layer0_out[10146] | layer0_out[10147]);
     layer1_out[11880] <= ~layer0_out[2948] | layer0_out[2949];
     layer1_out[11881] <= ~layer0_out[345] | layer0_out[344];
     layer1_out[11882] <= ~(layer0_out[10110] & layer0_out[10111]);
     layer1_out[11883] <= layer0_out[8317] & ~layer0_out[8318];
     layer1_out[11884] <= layer0_out[1163];
     layer1_out[11885] <= ~layer0_out[2089] | layer0_out[2088];
     layer1_out[11886] <= ~(layer0_out[11979] ^ layer0_out[11980]);
     layer1_out[11887] <= ~layer0_out[7863];
     layer1_out[11888] <= layer0_out[10278];
     layer1_out[11889] <= layer0_out[11957] & layer0_out[11958];
     layer1_out[11890] <= layer0_out[805] & layer0_out[806];
     layer1_out[11891] <= layer0_out[5858];
     layer1_out[11892] <= ~layer0_out[10484];
     layer1_out[11893] <= ~layer0_out[9710];
     layer1_out[11894] <= 1'b1;
     layer1_out[11895] <= layer0_out[7897];
     layer1_out[11896] <= layer0_out[8466];
     layer1_out[11897] <= ~layer0_out[8781];
     layer1_out[11898] <= layer0_out[6288];
     layer1_out[11899] <= ~layer0_out[9948];
     layer1_out[11900] <= layer0_out[3308] & ~layer0_out[3309];
     layer1_out[11901] <= ~layer0_out[11923];
     layer1_out[11902] <= layer0_out[4646] & ~layer0_out[4647];
     layer1_out[11903] <= ~(layer0_out[8309] | layer0_out[8310]);
     layer1_out[11904] <= layer0_out[224] & ~layer0_out[225];
     layer1_out[11905] <= layer0_out[7892] & ~layer0_out[7893];
     layer1_out[11906] <= layer0_out[1731] | layer0_out[1732];
     layer1_out[11907] <= ~(layer0_out[10182] & layer0_out[10183]);
     layer1_out[11908] <= ~layer0_out[5372];
     layer1_out[11909] <= layer0_out[6836];
     layer1_out[11910] <= ~layer0_out[5307] | layer0_out[5306];
     layer1_out[11911] <= layer0_out[5495] & layer0_out[5496];
     layer1_out[11912] <= ~(layer0_out[98] | layer0_out[99]);
     layer1_out[11913] <= 1'b0;
     layer1_out[11914] <= layer0_out[7404] | layer0_out[7405];
     layer1_out[11915] <= ~(layer0_out[10972] | layer0_out[10973]);
     layer1_out[11916] <= ~layer0_out[4647] | layer0_out[4648];
     layer1_out[11917] <= layer0_out[10491];
     layer1_out[11918] <= layer0_out[10059];
     layer1_out[11919] <= layer0_out[2824];
     layer1_out[11920] <= layer0_out[4123] | layer0_out[4124];
     layer1_out[11921] <= layer0_out[8924] & layer0_out[8925];
     layer1_out[11922] <= layer0_out[2919] | layer0_out[2920];
     layer1_out[11923] <= ~layer0_out[384] | layer0_out[385];
     layer1_out[11924] <= ~layer0_out[10262] | layer0_out[10263];
     layer1_out[11925] <= layer0_out[3568] & ~layer0_out[3567];
     layer1_out[11926] <= ~layer0_out[10831];
     layer1_out[11927] <= ~layer0_out[4332] | layer0_out[4333];
     layer1_out[11928] <= layer0_out[10672] | layer0_out[10673];
     layer1_out[11929] <= ~layer0_out[1652] | layer0_out[1651];
     layer1_out[11930] <= ~(layer0_out[4350] ^ layer0_out[4351]);
     layer1_out[11931] <= ~layer0_out[6248];
     layer1_out[11932] <= ~layer0_out[2981] | layer0_out[2980];
     layer1_out[11933] <= layer0_out[11480] & ~layer0_out[11481];
     layer1_out[11934] <= layer0_out[4207];
     layer1_out[11935] <= ~layer0_out[735];
     layer1_out[11936] <= layer0_out[2702];
     layer1_out[11937] <= layer0_out[11160] & ~layer0_out[11159];
     layer1_out[11938] <= layer0_out[4602] & ~layer0_out[4603];
     layer1_out[11939] <= layer0_out[6694] & ~layer0_out[6695];
     layer1_out[11940] <= layer0_out[10806] & ~layer0_out[10807];
     layer1_out[11941] <= ~layer0_out[7012];
     layer1_out[11942] <= layer0_out[7900] & layer0_out[7901];
     layer1_out[11943] <= layer0_out[4820] | layer0_out[4821];
     layer1_out[11944] <= layer0_out[8622] ^ layer0_out[8623];
     layer1_out[11945] <= layer0_out[9149];
     layer1_out[11946] <= ~layer0_out[4154] | layer0_out[4155];
     layer1_out[11947] <= layer0_out[11967];
     layer1_out[11948] <= layer0_out[2705];
     layer1_out[11949] <= ~(layer0_out[10450] ^ layer0_out[10451]);
     layer1_out[11950] <= 1'b1;
     layer1_out[11951] <= ~layer0_out[10337];
     layer1_out[11952] <= ~layer0_out[6214] | layer0_out[6215];
     layer1_out[11953] <= layer0_out[4562] & ~layer0_out[4563];
     layer1_out[11954] <= ~(layer0_out[8886] ^ layer0_out[8887]);
     layer1_out[11955] <= layer0_out[6315] ^ layer0_out[6316];
     layer1_out[11956] <= layer0_out[1602] | layer0_out[1603];
     layer1_out[11957] <= layer0_out[10862] ^ layer0_out[10863];
     layer1_out[11958] <= layer0_out[2280];
     layer1_out[11959] <= ~layer0_out[8176];
     layer1_out[11960] <= ~layer0_out[5276];
     layer1_out[11961] <= ~(layer0_out[2600] ^ layer0_out[2601]);
     layer1_out[11962] <= ~(layer0_out[9959] | layer0_out[9960]);
     layer1_out[11963] <= ~layer0_out[9450];
     layer1_out[11964] <= 1'b0;
     layer1_out[11965] <= ~layer0_out[3844];
     layer1_out[11966] <= layer0_out[3785];
     layer1_out[11967] <= ~layer0_out[4249] | layer0_out[4248];
     layer1_out[11968] <= ~layer0_out[6859];
     layer1_out[11969] <= ~layer0_out[4980] | layer0_out[4981];
     layer1_out[11970] <= ~(layer0_out[5967] & layer0_out[5968]);
     layer1_out[11971] <= layer0_out[10519] & ~layer0_out[10518];
     layer1_out[11972] <= ~layer0_out[137];
     layer1_out[11973] <= ~layer0_out[4020];
     layer1_out[11974] <= layer0_out[9328];
     layer1_out[11975] <= ~layer0_out[376];
     layer1_out[11976] <= ~layer0_out[10148] | layer0_out[10149];
     layer1_out[11977] <= ~layer0_out[4470];
     layer1_out[11978] <= ~(layer0_out[4768] | layer0_out[4769]);
     layer1_out[11979] <= ~layer0_out[7014] | layer0_out[7013];
     layer1_out[11980] <= layer0_out[8799] | layer0_out[8800];
     layer1_out[11981] <= ~layer0_out[4534] | layer0_out[4533];
     layer1_out[11982] <= ~(layer0_out[9706] ^ layer0_out[9707]);
     layer1_out[11983] <= ~(layer0_out[9046] ^ layer0_out[9047]);
     layer1_out[11984] <= ~layer0_out[6280];
     layer1_out[11985] <= layer0_out[5222] & ~layer0_out[5221];
     layer1_out[11986] <= layer0_out[11207] & layer0_out[11208];
     layer1_out[11987] <= layer0_out[4546] & ~layer0_out[4547];
     layer1_out[11988] <= 1'b0;
     layer1_out[11989] <= ~layer0_out[10534] | layer0_out[10535];
     layer1_out[11990] <= layer0_out[4706];
     layer1_out[11991] <= ~layer0_out[2143] | layer0_out[2142];
     layer1_out[11992] <= layer0_out[1627];
     layer1_out[11993] <= ~layer0_out[1464];
     layer1_out[11994] <= ~layer0_out[8045];
     layer1_out[11995] <= layer0_out[5504] & layer0_out[5505];
     layer1_out[11996] <= layer0_out[9201] & ~layer0_out[9202];
     layer1_out[11997] <= ~layer0_out[1524] | layer0_out[1523];
     layer1_out[11998] <= ~layer0_out[6737];
     layer1_out[11999] <= layer0_out[8684] & ~layer0_out[8683];
     layer2_out[0] <= ~(layer1_out[6307] ^ layer1_out[6308]);
     layer2_out[1] <= layer1_out[3669];
     layer2_out[2] <= ~layer1_out[3752];
     layer2_out[3] <= layer1_out[1597] & ~layer1_out[1598];
     layer2_out[4] <= layer1_out[3984];
     layer2_out[5] <= layer1_out[1590];
     layer2_out[6] <= layer1_out[4017] & ~layer1_out[4018];
     layer2_out[7] <= layer1_out[11424] & layer1_out[11425];
     layer2_out[8] <= ~(layer1_out[8480] | layer1_out[8481]);
     layer2_out[9] <= layer1_out[2389];
     layer2_out[10] <= ~(layer1_out[11519] & layer1_out[11520]);
     layer2_out[11] <= ~layer1_out[495] | layer1_out[496];
     layer2_out[12] <= 1'b0;
     layer2_out[13] <= layer1_out[3024];
     layer2_out[14] <= ~layer1_out[4859];
     layer2_out[15] <= layer1_out[4794] & layer1_out[4795];
     layer2_out[16] <= ~(layer1_out[6530] & layer1_out[6531]);
     layer2_out[17] <= ~layer1_out[10469] | layer1_out[10468];
     layer2_out[18] <= layer1_out[6892] ^ layer1_out[6893];
     layer2_out[19] <= layer1_out[9993] & layer1_out[9994];
     layer2_out[20] <= ~layer1_out[7579] | layer1_out[7578];
     layer2_out[21] <= layer1_out[3351] & ~layer1_out[3350];
     layer2_out[22] <= layer1_out[11447] & layer1_out[11448];
     layer2_out[23] <= layer1_out[7400] | layer1_out[7401];
     layer2_out[24] <= ~(layer1_out[6953] & layer1_out[6954]);
     layer2_out[25] <= layer1_out[419];
     layer2_out[26] <= ~layer1_out[8009] | layer1_out[8008];
     layer2_out[27] <= ~layer1_out[6252] | layer1_out[6253];
     layer2_out[28] <= layer1_out[10788] | layer1_out[10789];
     layer2_out[29] <= ~(layer1_out[7600] | layer1_out[7601]);
     layer2_out[30] <= layer1_out[273] & layer1_out[274];
     layer2_out[31] <= layer1_out[5864];
     layer2_out[32] <= layer1_out[689];
     layer2_out[33] <= ~layer1_out[9257];
     layer2_out[34] <= layer1_out[3970] | layer1_out[3971];
     layer2_out[35] <= ~(layer1_out[5190] ^ layer1_out[5191]);
     layer2_out[36] <= layer1_out[11113] & layer1_out[11114];
     layer2_out[37] <= layer1_out[4557];
     layer2_out[38] <= ~(layer1_out[7655] ^ layer1_out[7656]);
     layer2_out[39] <= ~layer1_out[9010];
     layer2_out[40] <= ~(layer1_out[10455] | layer1_out[10456]);
     layer2_out[41] <= layer1_out[8094] ^ layer1_out[8095];
     layer2_out[42] <= layer1_out[4258];
     layer2_out[43] <= layer1_out[5399];
     layer2_out[44] <= ~layer1_out[9864] | layer1_out[9865];
     layer2_out[45] <= layer1_out[10173] & ~layer1_out[10174];
     layer2_out[46] <= ~layer1_out[10265] | layer1_out[10266];
     layer2_out[47] <= layer1_out[10010] & layer1_out[10011];
     layer2_out[48] <= layer1_out[6039];
     layer2_out[49] <= layer1_out[7759] & layer1_out[7760];
     layer2_out[50] <= layer1_out[4734] & ~layer1_out[4735];
     layer2_out[51] <= layer1_out[6317];
     layer2_out[52] <= layer1_out[11488] | layer1_out[11489];
     layer2_out[53] <= layer1_out[6545] ^ layer1_out[6546];
     layer2_out[54] <= 1'b0;
     layer2_out[55] <= ~(layer1_out[556] & layer1_out[557]);
     layer2_out[56] <= layer1_out[1436];
     layer2_out[57] <= ~(layer1_out[5381] | layer1_out[5382]);
     layer2_out[58] <= 1'b0;
     layer2_out[59] <= layer1_out[4515];
     layer2_out[60] <= layer1_out[11546] & layer1_out[11547];
     layer2_out[61] <= ~layer1_out[8145];
     layer2_out[62] <= layer1_out[11124] & ~layer1_out[11125];
     layer2_out[63] <= layer1_out[5120] & ~layer1_out[5121];
     layer2_out[64] <= 1'b1;
     layer2_out[65] <= layer1_out[4649];
     layer2_out[66] <= ~(layer1_out[2109] ^ layer1_out[2110]);
     layer2_out[67] <= ~(layer1_out[97] | layer1_out[98]);
     layer2_out[68] <= ~(layer1_out[5074] | layer1_out[5075]);
     layer2_out[69] <= ~(layer1_out[8142] ^ layer1_out[8143]);
     layer2_out[70] <= layer1_out[2073] & ~layer1_out[2074];
     layer2_out[71] <= ~layer1_out[10847] | layer1_out[10846];
     layer2_out[72] <= layer1_out[6638];
     layer2_out[73] <= layer1_out[3922] & ~layer1_out[3923];
     layer2_out[74] <= layer1_out[10407] ^ layer1_out[10408];
     layer2_out[75] <= ~layer1_out[4790];
     layer2_out[76] <= ~(layer1_out[7335] & layer1_out[7336]);
     layer2_out[77] <= layer1_out[11077] & ~layer1_out[11078];
     layer2_out[78] <= layer1_out[1485] & ~layer1_out[1486];
     layer2_out[79] <= ~layer1_out[3388];
     layer2_out[80] <= ~(layer1_out[11245] & layer1_out[11246]);
     layer2_out[81] <= ~layer1_out[3780];
     layer2_out[82] <= ~layer1_out[2492];
     layer2_out[83] <= ~(layer1_out[3077] & layer1_out[3078]);
     layer2_out[84] <= ~layer1_out[1871] | layer1_out[1870];
     layer2_out[85] <= layer1_out[8635] & ~layer1_out[8636];
     layer2_out[86] <= layer1_out[11070] & layer1_out[11071];
     layer2_out[87] <= ~(layer1_out[4264] & layer1_out[4265]);
     layer2_out[88] <= layer1_out[8819];
     layer2_out[89] <= layer1_out[3540];
     layer2_out[90] <= layer1_out[1776] & ~layer1_out[1775];
     layer2_out[91] <= layer1_out[10543] & ~layer1_out[10544];
     layer2_out[92] <= layer1_out[8628];
     layer2_out[93] <= layer1_out[5260] | layer1_out[5261];
     layer2_out[94] <= layer1_out[6975] | layer1_out[6976];
     layer2_out[95] <= layer1_out[9190] & ~layer1_out[9189];
     layer2_out[96] <= ~layer1_out[4094];
     layer2_out[97] <= ~layer1_out[5132];
     layer2_out[98] <= ~(layer1_out[3231] ^ layer1_out[3232]);
     layer2_out[99] <= layer1_out[7874] | layer1_out[7875];
     layer2_out[100] <= layer1_out[7587] | layer1_out[7588];
     layer2_out[101] <= layer1_out[8285] | layer1_out[8286];
     layer2_out[102] <= ~layer1_out[9341];
     layer2_out[103] <= ~(layer1_out[3878] ^ layer1_out[3879]);
     layer2_out[104] <= layer1_out[6067];
     layer2_out[105] <= ~(layer1_out[10615] & layer1_out[10616]);
     layer2_out[106] <= ~layer1_out[5910] | layer1_out[5909];
     layer2_out[107] <= ~(layer1_out[5688] & layer1_out[5689]);
     layer2_out[108] <= layer1_out[10991];
     layer2_out[109] <= layer1_out[9271] & ~layer1_out[9272];
     layer2_out[110] <= layer1_out[9320];
     layer2_out[111] <= ~layer1_out[8923] | layer1_out[8924];
     layer2_out[112] <= ~(layer1_out[11964] & layer1_out[11965]);
     layer2_out[113] <= layer1_out[2420];
     layer2_out[114] <= ~(layer1_out[5299] | layer1_out[5300]);
     layer2_out[115] <= ~layer1_out[3384] | layer1_out[3385];
     layer2_out[116] <= ~layer1_out[11776];
     layer2_out[117] <= ~layer1_out[2060] | layer1_out[2059];
     layer2_out[118] <= ~layer1_out[6517] | layer1_out[6516];
     layer2_out[119] <= ~(layer1_out[10977] & layer1_out[10978]);
     layer2_out[120] <= ~layer1_out[8274] | layer1_out[8275];
     layer2_out[121] <= layer1_out[4987];
     layer2_out[122] <= layer1_out[2812];
     layer2_out[123] <= layer1_out[7904];
     layer2_out[124] <= layer1_out[9059] & ~layer1_out[9058];
     layer2_out[125] <= ~(layer1_out[11463] & layer1_out[11464]);
     layer2_out[126] <= ~layer1_out[5110];
     layer2_out[127] <= layer1_out[1634] & ~layer1_out[1635];
     layer2_out[128] <= ~layer1_out[11398];
     layer2_out[129] <= layer1_out[4290] ^ layer1_out[4291];
     layer2_out[130] <= layer1_out[6369] & ~layer1_out[6368];
     layer2_out[131] <= ~(layer1_out[9752] | layer1_out[9753]);
     layer2_out[132] <= layer1_out[7446] | layer1_out[7447];
     layer2_out[133] <= ~layer1_out[5593];
     layer2_out[134] <= layer1_out[175];
     layer2_out[135] <= layer1_out[2924] | layer1_out[2925];
     layer2_out[136] <= ~layer1_out[4203] | layer1_out[4204];
     layer2_out[137] <= layer1_out[2692] | layer1_out[2693];
     layer2_out[138] <= layer1_out[8853];
     layer2_out[139] <= layer1_out[9053];
     layer2_out[140] <= ~(layer1_out[5345] & layer1_out[5346]);
     layer2_out[141] <= layer1_out[3231] & ~layer1_out[3230];
     layer2_out[142] <= layer1_out[122] | layer1_out[123];
     layer2_out[143] <= ~layer1_out[1395] | layer1_out[1394];
     layer2_out[144] <= layer1_out[1602] ^ layer1_out[1603];
     layer2_out[145] <= ~(layer1_out[11700] & layer1_out[11701]);
     layer2_out[146] <= ~layer1_out[778] | layer1_out[777];
     layer2_out[147] <= ~layer1_out[4143];
     layer2_out[148] <= layer1_out[8999] & ~layer1_out[8998];
     layer2_out[149] <= ~layer1_out[1630];
     layer2_out[150] <= 1'b1;
     layer2_out[151] <= layer1_out[6287];
     layer2_out[152] <= layer1_out[8975] | layer1_out[8976];
     layer2_out[153] <= ~layer1_out[988] | layer1_out[987];
     layer2_out[154] <= ~(layer1_out[10848] | layer1_out[10849]);
     layer2_out[155] <= layer1_out[2892] & ~layer1_out[2893];
     layer2_out[156] <= layer1_out[3142] & layer1_out[3143];
     layer2_out[157] <= layer1_out[2075] & ~layer1_out[2076];
     layer2_out[158] <= ~layer1_out[10226] | layer1_out[10227];
     layer2_out[159] <= 1'b1;
     layer2_out[160] <= layer1_out[2861] & layer1_out[2862];
     layer2_out[161] <= layer1_out[1446] & layer1_out[1447];
     layer2_out[162] <= layer1_out[2695] & ~layer1_out[2694];
     layer2_out[163] <= layer1_out[9324] & ~layer1_out[9323];
     layer2_out[164] <= ~(layer1_out[6674] & layer1_out[6675]);
     layer2_out[165] <= layer1_out[11238] & ~layer1_out[11237];
     layer2_out[166] <= ~layer1_out[5214];
     layer2_out[167] <= layer1_out[2822] | layer1_out[2823];
     layer2_out[168] <= ~layer1_out[11729];
     layer2_out[169] <= layer1_out[11145] ^ layer1_out[11146];
     layer2_out[170] <= ~(layer1_out[7264] | layer1_out[7265]);
     layer2_out[171] <= ~layer1_out[1962];
     layer2_out[172] <= layer1_out[8643] & ~layer1_out[8644];
     layer2_out[173] <= ~layer1_out[11890] | layer1_out[11891];
     layer2_out[174] <= layer1_out[4367];
     layer2_out[175] <= layer1_out[11827] | layer1_out[11828];
     layer2_out[176] <= ~layer1_out[718] | layer1_out[719];
     layer2_out[177] <= layer1_out[1838] ^ layer1_out[1839];
     layer2_out[178] <= ~(layer1_out[8494] | layer1_out[8495]);
     layer2_out[179] <= ~layer1_out[8865];
     layer2_out[180] <= layer1_out[10776];
     layer2_out[181] <= ~(layer1_out[6089] ^ layer1_out[6090]);
     layer2_out[182] <= ~(layer1_out[4909] ^ layer1_out[4910]);
     layer2_out[183] <= layer1_out[7010] | layer1_out[7011];
     layer2_out[184] <= ~layer1_out[7432];
     layer2_out[185] <= ~(layer1_out[147] | layer1_out[148]);
     layer2_out[186] <= layer1_out[3223];
     layer2_out[187] <= layer1_out[4226];
     layer2_out[188] <= ~layer1_out[8879];
     layer2_out[189] <= layer1_out[9132];
     layer2_out[190] <= ~(layer1_out[11068] & layer1_out[11069]);
     layer2_out[191] <= ~layer1_out[2225];
     layer2_out[192] <= ~layer1_out[6690];
     layer2_out[193] <= layer1_out[6408] & layer1_out[6409];
     layer2_out[194] <= layer1_out[197];
     layer2_out[195] <= layer1_out[2169] | layer1_out[2170];
     layer2_out[196] <= layer1_out[3334] ^ layer1_out[3335];
     layer2_out[197] <= layer1_out[4222];
     layer2_out[198] <= ~layer1_out[2327] | layer1_out[2328];
     layer2_out[199] <= layer1_out[413];
     layer2_out[200] <= layer1_out[4190] & layer1_out[4191];
     layer2_out[201] <= layer1_out[7691];
     layer2_out[202] <= ~layer1_out[10430];
     layer2_out[203] <= layer1_out[64] ^ layer1_out[65];
     layer2_out[204] <= layer1_out[9758] & ~layer1_out[9757];
     layer2_out[205] <= ~layer1_out[9309];
     layer2_out[206] <= ~layer1_out[947];
     layer2_out[207] <= layer1_out[3222] & ~layer1_out[3221];
     layer2_out[208] <= layer1_out[1527] & ~layer1_out[1528];
     layer2_out[209] <= ~layer1_out[1536];
     layer2_out[210] <= layer1_out[3994];
     layer2_out[211] <= layer1_out[8701];
     layer2_out[212] <= layer1_out[5387] | layer1_out[5388];
     layer2_out[213] <= ~layer1_out[9485] | layer1_out[9484];
     layer2_out[214] <= layer1_out[2512];
     layer2_out[215] <= layer1_out[1102] & layer1_out[1103];
     layer2_out[216] <= ~layer1_out[10292] | layer1_out[10291];
     layer2_out[217] <= ~layer1_out[3499];
     layer2_out[218] <= ~(layer1_out[1844] ^ layer1_out[1845]);
     layer2_out[219] <= 1'b0;
     layer2_out[220] <= ~layer1_out[9192] | layer1_out[9193];
     layer2_out[221] <= ~(layer1_out[1583] | layer1_out[1584]);
     layer2_out[222] <= layer1_out[6223];
     layer2_out[223] <= ~layer1_out[455];
     layer2_out[224] <= layer1_out[4525];
     layer2_out[225] <= layer1_out[11186] & layer1_out[11187];
     layer2_out[226] <= ~(layer1_out[3997] ^ layer1_out[3998]);
     layer2_out[227] <= layer1_out[11608] ^ layer1_out[11609];
     layer2_out[228] <= ~(layer1_out[8549] | layer1_out[8550]);
     layer2_out[229] <= ~(layer1_out[6086] | layer1_out[6087]);
     layer2_out[230] <= layer1_out[1772];
     layer2_out[231] <= ~(layer1_out[9115] ^ layer1_out[9116]);
     layer2_out[232] <= ~(layer1_out[1143] & layer1_out[1144]);
     layer2_out[233] <= ~layer1_out[8987];
     layer2_out[234] <= ~layer1_out[8533] | layer1_out[8532];
     layer2_out[235] <= ~(layer1_out[4076] | layer1_out[4077]);
     layer2_out[236] <= ~layer1_out[3301];
     layer2_out[237] <= ~(layer1_out[229] & layer1_out[230]);
     layer2_out[238] <= ~layer1_out[11637] | layer1_out[11638];
     layer2_out[239] <= layer1_out[8924] & layer1_out[8925];
     layer2_out[240] <= layer1_out[3357] ^ layer1_out[3358];
     layer2_out[241] <= layer1_out[9590] & layer1_out[9591];
     layer2_out[242] <= ~layer1_out[5800];
     layer2_out[243] <= layer1_out[4270];
     layer2_out[244] <= layer1_out[6950] & layer1_out[6951];
     layer2_out[245] <= ~(layer1_out[7479] ^ layer1_out[7480]);
     layer2_out[246] <= ~layer1_out[10757] | layer1_out[10756];
     layer2_out[247] <= layer1_out[3809] & ~layer1_out[3808];
     layer2_out[248] <= ~layer1_out[2356];
     layer2_out[249] <= ~layer1_out[8983];
     layer2_out[250] <= ~layer1_out[3092];
     layer2_out[251] <= layer1_out[6516];
     layer2_out[252] <= ~(layer1_out[5533] ^ layer1_out[5534]);
     layer2_out[253] <= ~(layer1_out[4098] & layer1_out[4099]);
     layer2_out[254] <= layer1_out[6885] & ~layer1_out[6884];
     layer2_out[255] <= ~(layer1_out[162] | layer1_out[163]);
     layer2_out[256] <= ~layer1_out[10711];
     layer2_out[257] <= ~(layer1_out[5116] | layer1_out[5117]);
     layer2_out[258] <= layer1_out[3753] & layer1_out[3754];
     layer2_out[259] <= ~layer1_out[6012] | layer1_out[6013];
     layer2_out[260] <= ~(layer1_out[11528] | layer1_out[11529]);
     layer2_out[261] <= ~layer1_out[9176] | layer1_out[9175];
     layer2_out[262] <= layer1_out[10013];
     layer2_out[263] <= ~layer1_out[4059];
     layer2_out[264] <= layer1_out[11436] ^ layer1_out[11437];
     layer2_out[265] <= ~layer1_out[1581];
     layer2_out[266] <= ~layer1_out[3495] | layer1_out[3496];
     layer2_out[267] <= ~layer1_out[711];
     layer2_out[268] <= layer1_out[5013] & ~layer1_out[5014];
     layer2_out[269] <= layer1_out[6738];
     layer2_out[270] <= layer1_out[8164] & ~layer1_out[8163];
     layer2_out[271] <= layer1_out[7066];
     layer2_out[272] <= ~layer1_out[4755];
     layer2_out[273] <= layer1_out[3433] & ~layer1_out[3434];
     layer2_out[274] <= ~(layer1_out[5602] & layer1_out[5603]);
     layer2_out[275] <= layer1_out[3164];
     layer2_out[276] <= layer1_out[10581];
     layer2_out[277] <= layer1_out[7579] | layer1_out[7580];
     layer2_out[278] <= ~layer1_out[8820] | layer1_out[8821];
     layer2_out[279] <= ~layer1_out[5561];
     layer2_out[280] <= layer1_out[6306] & ~layer1_out[6307];
     layer2_out[281] <= layer1_out[6551];
     layer2_out[282] <= layer1_out[2231] & layer1_out[2232];
     layer2_out[283] <= layer1_out[11523];
     layer2_out[284] <= layer1_out[2930] | layer1_out[2931];
     layer2_out[285] <= ~layer1_out[4012];
     layer2_out[286] <= layer1_out[9862];
     layer2_out[287] <= ~layer1_out[813];
     layer2_out[288] <= layer1_out[10428] | layer1_out[10429];
     layer2_out[289] <= layer1_out[9370] | layer1_out[9371];
     layer2_out[290] <= layer1_out[7157];
     layer2_out[291] <= layer1_out[6646];
     layer2_out[292] <= ~(layer1_out[11252] ^ layer1_out[11253]);
     layer2_out[293] <= ~(layer1_out[975] & layer1_out[976]);
     layer2_out[294] <= layer1_out[3889];
     layer2_out[295] <= layer1_out[2172];
     layer2_out[296] <= layer1_out[26] ^ layer1_out[27];
     layer2_out[297] <= ~layer1_out[9058];
     layer2_out[298] <= layer1_out[9729] & ~layer1_out[9730];
     layer2_out[299] <= layer1_out[5576];
     layer2_out[300] <= ~layer1_out[530];
     layer2_out[301] <= layer1_out[2743];
     layer2_out[302] <= ~(layer1_out[9803] & layer1_out[9804]);
     layer2_out[303] <= ~(layer1_out[1857] & layer1_out[1858]);
     layer2_out[304] <= layer1_out[5053] | layer1_out[5054];
     layer2_out[305] <= ~layer1_out[4618] | layer1_out[4619];
     layer2_out[306] <= ~layer1_out[1279];
     layer2_out[307] <= ~(layer1_out[6062] & layer1_out[6063]);
     layer2_out[308] <= layer1_out[9553];
     layer2_out[309] <= layer1_out[10964] & ~layer1_out[10965];
     layer2_out[310] <= ~layer1_out[6808];
     layer2_out[311] <= ~layer1_out[8977];
     layer2_out[312] <= layer1_out[6709] & layer1_out[6710];
     layer2_out[313] <= ~(layer1_out[1431] & layer1_out[1432]);
     layer2_out[314] <= layer1_out[11226] | layer1_out[11227];
     layer2_out[315] <= layer1_out[1070];
     layer2_out[316] <= layer1_out[6957] & ~layer1_out[6958];
     layer2_out[317] <= ~(layer1_out[4738] | layer1_out[4739]);
     layer2_out[318] <= ~layer1_out[7542];
     layer2_out[319] <= ~layer1_out[8009] | layer1_out[8010];
     layer2_out[320] <= layer1_out[8335] & layer1_out[8336];
     layer2_out[321] <= layer1_out[4361] & layer1_out[4362];
     layer2_out[322] <= layer1_out[464];
     layer2_out[323] <= ~(layer1_out[2452] ^ layer1_out[2453]);
     layer2_out[324] <= layer1_out[200];
     layer2_out[325] <= ~layer1_out[5372];
     layer2_out[326] <= ~layer1_out[3184];
     layer2_out[327] <= layer1_out[8990] & ~layer1_out[8991];
     layer2_out[328] <= layer1_out[6695] & ~layer1_out[6696];
     layer2_out[329] <= ~layer1_out[3323];
     layer2_out[330] <= ~(layer1_out[506] | layer1_out[507]);
     layer2_out[331] <= ~layer1_out[9521];
     layer2_out[332] <= ~(layer1_out[4405] | layer1_out[4406]);
     layer2_out[333] <= layer1_out[2526] & ~layer1_out[2525];
     layer2_out[334] <= layer1_out[7931] | layer1_out[7932];
     layer2_out[335] <= layer1_out[10840];
     layer2_out[336] <= layer1_out[8170];
     layer2_out[337] <= ~layer1_out[3070];
     layer2_out[338] <= 1'b1;
     layer2_out[339] <= ~(layer1_out[4955] & layer1_out[4956]);
     layer2_out[340] <= ~(layer1_out[1916] & layer1_out[1917]);
     layer2_out[341] <= layer1_out[2079] ^ layer1_out[2080];
     layer2_out[342] <= layer1_out[10008];
     layer2_out[343] <= layer1_out[10753];
     layer2_out[344] <= layer1_out[2409] & ~layer1_out[2408];
     layer2_out[345] <= ~(layer1_out[5952] & layer1_out[5953]);
     layer2_out[346] <= layer1_out[2907];
     layer2_out[347] <= ~(layer1_out[9769] & layer1_out[9770]);
     layer2_out[348] <= layer1_out[359];
     layer2_out[349] <= layer1_out[8758] & ~layer1_out[8759];
     layer2_out[350] <= ~layer1_out[2048];
     layer2_out[351] <= layer1_out[5469] & ~layer1_out[5470];
     layer2_out[352] <= layer1_out[2385] ^ layer1_out[2386];
     layer2_out[353] <= layer1_out[10357];
     layer2_out[354] <= layer1_out[568] & ~layer1_out[567];
     layer2_out[355] <= ~layer1_out[2205] | layer1_out[2206];
     layer2_out[356] <= layer1_out[8725] ^ layer1_out[8726];
     layer2_out[357] <= layer1_out[9218];
     layer2_out[358] <= ~(layer1_out[3719] | layer1_out[3720]);
     layer2_out[359] <= ~layer1_out[1151];
     layer2_out[360] <= ~(layer1_out[5407] | layer1_out[5408]);
     layer2_out[361] <= layer1_out[1364] | layer1_out[1365];
     layer2_out[362] <= layer1_out[5596];
     layer2_out[363] <= ~layer1_out[6136];
     layer2_out[364] <= layer1_out[454] ^ layer1_out[455];
     layer2_out[365] <= ~layer1_out[10497];
     layer2_out[366] <= ~(layer1_out[2830] ^ layer1_out[2831]);
     layer2_out[367] <= layer1_out[10679];
     layer2_out[368] <= ~(layer1_out[4611] | layer1_out[4612]);
     layer2_out[369] <= ~layer1_out[8141];
     layer2_out[370] <= layer1_out[5845] | layer1_out[5846];
     layer2_out[371] <= layer1_out[1738] | layer1_out[1739];
     layer2_out[372] <= layer1_out[5251] & ~layer1_out[5252];
     layer2_out[373] <= ~layer1_out[11563] | layer1_out[11564];
     layer2_out[374] <= layer1_out[3264];
     layer2_out[375] <= ~(layer1_out[8397] | layer1_out[8398]);
     layer2_out[376] <= layer1_out[9317] & layer1_out[9318];
     layer2_out[377] <= ~layer1_out[5734] | layer1_out[5733];
     layer2_out[378] <= layer1_out[9867] | layer1_out[9868];
     layer2_out[379] <= ~(layer1_out[10397] | layer1_out[10398]);
     layer2_out[380] <= ~(layer1_out[2128] & layer1_out[2129]);
     layer2_out[381] <= ~layer1_out[7599];
     layer2_out[382] <= layer1_out[1731] ^ layer1_out[1732];
     layer2_out[383] <= ~(layer1_out[11975] ^ layer1_out[11976]);
     layer2_out[384] <= layer1_out[11229];
     layer2_out[385] <= ~(layer1_out[6654] & layer1_out[6655]);
     layer2_out[386] <= ~layer1_out[11464];
     layer2_out[387] <= ~layer1_out[4770] | layer1_out[4769];
     layer2_out[388] <= ~layer1_out[9798];
     layer2_out[389] <= layer1_out[11125] & layer1_out[11126];
     layer2_out[390] <= ~layer1_out[10709];
     layer2_out[391] <= layer1_out[7234] & layer1_out[7235];
     layer2_out[392] <= ~layer1_out[11394];
     layer2_out[393] <= ~(layer1_out[10061] | layer1_out[10062]);
     layer2_out[394] <= ~(layer1_out[8609] & layer1_out[8610]);
     layer2_out[395] <= layer1_out[8606] | layer1_out[8607];
     layer2_out[396] <= ~(layer1_out[10686] & layer1_out[10687]);
     layer2_out[397] <= ~layer1_out[4321];
     layer2_out[398] <= ~layer1_out[4032];
     layer2_out[399] <= ~(layer1_out[7612] | layer1_out[7613]);
     layer2_out[400] <= 1'b0;
     layer2_out[401] <= ~(layer1_out[10687] & layer1_out[10688]);
     layer2_out[402] <= layer1_out[2218];
     layer2_out[403] <= layer1_out[1901] | layer1_out[1902];
     layer2_out[404] <= layer1_out[9509];
     layer2_out[405] <= layer1_out[9140];
     layer2_out[406] <= layer1_out[6371];
     layer2_out[407] <= layer1_out[5652] & layer1_out[5653];
     layer2_out[408] <= layer1_out[7770];
     layer2_out[409] <= layer1_out[2594];
     layer2_out[410] <= ~(layer1_out[6776] | layer1_out[6777]);
     layer2_out[411] <= layer1_out[5542] | layer1_out[5543];
     layer2_out[412] <= layer1_out[4629];
     layer2_out[413] <= ~layer1_out[4408];
     layer2_out[414] <= layer1_out[173];
     layer2_out[415] <= ~layer1_out[10045];
     layer2_out[416] <= ~layer1_out[10691];
     layer2_out[417] <= ~layer1_out[6926] | layer1_out[6925];
     layer2_out[418] <= ~layer1_out[4522];
     layer2_out[419] <= layer1_out[3168] & layer1_out[3169];
     layer2_out[420] <= layer1_out[1060];
     layer2_out[421] <= layer1_out[1895] & layer1_out[1896];
     layer2_out[422] <= ~(layer1_out[10688] & layer1_out[10689]);
     layer2_out[423] <= ~layer1_out[9202];
     layer2_out[424] <= ~(layer1_out[4634] | layer1_out[4635]);
     layer2_out[425] <= ~layer1_out[1843];
     layer2_out[426] <= layer1_out[7905];
     layer2_out[427] <= layer1_out[11038] | layer1_out[11039];
     layer2_out[428] <= ~layer1_out[3095];
     layer2_out[429] <= layer1_out[8265] | layer1_out[8266];
     layer2_out[430] <= ~layer1_out[10717];
     layer2_out[431] <= layer1_out[5277] | layer1_out[5278];
     layer2_out[432] <= layer1_out[3901];
     layer2_out[433] <= ~layer1_out[10671];
     layer2_out[434] <= layer1_out[3983] & layer1_out[3984];
     layer2_out[435] <= layer1_out[11527];
     layer2_out[436] <= ~layer1_out[6766] | layer1_out[6767];
     layer2_out[437] <= layer1_out[9710] & ~layer1_out[9711];
     layer2_out[438] <= layer1_out[5061] ^ layer1_out[5062];
     layer2_out[439] <= layer1_out[4108] ^ layer1_out[4109];
     layer2_out[440] <= layer1_out[10815] & layer1_out[10816];
     layer2_out[441] <= layer1_out[6652] ^ layer1_out[6653];
     layer2_out[442] <= ~layer1_out[8535];
     layer2_out[443] <= ~layer1_out[1900] | layer1_out[1899];
     layer2_out[444] <= ~layer1_out[2149];
     layer2_out[445] <= ~(layer1_out[10327] | layer1_out[10328]);
     layer2_out[446] <= layer1_out[8036];
     layer2_out[447] <= layer1_out[7199] & ~layer1_out[7198];
     layer2_out[448] <= ~layer1_out[10820];
     layer2_out[449] <= ~layer1_out[2130] | layer1_out[2131];
     layer2_out[450] <= ~(layer1_out[701] & layer1_out[702]);
     layer2_out[451] <= ~(layer1_out[4599] & layer1_out[4600]);
     layer2_out[452] <= layer1_out[10210] & ~layer1_out[10209];
     layer2_out[453] <= 1'b0;
     layer2_out[454] <= ~layer1_out[2181];
     layer2_out[455] <= layer1_out[6529];
     layer2_out[456] <= layer1_out[5669];
     layer2_out[457] <= layer1_out[4889];
     layer2_out[458] <= ~layer1_out[8401] | layer1_out[8402];
     layer2_out[459] <= ~layer1_out[9645] | layer1_out[9644];
     layer2_out[460] <= layer1_out[4915];
     layer2_out[461] <= layer1_out[4040] & layer1_out[4041];
     layer2_out[462] <= layer1_out[770] & ~layer1_out[769];
     layer2_out[463] <= layer1_out[10980] & layer1_out[10981];
     layer2_out[464] <= layer1_out[11577];
     layer2_out[465] <= layer1_out[11474];
     layer2_out[466] <= ~(layer1_out[6547] ^ layer1_out[6548]);
     layer2_out[467] <= ~layer1_out[6431] | layer1_out[6430];
     layer2_out[468] <= layer1_out[6540] & ~layer1_out[6541];
     layer2_out[469] <= 1'b0;
     layer2_out[470] <= layer1_out[5294];
     layer2_out[471] <= ~(layer1_out[9194] | layer1_out[9195]);
     layer2_out[472] <= ~layer1_out[11883];
     layer2_out[473] <= layer1_out[1644];
     layer2_out[474] <= layer1_out[6031] | layer1_out[6032];
     layer2_out[475] <= ~(layer1_out[5736] & layer1_out[5737]);
     layer2_out[476] <= layer1_out[10778];
     layer2_out[477] <= layer1_out[10597] & ~layer1_out[10598];
     layer2_out[478] <= ~layer1_out[1653];
     layer2_out[479] <= ~(layer1_out[4798] | layer1_out[4799]);
     layer2_out[480] <= 1'b1;
     layer2_out[481] <= layer1_out[8168] & ~layer1_out[8169];
     layer2_out[482] <= ~(layer1_out[11348] & layer1_out[11349]);
     layer2_out[483] <= ~layer1_out[1676] | layer1_out[1677];
     layer2_out[484] <= ~layer1_out[11304];
     layer2_out[485] <= layer1_out[9777];
     layer2_out[486] <= ~layer1_out[5309] | layer1_out[5308];
     layer2_out[487] <= layer1_out[10278];
     layer2_out[488] <= ~(layer1_out[5314] & layer1_out[5315]);
     layer2_out[489] <= ~layer1_out[3313];
     layer2_out[490] <= layer1_out[3107] | layer1_out[3108];
     layer2_out[491] <= layer1_out[9567];
     layer2_out[492] <= layer1_out[766] & layer1_out[767];
     layer2_out[493] <= layer1_out[10435] & layer1_out[10436];
     layer2_out[494] <= layer1_out[9981];
     layer2_out[495] <= layer1_out[3516] ^ layer1_out[3517];
     layer2_out[496] <= ~layer1_out[4221];
     layer2_out[497] <= layer1_out[4778];
     layer2_out[498] <= ~layer1_out[10273];
     layer2_out[499] <= layer1_out[10680] ^ layer1_out[10681];
     layer2_out[500] <= layer1_out[9698] ^ layer1_out[9699];
     layer2_out[501] <= layer1_out[6655] & layer1_out[6656];
     layer2_out[502] <= ~layer1_out[9709];
     layer2_out[503] <= layer1_out[2974];
     layer2_out[504] <= ~layer1_out[3685];
     layer2_out[505] <= layer1_out[7786] ^ layer1_out[7787];
     layer2_out[506] <= ~(layer1_out[9380] ^ layer1_out[9381]);
     layer2_out[507] <= layer1_out[10499];
     layer2_out[508] <= layer1_out[1476];
     layer2_out[509] <= layer1_out[5259] | layer1_out[5260];
     layer2_out[510] <= layer1_out[551];
     layer2_out[511] <= ~(layer1_out[11878] ^ layer1_out[11879]);
     layer2_out[512] <= ~layer1_out[1054];
     layer2_out[513] <= layer1_out[6349];
     layer2_out[514] <= layer1_out[3616] | layer1_out[3617];
     layer2_out[515] <= ~(layer1_out[11672] | layer1_out[11673]);
     layer2_out[516] <= ~layer1_out[1373] | layer1_out[1374];
     layer2_out[517] <= layer1_out[11820] ^ layer1_out[11821];
     layer2_out[518] <= ~layer1_out[11289];
     layer2_out[519] <= ~(layer1_out[5166] & layer1_out[5167]);
     layer2_out[520] <= layer1_out[8757] | layer1_out[8758];
     layer2_out[521] <= ~layer1_out[8199];
     layer2_out[522] <= ~layer1_out[9732] | layer1_out[9731];
     layer2_out[523] <= ~layer1_out[5743];
     layer2_out[524] <= layer1_out[2006] & ~layer1_out[2007];
     layer2_out[525] <= layer1_out[3862];
     layer2_out[526] <= ~layer1_out[10966];
     layer2_out[527] <= layer1_out[11982] & ~layer1_out[11983];
     layer2_out[528] <= ~layer1_out[4849] | layer1_out[4848];
     layer2_out[529] <= layer1_out[3915] ^ layer1_out[3916];
     layer2_out[530] <= ~(layer1_out[8694] | layer1_out[8695]);
     layer2_out[531] <= layer1_out[7315] & ~layer1_out[7316];
     layer2_out[532] <= layer1_out[4158] ^ layer1_out[4159];
     layer2_out[533] <= layer1_out[10490];
     layer2_out[534] <= layer1_out[8254] & ~layer1_out[8255];
     layer2_out[535] <= ~(layer1_out[11903] | layer1_out[11904]);
     layer2_out[536] <= layer1_out[10112] & ~layer1_out[10111];
     layer2_out[537] <= ~layer1_out[6744] | layer1_out[6745];
     layer2_out[538] <= ~layer1_out[6778];
     layer2_out[539] <= ~(layer1_out[8496] | layer1_out[8497]);
     layer2_out[540] <= 1'b1;
     layer2_out[541] <= layer1_out[2507];
     layer2_out[542] <= ~layer1_out[8599];
     layer2_out[543] <= ~layer1_out[2761] | layer1_out[2760];
     layer2_out[544] <= ~(layer1_out[11684] ^ layer1_out[11685]);
     layer2_out[545] <= ~layer1_out[11660];
     layer2_out[546] <= ~layer1_out[6734];
     layer2_out[547] <= ~layer1_out[2827];
     layer2_out[548] <= ~(layer1_out[8037] & layer1_out[8038]);
     layer2_out[549] <= layer1_out[6875];
     layer2_out[550] <= layer1_out[3424];
     layer2_out[551] <= ~layer1_out[2679] | layer1_out[2680];
     layer2_out[552] <= ~(layer1_out[2285] & layer1_out[2286]);
     layer2_out[553] <= ~layer1_out[11178];
     layer2_out[554] <= layer1_out[7906] | layer1_out[7907];
     layer2_out[555] <= layer1_out[10138];
     layer2_out[556] <= ~(layer1_out[9554] | layer1_out[9555]);
     layer2_out[557] <= layer1_out[6421];
     layer2_out[558] <= layer1_out[1252];
     layer2_out[559] <= layer1_out[9855] & ~layer1_out[9856];
     layer2_out[560] <= layer1_out[1235] & ~layer1_out[1236];
     layer2_out[561] <= layer1_out[10211];
     layer2_out[562] <= layer1_out[3037];
     layer2_out[563] <= layer1_out[11819];
     layer2_out[564] <= ~layer1_out[4354];
     layer2_out[565] <= ~(layer1_out[8622] | layer1_out[8623]);
     layer2_out[566] <= ~layer1_out[8631];
     layer2_out[567] <= layer1_out[11816];
     layer2_out[568] <= layer1_out[5350];
     layer2_out[569] <= ~(layer1_out[3364] ^ layer1_out[3365]);
     layer2_out[570] <= ~(layer1_out[1320] & layer1_out[1321]);
     layer2_out[571] <= ~layer1_out[2967] | layer1_out[2966];
     layer2_out[572] <= layer1_out[3027] & ~layer1_out[3026];
     layer2_out[573] <= ~(layer1_out[5362] | layer1_out[5363]);
     layer2_out[574] <= ~layer1_out[8848];
     layer2_out[575] <= ~layer1_out[3597];
     layer2_out[576] <= layer1_out[11011] & ~layer1_out[11010];
     layer2_out[577] <= ~(layer1_out[7305] & layer1_out[7306]);
     layer2_out[578] <= ~(layer1_out[6003] & layer1_out[6004]);
     layer2_out[579] <= layer1_out[3181];
     layer2_out[580] <= layer1_out[9468];
     layer2_out[581] <= ~(layer1_out[8794] & layer1_out[8795]);
     layer2_out[582] <= ~(layer1_out[1472] ^ layer1_out[1473]);
     layer2_out[583] <= ~layer1_out[3468];
     layer2_out[584] <= layer1_out[1318] & ~layer1_out[1317];
     layer2_out[585] <= layer1_out[5779] & ~layer1_out[5778];
     layer2_out[586] <= layer1_out[3200] & ~layer1_out[3199];
     layer2_out[587] <= layer1_out[383];
     layer2_out[588] <= ~layer1_out[9418];
     layer2_out[589] <= layer1_out[9433] | layer1_out[9434];
     layer2_out[590] <= ~layer1_out[495];
     layer2_out[591] <= layer1_out[7071] & ~layer1_out[7072];
     layer2_out[592] <= layer1_out[8388];
     layer2_out[593] <= layer1_out[9862];
     layer2_out[594] <= ~layer1_out[10989];
     layer2_out[595] <= layer1_out[10208] | layer1_out[10209];
     layer2_out[596] <= ~layer1_out[1679] | layer1_out[1680];
     layer2_out[597] <= ~(layer1_out[9005] | layer1_out[9006]);
     layer2_out[598] <= ~(layer1_out[6865] | layer1_out[6866]);
     layer2_out[599] <= layer1_out[9577] | layer1_out[9578];
     layer2_out[600] <= ~layer1_out[4016];
     layer2_out[601] <= layer1_out[6873] & layer1_out[6874];
     layer2_out[602] <= layer1_out[4528] & ~layer1_out[4529];
     layer2_out[603] <= layer1_out[6332] & ~layer1_out[6331];
     layer2_out[604] <= layer1_out[1290] & layer1_out[1291];
     layer2_out[605] <= layer1_out[1017];
     layer2_out[606] <= ~layer1_out[9070];
     layer2_out[607] <= ~(layer1_out[974] | layer1_out[975]);
     layer2_out[608] <= layer1_out[3815];
     layer2_out[609] <= ~layer1_out[10450];
     layer2_out[610] <= ~layer1_out[5879];
     layer2_out[611] <= layer1_out[4091] | layer1_out[4092];
     layer2_out[612] <= layer1_out[2900];
     layer2_out[613] <= ~layer1_out[4855] | layer1_out[4856];
     layer2_out[614] <= ~(layer1_out[4333] | layer1_out[4334]);
     layer2_out[615] <= layer1_out[7029] | layer1_out[7030];
     layer2_out[616] <= ~(layer1_out[8630] & layer1_out[8631]);
     layer2_out[617] <= ~(layer1_out[7754] & layer1_out[7755]);
     layer2_out[618] <= ~layer1_out[11296];
     layer2_out[619] <= ~layer1_out[7428] | layer1_out[7427];
     layer2_out[620] <= ~layer1_out[1963];
     layer2_out[621] <= ~layer1_out[6816];
     layer2_out[622] <= ~layer1_out[6497] | layer1_out[6496];
     layer2_out[623] <= layer1_out[7231] & ~layer1_out[7230];
     layer2_out[624] <= layer1_out[11703] & layer1_out[11704];
     layer2_out[625] <= ~(layer1_out[9919] & layer1_out[9920]);
     layer2_out[626] <= ~layer1_out[3807];
     layer2_out[627] <= ~layer1_out[7753];
     layer2_out[628] <= ~(layer1_out[10554] ^ layer1_out[10555]);
     layer2_out[629] <= ~layer1_out[6704] | layer1_out[6705];
     layer2_out[630] <= ~layer1_out[5484];
     layer2_out[631] <= ~layer1_out[6759];
     layer2_out[632] <= layer1_out[3707];
     layer2_out[633] <= layer1_out[9475];
     layer2_out[634] <= ~layer1_out[4717];
     layer2_out[635] <= layer1_out[3369];
     layer2_out[636] <= layer1_out[11551] & ~layer1_out[11550];
     layer2_out[637] <= layer1_out[3659];
     layer2_out[638] <= ~layer1_out[626];
     layer2_out[639] <= layer1_out[3781] & layer1_out[3782];
     layer2_out[640] <= layer1_out[503] & ~layer1_out[502];
     layer2_out[641] <= ~(layer1_out[1504] & layer1_out[1505]);
     layer2_out[642] <= layer1_out[1412] & ~layer1_out[1413];
     layer2_out[643] <= ~layer1_out[1627];
     layer2_out[644] <= ~layer1_out[1368];
     layer2_out[645] <= layer1_out[5389];
     layer2_out[646] <= layer1_out[1710];
     layer2_out[647] <= ~(layer1_out[1218] | layer1_out[1219]);
     layer2_out[648] <= layer1_out[9161] ^ layer1_out[9162];
     layer2_out[649] <= layer1_out[3501] & layer1_out[3502];
     layer2_out[650] <= 1'b1;
     layer2_out[651] <= layer1_out[10234];
     layer2_out[652] <= layer1_out[11475] & ~layer1_out[11476];
     layer2_out[653] <= layer1_out[11673] | layer1_out[11674];
     layer2_out[654] <= layer1_out[3824];
     layer2_out[655] <= ~(layer1_out[150] | layer1_out[151]);
     layer2_out[656] <= layer1_out[3827] & ~layer1_out[3828];
     layer2_out[657] <= ~layer1_out[133];
     layer2_out[658] <= 1'b0;
     layer2_out[659] <= ~layer1_out[2917] | layer1_out[2916];
     layer2_out[660] <= ~layer1_out[1878] | layer1_out[1877];
     layer2_out[661] <= ~layer1_out[10086] | layer1_out[10087];
     layer2_out[662] <= ~(layer1_out[5700] | layer1_out[5701]);
     layer2_out[663] <= layer1_out[3353] & ~layer1_out[3352];
     layer2_out[664] <= ~layer1_out[7939] | layer1_out[7938];
     layer2_out[665] <= layer1_out[9044];
     layer2_out[666] <= ~layer1_out[3852] | layer1_out[3853];
     layer2_out[667] <= ~(layer1_out[4077] & layer1_out[4078]);
     layer2_out[668] <= layer1_out[10801] ^ layer1_out[10802];
     layer2_out[669] <= layer1_out[7914];
     layer2_out[670] <= ~(layer1_out[10089] | layer1_out[10090]);
     layer2_out[671] <= ~layer1_out[9872];
     layer2_out[672] <= ~layer1_out[4752] | layer1_out[4751];
     layer2_out[673] <= ~(layer1_out[7971] ^ layer1_out[7972]);
     layer2_out[674] <= ~layer1_out[1538];
     layer2_out[675] <= ~(layer1_out[2926] | layer1_out[2927]);
     layer2_out[676] <= layer1_out[2558];
     layer2_out[677] <= ~layer1_out[3827];
     layer2_out[678] <= layer1_out[9968] ^ layer1_out[9969];
     layer2_out[679] <= ~(layer1_out[7883] & layer1_out[7884]);
     layer2_out[680] <= ~layer1_out[760];
     layer2_out[681] <= layer1_out[8174] & ~layer1_out[8175];
     layer2_out[682] <= ~(layer1_out[6888] | layer1_out[6889]);
     layer2_out[683] <= layer1_out[1270] & layer1_out[1271];
     layer2_out[684] <= ~layer1_out[3061] | layer1_out[3060];
     layer2_out[685] <= layer1_out[7327] & layer1_out[7328];
     layer2_out[686] <= ~(layer1_out[3426] ^ layer1_out[3427]);
     layer2_out[687] <= layer1_out[9130];
     layer2_out[688] <= ~layer1_out[5383];
     layer2_out[689] <= layer1_out[3140] & layer1_out[3141];
     layer2_out[690] <= layer1_out[9792] | layer1_out[9793];
     layer2_out[691] <= layer1_out[2116] | layer1_out[2117];
     layer2_out[692] <= ~layer1_out[1932];
     layer2_out[693] <= ~layer1_out[10813] | layer1_out[10814];
     layer2_out[694] <= layer1_out[8455] & ~layer1_out[8456];
     layer2_out[695] <= layer1_out[333];
     layer2_out[696] <= layer1_out[7904] & ~layer1_out[7905];
     layer2_out[697] <= ~layer1_out[9446];
     layer2_out[698] <= ~(layer1_out[4712] | layer1_out[4713]);
     layer2_out[699] <= layer1_out[6794] | layer1_out[6795];
     layer2_out[700] <= layer1_out[9280] & ~layer1_out[9279];
     layer2_out[701] <= layer1_out[10838];
     layer2_out[702] <= layer1_out[4233] & ~layer1_out[4232];
     layer2_out[703] <= layer1_out[8326] & ~layer1_out[8327];
     layer2_out[704] <= ~layer1_out[2544] | layer1_out[2545];
     layer2_out[705] <= layer1_out[2210] ^ layer1_out[2211];
     layer2_out[706] <= layer1_out[4195] ^ layer1_out[4196];
     layer2_out[707] <= layer1_out[3807];
     layer2_out[708] <= layer1_out[1104] & ~layer1_out[1105];
     layer2_out[709] <= 1'b0;
     layer2_out[710] <= layer1_out[5457];
     layer2_out[711] <= layer1_out[3857];
     layer2_out[712] <= layer1_out[11340] | layer1_out[11341];
     layer2_out[713] <= layer1_out[4101] | layer1_out[4102];
     layer2_out[714] <= ~(layer1_out[9055] ^ layer1_out[9056]);
     layer2_out[715] <= ~layer1_out[3834];
     layer2_out[716] <= ~(layer1_out[6435] | layer1_out[6436]);
     layer2_out[717] <= ~(layer1_out[4166] & layer1_out[4167]);
     layer2_out[718] <= layer1_out[9347];
     layer2_out[719] <= ~layer1_out[8137];
     layer2_out[720] <= layer1_out[8757] & ~layer1_out[8756];
     layer2_out[721] <= layer1_out[1829] ^ layer1_out[1830];
     layer2_out[722] <= ~layer1_out[4573];
     layer2_out[723] <= layer1_out[7104] & layer1_out[7105];
     layer2_out[724] <= ~(layer1_out[3576] | layer1_out[3577]);
     layer2_out[725] <= ~(layer1_out[7034] | layer1_out[7035]);
     layer2_out[726] <= layer1_out[7548] & ~layer1_out[7549];
     layer2_out[727] <= layer1_out[7272];
     layer2_out[728] <= layer1_out[11014] & ~layer1_out[11013];
     layer2_out[729] <= ~layer1_out[9615];
     layer2_out[730] <= layer1_out[316] | layer1_out[317];
     layer2_out[731] <= layer1_out[3363] ^ layer1_out[3364];
     layer2_out[732] <= layer1_out[8833];
     layer2_out[733] <= layer1_out[4840] & layer1_out[4841];
     layer2_out[734] <= ~layer1_out[3774] | layer1_out[3773];
     layer2_out[735] <= layer1_out[5331];
     layer2_out[736] <= layer1_out[6044];
     layer2_out[737] <= layer1_out[6117] & ~layer1_out[6116];
     layer2_out[738] <= layer1_out[538];
     layer2_out[739] <= layer1_out[10486];
     layer2_out[740] <= ~layer1_out[9784] | layer1_out[9783];
     layer2_out[741] <= layer1_out[3653] ^ layer1_out[3654];
     layer2_out[742] <= ~layer1_out[4180];
     layer2_out[743] <= ~layer1_out[10938];
     layer2_out[744] <= ~(layer1_out[7077] | layer1_out[7078]);
     layer2_out[745] <= ~(layer1_out[650] ^ layer1_out[651]);
     layer2_out[746] <= ~layer1_out[8727];
     layer2_out[747] <= layer1_out[6027];
     layer2_out[748] <= layer1_out[2368];
     layer2_out[749] <= layer1_out[10386] & layer1_out[10387];
     layer2_out[750] <= ~layer1_out[11083] | layer1_out[11084];
     layer2_out[751] <= ~(layer1_out[2072] & layer1_out[2073]);
     layer2_out[752] <= ~layer1_out[2304] | layer1_out[2305];
     layer2_out[753] <= ~layer1_out[1268] | layer1_out[1267];
     layer2_out[754] <= ~layer1_out[10635];
     layer2_out[755] <= layer1_out[8870];
     layer2_out[756] <= layer1_out[3937];
     layer2_out[757] <= ~layer1_out[9096];
     layer2_out[758] <= layer1_out[10698] & layer1_out[10699];
     layer2_out[759] <= layer1_out[3648];
     layer2_out[760] <= layer1_out[8033];
     layer2_out[761] <= 1'b1;
     layer2_out[762] <= layer1_out[1069];
     layer2_out[763] <= ~layer1_out[9111] | layer1_out[9112];
     layer2_out[764] <= layer1_out[3614];
     layer2_out[765] <= ~layer1_out[10510] | layer1_out[10511];
     layer2_out[766] <= ~layer1_out[8399] | layer1_out[8398];
     layer2_out[767] <= ~(layer1_out[978] | layer1_out[979]);
     layer2_out[768] <= layer1_out[7671];
     layer2_out[769] <= ~(layer1_out[7451] ^ layer1_out[7452]);
     layer2_out[770] <= ~layer1_out[8914] | layer1_out[8913];
     layer2_out[771] <= layer1_out[11516] | layer1_out[11517];
     layer2_out[772] <= layer1_out[6928];
     layer2_out[773] <= ~layer1_out[9183];
     layer2_out[774] <= ~(layer1_out[2238] ^ layer1_out[2239]);
     layer2_out[775] <= ~(layer1_out[11201] | layer1_out[11202]);
     layer2_out[776] <= ~layer1_out[7430] | layer1_out[7429];
     layer2_out[777] <= layer1_out[3617] | layer1_out[3618];
     layer2_out[778] <= ~layer1_out[11746];
     layer2_out[779] <= layer1_out[1891];
     layer2_out[780] <= ~layer1_out[8556] | layer1_out[8557];
     layer2_out[781] <= ~(layer1_out[11308] & layer1_out[11309]);
     layer2_out[782] <= ~layer1_out[9233];
     layer2_out[783] <= layer1_out[3272] & ~layer1_out[3271];
     layer2_out[784] <= layer1_out[5525] & ~layer1_out[5526];
     layer2_out[785] <= layer1_out[3955];
     layer2_out[786] <= layer1_out[10050] & layer1_out[10051];
     layer2_out[787] <= layer1_out[3134] | layer1_out[3135];
     layer2_out[788] <= layer1_out[7726];
     layer2_out[789] <= layer1_out[3660] & ~layer1_out[3661];
     layer2_out[790] <= layer1_out[480] ^ layer1_out[481];
     layer2_out[791] <= ~layer1_out[2077] | layer1_out[2078];
     layer2_out[792] <= layer1_out[3768] & layer1_out[3769];
     layer2_out[793] <= ~layer1_out[7307] | layer1_out[7306];
     layer2_out[794] <= ~(layer1_out[11062] ^ layer1_out[11063]);
     layer2_out[795] <= ~layer1_out[5724];
     layer2_out[796] <= layer1_out[2789];
     layer2_out[797] <= layer1_out[7692] & layer1_out[7693];
     layer2_out[798] <= ~layer1_out[6678] | layer1_out[6677];
     layer2_out[799] <= ~layer1_out[6011];
     layer2_out[800] <= ~(layer1_out[1273] | layer1_out[1274]);
     layer2_out[801] <= layer1_out[9454] | layer1_out[9455];
     layer2_out[802] <= ~(layer1_out[397] | layer1_out[398]);
     layer2_out[803] <= ~layer1_out[6748];
     layer2_out[804] <= ~(layer1_out[1411] | layer1_out[1412]);
     layer2_out[805] <= layer1_out[8075] ^ layer1_out[8076];
     layer2_out[806] <= ~(layer1_out[6353] & layer1_out[6354]);
     layer2_out[807] <= layer1_out[11198];
     layer2_out[808] <= layer1_out[3094] & ~layer1_out[3093];
     layer2_out[809] <= ~layer1_out[6986];
     layer2_out[810] <= layer1_out[5360] & ~layer1_out[5361];
     layer2_out[811] <= ~(layer1_out[7939] & layer1_out[7940]);
     layer2_out[812] <= layer1_out[2813];
     layer2_out[813] <= ~layer1_out[8293] | layer1_out[8292];
     layer2_out[814] <= layer1_out[6477];
     layer2_out[815] <= layer1_out[10359] & ~layer1_out[10358];
     layer2_out[816] <= ~(layer1_out[1762] | layer1_out[1763]);
     layer2_out[817] <= layer1_out[621] & layer1_out[622];
     layer2_out[818] <= ~layer1_out[6641] | layer1_out[6642];
     layer2_out[819] <= ~layer1_out[10200];
     layer2_out[820] <= ~(layer1_out[1160] | layer1_out[1161]);
     layer2_out[821] <= layer1_out[7235] & ~layer1_out[7236];
     layer2_out[822] <= layer1_out[8644];
     layer2_out[823] <= ~(layer1_out[3542] & layer1_out[3543]);
     layer2_out[824] <= ~(layer1_out[1551] ^ layer1_out[1552]);
     layer2_out[825] <= layer1_out[2121] | layer1_out[2122];
     layer2_out[826] <= ~layer1_out[2186] | layer1_out[2185];
     layer2_out[827] <= layer1_out[4447] & ~layer1_out[4448];
     layer2_out[828] <= layer1_out[8315] & layer1_out[8316];
     layer2_out[829] <= layer1_out[4994] & ~layer1_out[4995];
     layer2_out[830] <= layer1_out[2618];
     layer2_out[831] <= layer1_out[9299] ^ layer1_out[9300];
     layer2_out[832] <= ~layer1_out[11166] | layer1_out[11167];
     layer2_out[833] <= ~(layer1_out[1328] & layer1_out[1329]);
     layer2_out[834] <= ~(layer1_out[7465] & layer1_out[7466]);
     layer2_out[835] <= layer1_out[2644];
     layer2_out[836] <= layer1_out[3873];
     layer2_out[837] <= ~layer1_out[4069] | layer1_out[4070];
     layer2_out[838] <= ~layer1_out[6579] | layer1_out[6580];
     layer2_out[839] <= layer1_out[7153];
     layer2_out[840] <= layer1_out[775] ^ layer1_out[776];
     layer2_out[841] <= layer1_out[10997];
     layer2_out[842] <= layer1_out[485] & ~layer1_out[486];
     layer2_out[843] <= layer1_out[1152] & layer1_out[1153];
     layer2_out[844] <= ~(layer1_out[7776] & layer1_out[7777]);
     layer2_out[845] <= layer1_out[2426] & ~layer1_out[2427];
     layer2_out[846] <= layer1_out[2230];
     layer2_out[847] <= layer1_out[9470] | layer1_out[9471];
     layer2_out[848] <= layer1_out[9894] | layer1_out[9895];
     layer2_out[849] <= layer1_out[6517] & layer1_out[6518];
     layer2_out[850] <= ~layer1_out[8245] | layer1_out[8246];
     layer2_out[851] <= ~(layer1_out[11943] ^ layer1_out[11944]);
     layer2_out[852] <= layer1_out[4617] & ~layer1_out[4618];
     layer2_out[853] <= ~layer1_out[4762] | layer1_out[4763];
     layer2_out[854] <= ~layer1_out[589];
     layer2_out[855] <= layer1_out[10884] & ~layer1_out[10885];
     layer2_out[856] <= 1'b0;
     layer2_out[857] <= layer1_out[8478] & layer1_out[8479];
     layer2_out[858] <= ~(layer1_out[2085] ^ layer1_out[2086]);
     layer2_out[859] <= ~layer1_out[4897] | layer1_out[4898];
     layer2_out[860] <= layer1_out[3778] & ~layer1_out[3779];
     layer2_out[861] <= ~(layer1_out[2140] ^ layer1_out[2141]);
     layer2_out[862] <= ~layer1_out[5492];
     layer2_out[863] <= layer1_out[1180];
     layer2_out[864] <= ~layer1_out[11042] | layer1_out[11043];
     layer2_out[865] <= ~(layer1_out[9219] ^ layer1_out[9220]);
     layer2_out[866] <= ~(layer1_out[5257] & layer1_out[5258]);
     layer2_out[867] <= ~layer1_out[9506];
     layer2_out[868] <= ~layer1_out[10426];
     layer2_out[869] <= layer1_out[9366];
     layer2_out[870] <= layer1_out[7] ^ layer1_out[8];
     layer2_out[871] <= layer1_out[4583];
     layer2_out[872] <= ~(layer1_out[747] & layer1_out[748]);
     layer2_out[873] <= layer1_out[6416] | layer1_out[6417];
     layer2_out[874] <= ~layer1_out[10835];
     layer2_out[875] <= layer1_out[2771] & ~layer1_out[2772];
     layer2_out[876] <= ~layer1_out[7582] | layer1_out[7581];
     layer2_out[877] <= layer1_out[10723] & ~layer1_out[10722];
     layer2_out[878] <= layer1_out[2890] & ~layer1_out[2891];
     layer2_out[879] <= ~layer1_out[4407];
     layer2_out[880] <= ~(layer1_out[11979] & layer1_out[11980]);
     layer2_out[881] <= layer1_out[9];
     layer2_out[882] <= ~(layer1_out[707] & layer1_out[708]);
     layer2_out[883] <= ~(layer1_out[6498] | layer1_out[6499]);
     layer2_out[884] <= layer1_out[8938];
     layer2_out[885] <= ~layer1_out[1174] | layer1_out[1175];
     layer2_out[886] <= ~layer1_out[4778] | layer1_out[4777];
     layer2_out[887] <= ~layer1_out[9661];
     layer2_out[888] <= ~layer1_out[6121];
     layer2_out[889] <= ~layer1_out[2419];
     layer2_out[890] <= ~layer1_out[4945] | layer1_out[4946];
     layer2_out[891] <= layer1_out[11995] ^ layer1_out[11996];
     layer2_out[892] <= ~layer1_out[5346] | layer1_out[5347];
     layer2_out[893] <= layer1_out[9493] ^ layer1_out[9494];
     layer2_out[894] <= ~layer1_out[11221] | layer1_out[11220];
     layer2_out[895] <= ~layer1_out[6942];
     layer2_out[896] <= ~layer1_out[1220];
     layer2_out[897] <= layer1_out[7500];
     layer2_out[898] <= layer1_out[6137] | layer1_out[6138];
     layer2_out[899] <= layer1_out[1824] ^ layer1_out[1825];
     layer2_out[900] <= ~(layer1_out[5529] ^ layer1_out[5530]);
     layer2_out[901] <= layer1_out[9693];
     layer2_out[902] <= ~layer1_out[9406];
     layer2_out[903] <= layer1_out[10188];
     layer2_out[904] <= layer1_out[11971] ^ layer1_out[11972];
     layer2_out[905] <= layer1_out[6981] & ~layer1_out[6980];
     layer2_out[906] <= ~(layer1_out[2484] | layer1_out[2485]);
     layer2_out[907] <= ~layer1_out[381] | layer1_out[382];
     layer2_out[908] <= layer1_out[2248] & layer1_out[2249];
     layer2_out[909] <= layer1_out[1865];
     layer2_out[910] <= layer1_out[8339];
     layer2_out[911] <= layer1_out[10755] ^ layer1_out[10756];
     layer2_out[912] <= layer1_out[5715];
     layer2_out[913] <= layer1_out[1208];
     layer2_out[914] <= ~layer1_out[6526];
     layer2_out[915] <= ~layer1_out[8302] | layer1_out[8303];
     layer2_out[916] <= ~layer1_out[2137];
     layer2_out[917] <= layer1_out[7076] | layer1_out[7077];
     layer2_out[918] <= layer1_out[192];
     layer2_out[919] <= layer1_out[906] & ~layer1_out[907];
     layer2_out[920] <= ~layer1_out[9062];
     layer2_out[921] <= ~(layer1_out[7160] ^ layer1_out[7161]);
     layer2_out[922] <= layer1_out[6426];
     layer2_out[923] <= ~(layer1_out[8778] & layer1_out[8779]);
     layer2_out[924] <= layer1_out[9938];
     layer2_out[925] <= 1'b0;
     layer2_out[926] <= layer1_out[9156];
     layer2_out[927] <= layer1_out[3615] | layer1_out[3616];
     layer2_out[928] <= layer1_out[2182];
     layer2_out[929] <= ~(layer1_out[10797] | layer1_out[10798]);
     layer2_out[930] <= ~(layer1_out[3] & layer1_out[4]);
     layer2_out[931] <= layer1_out[11322] & ~layer1_out[11321];
     layer2_out[932] <= ~layer1_out[11698];
     layer2_out[933] <= ~(layer1_out[5222] & layer1_out[5223]);
     layer2_out[934] <= layer1_out[2913] | layer1_out[2914];
     layer2_out[935] <= ~layer1_out[9467] | layer1_out[9466];
     layer2_out[936] <= layer1_out[9365] & ~layer1_out[9364];
     layer2_out[937] <= ~(layer1_out[8293] ^ layer1_out[8294]);
     layer2_out[938] <= layer1_out[5379];
     layer2_out[939] <= ~layer1_out[10308];
     layer2_out[940] <= layer1_out[5651] | layer1_out[5652];
     layer2_out[941] <= ~layer1_out[199] | layer1_out[200];
     layer2_out[942] <= layer1_out[10767] & layer1_out[10768];
     layer2_out[943] <= 1'b1;
     layer2_out[944] <= layer1_out[7506];
     layer2_out[945] <= layer1_out[10014];
     layer2_out[946] <= ~(layer1_out[1404] | layer1_out[1405]);
     layer2_out[947] <= ~layer1_out[1648];
     layer2_out[948] <= ~layer1_out[6574] | layer1_out[6573];
     layer2_out[949] <= layer1_out[11048] ^ layer1_out[11049];
     layer2_out[950] <= layer1_out[11582] & ~layer1_out[11583];
     layer2_out[951] <= layer1_out[6807];
     layer2_out[952] <= ~layer1_out[2825];
     layer2_out[953] <= ~(layer1_out[3446] ^ layer1_out[3447]);
     layer2_out[954] <= layer1_out[7332] & ~layer1_out[7333];
     layer2_out[955] <= ~layer1_out[7408];
     layer2_out[956] <= layer1_out[11219];
     layer2_out[957] <= layer1_out[6633];
     layer2_out[958] <= ~(layer1_out[2532] | layer1_out[2533]);
     layer2_out[959] <= layer1_out[8282];
     layer2_out[960] <= layer1_out[8210] & ~layer1_out[8209];
     layer2_out[961] <= 1'b1;
     layer2_out[962] <= ~layer1_out[9292];
     layer2_out[963] <= layer1_out[147];
     layer2_out[964] <= ~(layer1_out[4832] | layer1_out[4833]);
     layer2_out[965] <= layer1_out[6970] & ~layer1_out[6971];
     layer2_out[966] <= ~layer1_out[3284] | layer1_out[3285];
     layer2_out[967] <= layer1_out[8097] | layer1_out[8098];
     layer2_out[968] <= layer1_out[10840];
     layer2_out[969] <= layer1_out[4334] & layer1_out[4335];
     layer2_out[970] <= layer1_out[8410] ^ layer1_out[8411];
     layer2_out[971] <= 1'b0;
     layer2_out[972] <= layer1_out[984] & ~layer1_out[983];
     layer2_out[973] <= layer1_out[11897] ^ layer1_out[11898];
     layer2_out[974] <= ~(layer1_out[9060] ^ layer1_out[9061]);
     layer2_out[975] <= layer1_out[3822];
     layer2_out[976] <= layer1_out[8518] ^ layer1_out[8519];
     layer2_out[977] <= layer1_out[2663];
     layer2_out[978] <= ~layer1_out[5160];
     layer2_out[979] <= layer1_out[11832];
     layer2_out[980] <= ~(layer1_out[1116] & layer1_out[1117]);
     layer2_out[981] <= layer1_out[9899] | layer1_out[9900];
     layer2_out[982] <= layer1_out[8932];
     layer2_out[983] <= layer1_out[10713];
     layer2_out[984] <= layer1_out[3528];
     layer2_out[985] <= ~(layer1_out[3629] | layer1_out[3630]);
     layer2_out[986] <= layer1_out[1986];
     layer2_out[987] <= ~layer1_out[3210];
     layer2_out[988] <= ~layer1_out[11102];
     layer2_out[989] <= ~layer1_out[476];
     layer2_out[990] <= ~(layer1_out[7146] & layer1_out[7147]);
     layer2_out[991] <= ~layer1_out[6695] | layer1_out[6694];
     layer2_out[992] <= layer1_out[9217] ^ layer1_out[9218];
     layer2_out[993] <= layer1_out[9251] & ~layer1_out[9252];
     layer2_out[994] <= layer1_out[9637] & ~layer1_out[9638];
     layer2_out[995] <= layer1_out[2034] & layer1_out[2035];
     layer2_out[996] <= layer1_out[11917] & ~layer1_out[11918];
     layer2_out[997] <= ~layer1_out[1952];
     layer2_out[998] <= ~(layer1_out[10613] | layer1_out[10614]);
     layer2_out[999] <= ~layer1_out[9367];
     layer2_out[1000] <= layer1_out[8774] ^ layer1_out[8775];
     layer2_out[1001] <= layer1_out[6187] & layer1_out[6188];
     layer2_out[1002] <= ~(layer1_out[9540] ^ layer1_out[9541]);
     layer2_out[1003] <= ~layer1_out[8863] | layer1_out[8864];
     layer2_out[1004] <= ~layer1_out[11710];
     layer2_out[1005] <= ~layer1_out[8907] | layer1_out[8906];
     layer2_out[1006] <= layer1_out[7948];
     layer2_out[1007] <= ~(layer1_out[10085] & layer1_out[10086]);
     layer2_out[1008] <= layer1_out[8011] & layer1_out[8012];
     layer2_out[1009] <= layer1_out[7348] & ~layer1_out[7347];
     layer2_out[1010] <= layer1_out[3275] & ~layer1_out[3276];
     layer2_out[1011] <= layer1_out[1799] & layer1_out[1800];
     layer2_out[1012] <= ~(layer1_out[11183] ^ layer1_out[11184]);
     layer2_out[1013] <= layer1_out[8402];
     layer2_out[1014] <= ~layer1_out[2981];
     layer2_out[1015] <= ~(layer1_out[829] ^ layer1_out[830]);
     layer2_out[1016] <= layer1_out[5443];
     layer2_out[1017] <= layer1_out[859];
     layer2_out[1018] <= ~layer1_out[3214];
     layer2_out[1019] <= ~layer1_out[4051];
     layer2_out[1020] <= ~layer1_out[8800];
     layer2_out[1021] <= layer1_out[2702] & layer1_out[2703];
     layer2_out[1022] <= layer1_out[10337] & layer1_out[10338];
     layer2_out[1023] <= layer1_out[10198] | layer1_out[10199];
     layer2_out[1024] <= layer1_out[4821] & layer1_out[4822];
     layer2_out[1025] <= layer1_out[6381];
     layer2_out[1026] <= ~layer1_out[1665];
     layer2_out[1027] <= layer1_out[1742] & layer1_out[1743];
     layer2_out[1028] <= ~(layer1_out[5163] & layer1_out[5164]);
     layer2_out[1029] <= ~layer1_out[11415];
     layer2_out[1030] <= layer1_out[10812];
     layer2_out[1031] <= ~layer1_out[3518];
     layer2_out[1032] <= ~(layer1_out[6850] ^ layer1_out[6851]);
     layer2_out[1033] <= layer1_out[11174] ^ layer1_out[11175];
     layer2_out[1034] <= layer1_out[1512] ^ layer1_out[1513];
     layer2_out[1035] <= layer1_out[10581];
     layer2_out[1036] <= ~layer1_out[2685] | layer1_out[2684];
     layer2_out[1037] <= ~layer1_out[5732];
     layer2_out[1038] <= ~layer1_out[3759];
     layer2_out[1039] <= layer1_out[8650] & ~layer1_out[8651];
     layer2_out[1040] <= 1'b1;
     layer2_out[1041] <= layer1_out[6314];
     layer2_out[1042] <= ~layer1_out[5956] | layer1_out[5955];
     layer2_out[1043] <= layer1_out[2222];
     layer2_out[1044] <= ~layer1_out[2040];
     layer2_out[1045] <= ~layer1_out[2241] | layer1_out[2242];
     layer2_out[1046] <= layer1_out[5407];
     layer2_out[1047] <= 1'b0;
     layer2_out[1048] <= layer1_out[8777] & ~layer1_out[8778];
     layer2_out[1049] <= layer1_out[5614] | layer1_out[5615];
     layer2_out[1050] <= layer1_out[4681];
     layer2_out[1051] <= ~layer1_out[3659] | layer1_out[3660];
     layer2_out[1052] <= ~(layer1_out[7382] | layer1_out[7383]);
     layer2_out[1053] <= ~layer1_out[6601] | layer1_out[6602];
     layer2_out[1054] <= layer1_out[10919];
     layer2_out[1055] <= ~layer1_out[11170];
     layer2_out[1056] <= ~(layer1_out[3742] | layer1_out[3743]);
     layer2_out[1057] <= layer1_out[9583];
     layer2_out[1058] <= layer1_out[2541] ^ layer1_out[2542];
     layer2_out[1059] <= layer1_out[9079] | layer1_out[9080];
     layer2_out[1060] <= layer1_out[2378];
     layer2_out[1061] <= layer1_out[9017] & layer1_out[9018];
     layer2_out[1062] <= ~(layer1_out[10922] | layer1_out[10923]);
     layer2_out[1063] <= layer1_out[10335];
     layer2_out[1064] <= ~layer1_out[753];
     layer2_out[1065] <= ~layer1_out[4169];
     layer2_out[1066] <= ~(layer1_out[8544] ^ layer1_out[8545]);
     layer2_out[1067] <= ~(layer1_out[3296] & layer1_out[3297]);
     layer2_out[1068] <= ~(layer1_out[6676] ^ layer1_out[6677]);
     layer2_out[1069] <= layer1_out[10284];
     layer2_out[1070] <= ~layer1_out[315];
     layer2_out[1071] <= 1'b1;
     layer2_out[1072] <= ~(layer1_out[4373] & layer1_out[4374]);
     layer2_out[1073] <= ~layer1_out[231];
     layer2_out[1074] <= layer1_out[6683] ^ layer1_out[6684];
     layer2_out[1075] <= layer1_out[1813];
     layer2_out[1076] <= ~layer1_out[11576];
     layer2_out[1077] <= ~(layer1_out[3000] & layer1_out[3001]);
     layer2_out[1078] <= layer1_out[1356] | layer1_out[1357];
     layer2_out[1079] <= layer1_out[5430] | layer1_out[5431];
     layer2_out[1080] <= layer1_out[9190] & layer1_out[9191];
     layer2_out[1081] <= ~(layer1_out[2638] & layer1_out[2639]);
     layer2_out[1082] <= ~layer1_out[6346];
     layer2_out[1083] <= layer1_out[11149];
     layer2_out[1084] <= ~layer1_out[11342];
     layer2_out[1085] <= ~layer1_out[5130] | layer1_out[5129];
     layer2_out[1086] <= ~(layer1_out[7698] | layer1_out[7699]);
     layer2_out[1087] <= ~(layer1_out[7584] | layer1_out[7585]);
     layer2_out[1088] <= layer1_out[10163];
     layer2_out[1089] <= layer1_out[11064];
     layer2_out[1090] <= ~(layer1_out[10502] & layer1_out[10503]);
     layer2_out[1091] <= ~layer1_out[10345];
     layer2_out[1092] <= layer1_out[2791];
     layer2_out[1093] <= ~(layer1_out[3513] ^ layer1_out[3514]);
     layer2_out[1094] <= layer1_out[2327];
     layer2_out[1095] <= layer1_out[9818];
     layer2_out[1096] <= layer1_out[1568];
     layer2_out[1097] <= layer1_out[3531];
     layer2_out[1098] <= ~layer1_out[6540] | layer1_out[6539];
     layer2_out[1099] <= layer1_out[2881] | layer1_out[2882];
     layer2_out[1100] <= ~layer1_out[1237];
     layer2_out[1101] <= layer1_out[32];
     layer2_out[1102] <= layer1_out[4259] & layer1_out[4260];
     layer2_out[1103] <= layer1_out[3702];
     layer2_out[1104] <= ~layer1_out[10648];
     layer2_out[1105] <= layer1_out[6075];
     layer2_out[1106] <= layer1_out[2305] & ~layer1_out[2306];
     layer2_out[1107] <= ~(layer1_out[11908] | layer1_out[11909]);
     layer2_out[1108] <= layer1_out[4635] & ~layer1_out[4636];
     layer2_out[1109] <= layer1_out[11814] | layer1_out[11815];
     layer2_out[1110] <= layer1_out[6236];
     layer2_out[1111] <= layer1_out[291] | layer1_out[292];
     layer2_out[1112] <= ~(layer1_out[5331] ^ layer1_out[5332]);
     layer2_out[1113] <= ~(layer1_out[11595] & layer1_out[11596]);
     layer2_out[1114] <= ~layer1_out[5559];
     layer2_out[1115] <= layer1_out[7399] & ~layer1_out[7398];
     layer2_out[1116] <= ~layer1_out[10468];
     layer2_out[1117] <= ~(layer1_out[5738] | layer1_out[5739]);
     layer2_out[1118] <= layer1_out[5285];
     layer2_out[1119] <= layer1_out[3383];
     layer2_out[1120] <= ~(layer1_out[7970] ^ layer1_out[7971]);
     layer2_out[1121] <= ~layer1_out[7362];
     layer2_out[1122] <= layer1_out[4716];
     layer2_out[1123] <= ~layer1_out[3120] | layer1_out[3121];
     layer2_out[1124] <= ~layer1_out[1573];
     layer2_out[1125] <= layer1_out[3873] & ~layer1_out[3874];
     layer2_out[1126] <= layer1_out[3177];
     layer2_out[1127] <= layer1_out[2710];
     layer2_out[1128] <= layer1_out[8707];
     layer2_out[1129] <= layer1_out[2763] | layer1_out[2764];
     layer2_out[1130] <= layer1_out[768] & ~layer1_out[769];
     layer2_out[1131] <= layer1_out[4873] | layer1_out[4874];
     layer2_out[1132] <= layer1_out[10985];
     layer2_out[1133] <= 1'b0;
     layer2_out[1134] <= layer1_out[511] & ~layer1_out[512];
     layer2_out[1135] <= ~layer1_out[9756];
     layer2_out[1136] <= layer1_out[344];
     layer2_out[1137] <= layer1_out[5382] ^ layer1_out[5383];
     layer2_out[1138] <= ~layer1_out[10798] | layer1_out[10799];
     layer2_out[1139] <= layer1_out[837] ^ layer1_out[838];
     layer2_out[1140] <= ~layer1_out[4119];
     layer2_out[1141] <= layer1_out[4926] | layer1_out[4927];
     layer2_out[1142] <= layer1_out[7038] | layer1_out[7039];
     layer2_out[1143] <= layer1_out[8312];
     layer2_out[1144] <= layer1_out[6297] & ~layer1_out[6296];
     layer2_out[1145] <= layer1_out[4487] | layer1_out[4488];
     layer2_out[1146] <= ~layer1_out[5104];
     layer2_out[1147] <= layer1_out[1610] & ~layer1_out[1609];
     layer2_out[1148] <= ~(layer1_out[3177] & layer1_out[3178]);
     layer2_out[1149] <= layer1_out[4671];
     layer2_out[1150] <= ~layer1_out[11443];
     layer2_out[1151] <= ~(layer1_out[5990] | layer1_out[5991]);
     layer2_out[1152] <= layer1_out[2875];
     layer2_out[1153] <= ~layer1_out[8110] | layer1_out[8111];
     layer2_out[1154] <= layer1_out[4242] ^ layer1_out[4243];
     layer2_out[1155] <= layer1_out[1377] & ~layer1_out[1378];
     layer2_out[1156] <= layer1_out[9627];
     layer2_out[1157] <= ~layer1_out[2266] | layer1_out[2267];
     layer2_out[1158] <= layer1_out[246];
     layer2_out[1159] <= ~(layer1_out[553] & layer1_out[554]);
     layer2_out[1160] <= ~layer1_out[6824];
     layer2_out[1161] <= layer1_out[1188];
     layer2_out[1162] <= layer1_out[1478];
     layer2_out[1163] <= ~layer1_out[1612];
     layer2_out[1164] <= layer1_out[2456] ^ layer1_out[2457];
     layer2_out[1165] <= layer1_out[3982] & ~layer1_out[3983];
     layer2_out[1166] <= layer1_out[3309] | layer1_out[3310];
     layer2_out[1167] <= layer1_out[7723] & layer1_out[7724];
     layer2_out[1168] <= layer1_out[10247];
     layer2_out[1169] <= layer1_out[5476] & layer1_out[5477];
     layer2_out[1170] <= ~layer1_out[2243] | layer1_out[2244];
     layer2_out[1171] <= layer1_out[11606];
     layer2_out[1172] <= ~(layer1_out[8973] | layer1_out[8974]);
     layer2_out[1173] <= layer1_out[8584] & ~layer1_out[8585];
     layer2_out[1174] <= ~(layer1_out[3412] ^ layer1_out[3413]);
     layer2_out[1175] <= layer1_out[9103] & layer1_out[9104];
     layer2_out[1176] <= layer1_out[10979] & ~layer1_out[10980];
     layer2_out[1177] <= layer1_out[6803];
     layer2_out[1178] <= ~layer1_out[2755];
     layer2_out[1179] <= ~layer1_out[4673];
     layer2_out[1180] <= layer1_out[4357] & layer1_out[4358];
     layer2_out[1181] <= 1'b1;
     layer2_out[1182] <= layer1_out[4435];
     layer2_out[1183] <= layer1_out[4706] ^ layer1_out[4707];
     layer2_out[1184] <= layer1_out[11176] & layer1_out[11177];
     layer2_out[1185] <= ~(layer1_out[8871] & layer1_out[8872]);
     layer2_out[1186] <= layer1_out[10022] ^ layer1_out[10023];
     layer2_out[1187] <= layer1_out[7691];
     layer2_out[1188] <= layer1_out[1696];
     layer2_out[1189] <= ~layer1_out[689] | layer1_out[688];
     layer2_out[1190] <= ~layer1_out[5978];
     layer2_out[1191] <= layer1_out[341];
     layer2_out[1192] <= ~layer1_out[10375];
     layer2_out[1193] <= layer1_out[7312] ^ layer1_out[7313];
     layer2_out[1194] <= ~layer1_out[6069] | layer1_out[6070];
     layer2_out[1195] <= layer1_out[7477];
     layer2_out[1196] <= layer1_out[8588];
     layer2_out[1197] <= layer1_out[5056];
     layer2_out[1198] <= layer1_out[878] & ~layer1_out[879];
     layer2_out[1199] <= layer1_out[9714];
     layer2_out[1200] <= ~(layer1_out[7660] & layer1_out[7661]);
     layer2_out[1201] <= ~layer1_out[864];
     layer2_out[1202] <= ~layer1_out[4575] | layer1_out[4574];
     layer2_out[1203] <= layer1_out[11936];
     layer2_out[1204] <= layer1_out[9700] & ~layer1_out[9701];
     layer2_out[1205] <= ~layer1_out[4365] | layer1_out[4366];
     layer2_out[1206] <= layer1_out[6843];
     layer2_out[1207] <= ~(layer1_out[209] | layer1_out[210]);
     layer2_out[1208] <= ~layer1_out[10242];
     layer2_out[1209] <= layer1_out[10937];
     layer2_out[1210] <= ~(layer1_out[210] | layer1_out[211]);
     layer2_out[1211] <= ~(layer1_out[8470] ^ layer1_out[8471]);
     layer2_out[1212] <= layer1_out[5164] | layer1_out[5165];
     layer2_out[1213] <= layer1_out[10053];
     layer2_out[1214] <= layer1_out[4368];
     layer2_out[1215] <= layer1_out[10846];
     layer2_out[1216] <= ~layer1_out[6066] | layer1_out[6065];
     layer2_out[1217] <= ~layer1_out[131] | layer1_out[130];
     layer2_out[1218] <= layer1_out[191];
     layer2_out[1219] <= layer1_out[6119];
     layer2_out[1220] <= ~(layer1_out[9477] ^ layer1_out[9478]);
     layer2_out[1221] <= ~(layer1_out[9607] & layer1_out[9608]);
     layer2_out[1222] <= ~(layer1_out[2451] ^ layer1_out[2452]);
     layer2_out[1223] <= layer1_out[1068] & layer1_out[1069];
     layer2_out[1224] <= ~(layer1_out[4206] ^ layer1_out[4207]);
     layer2_out[1225] <= ~layer1_out[10405] | layer1_out[10406];
     layer2_out[1226] <= ~layer1_out[1165] | layer1_out[1164];
     layer2_out[1227] <= ~layer1_out[7694];
     layer2_out[1228] <= layer1_out[2530];
     layer2_out[1229] <= layer1_out[3126];
     layer2_out[1230] <= ~layer1_out[2045] | layer1_out[2046];
     layer2_out[1231] <= ~(layer1_out[2288] & layer1_out[2289]);
     layer2_out[1232] <= layer1_out[6505] | layer1_out[6506];
     layer2_out[1233] <= layer1_out[8159] | layer1_out[8160];
     layer2_out[1234] <= ~layer1_out[10475] | layer1_out[10474];
     layer2_out[1235] <= layer1_out[6577] ^ layer1_out[6578];
     layer2_out[1236] <= ~layer1_out[11064];
     layer2_out[1237] <= layer1_out[10444] | layer1_out[10445];
     layer2_out[1238] <= layer1_out[8127] & ~layer1_out[8128];
     layer2_out[1239] <= ~layer1_out[2535] | layer1_out[2534];
     layer2_out[1240] <= layer1_out[9321] | layer1_out[9322];
     layer2_out[1241] <= layer1_out[344];
     layer2_out[1242] <= layer1_out[1417];
     layer2_out[1243] <= layer1_out[3848];
     layer2_out[1244] <= layer1_out[4813] & ~layer1_out[4812];
     layer2_out[1245] <= layer1_out[3941] & ~layer1_out[3940];
     layer2_out[1246] <= ~(layer1_out[3094] | layer1_out[3095]);
     layer2_out[1247] <= ~layer1_out[1714] | layer1_out[1715];
     layer2_out[1248] <= layer1_out[4996];
     layer2_out[1249] <= layer1_out[4784];
     layer2_out[1250] <= ~(layer1_out[5502] | layer1_out[5503]);
     layer2_out[1251] <= layer1_out[6410] & ~layer1_out[6409];
     layer2_out[1252] <= ~layer1_out[10892] | layer1_out[10893];
     layer2_out[1253] <= layer1_out[1696] | layer1_out[1697];
     layer2_out[1254] <= layer1_out[7212] & ~layer1_out[7211];
     layer2_out[1255] <= layer1_out[8741];
     layer2_out[1256] <= 1'b1;
     layer2_out[1257] <= ~layer1_out[6687];
     layer2_out[1258] <= ~layer1_out[6699];
     layer2_out[1259] <= ~layer1_out[1532];
     layer2_out[1260] <= layer1_out[11758] & ~layer1_out[11757];
     layer2_out[1261] <= ~layer1_out[4370];
     layer2_out[1262] <= 1'b0;
     layer2_out[1263] <= layer1_out[2291] & layer1_out[2292];
     layer2_out[1264] <= ~layer1_out[3821] | layer1_out[3820];
     layer2_out[1265] <= layer1_out[7837] & ~layer1_out[7838];
     layer2_out[1266] <= ~layer1_out[4823];
     layer2_out[1267] <= ~layer1_out[6585] | layer1_out[6584];
     layer2_out[1268] <= layer1_out[9842];
     layer2_out[1269] <= layer1_out[3582] & ~layer1_out[3581];
     layer2_out[1270] <= ~(layer1_out[212] | layer1_out[213]);
     layer2_out[1271] <= layer1_out[7890] ^ layer1_out[7891];
     layer2_out[1272] <= ~layer1_out[1755] | layer1_out[1756];
     layer2_out[1273] <= layer1_out[4850] & layer1_out[4851];
     layer2_out[1274] <= ~layer1_out[7930] | layer1_out[7931];
     layer2_out[1275] <= ~layer1_out[1740];
     layer2_out[1276] <= ~layer1_out[3469];
     layer2_out[1277] <= layer1_out[774];
     layer2_out[1278] <= ~layer1_out[1303];
     layer2_out[1279] <= ~(layer1_out[10916] | layer1_out[10917]);
     layer2_out[1280] <= ~(layer1_out[6099] & layer1_out[6100]);
     layer2_out[1281] <= ~layer1_out[6832] | layer1_out[6831];
     layer2_out[1282] <= 1'b0;
     layer2_out[1283] <= ~layer1_out[2101] | layer1_out[2102];
     layer2_out[1284] <= ~layer1_out[1130] | layer1_out[1129];
     layer2_out[1285] <= layer1_out[2917] & layer1_out[2918];
     layer2_out[1286] <= layer1_out[6220] & layer1_out[6221];
     layer2_out[1287] <= layer1_out[9513] & ~layer1_out[9514];
     layer2_out[1288] <= ~(layer1_out[7154] | layer1_out[7155]);
     layer2_out[1289] <= ~(layer1_out[10270] & layer1_out[10271]);
     layer2_out[1290] <= ~layer1_out[2955];
     layer2_out[1291] <= layer1_out[2977] | layer1_out[2978];
     layer2_out[1292] <= layer1_out[4749];
     layer2_out[1293] <= layer1_out[5183];
     layer2_out[1294] <= ~layer1_out[11498];
     layer2_out[1295] <= ~layer1_out[10696];
     layer2_out[1296] <= layer1_out[11721];
     layer2_out[1297] <= layer1_out[2139] & ~layer1_out[2138];
     layer2_out[1298] <= layer1_out[10663] | layer1_out[10664];
     layer2_out[1299] <= layer1_out[4355] | layer1_out[4356];
     layer2_out[1300] <= ~layer1_out[1375] | layer1_out[1376];
     layer2_out[1301] <= layer1_out[3440] & layer1_out[3441];
     layer2_out[1302] <= layer1_out[6612] | layer1_out[6613];
     layer2_out[1303] <= ~layer1_out[5872] | layer1_out[5873];
     layer2_out[1304] <= ~layer1_out[10524];
     layer2_out[1305] <= layer1_out[5640];
     layer2_out[1306] <= ~layer1_out[6256] | layer1_out[6255];
     layer2_out[1307] <= ~layer1_out[1168];
     layer2_out[1308] <= layer1_out[4080];
     layer2_out[1309] <= ~layer1_out[1298] | layer1_out[1297];
     layer2_out[1310] <= layer1_out[4977] & layer1_out[4978];
     layer2_out[1311] <= ~layer1_out[6308] | layer1_out[6309];
     layer2_out[1312] <= layer1_out[187] | layer1_out[188];
     layer2_out[1313] <= layer1_out[7103] | layer1_out[7104];
     layer2_out[1314] <= layer1_out[11596] ^ layer1_out[11597];
     layer2_out[1315] <= ~layer1_out[9675];
     layer2_out[1316] <= ~layer1_out[1302];
     layer2_out[1317] <= ~(layer1_out[6941] ^ layer1_out[6942]);
     layer2_out[1318] <= layer1_out[5023] | layer1_out[5024];
     layer2_out[1319] <= ~(layer1_out[10278] ^ layer1_out[10279]);
     layer2_out[1320] <= ~layer1_out[7713];
     layer2_out[1321] <= ~layer1_out[2475];
     layer2_out[1322] <= layer1_out[11296];
     layer2_out[1323] <= ~(layer1_out[7414] & layer1_out[7415]);
     layer2_out[1324] <= layer1_out[5746] & layer1_out[5747];
     layer2_out[1325] <= layer1_out[7220];
     layer2_out[1326] <= layer1_out[11541] & ~layer1_out[11540];
     layer2_out[1327] <= layer1_out[6868];
     layer2_out[1328] <= layer1_out[4598] & layer1_out[4599];
     layer2_out[1329] <= layer1_out[7452] | layer1_out[7453];
     layer2_out[1330] <= ~(layer1_out[10471] ^ layer1_out[10472]);
     layer2_out[1331] <= 1'b1;
     layer2_out[1332] <= ~layer1_out[925];
     layer2_out[1333] <= ~layer1_out[7736] | layer1_out[7737];
     layer2_out[1334] <= layer1_out[59] ^ layer1_out[60];
     layer2_out[1335] <= ~(layer1_out[3529] ^ layer1_out[3530]);
     layer2_out[1336] <= layer1_out[9319];
     layer2_out[1337] <= ~(layer1_out[5475] & layer1_out[5476]);
     layer2_out[1338] <= ~layer1_out[10412] | layer1_out[10413];
     layer2_out[1339] <= ~(layer1_out[5069] ^ layer1_out[5070]);
     layer2_out[1340] <= layer1_out[1244] | layer1_out[1245];
     layer2_out[1341] <= ~(layer1_out[11559] | layer1_out[11560]);
     layer2_out[1342] <= layer1_out[446];
     layer2_out[1343] <= ~(layer1_out[11756] ^ layer1_out[11757]);
     layer2_out[1344] <= layer1_out[5649] | layer1_out[5650];
     layer2_out[1345] <= layer1_out[7717] & ~layer1_out[7716];
     layer2_out[1346] <= layer1_out[3882];
     layer2_out[1347] <= layer1_out[3766] ^ layer1_out[3767];
     layer2_out[1348] <= ~layer1_out[91] | layer1_out[90];
     layer2_out[1349] <= layer1_out[11205] & layer1_out[11206];
     layer2_out[1350] <= layer1_out[10960];
     layer2_out[1351] <= layer1_out[8070] | layer1_out[8071];
     layer2_out[1352] <= ~(layer1_out[195] & layer1_out[196]);
     layer2_out[1353] <= layer1_out[8026] & ~layer1_out[8027];
     layer2_out[1354] <= ~layer1_out[4424] | layer1_out[4425];
     layer2_out[1355] <= ~layer1_out[5985] | layer1_out[5984];
     layer2_out[1356] <= layer1_out[2310] | layer1_out[2311];
     layer2_out[1357] <= ~(layer1_out[3959] | layer1_out[3960]);
     layer2_out[1358] <= layer1_out[2510];
     layer2_out[1359] <= layer1_out[5212];
     layer2_out[1360] <= ~layer1_out[4463];
     layer2_out[1361] <= layer1_out[9709];
     layer2_out[1362] <= ~(layer1_out[4492] & layer1_out[4493]);
     layer2_out[1363] <= ~(layer1_out[4452] | layer1_out[4453]);
     layer2_out[1364] <= ~layer1_out[685] | layer1_out[686];
     layer2_out[1365] <= ~(layer1_out[10267] | layer1_out[10268]);
     layer2_out[1366] <= layer1_out[5352];
     layer2_out[1367] <= ~layer1_out[6250];
     layer2_out[1368] <= layer1_out[2325] & ~layer1_out[2326];
     layer2_out[1369] <= layer1_out[10488] & layer1_out[10489];
     layer2_out[1370] <= ~(layer1_out[9212] | layer1_out[9213]);
     layer2_out[1371] <= layer1_out[8200] & ~layer1_out[8199];
     layer2_out[1372] <= layer1_out[2574] & ~layer1_out[2573];
     layer2_out[1373] <= ~layer1_out[3797];
     layer2_out[1374] <= layer1_out[5607];
     layer2_out[1375] <= layer1_out[4750] | layer1_out[4751];
     layer2_out[1376] <= layer1_out[10420] & ~layer1_out[10421];
     layer2_out[1377] <= ~layer1_out[1334];
     layer2_out[1378] <= layer1_out[11248];
     layer2_out[1379] <= ~layer1_out[6326] | layer1_out[6325];
     layer2_out[1380] <= layer1_out[8987] | layer1_out[8988];
     layer2_out[1381] <= ~(layer1_out[6698] ^ layer1_out[6699]);
     layer2_out[1382] <= layer1_out[867] ^ layer1_out[868];
     layer2_out[1383] <= ~layer1_out[9323];
     layer2_out[1384] <= layer1_out[8782] & ~layer1_out[8783];
     layer2_out[1385] <= ~layer1_out[3869];
     layer2_out[1386] <= 1'b0;
     layer2_out[1387] <= layer1_out[5169] & ~layer1_out[5170];
     layer2_out[1388] <= layer1_out[8602] & ~layer1_out[8601];
     layer2_out[1389] <= ~(layer1_out[6165] | layer1_out[6166]);
     layer2_out[1390] <= ~layer1_out[5745] | layer1_out[5746];
     layer2_out[1391] <= layer1_out[9391] & ~layer1_out[9390];
     layer2_out[1392] <= layer1_out[9526];
     layer2_out[1393] <= layer1_out[1442];
     layer2_out[1394] <= layer1_out[1458];
     layer2_out[1395] <= layer1_out[11056] ^ layer1_out[11057];
     layer2_out[1396] <= ~layer1_out[2579];
     layer2_out[1397] <= ~layer1_out[8099] | layer1_out[8098];
     layer2_out[1398] <= layer1_out[8244];
     layer2_out[1399] <= layer1_out[1192] & layer1_out[1193];
     layer2_out[1400] <= ~layer1_out[3693];
     layer2_out[1401] <= layer1_out[93] & ~layer1_out[92];
     layer2_out[1402] <= ~layer1_out[4923];
     layer2_out[1403] <= ~(layer1_out[7658] & layer1_out[7659]);
     layer2_out[1404] <= ~layer1_out[3510];
     layer2_out[1405] <= layer1_out[8220] & layer1_out[8221];
     layer2_out[1406] <= 1'b0;
     layer2_out[1407] <= ~layer1_out[6586] | layer1_out[6585];
     layer2_out[1408] <= 1'b0;
     layer2_out[1409] <= ~(layer1_out[4524] | layer1_out[4525]);
     layer2_out[1410] <= layer1_out[10743] & layer1_out[10744];
     layer2_out[1411] <= layer1_out[5674] & ~layer1_out[5675];
     layer2_out[1412] <= layer1_out[2879] | layer1_out[2880];
     layer2_out[1413] <= ~layer1_out[8670];
     layer2_out[1414] <= layer1_out[7729];
     layer2_out[1415] <= ~(layer1_out[3115] | layer1_out[3116]);
     layer2_out[1416] <= layer1_out[3205];
     layer2_out[1417] <= layer1_out[5638];
     layer2_out[1418] <= layer1_out[2758] & ~layer1_out[2757];
     layer2_out[1419] <= ~layer1_out[6432];
     layer2_out[1420] <= layer1_out[7822];
     layer2_out[1421] <= ~(layer1_out[7790] | layer1_out[7791]);
     layer2_out[1422] <= ~layer1_out[4872] | layer1_out[4871];
     layer2_out[1423] <= ~(layer1_out[7979] & layer1_out[7980]);
     layer2_out[1424] <= ~layer1_out[8579];
     layer2_out[1425] <= ~layer1_out[10646];
     layer2_out[1426] <= layer1_out[2858];
     layer2_out[1427] <= layer1_out[4506];
     layer2_out[1428] <= layer1_out[4989] & ~layer1_out[4988];
     layer2_out[1429] <= ~layer1_out[7551] | layer1_out[7552];
     layer2_out[1430] <= layer1_out[8271];
     layer2_out[1431] <= ~layer1_out[1489];
     layer2_out[1432] <= ~layer1_out[11545] | layer1_out[11546];
     layer2_out[1433] <= layer1_out[4283] & ~layer1_out[4284];
     layer2_out[1434] <= ~layer1_out[3704];
     layer2_out[1435] <= ~(layer1_out[11583] ^ layer1_out[11584]);
     layer2_out[1436] <= layer1_out[2844] & ~layer1_out[2843];
     layer2_out[1437] <= layer1_out[5870] | layer1_out[5871];
     layer2_out[1438] <= ~layer1_out[4438];
     layer2_out[1439] <= layer1_out[6967] & ~layer1_out[6968];
     layer2_out[1440] <= ~(layer1_out[5125] & layer1_out[5126]);
     layer2_out[1441] <= layer1_out[8090] & ~layer1_out[8091];
     layer2_out[1442] <= ~(layer1_out[4433] ^ layer1_out[4434]);
     layer2_out[1443] <= layer1_out[1921] & ~layer1_out[1922];
     layer2_out[1444] <= ~(layer1_out[2216] & layer1_out[2217]);
     layer2_out[1445] <= ~(layer1_out[8378] | layer1_out[8379]);
     layer2_out[1446] <= layer1_out[6976] | layer1_out[6977];
     layer2_out[1447] <= ~layer1_out[4389];
     layer2_out[1448] <= layer1_out[6759];
     layer2_out[1449] <= ~(layer1_out[3693] & layer1_out[3694]);
     layer2_out[1450] <= layer1_out[1428];
     layer2_out[1451] <= ~layer1_out[1543];
     layer2_out[1452] <= layer1_out[5665];
     layer2_out[1453] <= layer1_out[7210] & ~layer1_out[7211];
     layer2_out[1454] <= ~layer1_out[10237];
     layer2_out[1455] <= ~layer1_out[4577] | layer1_out[4576];
     layer2_out[1456] <= layer1_out[6392];
     layer2_out[1457] <= ~(layer1_out[5485] | layer1_out[5486]);
     layer2_out[1458] <= ~layer1_out[10192];
     layer2_out[1459] <= ~layer1_out[6229] | layer1_out[6230];
     layer2_out[1460] <= layer1_out[6054] & ~layer1_out[6053];
     layer2_out[1461] <= layer1_out[41];
     layer2_out[1462] <= layer1_out[4145] & ~layer1_out[4144];
     layer2_out[1463] <= layer1_out[10121] & ~layer1_out[10122];
     layer2_out[1464] <= layer1_out[1510];
     layer2_out[1465] <= ~(layer1_out[4392] & layer1_out[4393]);
     layer2_out[1466] <= ~(layer1_out[10247] & layer1_out[10248]);
     layer2_out[1467] <= ~(layer1_out[3122] & layer1_out[3123]);
     layer2_out[1468] <= ~layer1_out[5234];
     layer2_out[1469] <= layer1_out[4949] & ~layer1_out[4950];
     layer2_out[1470] <= ~layer1_out[5519];
     layer2_out[1471] <= layer1_out[3964] & ~layer1_out[3963];
     layer2_out[1472] <= layer1_out[1117] & layer1_out[1118];
     layer2_out[1473] <= layer1_out[7731] ^ layer1_out[7732];
     layer2_out[1474] <= layer1_out[1401];
     layer2_out[1475] <= layer1_out[8041] & layer1_out[8042];
     layer2_out[1476] <= layer1_out[2520];
     layer2_out[1477] <= layer1_out[8184] & layer1_out[8185];
     layer2_out[1478] <= layer1_out[7619];
     layer2_out[1479] <= layer1_out[6757] & layer1_out[6758];
     layer2_out[1480] <= layer1_out[365] & ~layer1_out[366];
     layer2_out[1481] <= ~(layer1_out[9837] ^ layer1_out[9838]);
     layer2_out[1482] <= layer1_out[2559];
     layer2_out[1483] <= layer1_out[7850] ^ layer1_out[7851];
     layer2_out[1484] <= ~(layer1_out[5010] & layer1_out[5011]);
     layer2_out[1485] <= layer1_out[5052];
     layer2_out[1486] <= ~layer1_out[1762];
     layer2_out[1487] <= layer1_out[6457] | layer1_out[6458];
     layer2_out[1488] <= layer1_out[1332] & ~layer1_out[1331];
     layer2_out[1489] <= layer1_out[9857] & ~layer1_out[9858];
     layer2_out[1490] <= layer1_out[6575];
     layer2_out[1491] <= ~layer1_out[10781];
     layer2_out[1492] <= ~layer1_out[10522];
     layer2_out[1493] <= ~(layer1_out[824] | layer1_out[825]);
     layer2_out[1494] <= ~(layer1_out[10895] & layer1_out[10896]);
     layer2_out[1495] <= layer1_out[8734] & ~layer1_out[8733];
     layer2_out[1496] <= ~(layer1_out[1418] | layer1_out[1419]);
     layer2_out[1497] <= layer1_out[10071] & ~layer1_out[10072];
     layer2_out[1498] <= ~(layer1_out[1743] ^ layer1_out[1744]);
     layer2_out[1499] <= ~layer1_out[28];
     layer2_out[1500] <= layer1_out[9129] & ~layer1_out[9128];
     layer2_out[1501] <= ~layer1_out[7368];
     layer2_out[1502] <= layer1_out[1764] | layer1_out[1765];
     layer2_out[1503] <= ~layer1_out[7778];
     layer2_out[1504] <= layer1_out[1505] | layer1_out[1506];
     layer2_out[1505] <= layer1_out[1444];
     layer2_out[1506] <= ~(layer1_out[11566] ^ layer1_out[11567]);
     layer2_out[1507] <= ~layer1_out[6528] | layer1_out[6527];
     layer2_out[1508] <= layer1_out[1948] ^ layer1_out[1949];
     layer2_out[1509] <= layer1_out[9953] | layer1_out[9954];
     layer2_out[1510] <= layer1_out[3251] ^ layer1_out[3252];
     layer2_out[1511] <= layer1_out[9371];
     layer2_out[1512] <= layer1_out[6456];
     layer2_out[1513] <= ~(layer1_out[386] | layer1_out[387]);
     layer2_out[1514] <= ~layer1_out[9976];
     layer2_out[1515] <= layer1_out[1945];
     layer2_out[1516] <= ~(layer1_out[8689] ^ layer1_out[8690]);
     layer2_out[1517] <= layer1_out[9529] & layer1_out[9530];
     layer2_out[1518] <= ~(layer1_out[5948] | layer1_out[5949]);
     layer2_out[1519] <= ~layer1_out[156];
     layer2_out[1520] <= ~layer1_out[7279] | layer1_out[7280];
     layer2_out[1521] <= layer1_out[11655];
     layer2_out[1522] <= layer1_out[5248] | layer1_out[5249];
     layer2_out[1523] <= layer1_out[6578] ^ layer1_out[6579];
     layer2_out[1524] <= layer1_out[10590] ^ layer1_out[10591];
     layer2_out[1525] <= ~(layer1_out[3638] | layer1_out[3639]);
     layer2_out[1526] <= ~layer1_out[9215];
     layer2_out[1527] <= layer1_out[11706];
     layer2_out[1528] <= layer1_out[1897] & ~layer1_out[1896];
     layer2_out[1529] <= ~(layer1_out[6715] | layer1_out[6716]);
     layer2_out[1530] <= layer1_out[6192] ^ layer1_out[6193];
     layer2_out[1531] <= layer1_out[10417] | layer1_out[10418];
     layer2_out[1532] <= ~layer1_out[5851] | layer1_out[5852];
     layer2_out[1533] <= layer1_out[2406];
     layer2_out[1534] <= ~(layer1_out[1556] ^ layer1_out[1557]);
     layer2_out[1535] <= ~layer1_out[2211];
     layer2_out[1536] <= layer1_out[2098];
     layer2_out[1537] <= ~layer1_out[7170];
     layer2_out[1538] <= ~layer1_out[2446];
     layer2_out[1539] <= layer1_out[134];
     layer2_out[1540] <= ~layer1_out[3603] | layer1_out[3604];
     layer2_out[1541] <= ~layer1_out[7922];
     layer2_out[1542] <= layer1_out[9874];
     layer2_out[1543] <= layer1_out[4655] & layer1_out[4656];
     layer2_out[1544] <= ~(layer1_out[10259] & layer1_out[10260]);
     layer2_out[1545] <= layer1_out[5281] | layer1_out[5282];
     layer2_out[1546] <= layer1_out[2997];
     layer2_out[1547] <= layer1_out[8856];
     layer2_out[1548] <= ~(layer1_out[8299] | layer1_out[8300]);
     layer2_out[1549] <= ~layer1_out[522];
     layer2_out[1550] <= layer1_out[8892] & layer1_out[8893];
     layer2_out[1551] <= ~(layer1_out[10239] | layer1_out[10240]);
     layer2_out[1552] <= layer1_out[9198] ^ layer1_out[9199];
     layer2_out[1553] <= ~layer1_out[3904] | layer1_out[3905];
     layer2_out[1554] <= ~layer1_out[2500];
     layer2_out[1555] <= ~(layer1_out[1401] ^ layer1_out[1402]);
     layer2_out[1556] <= layer1_out[4605] & layer1_out[4606];
     layer2_out[1557] <= layer1_out[4913] ^ layer1_out[4914];
     layer2_out[1558] <= layer1_out[1494] | layer1_out[1495];
     layer2_out[1559] <= ~layer1_out[9498];
     layer2_out[1560] <= ~layer1_out[773];
     layer2_out[1561] <= layer1_out[9996] ^ layer1_out[9997];
     layer2_out[1562] <= ~layer1_out[5061] | layer1_out[5060];
     layer2_out[1563] <= ~layer1_out[8877] | layer1_out[8878];
     layer2_out[1564] <= layer1_out[10625];
     layer2_out[1565] <= ~layer1_out[7389];
     layer2_out[1566] <= layer1_out[1781];
     layer2_out[1567] <= layer1_out[10833] | layer1_out[10834];
     layer2_out[1568] <= ~layer1_out[11684];
     layer2_out[1569] <= layer1_out[11387];
     layer2_out[1570] <= layer1_out[4148] & ~layer1_out[4147];
     layer2_out[1571] <= ~layer1_out[5137];
     layer2_out[1572] <= ~(layer1_out[11863] & layer1_out[11864]);
     layer2_out[1573] <= ~layer1_out[11003];
     layer2_out[1574] <= ~(layer1_out[8158] | layer1_out[8159]);
     layer2_out[1575] <= layer1_out[8409];
     layer2_out[1576] <= ~layer1_out[10852];
     layer2_out[1577] <= layer1_out[4319] | layer1_out[4320];
     layer2_out[1578] <= layer1_out[489];
     layer2_out[1579] <= layer1_out[7422] | layer1_out[7423];
     layer2_out[1580] <= ~(layer1_out[3755] | layer1_out[3756]);
     layer2_out[1581] <= ~(layer1_out[5105] ^ layer1_out[5106]);
     layer2_out[1582] <= layer1_out[8395] & ~layer1_out[8394];
     layer2_out[1583] <= layer1_out[1593] & ~layer1_out[1592];
     layer2_out[1584] <= ~layer1_out[9837] | layer1_out[9836];
     layer2_out[1585] <= ~layer1_out[4771];
     layer2_out[1586] <= ~(layer1_out[9696] & layer1_out[9697]);
     layer2_out[1587] <= ~(layer1_out[4339] & layer1_out[4340]);
     layer2_out[1588] <= layer1_out[4231] | layer1_out[4232];
     layer2_out[1589] <= layer1_out[9622] & ~layer1_out[9621];
     layer2_out[1590] <= layer1_out[7999];
     layer2_out[1591] <= ~(layer1_out[6927] | layer1_out[6928]);
     layer2_out[1592] <= layer1_out[1703] & layer1_out[1704];
     layer2_out[1593] <= ~layer1_out[4240] | layer1_out[4241];
     layer2_out[1594] <= ~(layer1_out[889] & layer1_out[890]);
     layer2_out[1595] <= ~layer1_out[7269];
     layer2_out[1596] <= ~(layer1_out[4676] & layer1_out[4677]);
     layer2_out[1597] <= ~layer1_out[11122];
     layer2_out[1598] <= ~layer1_out[549];
     layer2_out[1599] <= ~(layer1_out[5108] | layer1_out[5109]);
     layer2_out[1600] <= layer1_out[293] & ~layer1_out[294];
     layer2_out[1601] <= ~(layer1_out[6592] ^ layer1_out[6593]);
     layer2_out[1602] <= ~layer1_out[10693];
     layer2_out[1603] <= ~(layer1_out[5204] & layer1_out[5205]);
     layer2_out[1604] <= layer1_out[3436];
     layer2_out[1605] <= ~(layer1_out[4646] & layer1_out[4647]);
     layer2_out[1606] <= 1'b0;
     layer2_out[1607] <= layer1_out[7200];
     layer2_out[1608] <= layer1_out[1133];
     layer2_out[1609] <= layer1_out[6829] & layer1_out[6830];
     layer2_out[1610] <= layer1_out[1867] & ~layer1_out[1866];
     layer2_out[1611] <= layer1_out[10556] & layer1_out[10557];
     layer2_out[1612] <= layer1_out[9955];
     layer2_out[1613] <= ~layer1_out[211];
     layer2_out[1614] <= layer1_out[831] ^ layer1_out[832];
     layer2_out[1615] <= layer1_out[4288];
     layer2_out[1616] <= layer1_out[8361] & layer1_out[8362];
     layer2_out[1617] <= layer1_out[6125] & ~layer1_out[6126];
     layer2_out[1618] <= ~layer1_out[8996];
     layer2_out[1619] <= ~layer1_out[8927];
     layer2_out[1620] <= ~layer1_out[10214];
     layer2_out[1621] <= ~layer1_out[3783];
     layer2_out[1622] <= ~layer1_out[7177];
     layer2_out[1623] <= layer1_out[6004] & ~layer1_out[6005];
     layer2_out[1624] <= ~(layer1_out[3893] & layer1_out[3894]);
     layer2_out[1625] <= ~layer1_out[5809];
     layer2_out[1626] <= ~(layer1_out[7436] & layer1_out[7437]);
     layer2_out[1627] <= layer1_out[6784];
     layer2_out[1628] <= layer1_out[5115];
     layer2_out[1629] <= ~layer1_out[4079];
     layer2_out[1630] <= 1'b1;
     layer2_out[1631] <= layer1_out[1029] ^ layer1_out[1030];
     layer2_out[1632] <= layer1_out[11738];
     layer2_out[1633] <= layer1_out[5581] & ~layer1_out[5580];
     layer2_out[1634] <= ~layer1_out[10392];
     layer2_out[1635] <= ~(layer1_out[779] ^ layer1_out[780]);
     layer2_out[1636] <= ~(layer1_out[2449] ^ layer1_out[2450]);
     layer2_out[1637] <= ~(layer1_out[10830] ^ layer1_out[10831]);
     layer2_out[1638] <= layer1_out[6246];
     layer2_out[1639] <= ~(layer1_out[1840] ^ layer1_out[1841]);
     layer2_out[1640] <= layer1_out[2220];
     layer2_out[1641] <= layer1_out[9462] & ~layer1_out[9463];
     layer2_out[1642] <= layer1_out[875] | layer1_out[876];
     layer2_out[1643] <= ~layer1_out[1868] | layer1_out[1869];
     layer2_out[1644] <= layer1_out[10883];
     layer2_out[1645] <= ~layer1_out[9831];
     layer2_out[1646] <= layer1_out[4755] & layer1_out[4756];
     layer2_out[1647] <= ~layer1_out[5503];
     layer2_out[1648] <= layer1_out[3867] | layer1_out[3868];
     layer2_out[1649] <= layer1_out[1224];
     layer2_out[1650] <= layer1_out[4472] & ~layer1_out[4471];
     layer2_out[1651] <= ~layer1_out[10481];
     layer2_out[1652] <= ~(layer1_out[498] & layer1_out[499]);
     layer2_out[1653] <= ~layer1_out[5467] | layer1_out[5466];
     layer2_out[1654] <= ~layer1_out[1080] | layer1_out[1079];
     layer2_out[1655] <= layer1_out[3494];
     layer2_out[1656] <= layer1_out[6167] & ~layer1_out[6168];
     layer2_out[1657] <= layer1_out[6945] ^ layer1_out[6946];
     layer2_out[1658] <= ~(layer1_out[1607] & layer1_out[1608]);
     layer2_out[1659] <= ~layer1_out[2548] | layer1_out[2547];
     layer2_out[1660] <= layer1_out[395] ^ layer1_out[396];
     layer2_out[1661] <= layer1_out[514] ^ layer1_out[515];
     layer2_out[1662] <= 1'b0;
     layer2_out[1663] <= layer1_out[1882];
     layer2_out[1664] <= layer1_out[4080] & ~layer1_out[4079];
     layer2_out[1665] <= ~layer1_out[1103];
     layer2_out[1666] <= ~layer1_out[923];
     layer2_out[1667] <= layer1_out[9222];
     layer2_out[1668] <= ~(layer1_out[72] ^ layer1_out[73]);
     layer2_out[1669] <= ~layer1_out[7784];
     layer2_out[1670] <= layer1_out[11744] & layer1_out[11745];
     layer2_out[1671] <= layer1_out[7127] & layer1_out[7128];
     layer2_out[1672] <= ~(layer1_out[7543] ^ layer1_out[7544]);
     layer2_out[1673] <= ~(layer1_out[6360] | layer1_out[6361]);
     layer2_out[1674] <= layer1_out[4207] | layer1_out[4208];
     layer2_out[1675] <= ~layer1_out[5026];
     layer2_out[1676] <= ~layer1_out[4371];
     layer2_out[1677] <= layer1_out[6545] & ~layer1_out[6544];
     layer2_out[1678] <= layer1_out[7152] & ~layer1_out[7151];
     layer2_out[1679] <= ~layer1_out[11806];
     layer2_out[1680] <= ~(layer1_out[1875] & layer1_out[1876]);
     layer2_out[1681] <= ~layer1_out[11431];
     layer2_out[1682] <= layer1_out[2374] & ~layer1_out[2375];
     layer2_out[1683] <= layer1_out[8561];
     layer2_out[1684] <= layer1_out[9562];
     layer2_out[1685] <= ~layer1_out[4238];
     layer2_out[1686] <= ~layer1_out[10733];
     layer2_out[1687] <= layer1_out[3849] & ~layer1_out[3850];
     layer2_out[1688] <= layer1_out[9979] & layer1_out[9980];
     layer2_out[1689] <= ~layer1_out[11132] | layer1_out[11133];
     layer2_out[1690] <= layer1_out[3191] & ~layer1_out[3192];
     layer2_out[1691] <= layer1_out[3583] | layer1_out[3584];
     layer2_out[1692] <= layer1_out[11029];
     layer2_out[1693] <= ~(layer1_out[3990] ^ layer1_out[3991]);
     layer2_out[1694] <= 1'b1;
     layer2_out[1695] <= layer1_out[4042] & ~layer1_out[4043];
     layer2_out[1696] <= layer1_out[8176] & layer1_out[8177];
     layer2_out[1697] <= layer1_out[519] & ~layer1_out[520];
     layer2_out[1698] <= ~layer1_out[2848] | layer1_out[2847];
     layer2_out[1699] <= ~layer1_out[5763];
     layer2_out[1700] <= ~layer1_out[11679] | layer1_out[11678];
     layer2_out[1701] <= ~layer1_out[9086];
     layer2_out[1702] <= ~layer1_out[87];
     layer2_out[1703] <= ~(layer1_out[10981] & layer1_out[10982]);
     layer2_out[1704] <= ~(layer1_out[4070] | layer1_out[4071]);
     layer2_out[1705] <= layer1_out[4050] | layer1_out[4051];
     layer2_out[1706] <= ~layer1_out[1771];
     layer2_out[1707] <= layer1_out[10759];
     layer2_out[1708] <= layer1_out[10458];
     layer2_out[1709] <= ~(layer1_out[822] | layer1_out[823]);
     layer2_out[1710] <= layer1_out[8676] & layer1_out[8677];
     layer2_out[1711] <= ~layer1_out[7072];
     layer2_out[1712] <= ~(layer1_out[4325] & layer1_out[4326]);
     layer2_out[1713] <= ~layer1_out[813];
     layer2_out[1714] <= layer1_out[10428] & ~layer1_out[10427];
     layer2_out[1715] <= ~(layer1_out[5079] ^ layer1_out[5080]);
     layer2_out[1716] <= ~(layer1_out[10484] | layer1_out[10485]);
     layer2_out[1717] <= ~(layer1_out[10542] | layer1_out[10543]);
     layer2_out[1718] <= layer1_out[4251] | layer1_out[4252];
     layer2_out[1719] <= ~layer1_out[2319];
     layer2_out[1720] <= ~layer1_out[11127];
     layer2_out[1721] <= ~(layer1_out[4726] & layer1_out[4727]);
     layer2_out[1722] <= layer1_out[5287] & layer1_out[5288];
     layer2_out[1723] <= layer1_out[9611];
     layer2_out[1724] <= ~layer1_out[943];
     layer2_out[1725] <= layer1_out[11209];
     layer2_out[1726] <= layer1_out[6201];
     layer2_out[1727] <= layer1_out[3655] | layer1_out[3656];
     layer2_out[1728] <= ~layer1_out[9422] | layer1_out[9423];
     layer2_out[1729] <= ~layer1_out[2556] | layer1_out[2555];
     layer2_out[1730] <= ~layer1_out[11287];
     layer2_out[1731] <= layer1_out[11378];
     layer2_out[1732] <= layer1_out[10092] ^ layer1_out[10093];
     layer2_out[1733] <= ~layer1_out[4124];
     layer2_out[1734] <= layer1_out[10272] & layer1_out[10273];
     layer2_out[1735] <= layer1_out[11478] & ~layer1_out[11477];
     layer2_out[1736] <= layer1_out[1576] & ~layer1_out[1575];
     layer2_out[1737] <= ~layer1_out[6338];
     layer2_out[1738] <= ~layer1_out[11404];
     layer2_out[1739] <= layer1_out[11221] | layer1_out[11222];
     layer2_out[1740] <= ~(layer1_out[592] | layer1_out[593]);
     layer2_out[1741] <= layer1_out[10098];
     layer2_out[1742] <= layer1_out[5136] | layer1_out[5137];
     layer2_out[1743] <= ~layer1_out[5277];
     layer2_out[1744] <= ~layer1_out[11706] | layer1_out[11707];
     layer2_out[1745] <= ~layer1_out[11565];
     layer2_out[1746] <= layer1_out[4014];
     layer2_out[1747] <= ~(layer1_out[2661] & layer1_out[2662]);
     layer2_out[1748] <= layer1_out[11654] & ~layer1_out[11655];
     layer2_out[1749] <= ~(layer1_out[2606] ^ layer1_out[2607]);
     layer2_out[1750] <= layer1_out[1461] & layer1_out[1462];
     layer2_out[1751] <= layer1_out[422] & layer1_out[423];
     layer2_out[1752] <= layer1_out[11315];
     layer2_out[1753] <= layer1_out[3636] | layer1_out[3637];
     layer2_out[1754] <= layer1_out[5426];
     layer2_out[1755] <= ~(layer1_out[2984] & layer1_out[2985]);
     layer2_out[1756] <= ~(layer1_out[8384] ^ layer1_out[8385]);
     layer2_out[1757] <= layer1_out[10103] & ~layer1_out[10102];
     layer2_out[1758] <= layer1_out[9105];
     layer2_out[1759] <= layer1_out[6165] & ~layer1_out[6164];
     layer2_out[1760] <= layer1_out[9668] | layer1_out[9669];
     layer2_out[1761] <= ~layer1_out[10351];
     layer2_out[1762] <= ~layer1_out[4135] | layer1_out[4136];
     layer2_out[1763] <= ~layer1_out[2781];
     layer2_out[1764] <= ~layer1_out[8148] | layer1_out[8147];
     layer2_out[1765] <= layer1_out[10934] ^ layer1_out[10935];
     layer2_out[1766] <= layer1_out[2577] & ~layer1_out[2578];
     layer2_out[1767] <= layer1_out[5495] ^ layer1_out[5496];
     layer2_out[1768] <= layer1_out[2620];
     layer2_out[1769] <= layer1_out[2030] & ~layer1_out[2029];
     layer2_out[1770] <= layer1_out[9824] | layer1_out[9825];
     layer2_out[1771] <= layer1_out[9818];
     layer2_out[1772] <= layer1_out[4837] & ~layer1_out[4836];
     layer2_out[1773] <= ~(layer1_out[11619] | layer1_out[11620]);
     layer2_out[1774] <= layer1_out[2018] ^ layer1_out[2019];
     layer2_out[1775] <= ~layer1_out[10125] | layer1_out[10124];
     layer2_out[1776] <= ~layer1_out[6583];
     layer2_out[1777] <= layer1_out[11128] & layer1_out[11129];
     layer2_out[1778] <= ~layer1_out[8582];
     layer2_out[1779] <= ~(layer1_out[7840] & layer1_out[7841]);
     layer2_out[1780] <= ~(layer1_out[4534] | layer1_out[4535]);
     layer2_out[1781] <= ~(layer1_out[8059] | layer1_out[8060]);
     layer2_out[1782] <= layer1_out[4111];
     layer2_out[1783] <= ~layer1_out[9463];
     layer2_out[1784] <= layer1_out[4538] | layer1_out[4539];
     layer2_out[1785] <= layer1_out[2503];
     layer2_out[1786] <= ~layer1_out[3592];
     layer2_out[1787] <= layer1_out[8183] & ~layer1_out[8184];
     layer2_out[1788] <= ~layer1_out[2785] | layer1_out[2786];
     layer2_out[1789] <= ~layer1_out[3696] | layer1_out[3695];
     layer2_out[1790] <= ~(layer1_out[7748] ^ layer1_out[7749]);
     layer2_out[1791] <= layer1_out[1378];
     layer2_out[1792] <= layer1_out[11823] ^ layer1_out[11824];
     layer2_out[1793] <= ~(layer1_out[5814] ^ layer1_out[5815]);
     layer2_out[1794] <= layer1_out[3279] & ~layer1_out[3280];
     layer2_out[1795] <= layer1_out[3144];
     layer2_out[1796] <= ~(layer1_out[3843] & layer1_out[3844]);
     layer2_out[1797] <= layer1_out[4540];
     layer2_out[1798] <= layer1_out[747];
     layer2_out[1799] <= layer1_out[10868] & ~layer1_out[10867];
     layer2_out[1800] <= ~layer1_out[3825];
     layer2_out[1801] <= ~(layer1_out[3858] & layer1_out[3859]);
     layer2_out[1802] <= ~layer1_out[6385] | layer1_out[6386];
     layer2_out[1803] <= ~layer1_out[3474] | layer1_out[3475];
     layer2_out[1804] <= ~layer1_out[11359];
     layer2_out[1805] <= layer1_out[8585] ^ layer1_out[8586];
     layer2_out[1806] <= ~layer1_out[9241] | layer1_out[9240];
     layer2_out[1807] <= ~layer1_out[10872];
     layer2_out[1808] <= ~layer1_out[6748] | layer1_out[6749];
     layer2_out[1809] <= ~layer1_out[10762];
     layer2_out[1810] <= layer1_out[10363];
     layer2_out[1811] <= ~layer1_out[11232] | layer1_out[11233];
     layer2_out[1812] <= ~(layer1_out[10828] | layer1_out[10829]);
     layer2_out[1813] <= ~(layer1_out[11884] | layer1_out[11885]);
     layer2_out[1814] <= ~layer1_out[5325];
     layer2_out[1815] <= ~layer1_out[308] | layer1_out[309];
     layer2_out[1816] <= ~layer1_out[4480] | layer1_out[4481];
     layer2_out[1817] <= layer1_out[634];
     layer2_out[1818] <= ~layer1_out[5547];
     layer2_out[1819] <= layer1_out[7025] & ~layer1_out[7024];
     layer2_out[1820] <= ~layer1_out[1788];
     layer2_out[1821] <= ~layer1_out[6918] | layer1_out[6917];
     layer2_out[1822] <= layer1_out[4450] & ~layer1_out[4449];
     layer2_out[1823] <= ~(layer1_out[5573] | layer1_out[5574]);
     layer2_out[1824] <= ~(layer1_out[10439] ^ layer1_out[10440]);
     layer2_out[1825] <= ~layer1_out[9274];
     layer2_out[1826] <= layer1_out[9841];
     layer2_out[1827] <= ~layer1_out[3313] | layer1_out[3312];
     layer2_out[1828] <= ~layer1_out[3117] | layer1_out[3116];
     layer2_out[1829] <= layer1_out[776];
     layer2_out[1830] <= layer1_out[4514] & ~layer1_out[4515];
     layer2_out[1831] <= ~layer1_out[6037];
     layer2_out[1832] <= ~(layer1_out[10650] | layer1_out[10651]);
     layer2_out[1833] <= layer1_out[3305] & ~layer1_out[3306];
     layer2_out[1834] <= layer1_out[930] & ~layer1_out[929];
     layer2_out[1835] <= layer1_out[91] | layer1_out[92];
     layer2_out[1836] <= layer1_out[9012] | layer1_out[9013];
     layer2_out[1837] <= ~(layer1_out[11517] ^ layer1_out[11518]);
     layer2_out[1838] <= layer1_out[10495] ^ layer1_out[10496];
     layer2_out[1839] <= ~(layer1_out[2944] ^ layer1_out[2945]);
     layer2_out[1840] <= layer1_out[9495] & ~layer1_out[9494];
     layer2_out[1841] <= layer1_out[10149];
     layer2_out[1842] <= ~layer1_out[9876] | layer1_out[9877];
     layer2_out[1843] <= ~(layer1_out[1544] & layer1_out[1545]);
     layer2_out[1844] <= ~(layer1_out[2316] | layer1_out[2317]);
     layer2_out[1845] <= layer1_out[259] & layer1_out[260];
     layer2_out[1846] <= ~(layer1_out[11408] & layer1_out[11409]);
     layer2_out[1847] <= 1'b1;
     layer2_out[1848] <= layer1_out[5472];
     layer2_out[1849] <= ~layer1_out[431];
     layer2_out[1850] <= layer1_out[6588] ^ layer1_out[6589];
     layer2_out[1851] <= layer1_out[2207];
     layer2_out[1852] <= layer1_out[3223] & ~layer1_out[3224];
     layer2_out[1853] <= layer1_out[4870] & ~layer1_out[4869];
     layer2_out[1854] <= ~layer1_out[9904] | layer1_out[9903];
     layer2_out[1855] <= ~layer1_out[7591] | layer1_out[7590];
     layer2_out[1856] <= ~layer1_out[8257];
     layer2_out[1857] <= ~layer1_out[3568] | layer1_out[3569];
     layer2_out[1858] <= layer1_out[8518] & ~layer1_out[8517];
     layer2_out[1859] <= ~layer1_out[6898];
     layer2_out[1860] <= layer1_out[7537];
     layer2_out[1861] <= ~layer1_out[7568];
     layer2_out[1862] <= ~(layer1_out[7087] & layer1_out[7088]);
     layer2_out[1863] <= layer1_out[3624];
     layer2_out[1864] <= layer1_out[723];
     layer2_out[1865] <= 1'b0;
     layer2_out[1866] <= layer1_out[6909];
     layer2_out[1867] <= ~layer1_out[8836] | layer1_out[8837];
     layer2_out[1868] <= layer1_out[3406] | layer1_out[3407];
     layer2_out[1869] <= layer1_out[9524] & layer1_out[9525];
     layer2_out[1870] <= layer1_out[11432] & ~layer1_out[11433];
     layer2_out[1871] <= layer1_out[6341] & ~layer1_out[6340];
     layer2_out[1872] <= layer1_out[1146] & ~layer1_out[1147];
     layer2_out[1873] <= ~(layer1_out[1195] | layer1_out[1196]);
     layer2_out[1874] <= 1'b1;
     layer2_out[1875] <= layer1_out[237] & layer1_out[238];
     layer2_out[1876] <= layer1_out[3481];
     layer2_out[1877] <= layer1_out[8995];
     layer2_out[1878] <= ~(layer1_out[298] ^ layer1_out[299]);
     layer2_out[1879] <= ~layer1_out[9908] | layer1_out[9909];
     layer2_out[1880] <= ~layer1_out[6294] | layer1_out[6293];
     layer2_out[1881] <= ~(layer1_out[10953] & layer1_out[10954]);
     layer2_out[1882] <= ~layer1_out[5375];
     layer2_out[1883] <= ~layer1_out[408];
     layer2_out[1884] <= ~(layer1_out[9951] | layer1_out[9952]);
     layer2_out[1885] <= ~layer1_out[11868] | layer1_out[11869];
     layer2_out[1886] <= layer1_out[1821] | layer1_out[1822];
     layer2_out[1887] <= ~(layer1_out[5840] & layer1_out[5841]);
     layer2_out[1888] <= layer1_out[11428] & ~layer1_out[11427];
     layer2_out[1889] <= layer1_out[10643] & ~layer1_out[10642];
     layer2_out[1890] <= ~layer1_out[11768];
     layer2_out[1891] <= ~(layer1_out[9591] & layer1_out[9592]);
     layer2_out[1892] <= layer1_out[10705] & ~layer1_out[10706];
     layer2_out[1893] <= layer1_out[3988];
     layer2_out[1894] <= ~layer1_out[3197];
     layer2_out[1895] <= layer1_out[2767] ^ layer1_out[2768];
     layer2_out[1896] <= layer1_out[2127] ^ layer1_out[2128];
     layer2_out[1897] <= ~layer1_out[4803];
     layer2_out[1898] <= ~(layer1_out[10611] ^ layer1_out[10612]);
     layer2_out[1899] <= ~layer1_out[3918];
     layer2_out[1900] <= layer1_out[5757] & ~layer1_out[5756];
     layer2_out[1901] <= layer1_out[10730] & ~layer1_out[10729];
     layer2_out[1902] <= ~layer1_out[3811];
     layer2_out[1903] <= ~layer1_out[9415];
     layer2_out[1904] <= layer1_out[5960] & layer1_out[5961];
     layer2_out[1905] <= layer1_out[4270];
     layer2_out[1906] <= ~(layer1_out[9159] & layer1_out[9160]);
     layer2_out[1907] <= layer1_out[4460];
     layer2_out[1908] <= ~layer1_out[10184];
     layer2_out[1909] <= ~layer1_out[2002];
     layer2_out[1910] <= ~layer1_out[6258];
     layer2_out[1911] <= layer1_out[7113] & layer1_out[7114];
     layer2_out[1912] <= ~layer1_out[4027];
     layer2_out[1913] <= layer1_out[7133];
     layer2_out[1914] <= layer1_out[3791] & layer1_out[3792];
     layer2_out[1915] <= ~(layer1_out[6912] ^ layer1_out[6913]);
     layer2_out[1916] <= ~layer1_out[7782];
     layer2_out[1917] <= ~layer1_out[995];
     layer2_out[1918] <= ~layer1_out[7772];
     layer2_out[1919] <= layer1_out[4693] | layer1_out[4694];
     layer2_out[1920] <= layer1_out[8029] & ~layer1_out[8030];
     layer2_out[1921] <= layer1_out[10158] | layer1_out[10159];
     layer2_out[1922] <= layer1_out[2195];
     layer2_out[1923] <= layer1_out[7088] | layer1_out[7089];
     layer2_out[1924] <= layer1_out[1967] & ~layer1_out[1966];
     layer2_out[1925] <= ~(layer1_out[4004] & layer1_out[4005]);
     layer2_out[1926] <= layer1_out[5170] | layer1_out[5171];
     layer2_out[1927] <= ~(layer1_out[10535] ^ layer1_out[10536]);
     layer2_out[1928] <= layer1_out[5793] & ~layer1_out[5792];
     layer2_out[1929] <= layer1_out[4472] & ~layer1_out[4473];
     layer2_out[1930] <= layer1_out[2586];
     layer2_out[1931] <= ~(layer1_out[10216] & layer1_out[10217]);
     layer2_out[1932] <= layer1_out[11055] | layer1_out[11056];
     layer2_out[1933] <= layer1_out[11026];
     layer2_out[1934] <= layer1_out[6436] & ~layer1_out[6437];
     layer2_out[1935] <= ~(layer1_out[1519] | layer1_out[1520]);
     layer2_out[1936] <= ~layer1_out[2904];
     layer2_out[1937] <= layer1_out[9596];
     layer2_out[1938] <= layer1_out[1123] & layer1_out[1124];
     layer2_out[1939] <= ~layer1_out[340] | layer1_out[339];
     layer2_out[1940] <= ~layer1_out[7232];
     layer2_out[1941] <= ~layer1_out[6205];
     layer2_out[1942] <= layer1_out[8861];
     layer2_out[1943] <= layer1_out[11941] & ~layer1_out[11942];
     layer2_out[1944] <= ~layer1_out[4717] | layer1_out[4718];
     layer2_out[1945] <= layer1_out[6600] | layer1_out[6601];
     layer2_out[1946] <= ~layer1_out[2383];
     layer2_out[1947] <= ~layer1_out[8060];
     layer2_out[1948] <= ~(layer1_out[8560] & layer1_out[8561]);
     layer2_out[1949] <= ~layer1_out[6098];
     layer2_out[1950] <= ~layer1_out[10594];
     layer2_out[1951] <= layer1_out[2465];
     layer2_out[1952] <= layer1_out[7487];
     layer2_out[1953] <= ~(layer1_out[6061] & layer1_out[6062]);
     layer2_out[1954] <= ~(layer1_out[1516] & layer1_out[1517]);
     layer2_out[1955] <= layer1_out[5557];
     layer2_out[1956] <= ~layer1_out[11853];
     layer2_out[1957] <= ~(layer1_out[10017] | layer1_out[10018]);
     layer2_out[1958] <= layer1_out[11002];
     layer2_out[1959] <= ~(layer1_out[8762] & layer1_out[8763]);
     layer2_out[1960] <= ~(layer1_out[10558] ^ layer1_out[10559]);
     layer2_out[1961] <= ~layer1_out[9998];
     layer2_out[1962] <= layer1_out[6129] & layer1_out[6130];
     layer2_out[1963] <= ~layer1_out[7136];
     layer2_out[1964] <= layer1_out[11961] & ~layer1_out[11960];
     layer2_out[1965] <= 1'b1;
     layer2_out[1966] <= layer1_out[3855] & ~layer1_out[3856];
     layer2_out[1967] <= ~layer1_out[6318];
     layer2_out[1968] <= layer1_out[696];
     layer2_out[1969] <= ~layer1_out[4845] | layer1_out[4846];
     layer2_out[1970] <= 1'b1;
     layer2_out[1971] <= ~(layer1_out[856] | layer1_out[857]);
     layer2_out[1972] <= layer1_out[4484] ^ layer1_out[4485];
     layer2_out[1973] <= layer1_out[25];
     layer2_out[1974] <= layer1_out[2531] & layer1_out[2532];
     layer2_out[1975] <= ~(layer1_out[5719] ^ layer1_out[5720]);
     layer2_out[1976] <= ~layer1_out[4963];
     layer2_out[1977] <= layer1_out[1613];
     layer2_out[1978] <= ~layer1_out[2617] | layer1_out[2616];
     layer2_out[1979] <= ~(layer1_out[7359] | layer1_out[7360]);
     layer2_out[1980] <= ~layer1_out[4331];
     layer2_out[1981] <= ~layer1_out[11951];
     layer2_out[1982] <= layer1_out[4878] ^ layer1_out[4879];
     layer2_out[1983] <= ~layer1_out[7977];
     layer2_out[1984] <= layer1_out[169] ^ layer1_out[170];
     layer2_out[1985] <= ~layer1_out[10534];
     layer2_out[1986] <= layer1_out[4398] ^ layer1_out[4399];
     layer2_out[1987] <= layer1_out[2870];
     layer2_out[1988] <= layer1_out[10276];
     layer2_out[1989] <= ~layer1_out[107];
     layer2_out[1990] <= ~(layer1_out[1426] ^ layer1_out[1427]);
     layer2_out[1991] <= ~layer1_out[6995];
     layer2_out[1992] <= ~layer1_out[8763] | layer1_out[8764];
     layer2_out[1993] <= ~layer1_out[9976];
     layer2_out[1994] <= layer1_out[2161] | layer1_out[2162];
     layer2_out[1995] <= ~layer1_out[8538] | layer1_out[8537];
     layer2_out[1996] <= layer1_out[4559] & ~layer1_out[4558];
     layer2_out[1997] <= ~(layer1_out[7807] ^ layer1_out[7808]);
     layer2_out[1998] <= layer1_out[4202] & layer1_out[4203];
     layer2_out[1999] <= ~layer1_out[1757] | layer1_out[1756];
     layer2_out[2000] <= ~layer1_out[2800];
     layer2_out[2001] <= ~(layer1_out[5032] & layer1_out[5033]);
     layer2_out[2002] <= ~(layer1_out[672] & layer1_out[673]);
     layer2_out[2003] <= 1'b0;
     layer2_out[2004] <= ~layer1_out[11399];
     layer2_out[2005] <= 1'b0;
     layer2_out[2006] <= layer1_out[9081] & ~layer1_out[9080];
     layer2_out[2007] <= ~layer1_out[3093];
     layer2_out[2008] <= ~layer1_out[788];
     layer2_out[2009] <= layer1_out[1393];
     layer2_out[2010] <= ~layer1_out[561] | layer1_out[560];
     layer2_out[2011] <= ~layer1_out[11259];
     layer2_out[2012] <= layer1_out[1976];
     layer2_out[2013] <= layer1_out[8715] ^ layer1_out[8716];
     layer2_out[2014] <= ~layer1_out[7481] | layer1_out[7480];
     layer2_out[2015] <= ~layer1_out[241];
     layer2_out[2016] <= ~layer1_out[8526];
     layer2_out[2017] <= layer1_out[5841] & layer1_out[5842];
     layer2_out[2018] <= layer1_out[8397];
     layer2_out[2019] <= ~(layer1_out[10834] ^ layer1_out[10835]);
     layer2_out[2020] <= layer1_out[10788];
     layer2_out[2021] <= layer1_out[9886];
     layer2_out[2022] <= ~layer1_out[6474];
     layer2_out[2023] <= ~layer1_out[10523] | layer1_out[10524];
     layer2_out[2024] <= layer1_out[7256] & ~layer1_out[7255];
     layer2_out[2025] <= layer1_out[4024];
     layer2_out[2026] <= ~layer1_out[5049];
     layer2_out[2027] <= layer1_out[6853];
     layer2_out[2028] <= layer1_out[815] & ~layer1_out[816];
     layer2_out[2029] <= layer1_out[2708];
     layer2_out[2030] <= layer1_out[6982];
     layer2_out[2031] <= layer1_out[2728] & ~layer1_out[2729];
     layer2_out[2032] <= layer1_out[8476] & ~layer1_out[8477];
     layer2_out[2033] <= ~layer1_out[11046] | layer1_out[11047];
     layer2_out[2034] <= layer1_out[10807];
     layer2_out[2035] <= ~layer1_out[7993] | layer1_out[7992];
     layer2_out[2036] <= layer1_out[8902] ^ layer1_out[8903];
     layer2_out[2037] <= layer1_out[3672];
     layer2_out[2038] <= ~layer1_out[2875];
     layer2_out[2039] <= ~layer1_out[6514];
     layer2_out[2040] <= ~(layer1_out[3901] | layer1_out[3902]);
     layer2_out[2041] <= ~layer1_out[10564] | layer1_out[10565];
     layer2_out[2042] <= ~layer1_out[9474];
     layer2_out[2043] <= layer1_out[3477] & ~layer1_out[3478];
     layer2_out[2044] <= layer1_out[604];
     layer2_out[2045] <= layer1_out[418];
     layer2_out[2046] <= layer1_out[7081] & ~layer1_out[7080];
     layer2_out[2047] <= layer1_out[2247];
     layer2_out[2048] <= layer1_out[3929];
     layer2_out[2049] <= ~(layer1_out[2993] & layer1_out[2994]);
     layer2_out[2050] <= layer1_out[9619] | layer1_out[9620];
     layer2_out[2051] <= layer1_out[7764] & ~layer1_out[7765];
     layer2_out[2052] <= 1'b0;
     layer2_out[2053] <= layer1_out[3127] | layer1_out[3128];
     layer2_out[2054] <= ~layer1_out[10370] | layer1_out[10371];
     layer2_out[2055] <= ~layer1_out[4742];
     layer2_out[2056] <= ~layer1_out[4730];
     layer2_out[2057] <= layer1_out[3463] & ~layer1_out[3464];
     layer2_out[2058] <= layer1_out[7800];
     layer2_out[2059] <= layer1_out[11549] & ~layer1_out[11550];
     layer2_out[2060] <= ~(layer1_out[9684] ^ layer1_out[9685]);
     layer2_out[2061] <= ~layer1_out[6366] | layer1_out[6367];
     layer2_out[2062] <= ~(layer1_out[2409] | layer1_out[2410]);
     layer2_out[2063] <= ~layer1_out[2151] | layer1_out[2152];
     layer2_out[2064] <= ~(layer1_out[10503] ^ layer1_out[10504]);
     layer2_out[2065] <= ~(layer1_out[509] & layer1_out[510]);
     layer2_out[2066] <= layer1_out[8972];
     layer2_out[2067] <= layer1_out[710] & ~layer1_out[709];
     layer2_out[2068] <= 1'b1;
     layer2_out[2069] <= ~layer1_out[10955] | layer1_out[10954];
     layer2_out[2070] <= ~layer1_out[7628];
     layer2_out[2071] <= layer1_out[926] | layer1_out[927];
     layer2_out[2072] <= layer1_out[363] | layer1_out[364];
     layer2_out[2073] <= ~(layer1_out[7617] & layer1_out[7618]);
     layer2_out[2074] <= ~(layer1_out[9854] ^ layer1_out[9855]);
     layer2_out[2075] <= 1'b0;
     layer2_out[2076] <= layer1_out[2110] | layer1_out[2111];
     layer2_out[2077] <= ~layer1_out[7738];
     layer2_out[2078] <= layer1_out[6842];
     layer2_out[2079] <= layer1_out[11012];
     layer2_out[2080] <= ~(layer1_out[4395] & layer1_out[4396]);
     layer2_out[2081] <= 1'b1;
     layer2_out[2082] <= ~layer1_out[220];
     layer2_out[2083] <= ~layer1_out[1619];
     layer2_out[2084] <= layer1_out[5588] & layer1_out[5589];
     layer2_out[2085] <= ~layer1_out[8804];
     layer2_out[2086] <= layer1_out[2574] & layer1_out[2575];
     layer2_out[2087] <= layer1_out[3267] & ~layer1_out[3266];
     layer2_out[2088] <= ~(layer1_out[5611] ^ layer1_out[5612]);
     layer2_out[2089] <= layer1_out[617];
     layer2_out[2090] <= ~layer1_out[6077] | layer1_out[6076];
     layer2_out[2091] <= layer1_out[9727];
     layer2_out[2092] <= ~(layer1_out[2298] | layer1_out[2299]);
     layer2_out[2093] <= ~layer1_out[8787] | layer1_out[8786];
     layer2_out[2094] <= 1'b0;
     layer2_out[2095] <= layer1_out[1257];
     layer2_out[2096] <= layer1_out[76] & ~layer1_out[77];
     layer2_out[2097] <= ~layer1_out[10738] | layer1_out[10739];
     layer2_out[2098] <= layer1_out[5636] & ~layer1_out[5635];
     layer2_out[2099] <= layer1_out[9158];
     layer2_out[2100] <= ~layer1_out[84];
     layer2_out[2101] <= layer1_out[7902] | layer1_out[7903];
     layer2_out[2102] <= ~(layer1_out[6916] | layer1_out[6917]);
     layer2_out[2103] <= layer1_out[618];
     layer2_out[2104] <= layer1_out[7475] & ~layer1_out[7476];
     layer2_out[2105] <= ~(layer1_out[6920] | layer1_out[6921]);
     layer2_out[2106] <= ~layer1_out[8761] | layer1_out[8760];
     layer2_out[2107] <= ~layer1_out[6406];
     layer2_out[2108] <= ~(layer1_out[11774] | layer1_out[11775]);
     layer2_out[2109] <= ~(layer1_out[9328] & layer1_out[9329]);
     layer2_out[2110] <= layer1_out[636] & ~layer1_out[637];
     layer2_out[2111] <= layer1_out[1872];
     layer2_out[2112] <= layer1_out[9432] | layer1_out[9433];
     layer2_out[2113] <= layer1_out[11763] ^ layer1_out[11764];
     layer2_out[2114] <= ~layer1_out[10606];
     layer2_out[2115] <= layer1_out[1891];
     layer2_out[2116] <= layer1_out[2564] | layer1_out[2565];
     layer2_out[2117] <= layer1_out[7717];
     layer2_out[2118] <= layer1_out[9004] | layer1_out[9005];
     layer2_out[2119] <= layer1_out[1350] | layer1_out[1351];
     layer2_out[2120] <= ~layer1_out[2855] | layer1_out[2856];
     layer2_out[2121] <= layer1_out[379] ^ layer1_out[380];
     layer2_out[2122] <= ~(layer1_out[1230] & layer1_out[1231]);
     layer2_out[2123] <= layer1_out[1518];
     layer2_out[2124] <= layer1_out[8573] & ~layer1_out[8572];
     layer2_out[2125] <= layer1_out[11294] & layer1_out[11295];
     layer2_out[2126] <= layer1_out[4638] ^ layer1_out[4639];
     layer2_out[2127] <= layer1_out[909];
     layer2_out[2128] <= layer1_out[11781];
     layer2_out[2129] <= layer1_out[9078];
     layer2_out[2130] <= ~(layer1_out[3782] ^ layer1_out[3783]);
     layer2_out[2131] <= layer1_out[3902];
     layer2_out[2132] <= layer1_out[9209] & ~layer1_out[9208];
     layer2_out[2133] <= layer1_out[704] ^ layer1_out[705];
     layer2_out[2134] <= layer1_out[83] & ~layer1_out[84];
     layer2_out[2135] <= layer1_out[6058] & ~layer1_out[6057];
     layer2_out[2136] <= layer1_out[10170] & ~layer1_out[10171];
     layer2_out[2137] <= layer1_out[7949];
     layer2_out[2138] <= ~(layer1_out[7094] | layer1_out[7095]);
     layer2_out[2139] <= layer1_out[7334] & layer1_out[7335];
     layer2_out[2140] <= layer1_out[11948] & ~layer1_out[11949];
     layer2_out[2141] <= layer1_out[1825];
     layer2_out[2142] <= ~layer1_out[6565] | layer1_out[6566];
     layer2_out[2143] <= layer1_out[6132] ^ layer1_out[6133];
     layer2_out[2144] <= layer1_out[1033] ^ layer1_out[1034];
     layer2_out[2145] <= ~(layer1_out[5947] | layer1_out[5948]);
     layer2_out[2146] <= layer1_out[7577] & ~layer1_out[7576];
     layer2_out[2147] <= layer1_out[1717] & ~layer1_out[1716];
     layer2_out[2148] <= layer1_out[10577] & ~layer1_out[10578];
     layer2_out[2149] <= layer1_out[8358];
     layer2_out[2150] <= ~layer1_out[11246];
     layer2_out[2151] <= layer1_out[10891];
     layer2_out[2152] <= layer1_out[8719] ^ layer1_out[8720];
     layer2_out[2153] <= ~(layer1_out[1477] | layer1_out[1478]);
     layer2_out[2154] <= layer1_out[1793];
     layer2_out[2155] <= ~(layer1_out[8366] ^ layer1_out[8367]);
     layer2_out[2156] <= ~layer1_out[4724];
     layer2_out[2157] <= layer1_out[2395];
     layer2_out[2158] <= ~(layer1_out[5977] ^ layer1_out[5978]);
     layer2_out[2159] <= layer1_out[7100] & layer1_out[7101];
     layer2_out[2160] <= layer1_out[11217];
     layer2_out[2161] <= ~layer1_out[7140] | layer1_out[7139];
     layer2_out[2162] <= ~layer1_out[4696];
     layer2_out[2163] <= ~layer1_out[11250];
     layer2_out[2164] <= ~layer1_out[11380];
     layer2_out[2165] <= layer1_out[2811];
     layer2_out[2166] <= layer1_out[10711] & ~layer1_out[10712];
     layer2_out[2167] <= ~layer1_out[4630];
     layer2_out[2168] <= layer1_out[7150] | layer1_out[7151];
     layer2_out[2169] <= ~layer1_out[6896] | layer1_out[6895];
     layer2_out[2170] <= layer1_out[11847] & ~layer1_out[11846];
     layer2_out[2171] <= layer1_out[10320] & ~layer1_out[10319];
     layer2_out[2172] <= ~layer1_out[8743];
     layer2_out[2173] <= ~layer1_out[2003];
     layer2_out[2174] <= layer1_out[1048];
     layer2_out[2175] <= ~(layer1_out[39] | layer1_out[40]);
     layer2_out[2176] <= ~(layer1_out[11891] | layer1_out[11892]);
     layer2_out[2177] <= layer1_out[5318];
     layer2_out[2178] <= ~layer1_out[2430] | layer1_out[2431];
     layer2_out[2179] <= layer1_out[11789] & ~layer1_out[11790];
     layer2_out[2180] <= layer1_out[1633] ^ layer1_out[1634];
     layer2_out[2181] <= ~layer1_out[9978];
     layer2_out[2182] <= layer1_out[1720];
     layer2_out[2183] <= ~layer1_out[4516];
     layer2_out[2184] <= layer1_out[2637] ^ layer1_out[2638];
     layer2_out[2185] <= layer1_out[3366];
     layer2_out[2186] <= ~(layer1_out[9938] | layer1_out[9939]);
     layer2_out[2187] <= layer1_out[934] | layer1_out[935];
     layer2_out[2188] <= ~layer1_out[5230] | layer1_out[5229];
     layer2_out[2189] <= ~layer1_out[6703] | layer1_out[6704];
     layer2_out[2190] <= layer1_out[5920];
     layer2_out[2191] <= ~(layer1_out[7473] | layer1_out[7474]);
     layer2_out[2192] <= ~(layer1_out[9092] | layer1_out[9093]);
     layer2_out[2193] <= ~layer1_out[2818];
     layer2_out[2194] <= layer1_out[5122] & ~layer1_out[5123];
     layer2_out[2195] <= layer1_out[11882];
     layer2_out[2196] <= ~layer1_out[6119];
     layer2_out[2197] <= layer1_out[6148];
     layer2_out[2198] <= ~layer1_out[5356] | layer1_out[5355];
     layer2_out[2199] <= ~layer1_out[7879];
     layer2_out[2200] <= layer1_out[11665] & ~layer1_out[11664];
     layer2_out[2201] <= ~layer1_out[5555];
     layer2_out[2202] <= 1'b0;
     layer2_out[2203] <= layer1_out[4192] & layer1_out[4193];
     layer2_out[2204] <= ~(layer1_out[11390] | layer1_out[11391]);
     layer2_out[2205] <= layer1_out[11388];
     layer2_out[2206] <= ~layer1_out[7456];
     layer2_out[2207] <= layer1_out[1621] & ~layer1_out[1622];
     layer2_out[2208] <= ~(layer1_out[6662] | layer1_out[6663]);
     layer2_out[2209] <= ~layer1_out[10603];
     layer2_out[2210] <= layer1_out[5562];
     layer2_out[2211] <= layer1_out[1194];
     layer2_out[2212] <= ~(layer1_out[9071] & layer1_out[9072]);
     layer2_out[2213] <= ~(layer1_out[8755] & layer1_out[8756]);
     layer2_out[2214] <= ~layer1_out[9376];
     layer2_out[2215] <= ~layer1_out[3039];
     layer2_out[2216] <= layer1_out[2649];
     layer2_out[2217] <= layer1_out[11687] & layer1_out[11688];
     layer2_out[2218] <= layer1_out[5722];
     layer2_out[2219] <= layer1_out[8134] & ~layer1_out[8135];
     layer2_out[2220] <= layer1_out[7855];
     layer2_out[2221] <= layer1_out[10128] & layer1_out[10129];
     layer2_out[2222] <= layer1_out[8709] & ~layer1_out[8708];
     layer2_out[2223] <= ~(layer1_out[6858] ^ layer1_out[6859]);
     layer2_out[2224] <= layer1_out[23] & layer1_out[24];
     layer2_out[2225] <= layer1_out[10194] & ~layer1_out[10195];
     layer2_out[2226] <= layer1_out[8315];
     layer2_out[2227] <= ~layer1_out[10070];
     layer2_out[2228] <= ~layer1_out[2039];
     layer2_out[2229] <= layer1_out[3567];
     layer2_out[2230] <= layer1_out[4616] | layer1_out[4617];
     layer2_out[2231] <= layer1_out[3965] | layer1_out[3966];
     layer2_out[2232] <= ~(layer1_out[10667] ^ layer1_out[10668]);
     layer2_out[2233] <= layer1_out[7591];
     layer2_out[2234] <= ~layer1_out[11333] | layer1_out[11334];
     layer2_out[2235] <= ~(layer1_out[7966] ^ layer1_out[7967]);
     layer2_out[2236] <= layer1_out[2287];
     layer2_out[2237] <= ~layer1_out[9663] | layer1_out[9664];
     layer2_out[2238] <= layer1_out[3356] & ~layer1_out[3355];
     layer2_out[2239] <= ~layer1_out[7544];
     layer2_out[2240] <= layer1_out[8874] & layer1_out[8875];
     layer2_out[2241] <= layer1_out[4275];
     layer2_out[2242] <= ~layer1_out[4563];
     layer2_out[2243] <= layer1_out[9353];
     layer2_out[2244] <= ~layer1_out[1431];
     layer2_out[2245] <= layer1_out[1646] & ~layer1_out[1647];
     layer2_out[2246] <= ~layer1_out[6381] | layer1_out[6380];
     layer2_out[2247] <= ~(layer1_out[3083] | layer1_out[3084]);
     layer2_out[2248] <= layer1_out[5243] | layer1_out[5244];
     layer2_out[2249] <= ~layer1_out[5950];
     layer2_out[2250] <= layer1_out[6445];
     layer2_out[2251] <= layer1_out[8626];
     layer2_out[2252] <= layer1_out[2754] | layer1_out[2755];
     layer2_out[2253] <= layer1_out[5761] & layer1_out[5762];
     layer2_out[2254] <= ~(layer1_out[841] | layer1_out[842]);
     layer2_out[2255] <= layer1_out[1415] & layer1_out[1416];
     layer2_out[2256] <= ~layer1_out[708] | layer1_out[709];
     layer2_out[2257] <= layer1_out[11539] & ~layer1_out[11540];
     layer2_out[2258] <= ~layer1_out[1791] | layer1_out[1792];
     layer2_out[2259] <= layer1_out[5175];
     layer2_out[2260] <= ~layer1_out[9841] | layer1_out[9842];
     layer2_out[2261] <= ~layer1_out[4708];
     layer2_out[2262] <= layer1_out[9584] ^ layer1_out[9585];
     layer2_out[2263] <= layer1_out[272];
     layer2_out[2264] <= layer1_out[2163] & layer1_out[2164];
     layer2_out[2265] <= ~layer1_out[4521] | layer1_out[4520];
     layer2_out[2266] <= layer1_out[1893] ^ layer1_out[1894];
     layer2_out[2267] <= layer1_out[1367];
     layer2_out[2268] <= layer1_out[9353];
     layer2_out[2269] <= 1'b0;
     layer2_out[2270] <= ~layer1_out[9671] | layer1_out[9670];
     layer2_out[2271] <= layer1_out[4967] & ~layer1_out[4966];
     layer2_out[2272] <= ~layer1_out[9674];
     layer2_out[2273] <= ~layer1_out[2517];
     layer2_out[2274] <= ~layer1_out[6987];
     layer2_out[2275] <= layer1_out[857];
     layer2_out[2276] <= layer1_out[1660];
     layer2_out[2277] <= ~layer1_out[11697];
     layer2_out[2278] <= ~layer1_out[7643];
     layer2_out[2279] <= ~layer1_out[10629];
     layer2_out[2280] <= ~layer1_out[7997];
     layer2_out[2281] <= layer1_out[3891];
     layer2_out[2282] <= layer1_out[11006];
     layer2_out[2283] <= ~(layer1_out[10373] & layer1_out[10374]);
     layer2_out[2284] <= ~(layer1_out[9288] & layer1_out[9289]);
     layer2_out[2285] <= layer1_out[2404] & ~layer1_out[2405];
     layer2_out[2286] <= layer1_out[5181] & ~layer1_out[5180];
     layer2_out[2287] <= ~(layer1_out[6144] & layer1_out[6145]);
     layer2_out[2288] <= ~layer1_out[5218];
     layer2_out[2289] <= ~layer1_out[3838];
     layer2_out[2290] <= layer1_out[2482] & ~layer1_out[2481];
     layer2_out[2291] <= ~(layer1_out[2129] & layer1_out[2130]);
     layer2_out[2292] <= layer1_out[3710] & ~layer1_out[3711];
     layer2_out[2293] <= ~layer1_out[2097] | layer1_out[2096];
     layer2_out[2294] <= ~layer1_out[7341];
     layer2_out[2295] <= ~(layer1_out[11865] & layer1_out[11866]);
     layer2_out[2296] <= ~(layer1_out[4417] ^ layer1_out[4418]);
     layer2_out[2297] <= layer1_out[9416] & layer1_out[9417];
     layer2_out[2298] <= layer1_out[9884];
     layer2_out[2299] <= layer1_out[918];
     layer2_out[2300] <= layer1_out[10156];
     layer2_out[2301] <= layer1_out[7712] ^ layer1_out[7713];
     layer2_out[2302] <= layer1_out[6939] & layer1_out[6940];
     layer2_out[2303] <= layer1_out[631];
     layer2_out[2304] <= layer1_out[7233];
     layer2_out[2305] <= ~layer1_out[9170];
     layer2_out[2306] <= ~(layer1_out[6232] & layer1_out[6233]);
     layer2_out[2307] <= ~(layer1_out[9325] ^ layer1_out[9326]);
     layer2_out[2308] <= layer1_out[6254] | layer1_out[6255];
     layer2_out[2309] <= layer1_out[6347] & layer1_out[6348];
     layer2_out[2310] <= ~layer1_out[6938];
     layer2_out[2311] <= layer1_out[4496];
     layer2_out[2312] <= layer1_out[11186];
     layer2_out[2313] <= layer1_out[5159] ^ layer1_out[5160];
     layer2_out[2314] <= 1'b0;
     layer2_out[2315] <= layer1_out[1032] & layer1_out[1033];
     layer2_out[2316] <= ~(layer1_out[2370] & layer1_out[2371]);
     layer2_out[2317] <= ~layer1_out[9680];
     layer2_out[2318] <= layer1_out[11263] | layer1_out[11264];
     layer2_out[2319] <= layer1_out[2499];
     layer2_out[2320] <= ~layer1_out[7302];
     layer2_out[2321] <= ~layer1_out[2182];
     layer2_out[2322] <= layer1_out[82] & ~layer1_out[83];
     layer2_out[2323] <= layer1_out[11592] & ~layer1_out[11593];
     layer2_out[2324] <= ~(layer1_out[3789] ^ layer1_out[3790]);
     layer2_out[2325] <= 1'b0;
     layer2_out[2326] <= layer1_out[9297] ^ layer1_out[9298];
     layer2_out[2327] <= layer1_out[8767] & ~layer1_out[8766];
     layer2_out[2328] <= ~(layer1_out[11059] | layer1_out[11060]);
     layer2_out[2329] <= layer1_out[3385] | layer1_out[3386];
     layer2_out[2330] <= layer1_out[7553] & ~layer1_out[7552];
     layer2_out[2331] <= layer1_out[6107] | layer1_out[6108];
     layer2_out[2332] <= layer1_out[5895];
     layer2_out[2333] <= layer1_out[10780] & layer1_out[10781];
     layer2_out[2334] <= layer1_out[610];
     layer2_out[2335] <= ~(layer1_out[11214] ^ layer1_out[11215]);
     layer2_out[2336] <= ~layer1_out[10823] | layer1_out[10824];
     layer2_out[2337] <= layer1_out[9774];
     layer2_out[2338] <= layer1_out[788];
     layer2_out[2339] <= layer1_out[9312] & ~layer1_out[9311];
     layer2_out[2340] <= layer1_out[303];
     layer2_out[2341] <= layer1_out[8880];
     layer2_out[2342] <= ~layer1_out[8483];
     layer2_out[2343] <= layer1_out[7295] & ~layer1_out[7294];
     layer2_out[2344] <= ~layer1_out[5773];
     layer2_out[2345] <= layer1_out[1059];
     layer2_out[2346] <= ~layer1_out[8661];
     layer2_out[2347] <= 1'b0;
     layer2_out[2348] <= layer1_out[8345] & layer1_out[8346];
     layer2_out[2349] <= ~layer1_out[6182] | layer1_out[6183];
     layer2_out[2350] <= ~layer1_out[338] | layer1_out[337];
     layer2_out[2351] <= layer1_out[4303] & ~layer1_out[4304];
     layer2_out[2352] <= ~(layer1_out[11714] | layer1_out[11715]);
     layer2_out[2353] <= ~layer1_out[11645];
     layer2_out[2354] <= layer1_out[3376] & ~layer1_out[3375];
     layer2_out[2355] <= ~(layer1_out[8454] & layer1_out[8455]);
     layer2_out[2356] <= 1'b0;
     layer2_out[2357] <= layer1_out[7257];
     layer2_out[2358] <= layer1_out[736] | layer1_out[737];
     layer2_out[2359] <= ~layer1_out[3726] | layer1_out[3727];
     layer2_out[2360] <= layer1_out[5955];
     layer2_out[2361] <= layer1_out[7324];
     layer2_out[2362] <= ~layer1_out[9669] | layer1_out[9670];
     layer2_out[2363] <= layer1_out[11343] & ~layer1_out[11344];
     layer2_out[2364] <= layer1_out[4146];
     layer2_out[2365] <= ~layer1_out[4190] | layer1_out[4189];
     layer2_out[2366] <= 1'b1;
     layer2_out[2367] <= ~(layer1_out[10016] & layer1_out[10017]);
     layer2_out[2368] <= ~(layer1_out[3973] ^ layer1_out[3974]);
     layer2_out[2369] <= ~(layer1_out[5368] & layer1_out[5369]);
     layer2_out[2370] <= ~layer1_out[6512];
     layer2_out[2371] <= ~(layer1_out[11110] | layer1_out[11111]);
     layer2_out[2372] <= ~layer1_out[8251] | layer1_out[8250];
     layer2_out[2373] <= layer1_out[10480] & ~layer1_out[10481];
     layer2_out[2374] <= layer1_out[7687];
     layer2_out[2375] <= ~(layer1_out[835] & layer1_out[836]);
     layer2_out[2376] <= layer1_out[8815] & ~layer1_out[8816];
     layer2_out[2377] <= ~(layer1_out[4790] ^ layer1_out[4791]);
     layer2_out[2378] <= layer1_out[7202] | layer1_out[7203];
     layer2_out[2379] <= ~layer1_out[2766];
     layer2_out[2380] <= ~layer1_out[2193];
     layer2_out[2381] <= ~(layer1_out[2844] & layer1_out[2845]);
     layer2_out[2382] <= ~layer1_out[4668];
     layer2_out[2383] <= ~(layer1_out[7633] | layer1_out[7634]);
     layer2_out[2384] <= layer1_out[2134] & ~layer1_out[2135];
     layer2_out[2385] <= layer1_out[7653] | layer1_out[7654];
     layer2_out[2386] <= ~layer1_out[10407] | layer1_out[10406];
     layer2_out[2387] <= layer1_out[1263] & ~layer1_out[1264];
     layer2_out[2388] <= ~layer1_out[10639];
     layer2_out[2389] <= ~layer1_out[2025];
     layer2_out[2390] <= ~layer1_out[9259];
     layer2_out[2391] <= ~(layer1_out[176] ^ layer1_out[177]);
     layer2_out[2392] <= ~layer1_out[3737] | layer1_out[3738];
     layer2_out[2393] <= ~layer1_out[5446] | layer1_out[5447];
     layer2_out[2394] <= layer1_out[7289] ^ layer1_out[7290];
     layer2_out[2395] <= ~layer1_out[8180];
     layer2_out[2396] <= layer1_out[5743];
     layer2_out[2397] <= ~layer1_out[5478];
     layer2_out[2398] <= ~layer1_out[3670];
     layer2_out[2399] <= layer1_out[3864] ^ layer1_out[3865];
     layer2_out[2400] <= layer1_out[3084] ^ layer1_out[3085];
     layer2_out[2401] <= ~layer1_out[1775] | layer1_out[1774];
     layer2_out[2402] <= layer1_out[9337] & ~layer1_out[9338];
     layer2_out[2403] <= 1'b1;
     layer2_out[2404] <= ~(layer1_out[2733] & layer1_out[2734]);
     layer2_out[2405] <= layer1_out[7909] & layer1_out[7910];
     layer2_out[2406] <= ~layer1_out[1101];
     layer2_out[2407] <= layer1_out[2228] & layer1_out[2229];
     layer2_out[2408] <= ~layer1_out[10370] | layer1_out[10369];
     layer2_out[2409] <= layer1_out[164];
     layer2_out[2410] <= layer1_out[1823] & layer1_out[1824];
     layer2_out[2411] <= ~(layer1_out[5176] ^ layer1_out[5177]);
     layer2_out[2412] <= ~(layer1_out[8010] | layer1_out[8011]);
     layer2_out[2413] <= ~(layer1_out[8456] | layer1_out[8457]);
     layer2_out[2414] <= ~layer1_out[7393];
     layer2_out[2415] <= ~layer1_out[5967];
     layer2_out[2416] <= layer1_out[4663] & layer1_out[4664];
     layer2_out[2417] <= ~(layer1_out[9067] ^ layer1_out[9068]);
     layer2_out[2418] <= ~layer1_out[6042] | layer1_out[6043];
     layer2_out[2419] <= layer1_out[4545] & ~layer1_out[4546];
     layer2_out[2420] <= ~layer1_out[6104];
     layer2_out[2421] <= layer1_out[7129] & layer1_out[7130];
     layer2_out[2422] <= layer1_out[5524] ^ layer1_out[5525];
     layer2_out[2423] <= layer1_out[10727] & layer1_out[10728];
     layer2_out[2424] <= ~layer1_out[5739];
     layer2_out[2425] <= 1'b1;
     layer2_out[2426] <= layer1_out[7342] & layer1_out[7343];
     layer2_out[2427] <= ~(layer1_out[3492] ^ layer1_out[3493]);
     layer2_out[2428] <= layer1_out[11180] & ~layer1_out[11181];
     layer2_out[2429] <= ~(layer1_out[3105] & layer1_out[3106]);
     layer2_out[2430] <= ~(layer1_out[3919] & layer1_out[3920]);
     layer2_out[2431] <= 1'b0;
     layer2_out[2432] <= layer1_out[7102] & ~layer1_out[7101];
     layer2_out[2433] <= layer1_out[9701] & layer1_out[9702];
     layer2_out[2434] <= ~(layer1_out[3836] ^ layer1_out[3837]);
     layer2_out[2435] <= layer1_out[10134];
     layer2_out[2436] <= ~layer1_out[799] | layer1_out[798];
     layer2_out[2437] <= ~layer1_out[1265];
     layer2_out[2438] <= ~layer1_out[2647] | layer1_out[2646];
     layer2_out[2439] <= layer1_out[5086] & layer1_out[5087];
     layer2_out[2440] <= layer1_out[6150];
     layer2_out[2441] <= ~layer1_out[3197];
     layer2_out[2442] <= layer1_out[164];
     layer2_out[2443] <= ~layer1_out[3681] | layer1_out[3682];
     layer2_out[2444] <= ~(layer1_out[1686] ^ layer1_out[1687]);
     layer2_out[2445] <= ~(layer1_out[4980] & layer1_out[4981]);
     layer2_out[2446] <= layer1_out[8193] | layer1_out[8194];
     layer2_out[2447] <= layer1_out[11337] | layer1_out[11338];
     layer2_out[2448] <= ~layer1_out[8034];
     layer2_out[2449] <= layer1_out[1546] | layer1_out[1547];
     layer2_out[2450] <= ~layer1_out[250] | layer1_out[249];
     layer2_out[2451] <= ~layer1_out[5270];
     layer2_out[2452] <= ~layer1_out[283];
     layer2_out[2453] <= ~(layer1_out[3913] | layer1_out[3914]);
     layer2_out[2454] <= layer1_out[5931] | layer1_out[5932];
     layer2_out[2455] <= ~layer1_out[11424] | layer1_out[11423];
     layer2_out[2456] <= 1'b1;
     layer2_out[2457] <= ~(layer1_out[9807] | layer1_out[9808]);
     layer2_out[2458] <= layer1_out[3965];
     layer2_out[2459] <= ~layer1_out[1835] | layer1_out[1834];
     layer2_out[2460] <= ~(layer1_out[3602] & layer1_out[3603]);
     layer2_out[2461] <= ~layer1_out[10117];
     layer2_out[2462] <= layer1_out[8304];
     layer2_out[2463] <= layer1_out[1231] ^ layer1_out[1232];
     layer2_out[2464] <= ~layer1_out[825];
     layer2_out[2465] <= ~layer1_out[2232];
     layer2_out[2466] <= ~(layer1_out[355] ^ layer1_out[356]);
     layer2_out[2467] <= ~(layer1_out[7695] | layer1_out[7696]);
     layer2_out[2468] <= ~layer1_out[1428] | layer1_out[1429];
     layer2_out[2469] <= layer1_out[7877];
     layer2_out[2470] <= ~(layer1_out[880] | layer1_out[881]);
     layer2_out[2471] <= layer1_out[8784] & layer1_out[8785];
     layer2_out[2472] <= layer1_out[1881] & ~layer1_out[1880];
     layer2_out[2473] <= ~(layer1_out[3152] & layer1_out[3153]);
     layer2_out[2474] <= layer1_out[4186] & ~layer1_out[4185];
     layer2_out[2475] <= layer1_out[2793] & ~layer1_out[2794];
     layer2_out[2476] <= layer1_out[7810] | layer1_out[7811];
     layer2_out[2477] <= layer1_out[1988] | layer1_out[1989];
     layer2_out[2478] <= layer1_out[9922] & ~layer1_out[9923];
     layer2_out[2479] <= layer1_out[7705] & layer1_out[7706];
     layer2_out[2480] <= ~(layer1_out[11617] | layer1_out[11618]);
     layer2_out[2481] <= layer1_out[32] & ~layer1_out[33];
     layer2_out[2482] <= ~layer1_out[8232] | layer1_out[8233];
     layer2_out[2483] <= layer1_out[8852];
     layer2_out[2484] <= layer1_out[185] & layer1_out[186];
     layer2_out[2485] <= layer1_out[2667] & layer1_out[2668];
     layer2_out[2486] <= ~layer1_out[1605];
     layer2_out[2487] <= layer1_out[9757];
     layer2_out[2488] <= ~layer1_out[6439];
     layer2_out[2489] <= ~(layer1_out[2166] & layer1_out[2167]);
     layer2_out[2490] <= layer1_out[10804] ^ layer1_out[10805];
     layer2_out[2491] <= ~(layer1_out[8233] | layer1_out[8234]);
     layer2_out[2492] <= ~layer1_out[6529];
     layer2_out[2493] <= ~(layer1_out[2761] & layer1_out[2762]);
     layer2_out[2494] <= layer1_out[802] & ~layer1_out[801];
     layer2_out[2495] <= layer1_out[6726] & ~layer1_out[6727];
     layer2_out[2496] <= layer1_out[4533];
     layer2_out[2497] <= ~layer1_out[1650];
     layer2_out[2498] <= ~(layer1_out[10763] | layer1_out[10764]);
     layer2_out[2499] <= ~layer1_out[10992];
     layer2_out[2500] <= layer1_out[1582];
     layer2_out[2501] <= layer1_out[483] | layer1_out[484];
     layer2_out[2502] <= layer1_out[941];
     layer2_out[2503] <= ~(layer1_out[2299] ^ layer1_out[2300]);
     layer2_out[2504] <= ~layer1_out[7422];
     layer2_out[2505] <= ~layer1_out[686];
     layer2_out[2506] <= ~(layer1_out[3645] & layer1_out[3646]);
     layer2_out[2507] <= ~layer1_out[758];
     layer2_out[2508] <= ~layer1_out[3685];
     layer2_out[2509] <= ~layer1_out[5842] | layer1_out[5843];
     layer2_out[2510] <= layer1_out[7727];
     layer2_out[2511] <= layer1_out[8641];
     layer2_out[2512] <= layer1_out[9580];
     layer2_out[2513] <= ~(layer1_out[1500] & layer1_out[1501]);
     layer2_out[2514] <= layer1_out[4385] & ~layer1_out[4386];
     layer2_out[2515] <= ~layer1_out[6564] | layer1_out[6565];
     layer2_out[2516] <= ~layer1_out[1974];
     layer2_out[2517] <= ~(layer1_out[8212] & layer1_out[8213]);
     layer2_out[2518] <= layer1_out[2803] ^ layer1_out[2804];
     layer2_out[2519] <= ~(layer1_out[11620] | layer1_out[11621]);
     layer2_out[2520] <= layer1_out[8956] | layer1_out[8957];
     layer2_out[2521] <= layer1_out[505] & ~layer1_out[504];
     layer2_out[2522] <= layer1_out[1333];
     layer2_out[2523] <= ~(layer1_out[3439] & layer1_out[3440]);
     layer2_out[2524] <= layer1_out[2344] | layer1_out[2345];
     layer2_out[2525] <= layer1_out[4125];
     layer2_out[2526] <= ~layer1_out[7636] | layer1_out[7635];
     layer2_out[2527] <= layer1_out[6769];
     layer2_out[2528] <= layer1_out[4933] | layer1_out[4934];
     layer2_out[2529] <= layer1_out[1522] & ~layer1_out[1523];
     layer2_out[2530] <= layer1_out[2035] & ~layer1_out[2036];
     layer2_out[2531] <= layer1_out[1582] & layer1_out[1583];
     layer2_out[2532] <= layer1_out[4106] | layer1_out[4107];
     layer2_out[2533] <= ~layer1_out[1272] | layer1_out[1271];
     layer2_out[2534] <= layer1_out[10183];
     layer2_out[2535] <= layer1_out[4557];
     layer2_out[2536] <= layer1_out[905];
     layer2_out[2537] <= ~(layer1_out[5138] ^ layer1_out[5139]);
     layer2_out[2538] <= ~layer1_out[8826];
     layer2_out[2539] <= layer1_out[7574] & ~layer1_out[7573];
     layer2_out[2540] <= ~(layer1_out[5208] & layer1_out[5209]);
     layer2_out[2541] <= layer1_out[2209] & ~layer1_out[2210];
     layer2_out[2542] <= layer1_out[9551] & ~layer1_out[9550];
     layer2_out[2543] <= layer1_out[8611];
     layer2_out[2544] <= ~layer1_out[4132];
     layer2_out[2545] <= layer1_out[6400];
     layer2_out[2546] <= ~layer1_out[1816] | layer1_out[1817];
     layer2_out[2547] <= ~layer1_out[8197] | layer1_out[8196];
     layer2_out[2548] <= layer1_out[7188];
     layer2_out[2549] <= ~layer1_out[10968] | layer1_out[10969];
     layer2_out[2550] <= ~(layer1_out[6557] & layer1_out[6558]);
     layer2_out[2551] <= ~layer1_out[10661];
     layer2_out[2552] <= layer1_out[5403];
     layer2_out[2553] <= ~layer1_out[11082] | layer1_out[11081];
     layer2_out[2554] <= layer1_out[4925] & ~layer1_out[4924];
     layer2_out[2555] <= layer1_out[5816] | layer1_out[5817];
     layer2_out[2556] <= ~layer1_out[2411] | layer1_out[2412];
     layer2_out[2557] <= ~layer1_out[10365];
     layer2_out[2558] <= ~layer1_out[759];
     layer2_out[2559] <= layer1_out[6121] & ~layer1_out[6122];
     layer2_out[2560] <= ~layer1_out[1294];
     layer2_out[2561] <= layer1_out[3569] & ~layer1_out[3570];
     layer2_out[2562] <= layer1_out[11803] | layer1_out[11804];
     layer2_out[2563] <= layer1_out[10811];
     layer2_out[2564] <= ~layer1_out[8745];
     layer2_out[2565] <= 1'b1;
     layer2_out[2566] <= ~(layer1_out[714] & layer1_out[715]);
     layer2_out[2567] <= ~layer1_out[7621] | layer1_out[7622];
     layer2_out[2568] <= layer1_out[3813];
     layer2_out[2569] <= ~layer1_out[11733] | layer1_out[11734];
     layer2_out[2570] <= ~layer1_out[5844] | layer1_out[5845];
     layer2_out[2571] <= layer1_out[3228] | layer1_out[3229];
     layer2_out[2572] <= ~(layer1_out[8301] | layer1_out[8302]);
     layer2_out[2573] <= ~layer1_out[10431] | layer1_out[10432];
     layer2_out[2574] <= ~(layer1_out[1887] ^ layer1_out[1888]);
     layer2_out[2575] <= layer1_out[7995] | layer1_out[7996];
     layer2_out[2576] <= ~layer1_out[11491];
     layer2_out[2577] <= layer1_out[6414];
     layer2_out[2578] <= ~layer1_out[5695];
     layer2_out[2579] <= ~layer1_out[4523];
     layer2_out[2580] <= ~(layer1_out[4631] | layer1_out[4632]);
     layer2_out[2581] <= ~(layer1_out[1371] ^ layer1_out[1372]);
     layer2_out[2582] <= ~layer1_out[7380] | layer1_out[7379];
     layer2_out[2583] <= layer1_out[6375] ^ layer1_out[6376];
     layer2_out[2584] <= ~layer1_out[4931];
     layer2_out[2585] <= layer1_out[705] & ~layer1_out[706];
     layer2_out[2586] <= ~layer1_out[8330];
     layer2_out[2587] <= ~(layer1_out[7430] & layer1_out[7431]);
     layer2_out[2588] <= layer1_out[2108];
     layer2_out[2589] <= ~(layer1_out[1698] ^ layer1_out[1699]);
     layer2_out[2590] <= ~(layer1_out[3206] ^ layer1_out[3207]);
     layer2_out[2591] <= ~layer1_out[10860];
     layer2_out[2592] <= layer1_out[8497] | layer1_out[8498];
     layer2_out[2593] <= ~(layer1_out[1036] | layer1_out[1037]);
     layer2_out[2594] <= ~(layer1_out[11282] ^ layer1_out[11283]);
     layer2_out[2595] <= 1'b1;
     layer2_out[2596] <= layer1_out[8639] & ~layer1_out[8640];
     layer2_out[2597] <= layer1_out[2753];
     layer2_out[2598] <= ~layer1_out[525];
     layer2_out[2599] <= layer1_out[1010] & ~layer1_out[1011];
     layer2_out[2600] <= ~layer1_out[6520];
     layer2_out[2601] <= layer1_out[4520] & ~layer1_out[4519];
     layer2_out[2602] <= ~(layer1_out[637] & layer1_out[638]);
     layer2_out[2603] <= layer1_out[11948];
     layer2_out[2604] <= ~layer1_out[11766];
     layer2_out[2605] <= layer1_out[7067];
     layer2_out[2606] <= ~(layer1_out[11633] | layer1_out[11634]);
     layer2_out[2607] <= 1'b1;
     layer2_out[2608] <= ~layer1_out[5626];
     layer2_out[2609] <= ~layer1_out[10056] | layer1_out[10057];
     layer2_out[2610] <= ~(layer1_out[7628] | layer1_out[7629]);
     layer2_out[2611] <= ~(layer1_out[6358] ^ layer1_out[6359]);
     layer2_out[2612] <= ~layer1_out[10095];
     layer2_out[2613] <= layer1_out[643] & ~layer1_out[644];
     layer2_out[2614] <= ~(layer1_out[7719] ^ layer1_out[7720]);
     layer2_out[2615] <= layer1_out[10311];
     layer2_out[2616] <= layer1_out[5227] & layer1_out[5228];
     layer2_out[2617] <= ~(layer1_out[2272] ^ layer1_out[2273]);
     layer2_out[2618] <= layer1_out[967];
     layer2_out[2619] <= ~layer1_out[3921];
     layer2_out[2620] <= ~layer1_out[4507];
     layer2_out[2621] <= ~layer1_out[2813];
     layer2_out[2622] <= ~layer1_out[4414];
     layer2_out[2623] <= ~(layer1_out[8229] | layer1_out[8230]);
     layer2_out[2624] <= ~(layer1_out[9770] | layer1_out[9771]);
     layer2_out[2625] <= layer1_out[2852] & ~layer1_out[2853];
     layer2_out[2626] <= ~layer1_out[6936];
     layer2_out[2627] <= ~layer1_out[827] | layer1_out[826];
     layer2_out[2628] <= ~layer1_out[1980];
     layer2_out[2629] <= ~layer1_out[1439];
     layer2_out[2630] <= ~layer1_out[5998];
     layer2_out[2631] <= layer1_out[5076] | layer1_out[5077];
     layer2_out[2632] <= ~layer1_out[1983];
     layer2_out[2633] <= ~layer1_out[11675];
     layer2_out[2634] <= ~(layer1_out[11434] & layer1_out[11435]);
     layer2_out[2635] <= layer1_out[319] & layer1_out[320];
     layer2_out[2636] <= ~layer1_out[6387];
     layer2_out[2637] <= layer1_out[1353] & layer1_out[1354];
     layer2_out[2638] <= ~(layer1_out[2775] | layer1_out[2776]);
     layer2_out[2639] <= ~layer1_out[2674];
     layer2_out[2640] <= ~layer1_out[6366];
     layer2_out[2641] <= layer1_out[6906] | layer1_out[6907];
     layer2_out[2642] <= layer1_out[363];
     layer2_out[2643] <= layer1_out[9619];
     layer2_out[2644] <= layer1_out[9350];
     layer2_out[2645] <= layer1_out[5297];
     layer2_out[2646] <= 1'b1;
     layer2_out[2647] <= layer1_out[2380] ^ layer1_out[2381];
     layer2_out[2648] <= layer1_out[3335];
     layer2_out[2649] <= layer1_out[7320] | layer1_out[7321];
     layer2_out[2650] <= layer1_out[11027];
     layer2_out[2651] <= ~layer1_out[9262];
     layer2_out[2652] <= ~(layer1_out[11260] & layer1_out[11261]);
     layer2_out[2653] <= ~layer1_out[8929];
     layer2_out[2654] <= ~layer1_out[3776];
     layer2_out[2655] <= ~layer1_out[9167] | layer1_out[9166];
     layer2_out[2656] <= ~(layer1_out[3866] ^ layer1_out[3867]);
     layer2_out[2657] <= ~(layer1_out[7442] ^ layer1_out[7443]);
     layer2_out[2658] <= layer1_out[10997];
     layer2_out[2659] <= layer1_out[6340];
     layer2_out[2660] <= ~(layer1_out[7418] | layer1_out[7419]);
     layer2_out[2661] <= ~(layer1_out[3389] ^ layer1_out[3390]);
     layer2_out[2662] <= ~layer1_out[7075];
     layer2_out[2663] <= ~layer1_out[3718] | layer1_out[3719];
     layer2_out[2664] <= layer1_out[2790] | layer1_out[2791];
     layer2_out[2665] <= ~layer1_out[1619] | layer1_out[1618];
     layer2_out[2666] <= ~layer1_out[7119];
     layer2_out[2667] <= ~layer1_out[3434] | layer1_out[3435];
     layer2_out[2668] <= layer1_out[10635] & ~layer1_out[10634];
     layer2_out[2669] <= ~(layer1_out[2044] ^ layer1_out[2045]);
     layer2_out[2670] <= layer1_out[2907] | layer1_out[2908];
     layer2_out[2671] <= ~(layer1_out[10437] & layer1_out[10438]);
     layer2_out[2672] <= ~layer1_out[5865];
     layer2_out[2673] <= layer1_out[1514] & ~layer1_out[1513];
     layer2_out[2674] <= ~(layer1_out[6400] | layer1_out[6401]);
     layer2_out[2675] <= layer1_out[2630] & ~layer1_out[2631];
     layer2_out[2676] <= layer1_out[1392];
     layer2_out[2677] <= ~(layer1_out[7380] ^ layer1_out[7381]);
     layer2_out[2678] <= ~(layer1_out[9829] ^ layer1_out[9830]);
     layer2_out[2679] <= layer1_out[3380];
     layer2_out[2680] <= ~layer1_out[6030];
     layer2_out[2681] <= ~(layer1_out[4483] | layer1_out[4484]);
     layer2_out[2682] <= ~layer1_out[8577];
     layer2_out[2683] <= layer1_out[10656] ^ layer1_out[10657];
     layer2_out[2684] <= layer1_out[4882] & ~layer1_out[4881];
     layer2_out[2685] <= layer1_out[8353];
     layer2_out[2686] <= ~layer1_out[2170] | layer1_out[2171];
     layer2_out[2687] <= ~layer1_out[3379] | layer1_out[3380];
     layer2_out[2688] <= ~(layer1_out[7539] ^ layer1_out[7540]);
     layer2_out[2689] <= ~(layer1_out[4141] & layer1_out[4142]);
     layer2_out[2690] <= ~layer1_out[3522] | layer1_out[3521];
     layer2_out[2691] <= ~layer1_out[4935];
     layer2_out[2692] <= ~layer1_out[9335];
     layer2_out[2693] <= layer1_out[10630];
     layer2_out[2694] <= ~layer1_out[438] | layer1_out[437];
     layer2_out[2695] <= layer1_out[352] & ~layer1_out[351];
     layer2_out[2696] <= ~layer1_out[6990] | layer1_out[6989];
     layer2_out[2697] <= ~layer1_out[3244];
     layer2_out[2698] <= layer1_out[1614];
     layer2_out[2699] <= ~(layer1_out[8661] & layer1_out[8662]);
     layer2_out[2700] <= ~(layer1_out[6608] & layer1_out[6609]);
     layer2_out[2701] <= ~layer1_out[2273] | layer1_out[2274];
     layer2_out[2702] <= layer1_out[9706] | layer1_out[9707];
     layer2_out[2703] <= layer1_out[6161] & ~layer1_out[6162];
     layer2_out[2704] <= layer1_out[8104];
     layer2_out[2705] <= layer1_out[9565] | layer1_out[9566];
     layer2_out[2706] <= ~layer1_out[4762] | layer1_out[4761];
     layer2_out[2707] <= layer1_out[11778] ^ layer1_out[11779];
     layer2_out[2708] <= layer1_out[5638] & ~layer1_out[5639];
     layer2_out[2709] <= layer1_out[3924] & ~layer1_out[3923];
     layer2_out[2710] <= layer1_out[5032];
     layer2_out[2711] <= ~(layer1_out[6463] & layer1_out[6464]);
     layer2_out[2712] <= ~layer1_out[9792];
     layer2_out[2713] <= ~layer1_out[6722] | layer1_out[6723];
     layer2_out[2714] <= layer1_out[1299] & layer1_out[1300];
     layer2_out[2715] <= layer1_out[11614] | layer1_out[11615];
     layer2_out[2716] <= layer1_out[3721] ^ layer1_out[3722];
     layer2_out[2717] <= layer1_out[1847] & ~layer1_out[1846];
     layer2_out[2718] <= layer1_out[9502] & layer1_out[9503];
     layer2_out[2719] <= ~(layer1_out[10260] | layer1_out[10261]);
     layer2_out[2720] <= ~(layer1_out[1711] & layer1_out[1712]);
     layer2_out[2721] <= layer1_out[7319] ^ layer1_out[7320];
     layer2_out[2722] <= ~layer1_out[598];
     layer2_out[2723] <= layer1_out[8868];
     layer2_out[2724] <= layer1_out[2414] & ~layer1_out[2413];
     layer2_out[2725] <= layer1_out[5684] & ~layer1_out[5683];
     layer2_out[2726] <= ~layer1_out[10592] | layer1_out[10593];
     layer2_out[2727] <= ~layer1_out[8442];
     layer2_out[2728] <= layer1_out[2484];
     layer2_out[2729] <= layer1_out[8036] & ~layer1_out[8035];
     layer2_out[2730] <= ~(layer1_out[9106] & layer1_out[9107]);
     layer2_out[2731] <= ~layer1_out[6717];
     layer2_out[2732] <= ~layer1_out[149];
     layer2_out[2733] <= ~layer1_out[4137] | layer1_out[4136];
     layer2_out[2734] <= ~(layer1_out[2839] ^ layer1_out[2840]);
     layer2_out[2735] <= ~layer1_out[6903] | layer1_out[6904];
     layer2_out[2736] <= ~layer1_out[11544];
     layer2_out[2737] <= layer1_out[6374] ^ layer1_out[6375];
     layer2_out[2738] <= layer1_out[6383];
     layer2_out[2739] <= ~(layer1_out[118] ^ layer1_out[119]);
     layer2_out[2740] <= layer1_out[7266] & layer1_out[7267];
     layer2_out[2741] <= layer1_out[11510] | layer1_out[11511];
     layer2_out[2742] <= layer1_out[11473] & ~layer1_out[11472];
     layer2_out[2743] <= layer1_out[2183] | layer1_out[2184];
     layer2_out[2744] <= layer1_out[9975];
     layer2_out[2745] <= ~layer1_out[5145];
     layer2_out[2746] <= layer1_out[9452];
     layer2_out[2747] <= ~layer1_out[5905];
     layer2_out[2748] <= ~layer1_out[8515] | layer1_out[8514];
     layer2_out[2749] <= ~layer1_out[10331] | layer1_out[10332];
     layer2_out[2750] <= layer1_out[534];
     layer2_out[2751] <= layer1_out[8989] ^ layer1_out[8990];
     layer2_out[2752] <= layer1_out[1064] ^ layer1_out[1065];
     layer2_out[2753] <= layer1_out[8228] | layer1_out[8229];
     layer2_out[2754] <= layer1_out[421];
     layer2_out[2755] <= ~layer1_out[10256] | layer1_out[10255];
     layer2_out[2756] <= layer1_out[4454] & ~layer1_out[4453];
     layer2_out[2757] <= layer1_out[11165];
     layer2_out[2758] <= ~layer1_out[1783] | layer1_out[1784];
     layer2_out[2759] <= ~layer1_out[7590] | layer1_out[7589];
     layer2_out[2760] <= ~(layer1_out[10588] ^ layer1_out[10589]);
     layer2_out[2761] <= ~layer1_out[6110];
     layer2_out[2762] <= layer1_out[10469] & layer1_out[10470];
     layer2_out[2763] <= layer1_out[4102];
     layer2_out[2764] <= ~layer1_out[11440];
     layer2_out[2765] <= 1'b0;
     layer2_out[2766] <= layer1_out[5322] & ~layer1_out[5321];
     layer2_out[2767] <= layer1_out[5401] | layer1_out[5402];
     layer2_out[2768] <= ~(layer1_out[9521] | layer1_out[9522]);
     layer2_out[2769] <= layer1_out[9766] & layer1_out[9767];
     layer2_out[2770] <= layer1_out[1329] | layer1_out[1330];
     layer2_out[2771] <= layer1_out[6993] & ~layer1_out[6992];
     layer2_out[2772] <= layer1_out[410];
     layer2_out[2773] <= ~layer1_out[7593];
     layer2_out[2774] <= ~layer1_out[5655];
     layer2_out[2775] <= ~(layer1_out[111] | layer1_out[112]);
     layer2_out[2776] <= layer1_out[4894] & ~layer1_out[4895];
     layer2_out[2777] <= layer1_out[6543] & ~layer1_out[6542];
     layer2_out[2778] <= layer1_out[6196] ^ layer1_out[6197];
     layer2_out[2779] <= layer1_out[2037];
     layer2_out[2780] <= layer1_out[11526] & layer1_out[11527];
     layer2_out[2781] <= layer1_out[3784] & layer1_out[3785];
     layer2_out[2782] <= layer1_out[3805];
     layer2_out[2783] <= layer1_out[10299] | layer1_out[10300];
     layer2_out[2784] <= layer1_out[115] & ~layer1_out[116];
     layer2_out[2785] <= ~(layer1_out[1777] & layer1_out[1778]);
     layer2_out[2786] <= layer1_out[9237];
     layer2_out[2787] <= ~(layer1_out[5804] ^ layer1_out[5805]);
     layer2_out[2788] <= ~(layer1_out[6534] | layer1_out[6535]);
     layer2_out[2789] <= ~layer1_out[6693] | layer1_out[6694];
     layer2_out[2790] <= layer1_out[10707] & ~layer1_out[10706];
     layer2_out[2791] <= layer1_out[100] & ~layer1_out[101];
     layer2_out[2792] <= layer1_out[2379] | layer1_out[2380];
     layer2_out[2793] <= ~(layer1_out[5884] & layer1_out[5885]);
     layer2_out[2794] <= layer1_out[11318];
     layer2_out[2795] <= layer1_out[6196] & ~layer1_out[6195];
     layer2_out[2796] <= ~layer1_out[434];
     layer2_out[2797] <= ~(layer1_out[8840] ^ layer1_out[8841]);
     layer2_out[2798] <= ~layer1_out[9158] | layer1_out[9159];
     layer2_out[2799] <= ~(layer1_out[2470] ^ layer1_out[2471]);
     layer2_out[2800] <= ~layer1_out[2422];
     layer2_out[2801] <= ~layer1_out[11910];
     layer2_out[2802] <= layer1_out[7025] ^ layer1_out[7026];
     layer2_out[2803] <= layer1_out[7174] & ~layer1_out[7175];
     layer2_out[2804] <= ~layer1_out[8440];
     layer2_out[2805] <= ~layer1_out[5512];
     layer2_out[2806] <= ~(layer1_out[5998] & layer1_out[5999]);
     layer2_out[2807] <= ~(layer1_out[11666] | layer1_out[11667]);
     layer2_out[2808] <= layer1_out[5767] & ~layer1_out[5768];
     layer2_out[2809] <= ~layer1_out[5261];
     layer2_out[2810] <= layer1_out[10548];
     layer2_out[2811] <= layer1_out[5731];
     layer2_out[2812] <= layer1_out[2124] & ~layer1_out[2125];
     layer2_out[2813] <= ~layer1_out[10817];
     layer2_out[2814] <= ~(layer1_out[9777] | layer1_out[9778]);
     layer2_out[2815] <= ~layer1_out[4297];
     layer2_out[2816] <= ~layer1_out[601] | layer1_out[600];
     layer2_out[2817] <= layer1_out[6170];
     layer2_out[2818] <= layer1_out[8681] | layer1_out[8682];
     layer2_out[2819] <= ~(layer1_out[5718] & layer1_out[5719]);
     layer2_out[2820] <= ~(layer1_out[3002] | layer1_out[3003]);
     layer2_out[2821] <= layer1_out[6055] | layer1_out[6056];
     layer2_out[2822] <= ~layer1_out[1023] | layer1_out[1024];
     layer2_out[2823] <= layer1_out[10057] & layer1_out[10058];
     layer2_out[2824] <= layer1_out[6590];
     layer2_out[2825] <= layer1_out[3087] | layer1_out[3088];
     layer2_out[2826] <= layer1_out[4295];
     layer2_out[2827] <= layer1_out[5178];
     layer2_out[2828] <= ~(layer1_out[2795] | layer1_out[2796]);
     layer2_out[2829] <= ~(layer1_out[9988] | layer1_out[9989]);
     layer2_out[2830] <= ~(layer1_out[5365] | layer1_out[5366]);
     layer2_out[2831] <= ~(layer1_out[10034] & layer1_out[10035]);
     layer2_out[2832] <= ~(layer1_out[8473] | layer1_out[8474]);
     layer2_out[2833] <= ~layer1_out[675] | layer1_out[676];
     layer2_out[2834] <= layer1_out[5873] & layer1_out[5874];
     layer2_out[2835] <= 1'b1;
     layer2_out[2836] <= ~layer1_out[1013];
     layer2_out[2837] <= layer1_out[6616];
     layer2_out[2838] <= ~(layer1_out[4943] | layer1_out[4944]);
     layer2_out[2839] <= ~(layer1_out[11074] & layer1_out[11075]);
     layer2_out[2840] <= ~layer1_out[7868] | layer1_out[7869];
     layer2_out[2841] <= layer1_out[4064] ^ layer1_out[4065];
     layer2_out[2842] <= layer1_out[9197] & ~layer1_out[9198];
     layer2_out[2843] <= layer1_out[7356] & ~layer1_out[7357];
     layer2_out[2844] <= layer1_out[2987];
     layer2_out[2845] <= ~layer1_out[9712] | layer1_out[9711];
     layer2_out[2846] <= ~layer1_out[9998];
     layer2_out[2847] <= layer1_out[1023];
     layer2_out[2848] <= layer1_out[5301] & ~layer1_out[5300];
     layer2_out[2849] <= layer1_out[2698] & layer1_out[2699];
     layer2_out[2850] <= ~layer1_out[11098];
     layer2_out[2851] <= layer1_out[122];
     layer2_out[2852] <= ~layer1_out[11936];
     layer2_out[2853] <= ~layer1_out[3371];
     layer2_out[2854] <= layer1_out[5982];
     layer2_out[2855] <= ~(layer1_out[2897] & layer1_out[2898]);
     layer2_out[2856] <= ~layer1_out[6298] | layer1_out[6299];
     layer2_out[2857] <= ~layer1_out[7556];
     layer2_out[2858] <= ~(layer1_out[3730] | layer1_out[3731]);
     layer2_out[2859] <= layer1_out[8527] & layer1_out[8528];
     layer2_out[2860] <= layer1_out[8667];
     layer2_out[2861] <= ~(layer1_out[278] ^ layer1_out[279]);
     layer2_out[2862] <= ~(layer1_out[10511] ^ layer1_out[10512]);
     layer2_out[2863] <= layer1_out[9161];
     layer2_out[2864] <= layer1_out[4086] & layer1_out[4087];
     layer2_out[2865] <= ~(layer1_out[11212] | layer1_out[11213]);
     layer2_out[2866] <= layer1_out[3056];
     layer2_out[2867] <= layer1_out[5660];
     layer2_out[2868] <= ~layer1_out[3228];
     layer2_out[2869] <= ~(layer1_out[9118] ^ layer1_out[9119]);
     layer2_out[2870] <= layer1_out[8070] & ~layer1_out[8069];
     layer2_out[2871] <= layer1_out[8771];
     layer2_out[2872] <= layer1_out[842] ^ layer1_out[843];
     layer2_out[2873] <= layer1_out[3804];
     layer2_out[2874] <= layer1_out[10008] & layer1_out[10009];
     layer2_out[2875] <= ~layer1_out[6474];
     layer2_out[2876] <= layer1_out[9995];
     layer2_out[2877] <= ~layer1_out[10125];
     layer2_out[2878] <= ~layer1_out[9084] | layer1_out[9083];
     layer2_out[2879] <= layer1_out[1158];
     layer2_out[2880] <= ~(layer1_out[8341] & layer1_out[8342]);
     layer2_out[2881] <= ~(layer1_out[891] | layer1_out[892]);
     layer2_out[2882] <= layer1_out[4830] | layer1_out[4831];
     layer2_out[2883] <= layer1_out[7563] | layer1_out[7564];
     layer2_out[2884] <= ~layer1_out[6151] | layer1_out[6152];
     layer2_out[2885] <= layer1_out[3097];
     layer2_out[2886] <= ~layer1_out[9880];
     layer2_out[2887] <= layer1_out[7617] & ~layer1_out[7616];
     layer2_out[2888] <= layer1_out[7757];
     layer2_out[2889] <= ~(layer1_out[1626] & layer1_out[1627]);
     layer2_out[2890] <= ~layer1_out[6350];
     layer2_out[2891] <= layer1_out[4686];
     layer2_out[2892] <= layer1_out[11452] & layer1_out[11453];
     layer2_out[2893] <= ~layer1_out[4340];
     layer2_out[2894] <= ~layer1_out[5265];
     layer2_out[2895] <= ~layer1_out[8226];
     layer2_out[2896] <= layer1_out[1547] & ~layer1_out[1548];
     layer2_out[2897] <= ~(layer1_out[8785] & layer1_out[8786]);
     layer2_out[2898] <= ~(layer1_out[8360] ^ layer1_out[8361]);
     layer2_out[2899] <= 1'b0;
     layer2_out[2900] <= ~(layer1_out[1715] ^ layer1_out[1716]);
     layer2_out[2901] <= ~layer1_out[1908] | layer1_out[1909];
     layer2_out[2902] <= ~layer1_out[5979] | layer1_out[5980];
     layer2_out[2903] <= ~(layer1_out[8538] | layer1_out[8539]);
     layer2_out[2904] <= layer1_out[4200] & layer1_out[4201];
     layer2_out[2905] <= ~layer1_out[6442];
     layer2_out[2906] <= layer1_out[3347] & layer1_out[3348];
     layer2_out[2907] <= layer1_out[2786];
     layer2_out[2908] <= 1'b1;
     layer2_out[2909] <= layer1_out[4595] & ~layer1_out[4596];
     layer2_out[2910] <= ~layer1_out[10561] | layer1_out[10562];
     layer2_out[2911] <= ~layer1_out[3557];
     layer2_out[2912] <= ~(layer1_out[7687] & layer1_out[7688]);
     layer2_out[2913] <= ~(layer1_out[1354] & layer1_out[1355]);
     layer2_out[2914] <= ~layer1_out[2348];
     layer2_out[2915] <= ~layer1_out[6502];
     layer2_out[2916] <= ~layer1_out[9278] | layer1_out[9279];
     layer2_out[2917] <= layer1_out[3628] ^ layer1_out[3629];
     layer2_out[2918] <= layer1_out[6274] ^ layer1_out[6275];
     layer2_out[2919] <= layer1_out[11130] & ~layer1_out[11131];
     layer2_out[2920] <= ~layer1_out[11411] | layer1_out[11412];
     layer2_out[2921] <= ~(layer1_out[5099] | layer1_out[5100]);
     layer2_out[2922] <= ~(layer1_out[3011] & layer1_out[3012]);
     layer2_out[2923] <= layer1_out[9775] | layer1_out[9776];
     layer2_out[2924] <= ~layer1_out[9764] | layer1_out[9765];
     layer2_out[2925] <= layer1_out[3337] & ~layer1_out[3338];
     layer2_out[2926] <= layer1_out[2876] & ~layer1_out[2877];
     layer2_out[2927] <= ~layer1_out[2152] | layer1_out[2153];
     layer2_out[2928] <= layer1_out[4165] ^ layer1_out[4166];
     layer2_out[2929] <= ~layer1_out[1565];
     layer2_out[2930] <= layer1_out[8328];
     layer2_out[2931] <= ~layer1_out[1920];
     layer2_out[2932] <= layer1_out[5197];
     layer2_out[2933] <= layer1_out[8611] & ~layer1_out[8610];
     layer2_out[2934] <= ~layer1_out[4286] | layer1_out[4287];
     layer2_out[2935] <= ~layer1_out[11428];
     layer2_out[2936] <= ~layer1_out[9608];
     layer2_out[2937] <= layer1_out[5448];
     layer2_out[2938] <= ~layer1_out[2929];
     layer2_out[2939] <= layer1_out[8008] & ~layer1_out[8007];
     layer2_out[2940] <= layer1_out[1500];
     layer2_out[2941] <= layer1_out[9245];
     layer2_out[2942] <= ~layer1_out[1143];
     layer2_out[2943] <= ~layer1_out[924];
     layer2_out[2944] <= ~layer1_out[10457] | layer1_out[10458];
     layer2_out[2945] <= layer1_out[3348];
     layer2_out[2946] <= ~(layer1_out[10669] | layer1_out[10670]);
     layer2_out[2947] <= ~layer1_out[7943];
     layer2_out[2948] <= layer1_out[3258] & layer1_out[3259];
     layer2_out[2949] <= layer1_out[7453] & layer1_out[7454];
     layer2_out[2950] <= layer1_out[4781] & ~layer1_out[4782];
     layer2_out[2951] <= ~layer1_out[304];
     layer2_out[2952] <= layer1_out[8732] & ~layer1_out[8733];
     layer2_out[2953] <= layer1_out[2935] & layer1_out[2936];
     layer2_out[2954] <= ~layer1_out[658];
     layer2_out[2955] <= layer1_out[8067] & layer1_out[8068];
     layer2_out[2956] <= ~layer1_out[1989];
     layer2_out[2957] <= ~(layer1_out[10067] ^ layer1_out[10068]);
     layer2_out[2958] <= ~layer1_out[8283];
     layer2_out[2959] <= layer1_out[9393];
     layer2_out[2960] <= ~(layer1_out[5808] & layer1_out[5809]);
     layer2_out[2961] <= ~(layer1_out[6273] & layer1_out[6274]);
     layer2_out[2962] <= layer1_out[2524] & ~layer1_out[2523];
     layer2_out[2963] <= layer1_out[6762];
     layer2_out[2964] <= ~layer1_out[2788] | layer1_out[2789];
     layer2_out[2965] <= layer1_out[7925];
     layer2_out[2966] <= layer1_out[7036] & layer1_out[7037];
     layer2_out[2967] <= layer1_out[8749] & layer1_out[8750];
     layer2_out[2968] <= layer1_out[5976];
     layer2_out[2969] <= layer1_out[8025];
     layer2_out[2970] <= layer1_out[11244] ^ layer1_out[11245];
     layer2_out[2971] <= ~layer1_out[4400] | layer1_out[4401];
     layer2_out[2972] <= ~layer1_out[114] | layer1_out[115];
     layer2_out[2973] <= layer1_out[10941];
     layer2_out[2974] <= ~layer1_out[8691];
     layer2_out[2975] <= ~layer1_out[503];
     layer2_out[2976] <= layer1_out[11889] & ~layer1_out[11890];
     layer2_out[2977] <= layer1_out[11969];
     layer2_out[2978] <= ~layer1_out[10372] | layer1_out[10373];
     layer2_out[2979] <= layer1_out[11334] | layer1_out[11335];
     layer2_out[2980] <= ~layer1_out[52];
     layer2_out[2981] <= layer1_out[3537];
     layer2_out[2982] <= ~(layer1_out[3686] & layer1_out[3687]);
     layer2_out[2983] <= ~(layer1_out[1080] ^ layer1_out[1081]);
     layer2_out[2984] <= ~layer1_out[10694];
     layer2_out[2985] <= ~(layer1_out[1432] ^ layer1_out[1433]);
     layer2_out[2986] <= ~(layer1_out[10399] ^ layer1_out[10400]);
     layer2_out[2987] <= layer1_out[5688];
     layer2_out[2988] <= ~layer1_out[7137] | layer1_out[7136];
     layer2_out[2989] <= ~layer1_out[6996] | layer1_out[6997];
     layer2_out[2990] <= layer1_out[2731] & ~layer1_out[2730];
     layer2_out[2991] <= ~layer1_out[8533];
     layer2_out[2992] <= ~(layer1_out[10326] | layer1_out[10327]);
     layer2_out[2993] <= layer1_out[2424] & ~layer1_out[2425];
     layer2_out[2994] <= layer1_out[1240] & layer1_out[1241];
     layer2_out[2995] <= ~layer1_out[5749];
     layer2_out[2996] <= ~layer1_out[9667] | layer1_out[9668];
     layer2_out[2997] <= layer1_out[899] ^ layer1_out[900];
     layer2_out[2998] <= ~layer1_out[3148];
     layer2_out[2999] <= ~(layer1_out[3172] | layer1_out[3173]);
     layer2_out[3000] <= layer1_out[9231] | layer1_out[9232];
     layer2_out[3001] <= ~(layer1_out[3174] | layer1_out[3175]);
     layer2_out[3002] <= ~layer1_out[1078];
     layer2_out[3003] <= layer1_out[620];
     layer2_out[3004] <= layer1_out[4002] & layer1_out[4003];
     layer2_out[3005] <= layer1_out[9141] | layer1_out[9142];
     layer2_out[3006] <= ~(layer1_out[3268] & layer1_out[3269]);
     layer2_out[3007] <= layer1_out[11396];
     layer2_out[3008] <= layer1_out[11688];
     layer2_out[3009] <= layer1_out[9589] ^ layer1_out[9590];
     layer2_out[3010] <= ~(layer1_out[2197] | layer1_out[2198]);
     layer2_out[3011] <= ~layer1_out[6904] | layer1_out[6905];
     layer2_out[3012] <= layer1_out[9672] & layer1_out[9673];
     layer2_out[3013] <= ~layer1_out[6644];
     layer2_out[3014] <= layer1_out[3300];
     layer2_out[3015] <= layer1_out[1521] ^ layer1_out[1522];
     layer2_out[3016] <= ~layer1_out[2993];
     layer2_out[3017] <= layer1_out[11482];
     layer2_out[3018] <= layer1_out[6016] ^ layer1_out[6017];
     layer2_out[3019] <= ~layer1_out[6161] | layer1_out[6160];
     layer2_out[3020] <= layer1_out[6157] ^ layer1_out[6158];
     layer2_out[3021] <= ~(layer1_out[11384] ^ layer1_out[11385]);
     layer2_out[3022] <= ~layer1_out[1364] | layer1_out[1363];
     layer2_out[3023] <= layer1_out[11567] & layer1_out[11568];
     layer2_out[3024] <= layer1_out[5914];
     layer2_out[3025] <= ~layer1_out[1661];
     layer2_out[3026] <= layer1_out[1241] & ~layer1_out[1242];
     layer2_out[3027] <= layer1_out[10874] & ~layer1_out[10873];
     layer2_out[3028] <= layer1_out[3658] & ~layer1_out[3657];
     layer2_out[3029] <= ~(layer1_out[8411] | layer1_out[8412]);
     layer2_out[3030] <= ~(layer1_out[3584] | layer1_out[3585]);
     layer2_out[3031] <= layer1_out[8573] & layer1_out[8574];
     layer2_out[3032] <= layer1_out[123] | layer1_out[124];
     layer2_out[3033] <= layer1_out[4890];
     layer2_out[3034] <= ~layer1_out[7835] | layer1_out[7836];
     layer2_out[3035] <= ~layer1_out[4886];
     layer2_out[3036] <= ~layer1_out[1000] | layer1_out[1001];
     layer2_out[3037] <= ~layer1_out[11825];
     layer2_out[3038] <= ~layer1_out[9401];
     layer2_out[3039] <= ~(layer1_out[3059] ^ layer1_out[3060]);
     layer2_out[3040] <= layer1_out[9152] & ~layer1_out[9151];
     layer2_out[3041] <= layer1_out[5079] & ~layer1_out[5078];
     layer2_out[3042] <= ~layer1_out[11726];
     layer2_out[3043] <= layer1_out[4294];
     layer2_out[3044] <= layer1_out[11934];
     layer2_out[3045] <= layer1_out[2608] & layer1_out[2609];
     layer2_out[3046] <= ~layer1_out[7284] | layer1_out[7285];
     layer2_out[3047] <= ~layer1_out[1859] | layer1_out[1858];
     layer2_out[3048] <= ~(layer1_out[10748] | layer1_out[10749]);
     layer2_out[3049] <= ~layer1_out[1840];
     layer2_out[3050] <= layer1_out[2428];
     layer2_out[3051] <= layer1_out[4011];
     layer2_out[3052] <= ~layer1_out[5515] | layer1_out[5516];
     layer2_out[3053] <= layer1_out[6971] | layer1_out[6972];
     layer2_out[3054] <= layer1_out[5011];
     layer2_out[3055] <= layer1_out[2846] | layer1_out[2847];
     layer2_out[3056] <= layer1_out[11345] & ~layer1_out[11346];
     layer2_out[3057] <= 1'b0;
     layer2_out[3058] <= layer1_out[10335] ^ layer1_out[10336];
     layer2_out[3059] <= layer1_out[6533] & ~layer1_out[6532];
     layer2_out[3060] <= ~(layer1_out[10514] & layer1_out[10515]);
     layer2_out[3061] <= layer1_out[2857];
     layer2_out[3062] <= layer1_out[10314] & ~layer1_out[10315];
     layer2_out[3063] <= ~layer1_out[9502];
     layer2_out[3064] <= layer1_out[3217];
     layer2_out[3065] <= ~layer1_out[8663] | layer1_out[8662];
     layer2_out[3066] <= layer1_out[6533];
     layer2_out[3067] <= ~layer1_out[10248] | layer1_out[10249];
     layer2_out[3068] <= ~layer1_out[7991];
     layer2_out[3069] <= ~(layer1_out[9444] | layer1_out[9445]);
     layer2_out[3070] <= ~layer1_out[3797];
     layer2_out[3071] <= ~(layer1_out[2174] ^ layer1_out[2175]);
     layer2_out[3072] <= layer1_out[2979] & ~layer1_out[2978];
     layer2_out[3073] <= ~layer1_out[11365];
     layer2_out[3074] <= ~layer1_out[1849];
     layer2_out[3075] <= layer1_out[2666] & layer1_out[2667];
     layer2_out[3076] <= ~layer1_out[3441];
     layer2_out[3077] <= layer1_out[8876];
     layer2_out[3078] <= layer1_out[3302] & ~layer1_out[3303];
     layer2_out[3079] <= ~(layer1_out[7918] & layer1_out[7919]);
     layer2_out[3080] <= ~layer1_out[9034];
     layer2_out[3081] <= ~(layer1_out[6878] ^ layer1_out[6879]);
     layer2_out[3082] <= ~(layer1_out[6842] & layer1_out[6843]);
     layer2_out[3083] <= ~layer1_out[9972] | layer1_out[9971];
     layer2_out[3084] <= ~layer1_out[1787] | layer1_out[1788];
     layer2_out[3085] <= ~layer1_out[8452];
     layer2_out[3086] <= ~layer1_out[10890];
     layer2_out[3087] <= layer1_out[8373] | layer1_out[8374];
     layer2_out[3088] <= layer1_out[6101] | layer1_out[6102];
     layer2_out[3089] <= layer1_out[16];
     layer2_out[3090] <= ~layer1_out[5548] | layer1_out[5547];
     layer2_out[3091] <= layer1_out[1795];
     layer2_out[3092] <= ~layer1_out[3023];
     layer2_out[3093] <= layer1_out[11069] ^ layer1_out[11070];
     layer2_out[3094] <= layer1_out[3678] & ~layer1_out[3677];
     layer2_out[3095] <= layer1_out[8224];
     layer2_out[3096] <= ~layer1_out[3419] | layer1_out[3420];
     layer2_out[3097] <= ~layer1_out[11157];
     layer2_out[3098] <= layer1_out[4987];
     layer2_out[3099] <= layer1_out[5080] & layer1_out[5081];
     layer2_out[3100] <= layer1_out[3809] | layer1_out[3810];
     layer2_out[3101] <= 1'b0;
     layer2_out[3102] <= ~(layer1_out[9516] ^ layer1_out[9517]);
     layer2_out[3103] <= ~(layer1_out[7078] | layer1_out[7079]);
     layer2_out[3104] <= layer1_out[3153];
     layer2_out[3105] <= layer1_out[4917] ^ layer1_out[4918];
     layer2_out[3106] <= ~layer1_out[2087];
     layer2_out[3107] <= ~layer1_out[6725];
     layer2_out[3108] <= layer1_out[5991] & ~layer1_out[5992];
     layer2_out[3109] <= ~layer1_out[7287];
     layer2_out[3110] <= ~layer1_out[3547];
     layer2_out[3111] <= layer1_out[540] | layer1_out[541];
     layer2_out[3112] <= layer1_out[9171] & ~layer1_out[9170];
     layer2_out[3113] <= 1'b1;
     layer2_out[3114] <= layer1_out[11254];
     layer2_out[3115] <= ~layer1_out[8769];
     layer2_out[3116] <= layer1_out[8820] & ~layer1_out[8819];
     layer2_out[3117] <= ~layer1_out[4502] | layer1_out[4503];
     layer2_out[3118] <= ~(layer1_out[11976] & layer1_out[11977]);
     layer2_out[3119] <= layer1_out[7093];
     layer2_out[3120] <= layer1_out[10783];
     layer2_out[3121] <= ~layer1_out[3316];
     layer2_out[3122] <= layer1_out[8016];
     layer2_out[3123] <= ~layer1_out[2476] | layer1_out[2475];
     layer2_out[3124] <= ~layer1_out[1225] | layer1_out[1226];
     layer2_out[3125] <= layer1_out[6621] & ~layer1_out[6620];
     layer2_out[3126] <= layer1_out[6955] & ~layer1_out[6956];
     layer2_out[3127] <= ~layer1_out[6050];
     layer2_out[3128] <= layer1_out[10051];
     layer2_out[3129] <= layer1_out[11987];
     layer2_out[3130] <= ~(layer1_out[3772] & layer1_out[3773]);
     layer2_out[3131] <= layer1_out[6239];
     layer2_out[3132] <= ~(layer1_out[6667] | layer1_out[6668]);
     layer2_out[3133] <= ~layer1_out[9868];
     layer2_out[3134] <= ~layer1_out[300];
     layer2_out[3135] <= ~layer1_out[7884];
     layer2_out[3136] <= ~layer1_out[8160];
     layer2_out[3137] <= ~layer1_out[11837];
     layer2_out[3138] <= layer1_out[8668];
     layer2_out[3139] <= layer1_out[4842];
     layer2_out[3140] <= layer1_out[1426];
     layer2_out[3141] <= ~layer1_out[8697];
     layer2_out[3142] <= ~layer1_out[5565] | layer1_out[5566];
     layer2_out[3143] <= layer1_out[11923] & layer1_out[11924];
     layer2_out[3144] <= layer1_out[11047] ^ layer1_out[11048];
     layer2_out[3145] <= layer1_out[5523];
     layer2_out[3146] <= layer1_out[4021];
     layer2_out[3147] <= layer1_out[4074];
     layer2_out[3148] <= ~layer1_out[5039];
     layer2_out[3149] <= layer1_out[8015] & layer1_out[8016];
     layer2_out[3150] <= ~layer1_out[9483];
     layer2_out[3151] <= layer1_out[9735] & ~layer1_out[9734];
     layer2_out[3152] <= layer1_out[6510] ^ layer1_out[6511];
     layer2_out[3153] <= layer1_out[6659];
     layer2_out[3154] <= ~layer1_out[1587];
     layer2_out[3155] <= layer1_out[2798];
     layer2_out[3156] <= layer1_out[4609];
     layer2_out[3157] <= ~layer1_out[7515];
     layer2_out[3158] <= ~layer1_out[4153];
     layer2_out[3159] <= layer1_out[6629] | layer1_out[6630];
     layer2_out[3160] <= layer1_out[7420];
     layer2_out[3161] <= layer1_out[5239] ^ layer1_out[5240];
     layer2_out[3162] <= layer1_out[6256] & ~layer1_out[6257];
     layer2_out[3163] <= ~layer1_out[177];
     layer2_out[3164] <= ~(layer1_out[11159] & layer1_out[11160]);
     layer2_out[3165] <= layer1_out[1967] & ~layer1_out[1968];
     layer2_out[3166] <= ~(layer1_out[3911] & layer1_out[3912]);
     layer2_out[3167] <= ~(layer1_out[6093] ^ layer1_out[6094]);
     layer2_out[3168] <= ~layer1_out[2973];
     layer2_out[3169] <= layer1_out[4966];
     layer2_out[3170] <= ~(layer1_out[4314] ^ layer1_out[4315]);
     layer2_out[3171] <= layer1_out[1277] & ~layer1_out[1276];
     layer2_out[3172] <= ~layer1_out[4674];
     layer2_out[3173] <= ~(layer1_out[4536] ^ layer1_out[4537]);
     layer2_out[3174] <= ~layer1_out[6543];
     layer2_out[3175] <= ~layer1_out[11084] | layer1_out[11085];
     layer2_out[3176] <= layer1_out[10522];
     layer2_out[3177] <= layer1_out[11867];
     layer2_out[3178] <= ~layer1_out[5861];
     layer2_out[3179] <= layer1_out[9109] & ~layer1_out[9108];
     layer2_out[3180] <= ~layer1_out[232];
     layer2_out[3181] <= ~layer1_out[6379] | layer1_out[6378];
     layer2_out[3182] <= layer1_out[955] | layer1_out[956];
     layer2_out[3183] <= layer1_out[4817];
     layer2_out[3184] <= layer1_out[9623] & ~layer1_out[9622];
     layer2_out[3185] <= layer1_out[8195];
     layer2_out[3186] <= layer1_out[7494] | layer1_out[7495];
     layer2_out[3187] <= layer1_out[11813] & ~layer1_out[11812];
     layer2_out[3188] <= layer1_out[6503] & layer1_out[6504];
     layer2_out[3189] <= ~layer1_out[4160] | layer1_out[4161];
     layer2_out[3190] <= ~layer1_out[3253];
     layer2_out[3191] <= ~layer1_out[3952];
     layer2_out[3192] <= ~layer1_out[1330] | layer1_out[1331];
     layer2_out[3193] <= layer1_out[6272];
     layer2_out[3194] <= layer1_out[10694] & ~layer1_out[10693];
     layer2_out[3195] <= ~(layer1_out[3599] | layer1_out[3600]);
     layer2_out[3196] <= layer1_out[11902];
     layer2_out[3197] <= layer1_out[2146];
     layer2_out[3198] <= ~(layer1_out[9452] ^ layer1_out[9453]);
     layer2_out[3199] <= ~layer1_out[5552] | layer1_out[5553];
     layer2_out[3200] <= ~layer1_out[3450] | layer1_out[3451];
     layer2_out[3201] <= layer1_out[6795] ^ layer1_out[6796];
     layer2_out[3202] <= layer1_out[5134] | layer1_out[5135];
     layer2_out[3203] <= layer1_out[11717];
     layer2_out[3204] <= layer1_out[4275] & ~layer1_out[4276];
     layer2_out[3205] <= ~layer1_out[9795];
     layer2_out[3206] <= layer1_out[5162] ^ layer1_out[5163];
     layer2_out[3207] <= ~layer1_out[4773] | layer1_out[4772];
     layer2_out[3208] <= layer1_out[2994] & layer1_out[2995];
     layer2_out[3209] <= ~(layer1_out[4998] ^ layer1_out[4999]);
     layer2_out[3210] <= ~layer1_out[4857];
     layer2_out[3211] <= ~layer1_out[10184];
     layer2_out[3212] <= ~layer1_out[6181];
     layer2_out[3213] <= layer1_out[10613] & ~layer1_out[10612];
     layer2_out[3214] <= ~(layer1_out[9399] ^ layer1_out[9400]);
     layer2_out[3215] <= layer1_out[5918] | layer1_out[5919];
     layer2_out[3216] <= layer1_out[9992];
     layer2_out[3217] <= ~layer1_out[9784];
     layer2_out[3218] <= ~(layer1_out[2214] ^ layer1_out[2215]);
     layer2_out[3219] <= ~layer1_out[2350];
     layer2_out[3220] <= ~layer1_out[8577];
     layer2_out[3221] <= ~layer1_out[1923];
     layer2_out[3222] <= layer1_out[11759] & ~layer1_out[11758];
     layer2_out[3223] <= layer1_out[2642] & layer1_out[2643];
     layer2_out[3224] <= ~(layer1_out[11521] & layer1_out[11522]);
     layer2_out[3225] <= ~layer1_out[2878] | layer1_out[2877];
     layer2_out[3226] <= layer1_out[5296] & layer1_out[5297];
     layer2_out[3227] <= layer1_out[8249] & ~layer1_out[8250];
     layer2_out[3228] <= ~(layer1_out[3370] & layer1_out[3371]);
     layer2_out[3229] <= layer1_out[5713] & layer1_out[5714];
     layer2_out[3230] <= ~(layer1_out[7545] | layer1_out[7546]);
     layer2_out[3231] <= ~layer1_out[3151];
     layer2_out[3232] <= ~(layer1_out[5409] & layer1_out[5410]);
     layer2_out[3233] <= ~layer1_out[966];
     layer2_out[3234] <= layer1_out[6199];
     layer2_out[3235] <= layer1_out[404];
     layer2_out[3236] <= ~layer1_out[473];
     layer2_out[3237] <= layer1_out[537] & ~layer1_out[536];
     layer2_out[3238] <= ~layer1_out[6247];
     layer2_out[3239] <= layer1_out[1970] & ~layer1_out[1971];
     layer2_out[3240] <= ~(layer1_out[3515] ^ layer1_out[3516]);
     layer2_out[3241] <= ~layer1_out[7565] | layer1_out[7564];
     layer2_out[3242] <= ~(layer1_out[8457] & layer1_out[8458]);
     layer2_out[3243] <= layer1_out[7983] & layer1_out[7984];
     layer2_out[3244] <= ~layer1_out[5298] | layer1_out[5299];
     layer2_out[3245] <= ~(layer1_out[1213] | layer1_out[1214]);
     layer2_out[3246] <= ~(layer1_out[5723] ^ layer1_out[5724]);
     layer2_out[3247] <= ~layer1_out[2777] | layer1_out[2778];
     layer2_out[3248] <= layer1_out[9239] & ~layer1_out[9240];
     layer2_out[3249] <= ~(layer1_out[8709] | layer1_out[8710]);
     layer2_out[3250] <= layer1_out[3687] & ~layer1_out[3688];
     layer2_out[3251] <= layer1_out[7520];
     layer2_out[3252] <= ~(layer1_out[9185] | layer1_out[9186]);
     layer2_out[3253] <= layer1_out[11076] | layer1_out[11077];
     layer2_out[3254] <= ~layer1_out[4287];
     layer2_out[3255] <= ~layer1_out[8104] | layer1_out[8105];
     layer2_out[3256] <= layer1_out[5092];
     layer2_out[3257] <= ~layer1_out[3005];
     layer2_out[3258] <= layer1_out[4575];
     layer2_out[3259] <= layer1_out[11009] & ~layer1_out[11008];
     layer2_out[3260] <= ~layer1_out[8422];
     layer2_out[3261] <= ~layer1_out[659];
     layer2_out[3262] <= 1'b0;
     layer2_out[3263] <= ~(layer1_out[104] | layer1_out[105]);
     layer2_out[3264] <= layer1_out[7053];
     layer2_out[3265] <= layer1_out[4880] | layer1_out[4881];
     layer2_out[3266] <= 1'b0;
     layer2_out[3267] <= ~(layer1_out[8562] ^ layer1_out[8563]);
     layer2_out[3268] <= ~layer1_out[9959];
     layer2_out[3269] <= ~layer1_out[7742] | layer1_out[7743];
     layer2_out[3270] <= layer1_out[11369];
     layer2_out[3271] <= layer1_out[442] & layer1_out[443];
     layer2_out[3272] <= ~layer1_out[5786];
     layer2_out[3273] <= ~layer1_out[8130];
     layer2_out[3274] <= layer1_out[7203] ^ layer1_out[7204];
     layer2_out[3275] <= layer1_out[7081] ^ layer1_out[7082];
     layer2_out[3276] <= ~layer1_out[3817];
     layer2_out[3277] <= ~layer1_out[695] | layer1_out[694];
     layer2_out[3278] <= ~(layer1_out[9168] ^ layer1_out[9169]);
     layer2_out[3279] <= layer1_out[4216];
     layer2_out[3280] <= ~layer1_out[5450];
     layer2_out[3281] <= layer1_out[11613] & layer1_out[11614];
     layer2_out[3282] <= ~layer1_out[4430];
     layer2_out[3283] <= 1'b1;
     layer2_out[3284] <= ~layer1_out[2524] | layer1_out[2525];
     layer2_out[3285] <= layer1_out[2281] & ~layer1_out[2282];
     layer2_out[3286] <= layer1_out[5242] & ~layer1_out[5243];
     layer2_out[3287] <= ~(layer1_out[5319] | layer1_out[5320]);
     layer2_out[3288] <= ~(layer1_out[11636] | layer1_out[11637]);
     layer2_out[3289] <= ~layer1_out[2369];
     layer2_out[3290] <= ~(layer1_out[8466] ^ layer1_out[8467]);
     layer2_out[3291] <= ~layer1_out[10750];
     layer2_out[3292] <= layer1_out[1539] | layer1_out[1540];
     layer2_out[3293] <= ~layer1_out[2461] | layer1_out[2460];
     layer2_out[3294] <= layer1_out[5002];
     layer2_out[3295] <= layer1_out[9295] & ~layer1_out[9294];
     layer2_out[3296] <= ~(layer1_out[5958] | layer1_out[5959]);
     layer2_out[3297] <= layer1_out[6916] & ~layer1_out[6915];
     layer2_out[3298] <= layer1_out[4255];
     layer2_out[3299] <= layer1_out[8898] & ~layer1_out[8899];
     layer2_out[3300] <= ~layer1_out[1937];
     layer2_out[3301] <= ~layer1_out[5766] | layer1_out[5767];
     layer2_out[3302] <= layer1_out[30];
     layer2_out[3303] <= layer1_out[8479] | layer1_out[8480];
     layer2_out[3304] <= ~layer1_out[3762];
     layer2_out[3305] <= layer1_out[7391] & layer1_out[7392];
     layer2_out[3306] <= ~(layer1_out[11105] | layer1_out[11106]);
     layer2_out[3307] <= ~(layer1_out[77] ^ layer1_out[78]);
     layer2_out[3308] <= ~(layer1_out[6786] ^ layer1_out[6787]);
     layer2_out[3309] <= layer1_out[3289] | layer1_out[3290];
     layer2_out[3310] <= ~layer1_out[6037];
     layer2_out[3311] <= layer1_out[8280] & ~layer1_out[8279];
     layer2_out[3312] <= layer1_out[8897];
     layer2_out[3313] <= layer1_out[6247];
     layer2_out[3314] <= ~layer1_out[7085] | layer1_out[7086];
     layer2_out[3315] <= layer1_out[6330] & ~layer1_out[6329];
     layer2_out[3316] <= layer1_out[7387] & ~layer1_out[7386];
     layer2_out[3317] <= ~(layer1_out[1469] | layer1_out[1470]);
     layer2_out[3318] <= layer1_out[598] | layer1_out[599];
     layer2_out[3319] <= layer1_out[9630];
     layer2_out[3320] <= layer1_out[9048] | layer1_out[9049];
     layer2_out[3321] <= ~layer1_out[2463] | layer1_out[2464];
     layer2_out[3322] <= layer1_out[10689] & ~layer1_out[10690];
     layer2_out[3323] <= layer1_out[7074] & layer1_out[7075];
     layer2_out[3324] <= ~layer1_out[4623] | layer1_out[4622];
     layer2_out[3325] <= ~layer1_out[5168];
     layer2_out[3326] <= layer1_out[6361] & layer1_out[6362];
     layer2_out[3327] <= ~layer1_out[11274];
     layer2_out[3328] <= layer1_out[2336] & layer1_out[2337];
     layer2_out[3329] <= ~layer1_out[8178];
     layer2_out[3330] <= ~layer1_out[11088] | layer1_out[11089];
     layer2_out[3331] <= ~(layer1_out[2683] ^ layer1_out[2684]);
     layer2_out[3332] <= ~layer1_out[9409] | layer1_out[9410];
     layer2_out[3333] <= layer1_out[4940] & layer1_out[4941];
     layer2_out[3334] <= layer1_out[4560];
     layer2_out[3335] <= ~layer1_out[5209];
     layer2_out[3336] <= layer1_out[7145] & ~layer1_out[7144];
     layer2_out[3337] <= layer1_out[695] | layer1_out[696];
     layer2_out[3338] <= ~(layer1_out[3272] ^ layer1_out[3273]);
     layer2_out[3339] <= layer1_out[9954] & ~layer1_out[9955];
     layer2_out[3340] <= ~layer1_out[3389];
     layer2_out[3341] <= layer1_out[5751];
     layer2_out[3342] <= ~layer1_out[245];
     layer2_out[3343] <= layer1_out[155];
     layer2_out[3344] <= ~layer1_out[1269];
     layer2_out[3345] <= layer1_out[4032];
     layer2_out[3346] <= ~(layer1_out[6930] & layer1_out[6931]);
     layer2_out[3347] <= ~layer1_out[6941];
     layer2_out[3348] <= ~layer1_out[9787];
     layer2_out[3349] <= ~layer1_out[289] | layer1_out[288];
     layer2_out[3350] <= ~layer1_out[3233];
     layer2_out[3351] <= layer1_out[10093];
     layer2_out[3352] <= ~layer1_out[8796] | layer1_out[8795];
     layer2_out[3353] <= layer1_out[11544];
     layer2_out[3354] <= layer1_out[1405];
     layer2_out[3355] <= layer1_out[3548];
     layer2_out[3356] <= ~layer1_out[231];
     layer2_out[3357] <= layer1_out[8150] ^ layer1_out[8151];
     layer2_out[3358] <= layer1_out[9456];
     layer2_out[3359] <= ~(layer1_out[8437] | layer1_out[8438]);
     layer2_out[3360] <= layer1_out[1118] & layer1_out[1119];
     layer2_out[3361] <= layer1_out[7132] | layer1_out[7133];
     layer2_out[3362] <= ~layer1_out[11773] | layer1_out[11774];
     layer2_out[3363] <= layer1_out[10828];
     layer2_out[3364] <= ~(layer1_out[8526] ^ layer1_out[8527]);
     layer2_out[3365] <= ~layer1_out[5438] | layer1_out[5437];
     layer2_out[3366] <= layer1_out[7115];
     layer2_out[3367] <= layer1_out[6490] & layer1_out[6491];
     layer2_out[3368] <= ~layer1_out[5016] | layer1_out[5017];
     layer2_out[3369] <= ~layer1_out[6263] | layer1_out[6264];
     layer2_out[3370] <= ~layer1_out[6197] | layer1_out[6198];
     layer2_out[3371] <= ~layer1_out[6267];
     layer2_out[3372] <= ~layer1_out[4155];
     layer2_out[3373] <= ~layer1_out[607];
     layer2_out[3374] <= ~layer1_out[8216];
     layer2_out[3375] <= layer1_out[6264] & ~layer1_out[6265];
     layer2_out[3376] <= layer1_out[10655] & ~layer1_out[10656];
     layer2_out[3377] <= ~layer1_out[11323] | layer1_out[11322];
     layer2_out[3378] <= ~layer1_out[8163] | layer1_out[8162];
     layer2_out[3379] <= ~layer1_out[11164] | layer1_out[11163];
     layer2_out[3380] <= layer1_out[8738];
     layer2_out[3381] <= ~layer1_out[2902];
     layer2_out[3382] <= layer1_out[5987];
     layer2_out[3383] <= layer1_out[5278] | layer1_out[5279];
     layer2_out[3384] <= layer1_out[2861];
     layer2_out[3385] <= ~(layer1_out[7194] ^ layer1_out[7195]);
     layer2_out[3386] <= ~(layer1_out[2587] & layer1_out[2588]);
     layer2_out[3387] <= ~layer1_out[5706];
     layer2_out[3388] <= ~layer1_out[11253];
     layer2_out[3389] <= layer1_out[8680] & ~layer1_out[8681];
     layer2_out[3390] <= ~layer1_out[1408] | layer1_out[1407];
     layer2_out[3391] <= layer1_out[2345] & ~layer1_out[2346];
     layer2_out[3392] <= ~layer1_out[10352] | layer1_out[10353];
     layer2_out[3393] <= layer1_out[751] & ~layer1_out[750];
     layer2_out[3394] <= layer1_out[9212];
     layer2_out[3395] <= ~layer1_out[4140];
     layer2_out[3396] <= layer1_out[5364];
     layer2_out[3397] <= ~layer1_out[9164];
     layer2_out[3398] <= layer1_out[6067];
     layer2_out[3399] <= ~layer1_out[565];
     layer2_out[3400] <= ~layer1_out[1939] | layer1_out[1940];
     layer2_out[3401] <= ~layer1_out[11272];
     layer2_out[3402] <= layer1_out[3188] | layer1_out[3189];
     layer2_out[3403] <= layer1_out[10169];
     layer2_out[3404] <= ~layer1_out[738] | layer1_out[737];
     layer2_out[3405] <= layer1_out[4306];
     layer2_out[3406] <= layer1_out[9318] | layer1_out[9319];
     layer2_out[3407] <= layer1_out[4250] & ~layer1_out[4249];
     layer2_out[3408] <= ~(layer1_out[5966] ^ layer1_out[5967]);
     layer2_out[3409] <= ~layer1_out[6087] | layer1_out[6088];
     layer2_out[3410] <= ~layer1_out[10348];
     layer2_out[3411] <= ~(layer1_out[8765] | layer1_out[8766]);
     layer2_out[3412] <= ~layer1_out[5112];
     layer2_out[3413] <= ~layer1_out[5801] | layer1_out[5802];
     layer2_out[3414] <= ~layer1_out[5183];
     layer2_out[3415] <= ~layer1_out[10381];
     layer2_out[3416] <= layer1_out[3473] & layer1_out[3474];
     layer2_out[3417] <= layer1_out[8791] & ~layer1_out[8792];
     layer2_out[3418] <= layer1_out[11211] ^ layer1_out[11212];
     layer2_out[3419] <= ~layer1_out[5938];
     layer2_out[3420] <= ~layer1_out[9015] | layer1_out[9016];
     layer2_out[3421] <= ~layer1_out[6357];
     layer2_out[3422] <= layer1_out[8322];
     layer2_out[3423] <= layer1_out[9412];
     layer2_out[3424] <= ~(layer1_out[1321] | layer1_out[1322]);
     layer2_out[3425] <= ~layer1_out[11390];
     layer2_out[3426] <= ~layer1_out[305] | layer1_out[306];
     layer2_out[3427] <= 1'b1;
     layer2_out[3428] <= ~layer1_out[3392];
     layer2_out[3429] <= ~layer1_out[7164];
     layer2_out[3430] <= ~(layer1_out[2258] & layer1_out[2259]);
     layer2_out[3431] <= layer1_out[1312] & ~layer1_out[1311];
     layer2_out[3432] <= ~layer1_out[9628] | layer1_out[9629];
     layer2_out[3433] <= ~layer1_out[8156];
     layer2_out[3434] <= ~(layer1_out[8187] ^ layer1_out[8188]);
     layer2_out[3435] <= layer1_out[7098] ^ layer1_out[7099];
     layer2_out[3436] <= ~layer1_out[4299];
     layer2_out[3437] <= ~layer1_out[9045];
     layer2_out[3438] <= layer1_out[2736] & layer1_out[2737];
     layer2_out[3439] <= ~(layer1_out[1727] | layer1_out[1728]);
     layer2_out[3440] <= ~layer1_out[11961] | layer1_out[11962];
     layer2_out[3441] <= ~layer1_out[11092] | layer1_out[11091];
     layer2_out[3442] <= ~layer1_out[7280] | layer1_out[7281];
     layer2_out[3443] <= ~layer1_out[6684];
     layer2_out[3444] <= layer1_out[7485];
     layer2_out[3445] <= 1'b0;
     layer2_out[3446] <= ~layer1_out[9145];
     layer2_out[3447] <= ~layer1_out[8028] | layer1_out[8029];
     layer2_out[3448] <= ~(layer1_out[11264] | layer1_out[11265]);
     layer2_out[3449] <= layer1_out[2276];
     layer2_out[3450] <= layer1_out[261] & ~layer1_out[262];
     layer2_out[3451] <= ~layer1_out[9947];
     layer2_out[3452] <= layer1_out[5944] & ~layer1_out[5943];
     layer2_out[3453] <= layer1_out[9116] ^ layer1_out[9117];
     layer2_out[3454] <= layer1_out[5102] & ~layer1_out[5101];
     layer2_out[3455] <= layer1_out[7344] & ~layer1_out[7343];
     layer2_out[3456] <= layer1_out[8511];
     layer2_out[3457] <= layer1_out[4652] & layer1_out[4653];
     layer2_out[3458] <= ~(layer1_out[3007] ^ layer1_out[3008]);
     layer2_out[3459] <= layer1_out[3194] ^ layer1_out[3195];
     layer2_out[3460] <= layer1_out[9072];
     layer2_out[3461] <= layer1_out[976];
     layer2_out[3462] <= layer1_out[2200] & ~layer1_out[2201];
     layer2_out[3463] <= ~(layer1_out[7175] ^ layer1_out[7176]);
     layer2_out[3464] <= layer1_out[8970];
     layer2_out[3465] <= layer1_out[5154];
     layer2_out[3466] <= layer1_out[1386] & ~layer1_out[1387];
     layer2_out[3467] <= ~layer1_out[11954] | layer1_out[11953];
     layer2_out[3468] <= ~layer1_out[10385];
     layer2_out[3469] <= layer1_out[9806] & ~layer1_out[9805];
     layer2_out[3470] <= layer1_out[10999];
     layer2_out[3471] <= layer1_out[6834] & ~layer1_out[6835];
     layer2_out[3472] <= ~(layer1_out[5668] | layer1_out[5669]);
     layer2_out[3473] <= ~(layer1_out[9718] & layer1_out[9719]);
     layer2_out[3474] <= layer1_out[11871];
     layer2_out[3475] <= layer1_out[2603] & ~layer1_out[2602];
     layer2_out[3476] <= layer1_out[367];
     layer2_out[3477] <= ~layer1_out[2353] | layer1_out[2354];
     layer2_out[3478] <= layer1_out[7425] | layer1_out[7426];
     layer2_out[3479] <= ~(layer1_out[8970] & layer1_out[8971]);
     layer2_out[3480] <= ~layer1_out[8892];
     layer2_out[3481] <= ~layer1_out[8390];
     layer2_out[3482] <= ~(layer1_out[6427] | layer1_out[6428]);
     layer2_out[3483] <= layer1_out[2401] & layer1_out[2402];
     layer2_out[3484] <= ~layer1_out[10640];
     layer2_out[3485] <= ~layer1_out[7974] | layer1_out[7975];
     layer2_out[3486] <= ~layer1_out[1068];
     layer2_out[3487] <= ~layer1_out[2501] | layer1_out[2502];
     layer2_out[3488] <= layer1_out[4052] & ~layer1_out[4053];
     layer2_out[3489] <= ~layer1_out[188];
     layer2_out[3490] <= ~layer1_out[7374];
     layer2_out[3491] <= layer1_out[951];
     layer2_out[3492] <= layer1_out[2522] | layer1_out[2523];
     layer2_out[3493] <= ~layer1_out[7679];
     layer2_out[3494] <= layer1_out[10880] | layer1_out[10881];
     layer2_out[3495] <= ~(layer1_out[11535] ^ layer1_out[11536]);
     layer2_out[3496] <= layer1_out[11630] & ~layer1_out[11631];
     layer2_out[3497] <= ~layer1_out[5035] | layer1_out[5034];
     layer2_out[3498] <= layer1_out[10565] & layer1_out[10566];
     layer2_out[3499] <= ~layer1_out[9138];
     layer2_out[3500] <= layer1_out[11926] & ~layer1_out[11927];
     layer2_out[3501] <= layer1_out[1360] & ~layer1_out[1361];
     layer2_out[3502] <= ~(layer1_out[7197] | layer1_out[7198]);
     layer2_out[3503] <= layer1_out[11485];
     layer2_out[3504] <= layer1_out[6844] ^ layer1_out[6845];
     layer2_out[3505] <= layer1_out[8376];
     layer2_out[3506] <= ~layer1_out[6788] | layer1_out[6789];
     layer2_out[3507] <= layer1_out[253] | layer1_out[254];
     layer2_out[3508] <= ~layer1_out[10715] | layer1_out[10716];
     layer2_out[3509] <= layer1_out[850] & ~layer1_out[851];
     layer2_out[3510] <= ~layer1_out[2701];
     layer2_out[3511] <= ~layer1_out[144];
     layer2_out[3512] <= ~(layer1_out[1610] & layer1_out[1611]);
     layer2_out[3513] <= layer1_out[7935] & layer1_out[7936];
     layer2_out[3514] <= ~layer1_out[1687];
     layer2_out[3515] <= layer1_out[2752];
     layer2_out[3516] <= ~layer1_out[1792];
     layer2_out[3517] <= layer1_out[8919] & ~layer1_out[8918];
     layer2_out[3518] <= layer1_out[8032];
     layer2_out[3519] <= layer1_out[3863] | layer1_out[3864];
     layer2_out[3520] <= layer1_out[9344] & ~layer1_out[9345];
     layer2_out[3521] <= ~layer1_out[1337];
     layer2_out[3522] <= ~layer1_out[744] | layer1_out[743];
     layer2_out[3523] <= layer1_out[2895];
     layer2_out[3524] <= layer1_out[11199] & ~layer1_out[11200];
     layer2_out[3525] <= ~(layer1_out[6060] | layer1_out[6061]);
     layer2_out[3526] <= ~layer1_out[1854] | layer1_out[1855];
     layer2_out[3527] <= layer1_out[72];
     layer2_out[3528] <= ~(layer1_out[10048] | layer1_out[10049]);
     layer2_out[3529] <= ~layer1_out[4585] | layer1_out[4586];
     layer2_out[3530] <= ~layer1_out[361];
     layer2_out[3531] <= ~(layer1_out[6063] ^ layer1_out[6064]);
     layer2_out[3532] <= ~layer1_out[3454];
     layer2_out[3533] <= ~layer1_out[8930] | layer1_out[8931];
     layer2_out[3534] <= layer1_out[7091] | layer1_out[7092];
     layer2_out[3535] <= layer1_out[9678];
     layer2_out[3536] <= layer1_out[4131] & ~layer1_out[4130];
     layer2_out[3537] <= layer1_out[11487];
     layer2_out[3538] <= ~layer1_out[8917];
     layer2_out[3539] <= layer1_out[20] & ~layer1_out[21];
     layer2_out[3540] <= layer1_out[1287] & ~layer1_out[1286];
     layer2_out[3541] <= ~layer1_out[2833] | layer1_out[2834];
     layer2_out[3542] <= ~layer1_out[2614];
     layer2_out[3543] <= ~layer1_out[3130];
     layer2_out[3544] <= ~layer1_out[10256];
     layer2_out[3545] <= layer1_out[10223];
     layer2_out[3546] <= layer1_out[11433] & ~layer1_out[11434];
     layer2_out[3547] <= ~layer1_out[10320];
     layer2_out[3548] <= ~layer1_out[5064];
     layer2_out[3549] <= layer1_out[11795] | layer1_out[11796];
     layer2_out[3550] <= ~layer1_out[11783];
     layer2_out[3551] <= layer1_out[11801] | layer1_out[11802];
     layer2_out[3552] <= layer1_out[3798] & ~layer1_out[3799];
     layer2_out[3553] <= ~layer1_out[8963];
     layer2_out[3554] <= ~(layer1_out[1748] ^ layer1_out[1749]);
     layer2_out[3555] <= ~(layer1_out[9532] & layer1_out[9533]);
     layer2_out[3556] <= 1'b1;
     layer2_out[3557] <= ~layer1_out[11788] | layer1_out[11789];
     layer2_out[3558] <= ~layer1_out[7900];
     layer2_out[3559] <= ~layer1_out[10464];
     layer2_out[3560] <= ~(layer1_out[11877] ^ layer1_out[11878]);
     layer2_out[3561] <= ~layer1_out[6174];
     layer2_out[3562] <= ~(layer1_out[247] & layer1_out[248]);
     layer2_out[3563] <= ~layer1_out[10001];
     layer2_out[3564] <= layer1_out[2594] | layer1_out[2595];
     layer2_out[3565] <= ~layer1_out[3350];
     layer2_out[3566] <= layer1_out[10991] | layer1_out[10992];
     layer2_out[3567] <= layer1_out[7985] | layer1_out[7986];
     layer2_out[3568] <= layer1_out[10107] & ~layer1_out[10108];
     layer2_out[3569] <= ~layer1_out[2470] | layer1_out[2469];
     layer2_out[3570] <= ~layer1_out[3459] | layer1_out[3458];
     layer2_out[3571] <= layer1_out[497];
     layer2_out[3572] <= layer1_out[1019] & ~layer1_out[1020];
     layer2_out[3573] <= layer1_out[2055];
     layer2_out[3574] <= layer1_out[10897];
     layer2_out[3575] <= ~layer1_out[9204];
     layer2_out[3576] <= ~layer1_out[449];
     layer2_out[3577] <= ~layer1_out[2759] | layer1_out[2760];
     layer2_out[3578] <= ~(layer1_out[8485] | layer1_out[8486]);
     layer2_out[3579] <= layer1_out[8118] & ~layer1_out[8117];
     layer2_out[3580] <= ~(layer1_out[5491] ^ layer1_out[5492]);
     layer2_out[3581] <= ~layer1_out[2836] | layer1_out[2835];
     layer2_out[3582] <= layer1_out[1204] | layer1_out[1205];
     layer2_out[3583] <= layer1_out[5752];
     layer2_out[3584] <= layer1_out[6492];
     layer2_out[3585] <= layer1_out[2965] & ~layer1_out[2964];
     layer2_out[3586] <= ~layer1_out[10060];
     layer2_out[3587] <= ~layer1_out[11525] | layer1_out[11524];
     layer2_out[3588] <= layer1_out[871] & ~layer1_out[870];
     layer2_out[3589] <= 1'b0;
     layer2_out[3590] <= ~layer1_out[11920];
     layer2_out[3591] <= ~(layer1_out[5898] ^ layer1_out[5899]);
     layer2_out[3592] <= layer1_out[5336];
     layer2_out[3593] <= layer1_out[11642] & ~layer1_out[11643];
     layer2_out[3594] <= ~(layer1_out[5373] | layer1_out[5374]);
     layer2_out[3595] <= ~(layer1_out[4659] ^ layer1_out[4660]);
     layer2_out[3596] <= layer1_out[2674] & layer1_out[2675];
     layer2_out[3597] <= layer1_out[10602];
     layer2_out[3598] <= layer1_out[2809];
     layer2_out[3599] <= layer1_out[3202] | layer1_out[3203];
     layer2_out[3600] <= ~layer1_out[6410];
     layer2_out[3601] <= ~layer1_out[6629] | layer1_out[6628];
     layer2_out[3602] <= layer1_out[7601] | layer1_out[7602];
     layer2_out[3603] <= layer1_out[257];
     layer2_out[3604] <= layer1_out[5337] ^ layer1_out[5338];
     layer2_out[3605] <= ~layer1_out[8365];
     layer2_out[3606] <= ~(layer1_out[2070] ^ layer1_out[2071]);
     layer2_out[3607] <= ~layer1_out[9047];
     layer2_out[3608] <= ~layer1_out[7059];
     layer2_out[3609] <= ~(layer1_out[3831] | layer1_out[3832]);
     layer2_out[3610] <= layer1_out[2051];
     layer2_out[3611] <= layer1_out[10941];
     layer2_out[3612] <= ~layer1_out[10027];
     layer2_out[3613] <= ~(layer1_out[5813] ^ layer1_out[5814]);
     layer2_out[3614] <= layer1_out[11568] & layer1_out[11569];
     layer2_out[3615] <= layer1_out[778] & ~layer1_out[779];
     layer2_out[3616] <= ~(layer1_out[5332] & layer1_out[5333]);
     layer2_out[3617] <= ~(layer1_out[8726] | layer1_out[8727]);
     layer2_out[3618] <= layer1_out[11895];
     layer2_out[3619] <= ~layer1_out[1629];
     layer2_out[3620] <= ~(layer1_out[2049] | layer1_out[2050]);
     layer2_out[3621] <= ~(layer1_out[1075] & layer1_out[1076]);
     layer2_out[3622] <= ~(layer1_out[1732] & layer1_out[1733]);
     layer2_out[3623] <= ~(layer1_out[8253] & layer1_out[8254]);
     layer2_out[3624] <= layer1_out[3064] & layer1_out[3065];
     layer2_out[3625] <= ~layer1_out[3723] | layer1_out[3724];
     layer2_out[3626] <= layer1_out[6869] & layer1_out[6870];
     layer2_out[3627] <= layer1_out[3633] & layer1_out[3634];
     layer2_out[3628] <= ~layer1_out[2219] | layer1_out[2218];
     layer2_out[3629] <= ~layer1_out[3473];
     layer2_out[3630] <= ~layer1_out[3761] | layer1_out[3760];
     layer2_out[3631] <= layer1_out[5949];
     layer2_out[3632] <= layer1_out[4946];
     layer2_out[3633] <= layer1_out[11017] & ~layer1_out[11016];
     layer2_out[3634] <= layer1_out[7024] & ~layer1_out[7023];
     layer2_out[3635] <= layer1_out[3972];
     layer2_out[3636] <= layer1_out[5022];
     layer2_out[3637] <= ~layer1_out[7575];
     layer2_out[3638] <= layer1_out[2156] | layer1_out[2157];
     layer2_out[3639] <= layer1_out[11329] & ~layer1_out[11328];
     layer2_out[3640] <= layer1_out[2297] & layer1_out[2298];
     layer2_out[3641] <= ~layer1_out[6848];
     layer2_out[3642] <= layer1_out[8131] & ~layer1_out[8132];
     layer2_out[3643] <= ~layer1_out[8350];
     layer2_out[3644] <= layer1_out[3081];
     layer2_out[3645] <= layer1_out[7142];
     layer2_out[3646] <= ~layer1_out[3070];
     layer2_out[3647] <= layer1_out[6745];
     layer2_out[3648] <= layer1_out[4765];
     layer2_out[3649] <= ~(layer1_out[11842] ^ layer1_out[11843]);
     layer2_out[3650] <= ~layer1_out[770];
     layer2_out[3651] <= ~(layer1_out[1702] | layer1_out[1703]);
     layer2_out[3652] <= layer1_out[9648];
     layer2_out[3653] <= ~(layer1_out[1836] | layer1_out[1837]);
     layer2_out[3654] <= ~layer1_out[10318];
     layer2_out[3655] <= layer1_out[1221] & layer1_out[1222];
     layer2_out[3656] <= ~layer1_out[4163];
     layer2_out[3657] <= ~layer1_out[4296] | layer1_out[4297];
     layer2_out[3658] <= layer1_out[8648] & ~layer1_out[8649];
     layer2_out[3659] <= ~layer1_out[1133] | layer1_out[1134];
     layer2_out[3660] <= 1'b1;
     layer2_out[3661] <= ~(layer1_out[3393] & layer1_out[3394]);
     layer2_out[3662] <= ~layer1_out[9038];
     layer2_out[3663] <= ~(layer1_out[545] & layer1_out[546]);
     layer2_out[3664] <= layer1_out[7045] & ~layer1_out[7046];
     layer2_out[3665] <= ~layer1_out[6731];
     layer2_out[3666] <= layer1_out[3035];
     layer2_out[3667] <= ~layer1_out[3081];
     layer2_out[3668] <= layer1_out[5442];
     layer2_out[3669] <= layer1_out[5215] & layer1_out[5216];
     layer2_out[3670] <= layer1_out[1168] & ~layer1_out[1169];
     layer2_out[3671] <= ~layer1_out[2563];
     layer2_out[3672] <= ~(layer1_out[11980] ^ layer1_out[11981]);
     layer2_out[3673] <= ~layer1_out[11841];
     layer2_out[3674] <= ~layer1_out[8917] | layer1_out[8918];
     layer2_out[3675] <= ~(layer1_out[11173] & layer1_out[11174]);
     layer2_out[3676] <= layer1_out[1106] | layer1_out[1107];
     layer2_out[3677] <= ~(layer1_out[11051] & layer1_out[11052]);
     layer2_out[3678] <= ~layer1_out[5488] | layer1_out[5489];
     layer2_out[3679] <= layer1_out[1425] & ~layer1_out[1424];
     layer2_out[3680] <= 1'b0;
     layer2_out[3681] <= layer1_out[4097] & layer1_out[4098];
     layer2_out[3682] <= layer1_out[4496] | layer1_out[4497];
     layer2_out[3683] <= ~layer1_out[2899] | layer1_out[2898];
     layer2_out[3684] <= layer1_out[9238];
     layer2_out[3685] <= layer1_out[4807];
     layer2_out[3686] <= ~(layer1_out[7583] & layer1_out[7584]);
     layer2_out[3687] <= ~layer1_out[3236] | layer1_out[3235];
     layer2_out[3688] <= ~(layer1_out[3061] ^ layer1_out[3062]);
     layer2_out[3689] <= layer1_out[9728] & ~layer1_out[9727];
     layer2_out[3690] <= ~layer1_out[11140];
     layer2_out[3691] <= layer1_out[6262];
     layer2_out[3692] <= ~layer1_out[2583] | layer1_out[2582];
     layer2_out[3693] <= ~layer1_out[1365];
     layer2_out[3694] <= ~layer1_out[4458] | layer1_out[4457];
     layer2_out[3695] <= layer1_out[5341] | layer1_out[5342];
     layer2_out[3696] <= layer1_out[4720];
     layer2_out[3697] <= layer1_out[11967] & layer1_out[11968];
     layer2_out[3698] <= ~layer1_out[10569];
     layer2_out[3699] <= layer1_out[10294];
     layer2_out[3700] <= layer1_out[7014];
     layer2_out[3701] <= ~(layer1_out[8702] | layer1_out[8703]);
     layer2_out[3702] <= layer1_out[6853] | layer1_out[6854];
     layer2_out[3703] <= ~(layer1_out[4289] & layer1_out[4290]);
     layer2_out[3704] <= layer1_out[6390] & ~layer1_out[6389];
     layer2_out[3705] <= layer1_out[6861] ^ layer1_out[6862];
     layer2_out[3706] <= ~layer1_out[992] | layer1_out[993];
     layer2_out[3707] <= layer1_out[8125];
     layer2_out[3708] <= ~(layer1_out[10700] ^ layer1_out[10701]);
     layer2_out[3709] <= 1'b0;
     layer2_out[3710] <= ~layer1_out[9614] | layer1_out[9613];
     layer2_out[3711] <= 1'b0;
     layer2_out[3712] <= ~layer1_out[2933] | layer1_out[2934];
     layer2_out[3713] <= layer1_out[844] & layer1_out[845];
     layer2_out[3714] <= layer1_out[5020];
     layer2_out[3715] <= layer1_out[11242] & layer1_out[11243];
     layer2_out[3716] <= ~(layer1_out[4566] & layer1_out[4567]);
     layer2_out[3717] <= layer1_out[8208] & layer1_out[8209];
     layer2_out[3718] <= ~layer1_out[3368];
     layer2_out[3719] <= layer1_out[11367];
     layer2_out[3720] <= layer1_out[6075] & ~layer1_out[6076];
     layer2_out[3721] <= 1'b1;
     layer2_out[3722] <= layer1_out[5030] & ~layer1_out[5031];
     layer2_out[3723] <= layer1_out[517];
     layer2_out[3724] <= ~(layer1_out[11415] ^ layer1_out[11416]);
     layer2_out[3725] <= ~layer1_out[3845];
     layer2_out[3726] <= layer1_out[2245] & ~layer1_out[2244];
     layer2_out[3727] <= layer1_out[9046] & ~layer1_out[9045];
     layer2_out[3728] <= layer1_out[6438] & ~layer1_out[6437];
     layer2_out[3729] <= layer1_out[1248] | layer1_out[1249];
     layer2_out[3730] <= layer1_out[8985] | layer1_out[8986];
     layer2_out[3731] <= ~layer1_out[6708] | layer1_out[6709];
     layer2_out[3732] <= layer1_out[8616] & layer1_out[8617];
     layer2_out[3733] <= layer1_out[4825];
     layer2_out[3734] <= ~layer1_out[6482] | layer1_out[6483];
     layer2_out[3735] <= layer1_out[95] & ~layer1_out[94];
     layer2_out[3736] <= ~layer1_out[5570];
     layer2_out[3737] <= layer1_out[7506];
     layer2_out[3738] <= ~(layer1_out[183] & layer1_out[184]);
     layer2_out[3739] <= ~(layer1_out[9623] | layer1_out[9624]);
     layer2_out[3740] <= layer1_out[1999] & layer1_out[2000];
     layer2_out[3741] <= layer1_out[9109] ^ layer1_out[9110];
     layer2_out[3742] <= layer1_out[1964] & layer1_out[1965];
     layer2_out[3743] <= ~layer1_out[2310];
     layer2_out[3744] <= layer1_out[1834] & ~layer1_out[1833];
     layer2_out[3745] <= layer1_out[11865];
     layer2_out[3746] <= ~layer1_out[5569] | layer1_out[5568];
     layer2_out[3747] <= layer1_out[2063] | layer1_out[2064];
     layer2_out[3748] <= layer1_out[2933];
     layer2_out[3749] <= ~layer1_out[9397];
     layer2_out[3750] <= layer1_out[414];
     layer2_out[3751] <= layer1_out[1837];
     layer2_out[3752] <= ~layer1_out[10555];
     layer2_out[3753] <= layer1_out[7675];
     layer2_out[3754] <= layer1_out[1562] | layer1_out[1563];
     layer2_out[3755] <= layer1_out[10709];
     layer2_out[3756] <= ~layer1_out[10381];
     layer2_out[3757] <= ~layer1_out[3256];
     layer2_out[3758] <= ~(layer1_out[11742] & layer1_out[11743]);
     layer2_out[3759] <= layer1_out[4057] & ~layer1_out[4058];
     layer2_out[3760] <= layer1_out[416];
     layer2_out[3761] <= ~(layer1_out[4623] | layer1_out[4624]);
     layer2_out[3762] <= ~layer1_out[2654];
     layer2_out[3763] <= layer1_out[5534] & ~layer1_out[5535];
     layer2_out[3764] <= ~layer1_out[8712];
     layer2_out[3765] <= layer1_out[6612];
     layer2_out[3766] <= layer1_out[8063] & layer1_out[8064];
     layer2_out[3767] <= ~layer1_out[8652] | layer1_out[8653];
     layer2_out[3768] <= ~layer1_out[10200];
     layer2_out[3769] <= layer1_out[5617];
     layer2_out[3770] <= layer1_out[9134] & ~layer1_out[9133];
     layer2_out[3771] <= 1'b1;
     layer2_out[3772] <= layer1_out[10463] & ~layer1_out[10462];
     layer2_out[3773] <= ~layer1_out[10782] | layer1_out[10783];
     layer2_out[3774] <= ~layer1_out[8776];
     layer2_out[3775] <= ~layer1_out[11504];
     layer2_out[3776] <= ~layer1_out[4089] | layer1_out[4088];
     layer2_out[3777] <= layer1_out[2852];
     layer2_out[3778] <= layer1_out[7689] & ~layer1_out[7690];
     layer2_out[3779] <= ~layer1_out[5781];
     layer2_out[3780] <= ~layer1_out[7665] | layer1_out[7664];
     layer2_out[3781] <= layer1_out[1392] ^ layer1_out[1393];
     layer2_out[3782] <= ~layer1_out[11259];
     layer2_out[3783] <= layer1_out[2251] ^ layer1_out[2252];
     layer2_out[3784] <= layer1_out[8427] & ~layer1_out[8426];
     layer2_out[3785] <= layer1_out[2673];
     layer2_out[3786] <= ~layer1_out[9431];
     layer2_out[3787] <= layer1_out[1196] ^ layer1_out[1197];
     layer2_out[3788] <= layer1_out[8541] | layer1_out[8542];
     layer2_out[3789] <= layer1_out[2081];
     layer2_out[3790] <= layer1_out[2568] & ~layer1_out[2569];
     layer2_out[3791] <= ~layer1_out[11298] | layer1_out[11297];
     layer2_out[3792] <= layer1_out[4854] & layer1_out[4855];
     layer2_out[3793] <= layer1_out[9009] & ~layer1_out[9008];
     layer2_out[3794] <= ~layer1_out[4170];
     layer2_out[3795] <= ~layer1_out[3744] | layer1_out[3745];
     layer2_out[3796] <= layer1_out[285] | layer1_out[286];
     layer2_out[3797] <= ~layer1_out[8989];
     layer2_out[3798] <= ~layer1_out[2272] | layer1_out[2271];
     layer2_out[3799] <= ~layer1_out[2150] | layer1_out[2151];
     layer2_out[3800] <= ~layer1_out[9051] | layer1_out[9052];
     layer2_out[3801] <= layer1_out[5403] | layer1_out[5404];
     layer2_out[3802] <= ~layer1_out[7260];
     layer2_out[3803] <= layer1_out[684];
     layer2_out[3804] <= layer1_out[2549];
     layer2_out[3805] <= ~layer1_out[2265] | layer1_out[2264];
     layer2_out[3806] <= ~(layer1_out[11114] ^ layer1_out[11115]);
     layer2_out[3807] <= layer1_out[3010] & ~layer1_out[3009];
     layer2_out[3808] <= ~layer1_out[3280];
     layer2_out[3809] <= ~layer1_out[2159];
     layer2_out[3810] <= layer1_out[408] ^ layer1_out[409];
     layer2_out[3811] <= layer1_out[11214];
     layer2_out[3812] <= layer1_out[10066];
     layer2_out[3813] <= layer1_out[9411];
     layer2_out[3814] <= layer1_out[4744];
     layer2_out[3815] <= ~layer1_out[11040];
     layer2_out[3816] <= layer1_out[2671];
     layer2_out[3817] <= ~layer1_out[9928] | layer1_out[9929];
     layer2_out[3818] <= ~(layer1_out[5930] ^ layer1_out[5931]);
     layer2_out[3819] <= ~(layer1_out[5376] | layer1_out[5377]);
     layer2_out[3820] <= layer1_out[5393];
     layer2_out[3821] <= ~(layer1_out[491] & layer1_out[492]);
     layer2_out[3822] <= ~layer1_out[11454] | layer1_out[11455];
     layer2_out[3823] <= layer1_out[11101] | layer1_out[11102];
     layer2_out[3824] <= layer1_out[1397] | layer1_out[1398];
     layer2_out[3825] <= layer1_out[1338] ^ layer1_out[1339];
     layer2_out[3826] <= layer1_out[9640] ^ layer1_out[9641];
     layer2_out[3827] <= ~(layer1_out[10530] & layer1_out[10531]);
     layer2_out[3828] <= ~(layer1_out[11916] & layer1_out[11917]);
     layer2_out[3829] <= layer1_out[7229];
     layer2_out[3830] <= layer1_out[2804] ^ layer1_out[2805];
     layer2_out[3831] <= layer1_out[8213] | layer1_out[8214];
     layer2_out[3832] <= ~layer1_out[11034];
     layer2_out[3833] <= 1'b1;
     layer2_out[3834] <= layer1_out[9267] & layer1_out[9268];
     layer2_out[3835] <= layer1_out[7413];
     layer2_out[3836] <= ~layer1_out[1131] | layer1_out[1132];
     layer2_out[3837] <= ~(layer1_out[8790] & layer1_out[8791]);
     layer2_out[3838] <= ~(layer1_out[11826] ^ layer1_out[11827]);
     layer2_out[3839] <= ~(layer1_out[10545] & layer1_out[10546]);
     layer2_out[3840] <= ~(layer1_out[8194] | layer1_out[8195]);
     layer2_out[3841] <= layer1_out[2463];
     layer2_out[3842] <= layer1_out[8614];
     layer2_out[3843] <= ~(layer1_out[1374] | layer1_out[1375]);
     layer2_out[3844] <= layer1_out[8548] | layer1_out[8549];
     layer2_out[3845] <= layer1_out[11017] & layer1_out[11018];
     layer2_out[3846] <= layer1_out[5155];
     layer2_out[3847] <= ~layer1_out[4028];
     layer2_out[3848] <= layer1_out[8845];
     layer2_out[3849] <= ~layer1_out[35];
     layer2_out[3850] <= ~layer1_out[7168];
     layer2_out[3851] <= ~(layer1_out[9533] & layer1_out[9534]);
     layer2_out[3852] <= ~layer1_out[3275] | layer1_out[3274];
     layer2_out[3853] <= ~layer1_out[3929] | layer1_out[3930];
     layer2_out[3854] <= ~layer1_out[6965] | layer1_out[6964];
     layer2_out[3855] <= ~(layer1_out[3938] ^ layer1_out[3939]);
     layer2_out[3856] <= ~layer1_out[7946];
     layer2_out[3857] <= ~layer1_out[7193] | layer1_out[7192];
     layer2_out[3858] <= ~layer1_out[1713];
     layer2_out[3859] <= ~layer1_out[276];
     layer2_out[3860] <= ~layer1_out[7987];
     layer2_out[3861] <= layer1_out[9069];
     layer2_out[3862] <= ~layer1_out[10046];
     layer2_out[3863] <= ~layer1_out[10041];
     layer2_out[3864] <= ~layer1_out[3908];
     layer2_out[3865] <= layer1_out[6606];
     layer2_out[3866] <= layer1_out[927] & ~layer1_out[928];
     layer2_out[3867] <= layer1_out[4869];
     layer2_out[3868] <= layer1_out[9431];
     layer2_out[3869] <= layer1_out[9740];
     layer2_out[3870] <= layer1_out[863];
     layer2_out[3871] <= layer1_out[2912] ^ layer1_out[2913];
     layer2_out[3872] <= ~layer1_out[1097];
     layer2_out[3873] <= layer1_out[7759] & ~layer1_out[7758];
     layer2_out[3874] <= layer1_out[9903];
     layer2_out[3875] <= layer1_out[10488] & ~layer1_out[10487];
     layer2_out[3876] <= layer1_out[5899];
     layer2_out[3877] <= layer1_out[2455] & layer1_out[2456];
     layer2_out[3878] <= layer1_out[1736] & layer1_out[1737];
     layer2_out[3879] <= layer1_out[2545] & ~layer1_out[2546];
     layer2_out[3880] <= ~(layer1_out[8729] | layer1_out[8730]);
     layer2_out[3881] <= ~(layer1_out[7710] | layer1_out[7711]);
     layer2_out[3882] <= ~layer1_out[7770];
     layer2_out[3883] <= layer1_out[2076] | layer1_out[2077];
     layer2_out[3884] <= layer1_out[5390];
     layer2_out[3885] <= ~(layer1_out[7262] & layer1_out[7263]);
     layer2_out[3886] <= ~(layer1_out[6431] | layer1_out[6432]);
     layer2_out[3887] <= ~layer1_out[3471] | layer1_out[3472];
     layer2_out[3888] <= ~(layer1_out[11638] | layer1_out[11639]);
     layer2_out[3889] <= layer1_out[785];
     layer2_out[3890] <= ~layer1_out[3759] | layer1_out[3760];
     layer2_out[3891] <= layer1_out[7309] & ~layer1_out[7310];
     layer2_out[3892] <= layer1_out[6045];
     layer2_out[3893] <= ~layer1_out[11816];
     layer2_out[3894] <= ~(layer1_out[4022] & layer1_out[4023]);
     layer2_out[3895] <= ~layer1_out[4704];
     layer2_out[3896] <= 1'b0;
     layer2_out[3897] <= layer1_out[5441] & layer1_out[5442];
     layer2_out[3898] <= ~layer1_out[11113];
     layer2_out[3899] <= layer1_out[329] & layer1_out[330];
     layer2_out[3900] <= layer1_out[5600];
     layer2_out[3901] <= ~layer1_out[3417];
     layer2_out[3902] <= layer1_out[1268] | layer1_out[1269];
     layer2_out[3903] <= layer1_out[1493] & ~layer1_out[1494];
     layer2_out[3904] <= layer1_out[6172];
     layer2_out[3905] <= ~layer1_out[9956];
     layer2_out[3906] <= ~(layer1_out[9312] & layer1_out[9313]);
     layer2_out[3907] <= ~layer1_out[9603] | layer1_out[9604];
     layer2_out[3908] <= layer1_out[3248];
     layer2_out[3909] <= ~layer1_out[10568] | layer1_out[10567];
     layer2_out[3910] <= layer1_out[11375] | layer1_out[11376];
     layer2_out[3911] <= layer1_out[8750];
     layer2_out[3912] <= ~layer1_out[4789];
     layer2_out[3913] <= ~layer1_out[8730] | layer1_out[8731];
     layer2_out[3914] <= layer1_out[8520];
     layer2_out[3915] <= ~layer1_out[7933] | layer1_out[7932];
     layer2_out[3916] <= ~(layer1_out[1643] | layer1_out[1644]);
     layer2_out[3917] <= layer1_out[3756] & ~layer1_out[3757];
     layer2_out[3918] <= ~layer1_out[3764];
     layer2_out[3919] <= layer1_out[1255] & ~layer1_out[1256];
     layer2_out[3920] <= layer1_out[1483];
     layer2_out[3921] <= ~(layer1_out[7328] ^ layer1_out[7329]);
     layer2_out[3922] <= ~layer1_out[8901] | layer1_out[8900];
     layer2_out[3923] <= ~layer1_out[7115] | layer1_out[7116];
     layer2_out[3924] <= layer1_out[4364] & ~layer1_out[4365];
     layer2_out[3925] <= layer1_out[9035] | layer1_out[9036];
     layer2_out[3926] <= layer1_out[281] & ~layer1_out[280];
     layer2_out[3927] <= layer1_out[6676] & ~layer1_out[6675];
     layer2_out[3928] <= ~layer1_out[3110] | layer1_out[3111];
     layer2_out[3929] <= ~(layer1_out[3788] | layer1_out[3789]);
     layer2_out[3930] <= ~(layer1_out[9272] | layer1_out[9273]);
     layer2_out[3931] <= ~layer1_out[2458] | layer1_out[2457];
     layer2_out[3932] <= ~layer1_out[602];
     layer2_out[3933] <= ~layer1_out[4404] | layer1_out[4403];
     layer2_out[3934] <= ~layer1_out[6856];
     layer2_out[3935] <= ~layer1_out[1796];
     layer2_out[3936] <= layer1_out[11745] & ~layer1_out[11746];
     layer2_out[3937] <= layer1_out[10961] & ~layer1_out[10960];
     layer2_out[3938] <= layer1_out[9277] & ~layer1_out[9276];
     layer2_out[3939] <= ~layer1_out[6596] | layer1_out[6597];
     layer2_out[3940] <= layer1_out[297];
     layer2_out[3941] <= ~layer1_out[9145];
     layer2_out[3942] <= layer1_out[888] & ~layer1_out[889];
     layer2_out[3943] <= layer1_out[6057] & ~layer1_out[6056];
     layer2_out[3944] <= layer1_out[2986] & ~layer1_out[2985];
     layer2_out[3945] <= layer1_out[5685] & ~layer1_out[5686];
     layer2_out[3946] <= layer1_out[10456] | layer1_out[10457];
     layer2_out[3947] <= ~layer1_out[9812] | layer1_out[9813];
     layer2_out[3948] <= 1'b1;
     layer2_out[3949] <= ~layer1_out[1171] | layer1_out[1172];
     layer2_out[3950] <= layer1_out[11861] ^ layer1_out[11862];
     layer2_out[3951] <= ~(layer1_out[5607] & layer1_out[5608]);
     layer2_out[3952] <= layer1_out[8618] & layer1_out[8619];
     layer2_out[3953] <= layer1_out[3578] | layer1_out[3579];
     layer2_out[3954] <= ~(layer1_out[6524] | layer1_out[6525]);
     layer2_out[3955] <= layer1_out[7338] & ~layer1_out[7337];
     layer2_out[3956] <= ~layer1_out[10378];
     layer2_out[3957] <= layer1_out[7362];
     layer2_out[3958] <= ~layer1_out[6326] | layer1_out[6327];
     layer2_out[3959] <= layer1_out[8077] & ~layer1_out[8078];
     layer2_out[3960] <= layer1_out[6248] & ~layer1_out[6249];
     layer2_out[3961] <= ~layer1_out[10974] | layer1_out[10975];
     layer2_out[3962] <= ~(layer1_out[9631] & layer1_out[9632]);
     layer2_out[3963] <= ~layer1_out[7285];
     layer2_out[3964] <= layer1_out[7385];
     layer2_out[3965] <= layer1_out[8673];
     layer2_out[3966] <= layer1_out[9396] & ~layer1_out[9395];
     layer2_out[3967] <= layer1_out[4482] ^ layer1_out[4483];
     layer2_out[3968] <= ~(layer1_out[1831] ^ layer1_out[1832]);
     layer2_out[3969] <= ~layer1_out[10638] | layer1_out[10637];
     layer2_out[3970] <= layer1_out[606] & ~layer1_out[607];
     layer2_out[3971] <= ~(layer1_out[10978] | layer1_out[10979]);
     layer2_out[3972] <= ~(layer1_out[383] & layer1_out[384]);
     layer2_out[3973] <= layer1_out[6329];
     layer2_out[3974] <= layer1_out[8703];
     layer2_out[3975] <= layer1_out[1198] | layer1_out[1199];
     layer2_out[3976] <= layer1_out[5106];
     layer2_out[3977] <= ~layer1_out[1113] | layer1_out[1114];
     layer2_out[3978] <= ~(layer1_out[8558] & layer1_out[8559]);
     layer2_out[3979] <= layer1_out[10897] & ~layer1_out[10896];
     layer2_out[3980] <= layer1_out[8101];
     layer2_out[3981] <= layer1_out[2321];
     layer2_out[3982] <= layer1_out[6033];
     layer2_out[3983] <= layer1_out[7485] & layer1_out[7486];
     layer2_out[3984] <= ~layer1_out[6210];
     layer2_out[3985] <= layer1_out[7511];
     layer2_out[3986] <= ~layer1_out[7438];
     layer2_out[3987] <= layer1_out[3295];
     layer2_out[3988] <= ~layer1_out[5013];
     layer2_out[3989] <= layer1_out[11671];
     layer2_out[3990] <= layer1_out[11336] | layer1_out[11337];
     layer2_out[3991] <= ~layer1_out[7070];
     layer2_out[3992] <= layer1_out[9853] ^ layer1_out[9854];
     layer2_out[3993] <= ~layer1_out[1154];
     layer2_out[3994] <= layer1_out[1981];
     layer2_out[3995] <= layer1_out[7331] & layer1_out[7332];
     layer2_out[3996] <= layer1_out[558];
     layer2_out[3997] <= layer1_out[717];
     layer2_out[3998] <= ~layer1_out[8879];
     layer2_out[3999] <= layer1_out[1114] ^ layer1_out[1115];
     layer2_out[4000] <= ~(layer1_out[11283] | layer1_out[11284]);
     layer2_out[4001] <= ~layer1_out[1814] | layer1_out[1813];
     layer2_out[4002] <= layer1_out[5151] & ~layer1_out[5152];
     layer2_out[4003] <= ~layer1_out[5882];
     layer2_out[4004] <= ~layer1_out[7207] | layer1_out[7208];
     layer2_out[4005] <= ~layer1_out[3428] | layer1_out[3429];
     layer2_out[4006] <= ~layer1_out[8504] | layer1_out[8505];
     layer2_out[4007] <= layer1_out[8023] & layer1_out[8024];
     layer2_out[4008] <= ~layer1_out[7504] | layer1_out[7503];
     layer2_out[4009] <= ~layer1_out[4188];
     layer2_out[4010] <= ~layer1_out[10433];
     layer2_out[4011] <= ~(layer1_out[10707] ^ layer1_out[10708]);
     layer2_out[4012] <= ~layer1_out[5694];
     layer2_out[4013] <= ~layer1_out[4121] | layer1_out[4122];
     layer2_out[4014] <= ~layer1_out[2703] | layer1_out[2704];
     layer2_out[4015] <= ~(layer1_out[3944] ^ layer1_out[3945]);
     layer2_out[4016] <= ~layer1_out[9662];
     layer2_out[4017] <= ~layer1_out[9925];
     layer2_out[4018] <= ~(layer1_out[6819] ^ layer1_out[6820]);
     layer2_out[4019] <= ~layer1_out[11320];
     layer2_out[4020] <= layer1_out[3796] & ~layer1_out[3795];
     layer2_out[4021] <= ~layer1_out[8937];
     layer2_out[4022] <= ~layer1_out[5649] | layer1_out[5648];
     layer2_out[4023] <= layer1_out[6741] | layer1_out[6742];
     layer2_out[4024] <= layer1_out[4300];
     layer2_out[4025] <= layer1_out[9556] & ~layer1_out[9555];
     layer2_out[4026] <= layer1_out[3400] | layer1_out[3401];
     layer2_out[4027] <= layer1_out[7815];
     layer2_out[4028] <= ~(layer1_out[6728] & layer1_out[6729]);
     layer2_out[4029] <= ~layer1_out[1234];
     layer2_out[4030] <= layer1_out[5342];
     layer2_out[4031] <= layer1_out[8406] & ~layer1_out[8407];
     layer2_out[4032] <= ~layer1_out[4278];
     layer2_out[4033] <= ~layer1_out[5762];
     layer2_out[4034] <= ~layer1_out[2015] | layer1_out[2014];
     layer2_out[4035] <= layer1_out[7225];
     layer2_out[4036] <= layer1_out[3099] & ~layer1_out[3100];
     layer2_out[4037] <= layer1_out[10923] & ~layer1_out[10924];
     layer2_out[4038] <= layer1_out[3274];
     layer2_out[4039] <= layer1_out[2087] & ~layer1_out[2088];
     layer2_out[4040] <= ~layer1_out[3229] | layer1_out[3230];
     layer2_out[4041] <= layer1_out[8375] & layer1_out[8376];
     layer2_out[4042] <= layer1_out[11810];
     layer2_out[4043] <= ~(layer1_out[4332] & layer1_out[4333]);
     layer2_out[4044] <= layer1_out[10973];
     layer2_out[4045] <= ~layer1_out[2433] | layer1_out[2432];
     layer2_out[4046] <= layer1_out[9888] ^ layer1_out[9889];
     layer2_out[4047] <= layer1_out[2397] | layer1_out[2398];
     layer2_out[4048] <= layer1_out[4228] ^ layer1_out[4229];
     layer2_out[4049] <= ~layer1_out[9139];
     layer2_out[4050] <= layer1_out[1669] | layer1_out[1670];
     layer2_out[4051] <= ~(layer1_out[2670] & layer1_out[2671]);
     layer2_out[4052] <= ~(layer1_out[9788] ^ layer1_out[9789]);
     layer2_out[4053] <= layer1_out[10321] | layer1_out[10322];
     layer2_out[4054] <= ~(layer1_out[8564] ^ layer1_out[8565]);
     layer2_out[4055] <= 1'b0;
     layer2_out[4056] <= layer1_out[8072];
     layer2_out[4057] <= layer1_out[11708] & layer1_out[11709];
     layer2_out[4058] <= ~layer1_out[3219];
     layer2_out[4059] <= ~layer1_out[4089];
     layer2_out[4060] <= layer1_out[10446] | layer1_out[10447];
     layer2_out[4061] <= layer1_out[5770] | layer1_out[5771];
     layer2_out[4062] <= layer1_out[5700];
     layer2_out[4063] <= ~(layer1_out[1326] | layer1_out[1327]);
     layer2_out[4064] <= ~layer1_out[2496];
     layer2_out[4065] <= ~layer1_out[4997];
     layer2_out[4066] <= layer1_out[1285];
     layer2_out[4067] <= layer1_out[4260] & ~layer1_out[4261];
     layer2_out[4068] <= layer1_out[2454] & ~layer1_out[2455];
     layer2_out[4069] <= ~layer1_out[6873];
     layer2_out[4070] <= ~layer1_out[7871];
     layer2_out[4071] <= layer1_out[2286] & layer1_out[2287];
     layer2_out[4072] <= ~(layer1_out[4488] | layer1_out[4489]);
     layer2_out[4073] <= layer1_out[11521] & ~layer1_out[11520];
     layer2_out[4074] <= layer1_out[11845] ^ layer1_out[11846];
     layer2_out[4075] <= 1'b1;
     layer2_out[4076] <= ~layer1_out[9095];
     layer2_out[4077] <= ~(layer1_out[1758] & layer1_out[1759]);
     layer2_out[4078] <= layer1_out[224] & ~layer1_out[225];
     layer2_out[4079] <= layer1_out[5744];
     layer2_out[4080] <= layer1_out[10411];
     layer2_out[4081] <= layer1_out[5475];
     layer2_out[4082] <= ~layer1_out[4804];
     layer2_out[4083] <= ~layer1_out[986];
     layer2_out[4084] <= ~layer1_out[1557];
     layer2_out[4085] <= ~layer1_out[4110];
     layer2_out[4086] <= ~layer1_out[5952];
     layer2_out[4087] <= ~layer1_out[7516] | layer1_out[7517];
     layer2_out[4088] <= layer1_out[426];
     layer2_out[4089] <= layer1_out[2289] & layer1_out[2290];
     layer2_out[4090] <= ~layer1_out[4072] | layer1_out[4073];
     layer2_out[4091] <= layer1_out[3310] | layer1_out[3311];
     layer2_out[4092] <= layer1_out[5960];
     layer2_out[4093] <= layer1_out[1209] & layer1_out[1210];
     layer2_out[4094] <= layer1_out[8277] | layer1_out[8278];
     layer2_out[4095] <= ~layer1_out[7016];
     layer2_out[4096] <= ~layer1_out[7283];
     layer2_out[4097] <= ~layer1_out[5400];
     layer2_out[4098] <= layer1_out[11571] & layer1_out[11572];
     layer2_out[4099] <= ~layer1_out[11265];
     layer2_out[4100] <= ~(layer1_out[1066] | layer1_out[1067]);
     layer2_out[4101] <= ~layer1_out[4830] | layer1_out[4829];
     layer2_out[4102] <= layer1_out[2894] | layer1_out[2895];
     layer2_out[4103] <= layer1_out[10671] & layer1_out[10672];
     layer2_out[4104] <= ~(layer1_out[7908] & layer1_out[7909]);
     layer2_out[4105] <= ~layer1_out[11530];
     layer2_out[4106] <= layer1_out[971];
     layer2_out[4107] <= ~(layer1_out[3226] & layer1_out[3227]);
     layer2_out[4108] <= layer1_out[2093] ^ layer1_out[2094];
     layer2_out[4109] <= ~(layer1_out[9085] ^ layer1_out[9086]);
     layer2_out[4110] <= ~layer1_out[5711];
     layer2_out[4111] <= layer1_out[11165];
     layer2_out[4112] <= layer1_out[1667];
     layer2_out[4113] <= layer1_out[4827] | layer1_out[4828];
     layer2_out[4114] <= ~layer1_out[3648];
     layer2_out[4115] <= ~(layer1_out[9177] ^ layer1_out[9178]);
     layer2_out[4116] <= layer1_out[5702] & layer1_out[5703];
     layer2_out[4117] <= ~layer1_out[7614];
     layer2_out[4118] <= layer1_out[4036] | layer1_out[4037];
     layer2_out[4119] <= ~(layer1_out[45] & layer1_out[46]);
     layer2_out[4120] <= ~layer1_out[6007];
     layer2_out[4121] <= layer1_out[5019] & ~layer1_out[5018];
     layer2_out[4122] <= ~layer1_out[19];
     layer2_out[4123] <= layer1_out[8442] ^ layer1_out[8443];
     layer2_out[4124] <= layer1_out[7842] & layer1_out[7843];
     layer2_out[4125] <= layer1_out[7856];
     layer2_out[4126] <= layer1_out[8881] & ~layer1_out[8882];
     layer2_out[4127] <= layer1_out[11660] & layer1_out[11661];
     layer2_out[4128] <= ~(layer1_out[11498] & layer1_out[11499]);
     layer2_out[4129] <= layer1_out[8688] | layer1_out[8689];
     layer2_out[4130] <= ~(layer1_out[9666] & layer1_out[9667]);
     layer2_out[4131] <= ~layer1_out[7411];
     layer2_out[4132] <= ~layer1_out[7050];
     layer2_out[4133] <= layer1_out[8528] & ~layer1_out[8529];
     layer2_out[4134] <= layer1_out[3321];
     layer2_out[4135] <= layer1_out[11515];
     layer2_out[4136] <= layer1_out[6235] ^ layer1_out[6236];
     layer2_out[4137] <= layer1_out[7726];
     layer2_out[4138] <= layer1_out[6211] & ~layer1_out[6210];
     layer2_out[4139] <= layer1_out[2544];
     layer2_out[4140] <= layer1_out[82] & ~layer1_out[81];
     layer2_out[4141] <= ~(layer1_out[4728] | layer1_out[4729]);
     layer2_out[4142] <= ~layer1_out[8044];
     layer2_out[4143] <= ~(layer1_out[9136] & layer1_out[9137]);
     layer2_out[4144] <= ~(layer1_out[1533] & layer1_out[1534]);
     layer2_out[4145] <= layer1_out[8883];
     layer2_out[4146] <= ~layer1_out[3732];
     layer2_out[4147] <= ~layer1_out[7218];
     layer2_out[4148] <= layer1_out[10397];
     layer2_out[4149] <= layer1_out[2746] & ~layer1_out[2747];
     layer2_out[4150] <= layer1_out[6269] & ~layer1_out[6268];
     layer2_out[4151] <= ~layer1_out[3340] | layer1_out[3339];
     layer2_out[4152] <= ~layer1_out[5007];
     layer2_out[4153] <= layer1_out[5827];
     layer2_out[4154] <= layer1_out[2851] & ~layer1_out[2850];
     layer2_out[4155] <= ~layer1_out[4811];
     layer2_out[4156] <= ~(layer1_out[4809] & layer1_out[4810]);
     layer2_out[4157] <= layer1_out[2174];
     layer2_out[4158] <= ~layer1_out[1672] | layer1_out[1671];
     layer2_out[4159] <= layer1_out[43] | layer1_out[44];
     layer2_out[4160] <= layer1_out[6899] & ~layer1_out[6900];
     layer2_out[4161] <= layer1_out[11985] & layer1_out[11986];
     layer2_out[4162] <= ~layer1_out[3040];
     layer2_out[4163] <= layer1_out[10868] & layer1_out[10869];
     layer2_out[4164] <= layer1_out[7558] | layer1_out[7559];
     layer2_out[4165] <= ~layer1_out[2832];
     layer2_out[4166] <= ~layer1_out[9416] | layer1_out[9415];
     layer2_out[4167] <= layer1_out[4283] & ~layer1_out[4282];
     layer2_out[4168] <= ~(layer1_out[3506] & layer1_out[3507]);
     layer2_out[4169] <= layer1_out[7193];
     layer2_out[4170] <= layer1_out[369];
     layer2_out[4171] <= layer1_out[7785] & ~layer1_out[7784];
     layer2_out[4172] <= layer1_out[11662] | layer1_out[11663];
     layer2_out[4173] <= layer1_out[7803];
     layer2_out[4174] <= ~layer1_out[6736] | layer1_out[6735];
     layer2_out[4175] <= layer1_out[11352] | layer1_out[11353];
     layer2_out[4176] <= layer1_out[10195];
     layer2_out[4177] <= ~layer1_out[11274];
     layer2_out[4178] <= ~(layer1_out[6156] | layer1_out[6157]);
     layer2_out[4179] <= ~layer1_out[5807];
     layer2_out[4180] <= layer1_out[339];
     layer2_out[4181] <= layer1_out[5193] & layer1_out[5194];
     layer2_out[4182] <= layer1_out[11278];
     layer2_out[4183] <= ~layer1_out[2133];
     layer2_out[4184] <= layer1_out[7143];
     layer2_out[4185] <= ~layer1_out[3103] | layer1_out[3102];
     layer2_out[4186] <= layer1_out[7789];
     layer2_out[4187] <= ~layer1_out[10218];
     layer2_out[4188] <= ~layer1_out[10507];
     layer2_out[4189] <= ~layer1_out[7937] | layer1_out[7936];
     layer2_out[4190] <= ~layer1_out[1673];
     layer2_out[4191] <= ~layer1_out[5058];
     layer2_out[4192] <= layer1_out[4257];
     layer2_out[4193] <= ~layer1_out[10070];
     layer2_out[4194] <= ~layer1_out[9941];
     layer2_out[4195] <= layer1_out[9538];
     layer2_out[4196] <= layer1_out[11605] & ~layer1_out[11604];
     layer2_out[4197] <= layer1_out[7662] & ~layer1_out[7663];
     layer2_out[4198] <= layer1_out[9333];
     layer2_out[4199] <= ~(layer1_out[251] | layer1_out[252]);
     layer2_out[4200] <= layer1_out[11609] | layer1_out[11610];
     layer2_out[4201] <= ~layer1_out[10282] | layer1_out[10281];
     layer2_out[4202] <= ~layer1_out[6752] | layer1_out[6751];
     layer2_out[4203] <= ~(layer1_out[8189] ^ layer1_out[8190]);
     layer2_out[4204] <= ~(layer1_out[406] & layer1_out[407]);
     layer2_out[4205] <= ~layer1_out[4775] | layer1_out[4776];
     layer2_out[4206] <= layer1_out[8682];
     layer2_out[4207] <= layer1_out[10894];
     layer2_out[4208] <= 1'b0;
     layer2_out[4209] <= ~layer1_out[10219];
     layer2_out[4210] <= layer1_out[4697] & layer1_out[4698];
     layer2_out[4211] <= layer1_out[3225] ^ layer1_out[3226];
     layer2_out[4212] <= layer1_out[7817] ^ layer1_out[7818];
     layer2_out[4213] <= layer1_out[1466];
     layer2_out[4214] <= ~(layer1_out[3012] | layer1_out[3013]);
     layer2_out[4215] <= layer1_out[4164] ^ layer1_out[4165];
     layer2_out[4216] <= layer1_out[9925];
     layer2_out[4217] <= layer1_out[7586];
     layer2_out[4218] <= ~layer1_out[10823] | layer1_out[10822];
     layer2_out[4219] <= ~(layer1_out[5729] & layer1_out[5730]);
     layer2_out[4220] <= ~layer1_out[1247];
     layer2_out[4221] <= ~layer1_out[9227];
     layer2_out[4222] <= layer1_out[11012];
     layer2_out[4223] <= ~layer1_out[9849] | layer1_out[9848];
     layer2_out[4224] <= ~layer1_out[9809] | layer1_out[9808];
     layer2_out[4225] <= layer1_out[8559] ^ layer1_out[8560];
     layer2_out[4226] <= layer1_out[10059];
     layer2_out[4227] <= layer1_out[11625] | layer1_out[11626];
     layer2_out[4228] <= ~layer1_out[5921] | layer1_out[5922];
     layer2_out[4229] <= ~(layer1_out[10587] & layer1_out[10588]);
     layer2_out[4230] <= 1'b1;
     layer2_out[4231] <= layer1_out[5253];
     layer2_out[4232] <= layer1_out[2028] & ~layer1_out[2027];
     layer2_out[4233] <= layer1_out[1641];
     layer2_out[4234] <= ~(layer1_out[9457] ^ layer1_out[9458]);
     layer2_out[4235] <= layer1_out[3163] | layer1_out[3164];
     layer2_out[4236] <= layer1_out[8803];
     layer2_out[4237] <= ~layer1_out[4002];
     layer2_out[4238] <= ~layer1_out[2885] | layer1_out[2884];
     layer2_out[4239] <= layer1_out[393] ^ layer1_out[394];
     layer2_out[4240] <= layer1_out[10478] & layer1_out[10479];
     layer2_out[4241] <= ~layer1_out[6104];
     layer2_out[4242] <= layer1_out[694];
     layer2_out[4243] <= layer1_out[11906] | layer1_out[11907];
     layer2_out[4244] <= layer1_out[6983] ^ layer1_out[6984];
     layer2_out[4245] <= layer1_out[2650];
     layer2_out[4246] <= layer1_out[8487] & ~layer1_out[8486];
     layer2_out[4247] <= ~layer1_out[12];
     layer2_out[4248] <= ~(layer1_out[350] | layer1_out[351]);
     layer2_out[4249] <= layer1_out[4499];
     layer2_out[4250] <= layer1_out[4517] | layer1_out[4518];
     layer2_out[4251] <= layer1_out[9070];
     layer2_out[4252] <= ~(layer1_out[11752] & layer1_out[11753]);
     layer2_out[4253] <= layer1_out[2434];
     layer2_out[4254] <= ~layer1_out[410] | layer1_out[411];
     layer2_out[4255] <= layer1_out[1550] & ~layer1_out[1549];
     layer2_out[4256] <= ~(layer1_out[3444] ^ layer1_out[3445]);
     layer2_out[4257] <= ~layer1_out[9845];
     layer2_out[4258] <= layer1_out[166];
     layer2_out[4259] <= layer1_out[1916];
     layer2_out[4260] <= layer1_out[11354] | layer1_out[11355];
     layer2_out[4261] <= ~layer1_out[11622];
     layer2_out[4262] <= ~layer1_out[7940];
     layer2_out[4263] <= ~(layer1_out[11115] | layer1_out[11116]);
     layer2_out[4264] <= 1'b0;
     layer2_out[4265] <= layer1_out[4683];
     layer2_out[4266] <= layer1_out[3133] | layer1_out[3134];
     layer2_out[4267] <= ~layer1_out[6043];
     layer2_out[4268] <= layer1_out[2716];
     layer2_out[4269] <= ~(layer1_out[1790] ^ layer1_out[1791]);
     layer2_out[4270] <= layer1_out[6109] & ~layer1_out[6108];
     layer2_out[4271] <= layer1_out[8740] & ~layer1_out[8741];
     layer2_out[4272] <= layer1_out[4569] ^ layer1_out[4570];
     layer2_out[4273] <= layer1_out[5572];
     layer2_out[4274] <= ~(layer1_out[8275] ^ layer1_out[8276]);
     layer2_out[4275] <= layer1_out[4419];
     layer2_out[4276] <= ~layer1_out[4868];
     layer2_out[4277] <= layer1_out[1586] | layer1_out[1587];
     layer2_out[4278] <= ~layer1_out[10037];
     layer2_out[4279] <= ~(layer1_out[2893] | layer1_out[2894]);
     layer2_out[4280] <= layer1_out[2690] & ~layer1_out[2689];
     layer2_out[4281] <= ~layer1_out[10518];
     layer2_out[4282] <= ~layer1_out[11319];
     layer2_out[4283] <= ~layer1_out[10250];
     layer2_out[4284] <= ~layer1_out[8501] | layer1_out[8500];
     layer2_out[4285] <= ~layer1_out[245];
     layer2_out[4286] <= 1'b0;
     layer2_out[4287] <= ~layer1_out[332] | layer1_out[331];
     layer2_out[4288] <= layer1_out[8444];
     layer2_out[4289] <= layer1_out[10684] & ~layer1_out[10685];
     layer2_out[4290] <= ~(layer1_out[8434] & layer1_out[8435]);
     layer2_out[4291] <= layer1_out[2853] | layer1_out[2854];
     layer2_out[4292] <= ~layer1_out[5043];
     layer2_out[4293] <= ~layer1_out[7173] | layer1_out[7172];
     layer2_out[4294] <= layer1_out[11860] & layer1_out[11861];
     layer2_out[4295] <= ~layer1_out[10715];
     layer2_out[4296] <= layer1_out[7833] & ~layer1_out[7832];
     layer2_out[4297] <= ~(layer1_out[6166] | layer1_out[6167]);
     layer2_out[4298] <= layer1_out[8107] | layer1_out[8108];
     layer2_out[4299] <= layer1_out[6089];
     layer2_out[4300] <= ~layer1_out[9755] | layer1_out[9754];
     layer2_out[4301] <= layer1_out[3101] ^ layer1_out[3102];
     layer2_out[4302] <= ~layer1_out[4999] | layer1_out[5000];
     layer2_out[4303] <= layer1_out[6081] & ~layer1_out[6080];
     layer2_out[4304] <= layer1_out[2482] & ~layer1_out[2483];
     layer2_out[4305] <= ~(layer1_out[4604] & layer1_out[4605]);
     layer2_out[4306] <= layer1_out[4863];
     layer2_out[4307] <= layer1_out[2471] & layer1_out[2472];
     layer2_out[4308] <= layer1_out[10600] & layer1_out[10601];
     layer2_out[4309] <= layer1_out[8685] | layer1_out[8686];
     layer2_out[4310] <= ~(layer1_out[6485] | layer1_out[6486]);
     layer2_out[4311] <= layer1_out[5107] & layer1_out[5108];
     layer2_out[4312] <= layer1_out[3417] ^ layer1_out[3418];
     layer2_out[4313] <= ~layer1_out[6469];
     layer2_out[4314] <= ~layer1_out[2644];
     layer2_out[4315] <= ~layer1_out[11019];
     layer2_out[4316] <= ~(layer1_out[11896] ^ layer1_out[11897]);
     layer2_out[4317] <= layer1_out[4099] & layer1_out[4100];
     layer2_out[4318] <= layer1_out[6535];
     layer2_out[4319] <= ~(layer1_out[8231] ^ layer1_out[8232]);
     layer2_out[4320] <= layer1_out[639] & layer1_out[640];
     layer2_out[4321] <= layer1_out[4081];
     layer2_out[4322] <= ~layer1_out[6687];
     layer2_out[4323] <= ~layer1_out[4313];
     layer2_out[4324] <= ~layer1_out[9746] | layer1_out[9745];
     layer2_out[4325] <= layer1_out[1349];
     layer2_out[4326] <= ~layer1_out[4654];
     layer2_out[4327] <= ~layer1_out[10138];
     layer2_out[4328] <= ~layer1_out[10284] | layer1_out[10283];
     layer2_out[4329] <= layer1_out[10620] & ~layer1_out[10621];
     layer2_out[4330] <= layer1_out[8608] & ~layer1_out[8607];
     layer2_out[4331] <= layer1_out[8017];
     layer2_out[4332] <= layer1_out[1593] & ~layer1_out[1594];
     layer2_out[4333] <= layer1_out[7730] & ~layer1_out[7731];
     layer2_out[4334] <= ~(layer1_out[900] ^ layer1_out[901]);
     layer2_out[4335] <= ~layer1_out[2140];
     layer2_out[4336] <= ~(layer1_out[570] | layer1_out[571]);
     layer2_out[4337] <= ~layer1_out[9009];
     layer2_out[4338] <= ~layer1_out[4954];
     layer2_out[4339] <= ~(layer1_out[8377] ^ layer1_out[8378]);
     layer2_out[4340] <= ~layer1_out[8969];
     layer2_out[4341] <= ~(layer1_out[2315] & layer1_out[2316]);
     layer2_out[4342] <= layer1_out[6555];
     layer2_out[4343] <= ~layer1_out[10146];
     layer2_out[4344] <= layer1_out[4643];
     layer2_out[4345] <= ~layer1_out[9666];
     layer2_out[4346] <= layer1_out[7243];
     layer2_out[4347] <= ~layer1_out[610] | layer1_out[611];
     layer2_out[4348] <= layer1_out[9210];
     layer2_out[4349] <= ~layer1_out[7386] | layer1_out[7385];
     layer2_out[4350] <= ~layer1_out[1251] | layer1_out[1250];
     layer2_out[4351] <= ~layer1_out[10423];
     layer2_out[4352] <= ~layer1_out[1445];
     layer2_out[4353] <= layer1_out[7288];
     layer2_out[4354] <= ~layer1_out[5394];
     layer2_out[4355] <= layer1_out[2656];
     layer2_out[4356] <= layer1_out[2468] & ~layer1_out[2469];
     layer2_out[4357] <= layer1_out[9775];
     layer2_out[4358] <= layer1_out[2131] & layer1_out[2132];
     layer2_out[4359] <= layer1_out[5552];
     layer2_out[4360] <= ~(layer1_out[10982] ^ layer1_out[10983]);
     layer2_out[4361] <= layer1_out[9221];
     layer2_out[4362] <= ~layer1_out[11857];
     layer2_out[4363] <= layer1_out[396] | layer1_out[397];
     layer2_out[4364] <= ~layer1_out[6575] | layer1_out[6576];
     layer2_out[4365] <= ~layer1_out[4820];
     layer2_out[4366] <= layer1_out[8475] & ~layer1_out[8474];
     layer2_out[4367] <= layer1_out[6218] ^ layer1_out[6219];
     layer2_out[4368] <= layer1_out[10408] ^ layer1_out[10409];
     layer2_out[4369] <= ~layer1_out[3698] | layer1_out[3699];
     layer2_out[4370] <= ~layer1_out[7149];
     layer2_out[4371] <= ~(layer1_out[959] & layer1_out[960]);
     layer2_out[4372] <= ~layer1_out[404] | layer1_out[403];
     layer2_out[4373] <= ~(layer1_out[7028] ^ layer1_out[7029]);
     layer2_out[4374] <= 1'b0;
     layer2_out[4375] <= layer1_out[670];
     layer2_out[4376] <= layer1_out[5799];
     layer2_out[4377] <= ~(layer1_out[6716] & layer1_out[6717]);
     layer2_out[4378] <= ~layer1_out[9000];
     layer2_out[4379] <= ~layer1_out[4655];
     layer2_out[4380] <= layer1_out[1776] & ~layer1_out[1777];
     layer2_out[4381] <= layer1_out[9281] & ~layer1_out[9280];
     layer2_out[4382] <= ~(layer1_out[4146] & layer1_out[4147]);
     layer2_out[4383] <= ~(layer1_out[1044] ^ layer1_out[1045]);
     layer2_out[4384] <= ~layer1_out[1178];
     layer2_out[4385] <= ~layer1_out[6163];
     layer2_out[4386] <= ~layer1_out[1574];
     layer2_out[4387] <= ~layer1_out[9180] | layer1_out[9179];
     layer2_out[4388] <= ~layer1_out[6008];
     layer2_out[4389] <= layer1_out[3395] | layer1_out[3396];
     layer2_out[4390] <= layer1_out[2854] & layer1_out[2855];
     layer2_out[4391] <= ~layer1_out[9293];
     layer2_out[4392] <= ~(layer1_out[9772] ^ layer1_out[9773]);
     layer2_out[4393] <= layer1_out[8767];
     layer2_out[4394] <= ~layer1_out[3586];
     layer2_out[4395] <= layer1_out[5621] ^ layer1_out[5622];
     layer2_out[4396] <= ~(layer1_out[3451] | layer1_out[3452]);
     layer2_out[4397] <= layer1_out[10076] & ~layer1_out[10077];
     layer2_out[4398] <= layer1_out[5276];
     layer2_out[4399] <= layer1_out[10557] | layer1_out[10558];
     layer2_out[4400] <= layer1_out[10667];
     layer2_out[4401] <= layer1_out[9871] & layer1_out[9872];
     layer2_out[4402] <= ~layer1_out[3086];
     layer2_out[4403] <= ~layer1_out[4526];
     layer2_out[4404] <= ~(layer1_out[3403] & layer1_out[3404]);
     layer2_out[4405] <= layer1_out[1485];
     layer2_out[4406] <= layer1_out[9107] & ~layer1_out[9108];
     layer2_out[4407] <= ~layer1_out[8916] | layer1_out[8915];
     layer2_out[4408] <= layer1_out[7317] & ~layer1_out[7318];
     layer2_out[4409] <= ~(layer1_out[5775] ^ layer1_out[5776]);
     layer2_out[4410] <= layer1_out[10493];
     layer2_out[4411] <= layer1_out[1578] | layer1_out[1579];
     layer2_out[4412] <= ~layer1_out[4418];
     layer2_out[4413] <= layer1_out[1221] & ~layer1_out[1220];
     layer2_out[4414] <= layer1_out[10445] | layer1_out[10446];
     layer2_out[4415] <= layer1_out[7900];
     layer2_out[4416] <= ~layer1_out[2983];
     layer2_out[4417] <= ~layer1_out[10156];
     layer2_out[4418] <= ~(layer1_out[6813] | layer1_out[6814]);
     layer2_out[4419] <= ~layer1_out[11468];
     layer2_out[4420] <= ~(layer1_out[2167] & layer1_out[2168]);
     layer2_out[4421] <= ~layer1_out[8648] | layer1_out[8647];
     layer2_out[4422] <= layer1_out[2872] & layer1_out[2873];
     layer2_out[4423] <= layer1_out[5132];
     layer2_out[4424] <= layer1_out[5613];
     layer2_out[4425] <= layer1_out[478] & ~layer1_out[479];
     layer2_out[4426] <= layer1_out[4937] ^ layer1_out[4938];
     layer2_out[4427] <= ~(layer1_out[4745] | layer1_out[4746]);
     layer2_out[4428] <= layer1_out[10958] | layer1_out[10959];
     layer2_out[4429] <= ~layer1_out[6422] | layer1_out[6423];
     layer2_out[4430] <= ~layer1_out[7458] | layer1_out[7459];
     layer2_out[4431] <= ~(layer1_out[11993] ^ layer1_out[11994]);
     layer2_out[4432] <= ~layer1_out[5146];
     layer2_out[4433] <= layer1_out[3263];
     layer2_out[4434] <= layer1_out[9930] & layer1_out[9931];
     layer2_out[4435] <= ~layer1_out[2156] | layer1_out[2155];
     layer2_out[4436] <= ~(layer1_out[8735] | layer1_out[8736]);
     layer2_out[4437] <= layer1_out[4543];
     layer2_out[4438] <= ~layer1_out[9194];
     layer2_out[4439] <= ~(layer1_out[10418] ^ layer1_out[10419]);
     layer2_out[4440] <= layer1_out[2632];
     layer2_out[4441] <= ~layer1_out[11741] | layer1_out[11740];
     layer2_out[4442] <= ~layer1_out[1683] | layer1_out[1684];
     layer2_out[4443] <= layer1_out[9734];
     layer2_out[4444] <= layer1_out[6747] & ~layer1_out[6746];
     layer2_out[4445] <= ~layer1_out[5787];
     layer2_out[4446] <= layer1_out[1728] & layer1_out[1729];
     layer2_out[4447] <= layer1_out[764] ^ layer1_out[765];
     layer2_out[4448] <= layer1_out[8809] & ~layer1_out[8808];
     layer2_out[4449] <= layer1_out[7707];
     layer2_out[4450] <= layer1_out[8780];
     layer2_out[4451] <= layer1_out[3044] | layer1_out[3045];
     layer2_out[4452] <= layer1_out[5579] & ~layer1_out[5578];
     layer2_out[4453] <= ~layer1_out[1290] | layer1_out[1289];
     layer2_out[4454] <= layer1_out[4285];
     layer2_out[4455] <= ~(layer1_out[2669] & layer1_out[2670]);
     layer2_out[4456] <= layer1_out[3110] & ~layer1_out[3109];
     layer2_out[4457] <= ~(layer1_out[1480] & layer1_out[1481]);
     layer2_out[4458] <= ~layer1_out[11336];
     layer2_out[4459] <= layer1_out[6424] & layer1_out[6425];
     layer2_out[4460] <= ~(layer1_out[11570] & layer1_out[11571]);
     layer2_out[4461] <= layer1_out[11990];
     layer2_out[4462] <= ~layer1_out[6494];
     layer2_out[4463] <= ~layer1_out[2406] | layer1_out[2405];
     layer2_out[4464] <= ~(layer1_out[4877] ^ layer1_out[4878]);
     layer2_out[4465] <= layer1_out[7997];
     layer2_out[4466] <= layer1_out[1810];
     layer2_out[4467] <= ~layer1_out[9302];
     layer2_out[4468] <= layer1_out[11224] & layer1_out[11225];
     layer2_out[4469] <= ~(layer1_out[8602] ^ layer1_out[8603]);
     layer2_out[4470] <= layer1_out[37] & ~layer1_out[38];
     layer2_out[4471] <= layer1_out[8831] & ~layer1_out[8832];
     layer2_out[4472] <= ~layer1_out[6526];
     layer2_out[4473] <= ~layer1_out[11100] | layer1_out[11099];
     layer2_out[4474] <= layer1_out[7295] & ~layer1_out[7296];
     layer2_out[4475] <= layer1_out[8532];
     layer2_out[4476] <= ~layer1_out[5734];
     layer2_out[4477] <= ~layer1_out[1690] | layer1_out[1691];
     layer2_out[4478] <= ~(layer1_out[2112] | layer1_out[2113]);
     layer2_out[4479] <= ~(layer1_out[771] ^ layer1_out[772]);
     layer2_out[4480] <= layer1_out[5757] & layer1_out[5758];
     layer2_out[4481] <= layer1_out[3278] & ~layer1_out[3277];
     layer2_out[4482] <= ~layer1_out[6571] | layer1_out[6570];
     layer2_out[4483] <= layer1_out[5249];
     layer2_out[4484] <= ~layer1_out[6000];
     layer2_out[4485] <= layer1_out[9442];
     layer2_out[4486] <= layer1_out[3317];
     layer2_out[4487] <= ~layer1_out[7899];
     layer2_out[4488] <= 1'b1;
     layer2_out[4489] <= layer1_out[5601] | layer1_out[5602];
     layer2_out[4490] <= layer1_out[8958];
     layer2_out[4491] <= layer1_out[207] & ~layer1_out[206];
     layer2_out[4492] <= ~(layer1_out[5822] ^ layer1_out[5823]);
     layer2_out[4493] <= ~layer1_out[10851];
     layer2_out[4494] <= layer1_out[8131];
     layer2_out[4495] <= layer1_out[3485];
     layer2_out[4496] <= ~(layer1_out[5427] ^ layer1_out[5428]);
     layer2_out[4497] <= ~layer1_out[8523];
     layer2_out[4498] <= layer1_out[2787] ^ layer1_out[2788];
     layer2_out[4499] <= layer1_out[4892] | layer1_out[4893];
     layer2_out[4500] <= layer1_out[11073] & layer1_out[11074];
     layer2_out[4501] <= layer1_out[10055] & layer1_out[10056];
     layer2_out[4502] <= 1'b0;
     layer2_out[4503] <= layer1_out[2914] | layer1_out[2915];
     layer2_out[4504] <= ~layer1_out[1447];
     layer2_out[4505] <= layer1_out[6443] | layer1_out[6444];
     layer2_out[4506] <= layer1_out[643];
     layer2_out[4507] <= layer1_out[2665];
     layer2_out[4508] <= layer1_out[1804] | layer1_out[1805];
     layer2_out[4509] <= layer1_out[7870] ^ layer1_out[7871];
     layer2_out[4510] <= ~layer1_out[336];
     layer2_out[4511] <= layer1_out[5220] & ~layer1_out[5221];
     layer2_out[4512] <= ~layer1_out[10577];
     layer2_out[4513] <= layer1_out[1227];
     layer2_out[4514] <= ~layer1_out[7138] | layer1_out[7139];
     layer2_out[4515] <= ~layer1_out[6212];
     layer2_out[4516] <= ~(layer1_out[925] | layer1_out[926]);
     layer2_out[4517] <= layer1_out[10419] & ~layer1_out[10420];
     layer2_out[4518] <= ~layer1_out[10400] | layer1_out[10401];
     layer2_out[4519] <= 1'b0;
     layer2_out[4520] <= ~layer1_out[1273] | layer1_out[1272];
     layer2_out[4521] <= layer1_out[4460] | layer1_out[4461];
     layer2_out[4522] <= 1'b0;
     layer2_out[4523] <= layer1_out[8504];
     layer2_out[4524] <= ~(layer1_out[4600] ^ layer1_out[4601]);
     layer2_out[4525] <= layer1_out[2052] ^ layer1_out[2053];
     layer2_out[4526] <= ~(layer1_out[65] ^ layer1_out[66]);
     layer2_out[4527] <= layer1_out[6606] | layer1_out[6607];
     layer2_out[4528] <= ~layer1_out[1734] | layer1_out[1733];
     layer2_out[4529] <= layer1_out[6507] & layer1_out[6508];
     layer2_out[4530] <= ~(layer1_out[10799] | layer1_out[10800]);
     layer2_out[4531] <= layer1_out[9264];
     layer2_out[4532] <= layer1_out[4224] & layer1_out[4225];
     layer2_out[4533] <= ~layer1_out[441];
     layer2_out[4534] <= ~(layer1_out[8240] & layer1_out[8241]);
     layer2_out[4535] <= layer1_out[389];
     layer2_out[4536] <= layer1_out[10067];
     layer2_out[4537] <= layer1_out[745];
     layer2_out[4538] <= ~layer1_out[9528] | layer1_out[9527];
     layer2_out[4539] <= layer1_out[8297] & ~layer1_out[8296];
     layer2_out[4540] <= layer1_out[6952] | layer1_out[6953];
     layer2_out[4541] <= ~layer1_out[9233];
     layer2_out[4542] <= layer1_out[10444];
     layer2_out[4543] <= ~(layer1_out[2067] | layer1_out[2068]);
     layer2_out[4544] <= ~(layer1_out[6949] & layer1_out[6950]);
     layer2_out[4545] <= ~(layer1_out[1909] ^ layer1_out[1910]);
     layer2_out[4546] <= layer1_out[6642];
     layer2_out[4547] <= layer1_out[3057];
     layer2_out[4548] <= layer1_out[1095] & layer1_out[1096];
     layer2_out[4549] <= ~layer1_out[10963];
     layer2_out[4550] <= ~(layer1_out[2731] | layer1_out[2732]);
     layer2_out[4551] <= layer1_out[2677] & ~layer1_out[2678];
     layer2_out[4552] <= ~layer1_out[9676] | layer1_out[9677];
     layer2_out[4553] <= ~layer1_out[8684] | layer1_out[8683];
     layer2_out[4554] <= ~(layer1_out[3916] & layer1_out[3917]);
     layer2_out[4555] <= layer1_out[7185];
     layer2_out[4556] <= ~layer1_out[10092] | layer1_out[10091];
     layer2_out[4557] <= layer1_out[3525];
     layer2_out[4558] <= ~layer1_out[4666] | layer1_out[4667];
     layer2_out[4559] <= layer1_out[7204] & layer1_out[7205];
     layer2_out[4560] <= ~(layer1_out[60] | layer1_out[61]);
     layer2_out[4561] <= layer1_out[5494];
     layer2_out[4562] <= layer1_out[4475];
     layer2_out[4563] <= ~(layer1_out[9567] ^ layer1_out[9568]);
     layer2_out[4564] <= ~(layer1_out[1314] & layer1_out[1315]);
     layer2_out[4565] <= ~layer1_out[8524];
     layer2_out[4566] <= ~layer1_out[9867] | layer1_out[9866];
     layer2_out[4567] <= ~layer1_out[1865];
     layer2_out[4568] <= ~layer1_out[3247];
     layer2_out[4569] <= layer1_out[7973] & layer1_out[7974];
     layer2_out[4570] <= layer1_out[2504] ^ layer1_out[2505];
     layer2_out[4571] <= ~(layer1_out[10237] ^ layer1_out[10238]);
     layer2_out[4572] <= ~(layer1_out[3802] | layer1_out[3803]);
     layer2_out[4573] <= ~(layer1_out[2268] | layer1_out[2269]);
     layer2_out[4574] <= ~layer1_out[9600] | layer1_out[9601];
     layer2_out[4575] <= layer1_out[11686];
     layer2_out[4576] <= ~(layer1_out[11441] & layer1_out[11442]);
     layer2_out[4577] <= layer1_out[3884];
     layer2_out[4578] <= layer1_out[57] & ~layer1_out[56];
     layer2_out[4579] <= ~layer1_out[5988];
     layer2_out[4580] <= ~(layer1_out[10553] ^ layer1_out[10554]);
     layer2_out[4581] <= layer1_out[6970] & ~layer1_out[6969];
     layer2_out[4582] <= layer1_out[3381];
     layer2_out[4583] <= layer1_out[10026] & ~layer1_out[10025];
     layer2_out[4584] <= layer1_out[6657];
     layer2_out[4585] <= ~layer1_out[9916] | layer1_out[9917];
     layer2_out[4586] <= ~layer1_out[5139] | layer1_out[5140];
     layer2_out[4587] <= layer1_out[10720] | layer1_out[10721];
     layer2_out[4588] <= ~(layer1_out[3351] & layer1_out[3352]);
     layer2_out[4589] <= ~layer1_out[838];
     layer2_out[4590] <= layer1_out[9539] & ~layer1_out[9540];
     layer2_out[4591] <= ~layer1_out[3455];
     layer2_out[4592] <= ~layer1_out[7522];
     layer2_out[4593] <= ~layer1_out[2057];
     layer2_out[4594] <= ~(layer1_out[881] ^ layer1_out[882]);
     layer2_out[4595] <= layer1_out[3491];
     layer2_out[4596] <= layer1_out[7236] | layer1_out[7237];
     layer2_out[4597] <= layer1_out[9120];
     layer2_out[4598] <= ~layer1_out[8172];
     layer2_out[4599] <= ~(layer1_out[960] & layer1_out[961]);
     layer2_out[4600] <= ~layer1_out[5966];
     layer2_out[4601] <= ~(layer1_out[1564] ^ layer1_out[1565]);
     layer2_out[4602] <= ~layer1_out[2243];
     layer2_out[4603] <= 1'b0;
     layer2_out[4604] <= ~(layer1_out[9424] ^ layer1_out[9425]);
     layer2_out[4605] <= layer1_out[1507] & ~layer1_out[1506];
     layer2_out[4606] <= ~layer1_out[7844] | layer1_out[7845];
     layer2_out[4607] <= 1'b0;
     layer2_out[4608] <= layer1_out[651] & ~layer1_out[652];
     layer2_out[4609] <= layer1_out[460] & layer1_out[461];
     layer2_out[4610] <= ~layer1_out[3051] | layer1_out[3050];
     layer2_out[4611] <= layer1_out[1978];
     layer2_out[4612] <= ~layer1_out[8915] | layer1_out[8914];
     layer2_out[4613] <= layer1_out[9056] & layer1_out[9057];
     layer2_out[4614] <= layer1_out[4358] & layer1_out[4359];
     layer2_out[4615] <= layer1_out[6017] & ~layer1_out[6018];
     layer2_out[4616] <= ~layer1_out[4663];
     layer2_out[4617] <= layer1_out[9356];
     layer2_out[4618] <= layer1_out[2301] & ~layer1_out[2302];
     layer2_out[4619] <= ~(layer1_out[10875] | layer1_out[10876]);
     layer2_out[4620] <= ~layer1_out[9790];
     layer2_out[4621] <= layer1_out[43] & ~layer1_out[42];
     layer2_out[4622] <= layer1_out[11236];
     layer2_out[4623] <= layer1_out[5754] & ~layer1_out[5753];
     layer2_out[4624] <= layer1_out[7290] & layer1_out[7291];
     layer2_out[4625] <= layer1_out[10773] & layer1_out[10774];
     layer2_out[4626] <= layer1_out[10965] | layer1_out[10966];
     layer2_out[4627] <= layer1_out[2987];
     layer2_out[4628] <= layer1_out[1245] & ~layer1_out[1246];
     layer2_out[4629] <= ~(layer1_out[596] | layer1_out[597]);
     layer2_out[4630] <= layer1_out[3139] & ~layer1_out[3138];
     layer2_out[4631] <= ~(layer1_out[3722] & layer1_out[3723]);
     layer2_out[4632] <= ~(layer1_out[5926] | layer1_out[5927]);
     layer2_out[4633] <= ~layer1_out[8078];
     layer2_out[4634] <= ~(layer1_out[5581] | layer1_out[5582]);
     layer2_out[4635] <= ~layer1_out[5773] | layer1_out[5772];
     layer2_out[4636] <= layer1_out[6959];
     layer2_out[4637] <= layer1_out[9596];
     layer2_out[4638] <= layer1_out[4942];
     layer2_out[4639] <= layer1_out[1217];
     layer2_out[4640] <= ~layer1_out[7110] | layer1_out[7109];
     layer2_out[4641] <= layer1_out[3775];
     layer2_out[4642] <= layer1_out[304] & ~layer1_out[303];
     layer2_out[4643] <= layer1_out[6890] & layer1_out[6891];
     layer2_out[4644] <= layer1_out[4056];
     layer2_out[4645] <= ~layer1_out[434];
     layer2_out[4646] <= ~(layer1_out[7490] ^ layer1_out[7491]);
     layer2_out[4647] <= layer1_out[7398];
     layer2_out[4648] <= layer1_out[2514];
     layer2_out[4649] <= layer1_out[4744] & layer1_out[4745];
     layer2_out[4650] <= ~layer1_out[1390];
     layer2_out[4651] <= layer1_out[11886] & layer1_out[11887];
     layer2_out[4652] <= ~layer1_out[2165] | layer1_out[2166];
     layer2_out[4653] <= layer1_out[5531] & layer1_out[5532];
     layer2_out[4654] <= layer1_out[6441];
     layer2_out[4655] <= ~layer1_out[4213];
     layer2_out[4656] <= layer1_out[6809] & layer1_out[6810];
     layer2_out[4657] <= ~layer1_out[3633];
     layer2_out[4658] <= ~(layer1_out[1201] ^ layer1_out[1202]);
     layer2_out[4659] <= layer1_out[9843] | layer1_out[9844];
     layer2_out[4660] <= ~(layer1_out[6199] & layer1_out[6200]);
     layer2_out[4661] <= ~layer1_out[2340];
     layer2_out[4662] <= ~layer1_out[9760];
     layer2_out[4663] <= ~(layer1_out[10702] ^ layer1_out[10703]);
     layer2_out[4664] <= layer1_out[5161];
     layer2_out[4665] <= layer1_out[4565] & ~layer1_out[4564];
     layer2_out[4666] <= ~layer1_out[6512];
     layer2_out[4667] <= layer1_out[10785];
     layer2_out[4668] <= layer1_out[8695] & layer1_out[8696];
     layer2_out[4669] <= ~layer1_out[1021];
     layer2_out[4670] <= ~(layer1_out[9303] | layer1_out[9304]);
     layer2_out[4671] <= layer1_out[5219];
     layer2_out[4672] <= ~layer1_out[10047] | layer1_out[10046];
     layer2_out[4673] <= ~layer1_out[294];
     layer2_out[4674] <= layer1_out[8139] & layer1_out[8140];
     layer2_out[4675] <= layer1_out[9917];
     layer2_out[4676] <= layer1_out[5370] ^ layer1_out[5371];
     layer2_out[4677] <= ~layer1_out[1214];
     layer2_out[4678] <= layer1_out[1725] | layer1_out[1726];
     layer2_out[4679] <= ~layer1_out[8414];
     layer2_out[4680] <= ~(layer1_out[11837] | layer1_out[11838]);
     layer2_out[4681] <= 1'b0;
     layer2_out[4682] <= ~(layer1_out[8004] | layer1_out[8005]);
     layer2_out[4683] <= ~layer1_out[1308] | layer1_out[1307];
     layer2_out[4684] <= layer1_out[9537] & ~layer1_out[9536];
     layer2_out[4685] <= layer1_out[5186] & ~layer1_out[5185];
     layer2_out[4686] <= layer1_out[11776] & layer1_out[11777];
     layer2_out[4687] <= layer1_out[578];
     layer2_out[4688] <= ~layer1_out[2013];
     layer2_out[4689] <= ~layer1_out[8137] | layer1_out[8138];
     layer2_out[4690] <= ~layer1_out[3552];
     layer2_out[4691] <= ~layer1_out[5630];
     layer2_out[4692] <= layer1_out[560];
     layer2_out[4693] <= ~layer1_out[4384];
     layer2_out[4694] <= ~(layer1_out[10701] ^ layer1_out[10702]);
     layer2_out[4695] <= ~layer1_out[5397];
     layer2_out[4696] <= layer1_out[6363];
     layer2_out[4697] <= layer1_out[11523] & ~layer1_out[11524];
     layer2_out[4698] <= layer1_out[3338];
     layer2_out[4699] <= ~layer1_out[1681];
     layer2_out[4700] <= ~layer1_out[8380];
     layer2_out[4701] <= ~(layer1_out[10888] & layer1_out[10889]);
     layer2_out[4702] <= 1'b0;
     layer2_out[4703] <= layer1_out[6370];
     layer2_out[4704] <= layer1_out[4178] & ~layer1_out[4179];
     layer2_out[4705] <= ~layer1_out[2011] | layer1_out[2012];
     layer2_out[4706] <= ~(layer1_out[7130] & layer1_out[7131]);
     layer2_out[4707] <= layer1_out[2656] & layer1_out[2657];
     layer2_out[4708] <= layer1_out[2141] ^ layer1_out[2142];
     layer2_out[4709] <= layer1_out[1186];
     layer2_out[4710] <= layer1_out[3709] & layer1_out[3710];
     layer2_out[4711] <= ~layer1_out[7316];
     layer2_out[4712] <= ~(layer1_out[7167] & layer1_out[7168]);
     layer2_out[4713] <= layer1_out[3834] & ~layer1_out[3835];
     layer2_out[4714] <= ~layer1_out[11405] | layer1_out[11404];
     layer2_out[4715] <= layer1_out[7933] & layer1_out[7934];
     layer2_out[4716] <= layer1_out[10914];
     layer2_out[4717] <= layer1_out[11914];
     layer2_out[4718] <= ~layer1_out[9174] | layer1_out[9175];
     layer2_out[4719] <= layer1_out[2635];
     layer2_out[4720] <= layer1_out[190];
     layer2_out[4721] <= layer1_out[684];
     layer2_out[4722] <= layer1_out[8529];
     layer2_out[4723] <= layer1_out[7893] | layer1_out[7894];
     layer2_out[4724] <= layer1_out[515] ^ layer1_out[516];
     layer2_out[4725] <= layer1_out[3674] | layer1_out[3675];
     layer2_out[4726] <= ~(layer1_out[11078] ^ layer1_out[11079]);
     layer2_out[4727] <= ~(layer1_out[10898] & layer1_out[10899]);
     layer2_out[4728] <= layer1_out[345] & layer1_out[346];
     layer2_out[4729] <= ~(layer1_out[3028] & layer1_out[3029]);
     layer2_out[4730] <= layer1_out[6638] & ~layer1_out[6637];
     layer2_out[4731] <= ~layer1_out[5454];
     layer2_out[4732] <= ~layer1_out[7635];
     layer2_out[4733] <= layer1_out[3432];
     layer2_out[4734] <= layer1_out[3238] ^ layer1_out[3239];
     layer2_out[4735] <= layer1_out[8372] & ~layer1_out[8371];
     layer2_out[4736] <= layer1_out[7873] ^ layer1_out[7874];
     layer2_out[4737] <= ~layer1_out[1518] | layer1_out[1519];
     layer2_out[4738] <= ~layer1_out[350];
     layer2_out[4739] <= ~layer1_out[7470] | layer1_out[7471];
     layer2_out[4740] <= ~layer1_out[459] | layer1_out[458];
     layer2_out[4741] <= ~(layer1_out[11327] | layer1_out[11328]);
     layer2_out[4742] <= ~(layer1_out[287] ^ layer1_out[288]);
     layer2_out[4743] <= ~layer1_out[6155];
     layer2_out[4744] <= ~(layer1_out[8427] ^ layer1_out[8428]);
     layer2_out[4745] <= layer1_out[8492];
     layer2_out[4746] <= ~(layer1_out[11634] ^ layer1_out[11635]);
     layer2_out[4747] <= ~layer1_out[10096];
     layer2_out[4748] <= layer1_out[5030] & ~layer1_out[5029];
     layer2_out[4749] <= layer1_out[2333] & layer1_out[2334];
     layer2_out[4750] <= layer1_out[5917];
     layer2_out[4751] <= layer1_out[5082] & ~layer1_out[5083];
     layer2_out[4752] <= ~(layer1_out[1224] ^ layer1_out[1225]);
     layer2_out[4753] <= ~layer1_out[5497];
     layer2_out[4754] <= ~layer1_out[3661];
     layer2_out[4755] <= layer1_out[8478] & ~layer1_out[8477];
     layer2_out[4756] <= layer1_out[4082] & ~layer1_out[4083];
     layer2_out[4757] <= ~(layer1_out[3642] | layer1_out[3643]);
     layer2_out[4758] <= layer1_out[10544] & layer1_out[10545];
     layer2_out[4759] <= ~(layer1_out[1954] | layer1_out[1955]);
     layer2_out[4760] <= layer1_out[10949] & ~layer1_out[10948];
     layer2_out[4761] <= ~(layer1_out[5065] ^ layer1_out[5066]);
     layer2_out[4762] <= ~layer1_out[3880];
     layer2_out[4763] <= layer1_out[10063] & ~layer1_out[10064];
     layer2_out[4764] <= layer1_out[89] & ~layer1_out[90];
     layer2_out[4765] <= layer1_out[9948] | layer1_out[9949];
     layer2_out[4766] <= layer1_out[8311];
     layer2_out[4767] <= layer1_out[2910] | layer1_out[2911];
     layer2_out[4768] <= ~layer1_out[4305];
     layer2_out[4769] <= ~layer1_out[9249] | layer1_out[9250];
     layer2_out[4770] <= ~layer1_out[11595] | layer1_out[11594];
     layer2_out[4771] <= ~(layer1_out[1642] ^ layer1_out[1643]);
     layer2_out[4772] <= ~(layer1_out[6133] & layer1_out[6134]);
     layer2_out[4773] <= ~(layer1_out[8586] ^ layer1_out[8587]);
     layer2_out[4774] <= layer1_out[7443] & layer1_out[7444];
     layer2_out[4775] <= layer1_out[596];
     layer2_out[4776] <= layer1_out[6982] & layer1_out[6983];
     layer2_out[4777] <= ~(layer1_out[6140] | layer1_out[6141]);
     layer2_out[4778] <= 1'b0;
     layer2_out[4779] <= ~layer1_out[4150];
     layer2_out[4780] <= ~layer1_out[9905];
     layer2_out[4781] <= ~layer1_out[480];
     layer2_out[4782] <= layer1_out[3634] & layer1_out[3635];
     layer2_out[4783] <= ~layer1_out[4010] | layer1_out[4009];
     layer2_out[4784] <= layer1_out[348];
     layer2_out[4785] <= ~(layer1_out[5194] & layer1_out[5195]);
     layer2_out[4786] <= layer1_out[1323] | layer1_out[1324];
     layer2_out[4787] <= layer1_out[6277];
     layer2_out[4788] <= layer1_out[8973];
     layer2_out[4789] <= layer1_out[11694] & layer1_out[11695];
     layer2_out[4790] <= ~(layer1_out[8204] | layer1_out[8205]);
     layer2_out[4791] <= layer1_out[803];
     layer2_out[4792] <= layer1_out[3187] & ~layer1_out[3186];
     layer2_out[4793] <= layer1_out[5827];
     layer2_out[4794] <= layer1_out[7838] ^ layer1_out[7839];
     layer2_out[4795] <= layer1_out[108] & ~layer1_out[109];
     layer2_out[4796] <= ~(layer1_out[5322] | layer1_out[5323]);
     layer2_out[4797] <= layer1_out[11753] & ~layer1_out[11754];
     layer2_out[4798] <= layer1_out[9911];
     layer2_out[4799] <= ~layer1_out[3626] | layer1_out[3625];
     layer2_out[4800] <= ~(layer1_out[282] & layer1_out[283]);
     layer2_out[4801] <= layer1_out[10299];
     layer2_out[4802] <= ~(layer1_out[4208] | layer1_out[4209]);
     layer2_out[4803] <= ~layer1_out[8594];
     layer2_out[4804] <= ~(layer1_out[4780] | layer1_out[4781]);
     layer2_out[4805] <= ~layer1_out[4415];
     layer2_out[4806] <= layer1_out[6867];
     layer2_out[4807] <= layer1_out[11466] & layer1_out[11467];
     layer2_out[4808] <= ~(layer1_out[4759] ^ layer1_out[4760]);
     layer2_out[4809] <= ~layer1_out[5501];
     layer2_out[4810] <= ~(layer1_out[10379] ^ layer1_out[10380]);
     layer2_out[4811] <= layer1_out[9] & ~layer1_out[8];
     layer2_out[4812] <= ~layer1_out[11998];
     layer2_out[4813] <= layer1_out[1089];
     layer2_out[4814] <= ~(layer1_out[7959] & layer1_out[7960]);
     layer2_out[4815] <= layer1_out[9557];
     layer2_out[4816] <= ~layer1_out[6538];
     layer2_out[4817] <= layer1_out[2084] & layer1_out[2085];
     layer2_out[4818] <= ~layer1_out[6680] | layer1_out[6681];
     layer2_out[4819] <= ~(layer1_out[7449] ^ layer1_out[7450]);
     layer2_out[4820] <= ~layer1_out[6038];
     layer2_out[4821] <= layer1_out[198] & ~layer1_out[197];
     layer2_out[4822] <= ~layer1_out[9309] | layer1_out[9310];
     layer2_out[4823] <= ~(layer1_out[6114] | layer1_out[6115]);
     layer2_out[4824] <= ~layer1_out[3697] | layer1_out[3698];
     layer2_out[4825] <= layer1_out[5272] | layer1_out[5273];
     layer2_out[4826] <= layer1_out[469] ^ layer1_out[470];
     layer2_out[4827] <= layer1_out[734];
     layer2_out[4828] <= layer1_out[8674];
     layer2_out[4829] <= layer1_out[8463] & layer1_out[8464];
     layer2_out[4830] <= layer1_out[424] & ~layer1_out[423];
     layer2_out[4831] <= layer1_out[4217] & ~layer1_out[4218];
     layer2_out[4832] <= ~(layer1_out[3958] & layer1_out[3959]);
     layer2_out[4833] <= layer1_out[8125] ^ layer1_out[8126];
     layer2_out[4834] <= ~layer1_out[5364] | layer1_out[5363];
     layer2_out[4835] <= ~(layer1_out[11376] | layer1_out[11377]);
     layer2_out[4836] <= layer1_out[8269] & layer1_out[8270];
     layer2_out[4837] <= ~layer1_out[2626];
     layer2_out[4838] <= layer1_out[811] & ~layer1_out[810];
     layer2_out[4839] <= layer1_out[5004];
     layer2_out[4840] <= layer1_out[8759] | layer1_out[8760];
     layer2_out[4841] <= ~layer1_out[2884];
     layer2_out[4842] <= layer1_out[1994];
     layer2_out[4843] <= layer1_out[7829];
     layer2_out[4844] <= ~layer1_out[6874];
     layer2_out[4845] <= layer1_out[1206] & ~layer1_out[1205];
     layer2_out[4846] <= ~(layer1_out[10460] ^ layer1_out[10461]);
     layer2_out[4847] <= layer1_out[1942] | layer1_out[1943];
     layer2_out[4848] <= ~(layer1_out[5613] ^ layer1_out[5614]);
     layer2_out[4849] <= ~(layer1_out[1832] | layer1_out[1833]);
     layer2_out[4850] <= layer1_out[4188];
     layer2_out[4851] <= ~(layer1_out[7492] | layer1_out[7493]);
     layer2_out[4852] <= ~layer1_out[5812];
     layer2_out[4853] <= layer1_out[4049] & ~layer1_out[4048];
     layer2_out[4854] <= ~(layer1_out[1490] | layer1_out[1491]);
     layer2_out[4855] <= ~(layer1_out[7244] & layer1_out[7245]);
     layer2_out[4856] <= ~(layer1_out[5461] | layer1_out[5462]);
     layer2_out[4857] <= layer1_out[7942] ^ layer1_out[7943];
     layer2_out[4858] <= ~layer1_out[5585];
     layer2_out[4859] <= layer1_out[11957];
     layer2_out[4860] <= layer1_out[2459] ^ layer1_out[2460];
     layer2_out[4861] <= ~layer1_out[9162] | layer1_out[9163];
     layer2_out[4862] <= ~(layer1_out[2377] & layer1_out[2378]);
     layer2_out[4863] <= ~layer1_out[8542];
     layer2_out[4864] <= ~layer1_out[8874];
     layer2_out[4865] <= layer1_out[11360] ^ layer1_out[11361];
     layer2_out[4866] <= ~layer1_out[8416];
     layer2_out[4867] <= ~(layer1_out[7849] & layer1_out[7850]);
     layer2_out[4868] <= layer1_out[74];
     layer2_out[4869] <= ~layer1_out[11810] | layer1_out[11811];
     layer2_out[4870] <= ~(layer1_out[11005] & layer1_out[11006]);
     layer2_out[4871] <= layer1_out[3605];
     layer2_out[4872] <= layer1_out[2720] | layer1_out[2721];
     layer2_out[4873] <= layer1_out[11123];
     layer2_out[4874] <= layer1_out[8799] | layer1_out[8800];
     layer2_out[4875] <= ~layer1_out[2569];
     layer2_out[4876] <= layer1_out[7483] | layer1_out[7484];
     layer2_out[4877] <= ~(layer1_out[4818] | layer1_out[4819]);
     layer2_out[4878] <= layer1_out[3543];
     layer2_out[4879] <= ~(layer1_out[11187] & layer1_out[11188]);
     layer2_out[4880] <= ~layer1_out[2191];
     layer2_out[4881] <= layer1_out[3905] & layer1_out[3906];
     layer2_out[4882] <= ~layer1_out[3785];
     layer2_out[4883] <= ~layer1_out[375];
     layer2_out[4884] <= ~layer1_out[7372];
     layer2_out[4885] <= ~layer1_out[2068] | layer1_out[2069];
     layer2_out[4886] <= ~layer1_out[3215];
     layer2_out[4887] <= layer1_out[9653];
     layer2_out[4888] <= ~(layer1_out[7638] | layer1_out[7639]);
     layer2_out[4889] <= layer1_out[7631];
     layer2_out[4890] <= ~layer1_out[8462] | layer1_out[8463];
     layer2_out[4891] <= layer1_out[8169] & layer1_out[8170];
     layer2_out[4892] <= ~(layer1_out[8258] & layer1_out[8259]);
     layer2_out[4893] <= layer1_out[8862] & layer1_out[8863];
     layer2_out[4894] <= ~(layer1_out[2179] | layer1_out[2180]);
     layer2_out[4895] <= ~(layer1_out[4787] & layer1_out[4788]);
     layer2_out[4896] <= ~(layer1_out[583] | layer1_out[584]);
     layer2_out[4897] <= ~layer1_out[10617];
     layer2_out[4898] <= layer1_out[10308];
     layer2_out[4899] <= ~layer1_out[2132] | layer1_out[2133];
     layer2_out[4900] <= layer1_out[5963];
     layer2_out[4901] <= ~layer1_out[5397];
     layer2_out[4902] <= ~(layer1_out[11009] ^ layer1_out[11010]);
     layer2_out[4903] <= layer1_out[2175] | layer1_out[2176];
     layer2_out[4904] <= ~layer1_out[10955];
     layer2_out[4905] <= layer1_out[11873] & ~layer1_out[11874];
     layer2_out[4906] <= layer1_out[8788] | layer1_out[8789];
     layer2_out[4907] <= ~(layer1_out[5662] ^ layer1_out[5663]);
     layer2_out[4908] <= ~layer1_out[2401];
     layer2_out[4909] <= layer1_out[1210] | layer1_out[1211];
     layer2_out[4910] <= layer1_out[11602];
     layer2_out[4911] <= ~layer1_out[3946];
     layer2_out[4912] <= ~(layer1_out[7648] & layer1_out[7649]);
     layer2_out[4913] <= ~layer1_out[8419] | layer1_out[8418];
     layer2_out[4914] <= layer1_out[7737] | layer1_out[7738];
     layer2_out[4915] <= layer1_out[8493];
     layer2_out[4916] <= ~layer1_out[8071];
     layer2_out[4917] <= layer1_out[2615] | layer1_out[2616];
     layer2_out[4918] <= ~(layer1_out[4008] | layer1_out[4009]);
     layer2_out[4919] <= 1'b1;
     layer2_out[4920] <= ~layer1_out[1235];
     layer2_out[4921] <= ~layer1_out[6146];
     layer2_out[4922] <= ~layer1_out[3438] | layer1_out[3439];
     layer2_out[4923] <= layer1_out[4324] & layer1_out[4325];
     layer2_out[4924] <= layer1_out[9587] & ~layer1_out[9588];
     layer2_out[4925] <= ~layer1_out[9229];
     layer2_out[4926] <= layer1_out[1100] & layer1_out[1101];
     layer2_out[4927] <= layer1_out[8327];
     layer2_out[4928] <= layer1_out[2004];
     layer2_out[4929] <= layer1_out[2915] ^ layer1_out[2916];
     layer2_out[4930] <= layer1_out[1998];
     layer2_out[4931] <= ~layer1_out[11409] | layer1_out[11410];
     layer2_out[4932] <= ~layer1_out[7126];
     layer2_out[4933] <= layer1_out[5306] | layer1_out[5307];
     layer2_out[4934] <= ~layer1_out[506];
     layer2_out[4935] <= layer1_out[7206] & layer1_out[7207];
     layer2_out[4936] <= layer1_out[10893] | layer1_out[10894];
     layer2_out[4937] <= layer1_out[5250] & layer1_out[5251];
     layer2_out[4938] <= ~layer1_out[11446] | layer1_out[11445];
     layer2_out[4939] <= ~(layer1_out[8663] ^ layer1_out[8664]);
     layer2_out[4940] <= ~(layer1_out[7478] & layer1_out[7479]);
     layer2_out[4941] <= ~(layer1_out[390] ^ layer1_out[391]);
     layer2_out[4942] <= ~layer1_out[7022];
     layer2_out[4943] <= ~layer1_out[5370];
     layer2_out[4944] <= ~layer1_out[3193];
     layer2_out[4945] <= ~layer1_out[9378] | layer1_out[9379];
     layer2_out[4946] <= layer1_out[7489];
     layer2_out[4947] <= ~(layer1_out[8596] ^ layer1_out[8597]);
     layer2_out[4948] <= layer1_out[3101] & ~layer1_out[3100];
     layer2_out[4949] <= ~layer1_out[6979] | layer1_out[6978];
     layer2_out[4950] <= layer1_out[5900];
     layer2_out[4951] <= layer1_out[8655];
     layer2_out[4952] <= layer1_out[5758] | layer1_out[5759];
     layer2_out[4953] <= ~layer1_out[807] | layer1_out[806];
     layer2_out[4954] <= layer1_out[10306] & ~layer1_out[10307];
     layer2_out[4955] <= ~(layer1_out[6350] & layer1_out[6351]);
     layer2_out[4956] <= ~layer1_out[6305];
     layer2_out[4957] <= ~(layer1_out[1115] ^ layer1_out[1116]);
     layer2_out[4958] <= layer1_out[5353] ^ layer1_out[5354];
     layer2_out[4959] <= layer1_out[692];
     layer2_out[4960] <= ~(layer1_out[9909] | layer1_out[9910]);
     layer2_out[4961] <= ~(layer1_out[4041] & layer1_out[4042]);
     layer2_out[4962] <= ~layer1_out[8287];
     layer2_out[4963] <= ~layer1_out[9712];
     layer2_out[4964] <= ~layer1_out[9663];
     layer2_out[4965] <= layer1_out[1626];
     layer2_out[4966] <= layer1_out[11719] & ~layer1_out[11720];
     layer2_out[4967] <= ~layer1_out[9291] | layer1_out[9290];
     layer2_out[4968] <= layer1_out[249];
     layer2_out[4969] <= layer1_out[8605];
     layer2_out[4970] <= ~(layer1_out[4137] & layer1_out[4138]);
     layer2_out[4971] <= layer1_out[1355] ^ layer1_out[1356];
     layer2_out[4972] <= ~layer1_out[7957];
     layer2_out[4973] <= ~(layer1_out[10264] & layer1_out[10265]);
     layer2_out[4974] <= layer1_out[11735] & ~layer1_out[11736];
     layer2_out[4975] <= ~layer1_out[1550];
     layer2_out[4976] <= layer1_out[1053];
     layer2_out[4977] <= ~layer1_out[6234] | layer1_out[6233];
     layer2_out[4978] <= layer1_out[10967] ^ layer1_out[10968];
     layer2_out[4979] <= layer1_out[2519] & ~layer1_out[2520];
     layer2_out[4980] <= layer1_out[4591];
     layer2_out[4981] <= ~(layer1_out[2712] | layer1_out[2713]);
     layer2_out[4982] <= layer1_out[9762] & layer1_out[9763];
     layer2_out[4983] <= layer1_out[7857] ^ layer1_out[7858];
     layer2_out[4984] <= layer1_out[3948] & ~layer1_out[3949];
     layer2_out[4985] <= ~(layer1_out[4956] | layer1_out[4957]);
     layer2_out[4986] <= layer1_out[11435] & layer1_out[11436];
     layer2_out[4987] <= ~(layer1_out[1298] | layer1_out[1299]);
     layer2_out[4988] <= ~(layer1_out[11702] & layer1_out[11703]);
     layer2_out[4989] <= layer1_out[1281];
     layer2_out[4990] <= layer1_out[1333];
     layer2_out[4991] <= layer1_out[3967] & ~layer1_out[3966];
     layer2_out[4992] <= ~layer1_out[9208];
     layer2_out[4993] <= layer1_out[9167] | layer1_out[9168];
     layer2_out[4994] <= layer1_out[9340] & ~layer1_out[9339];
     layer2_out[4995] <= ~(layer1_out[5795] | layer1_out[5796]);
     layer2_out[4996] <= ~layer1_out[11943];
     layer2_out[4997] <= ~layer1_out[4725];
     layer2_out[4998] <= ~layer1_out[5027] | layer1_out[5026];
     layer2_out[4999] <= ~layer1_out[228] | layer1_out[227];
     layer2_out[5000] <= ~(layer1_out[1474] ^ layer1_out[1475]);
     layer2_out[5001] <= layer1_out[2468];
     layer2_out[5002] <= layer1_out[10796] & ~layer1_out[10797];
     layer2_out[5003] <= ~(layer1_out[7047] | layer1_out[7048]);
     layer2_out[5004] <= 1'b0;
     layer2_out[5005] <= layer1_out[11690];
     layer2_out[5006] <= layer1_out[5422] ^ layer1_out[5423];
     layer2_out[5007] <= ~layer1_out[2887];
     layer2_out[5008] <= layer1_out[5860];
     layer2_out[5009] <= layer1_out[5831] | layer1_out[5832];
     layer2_out[5010] <= ~layer1_out[2679] | layer1_out[2678];
     layer2_out[5011] <= ~(layer1_out[7131] ^ layer1_out[7132]);
     layer2_out[5012] <= ~layer1_out[8314] | layer1_out[8313];
     layer2_out[5013] <= ~layer1_out[8183];
     layer2_out[5014] <= ~(layer1_out[5970] | layer1_out[5971]);
     layer2_out[5015] <= ~layer1_out[10034] | layer1_out[10033];
     layer2_out[5016] <= layer1_out[5641];
     layer2_out[5017] <= layer1_out[2337] & ~layer1_out[2338];
     layer2_out[5018] <= ~(layer1_out[3315] ^ layer1_out[3316]);
     layer2_out[5019] <= layer1_out[4914] & ~layer1_out[4915];
     layer2_out[5020] <= layer1_out[7446];
     layer2_out[5021] <= ~(layer1_out[5219] & layer1_out[5220]);
     layer2_out[5022] <= ~layer1_out[4963];
     layer2_out[5023] <= ~(layer1_out[1911] | layer1_out[1912]);
     layer2_out[5024] <= ~layer1_out[8708];
     layer2_out[5025] <= layer1_out[7523];
     layer2_out[5026] <= ~(layer1_out[8950] | layer1_out[8951]);
     layer2_out[5027] <= ~layer1_out[4446];
     layer2_out[5028] <= layer1_out[8563] & ~layer1_out[8564];
     layer2_out[5029] <= ~(layer1_out[10185] & layer1_out[10186]);
     layer2_out[5030] <= layer1_out[4976] & layer1_out[4977];
     layer2_out[5031] <= layer1_out[10461];
     layer2_out[5032] <= ~layer1_out[55];
     layer2_out[5033] <= layer1_out[1829] & ~layer1_out[1828];
     layer2_out[5034] <= ~layer1_out[2021] | layer1_out[2022];
     layer2_out[5035] <= ~layer1_out[7641];
     layer2_out[5036] <= layer1_out[5230];
     layer2_out[5037] <= layer1_out[2195] ^ layer1_out[2196];
     layer2_out[5038] <= layer1_out[7503];
     layer2_out[5039] <= ~(layer1_out[11934] & layer1_out[11935]);
     layer2_out[5040] <= ~layer1_out[1303] | layer1_out[1302];
     layer2_out[5041] <= ~layer1_out[5045] | layer1_out[5044];
     layer2_out[5042] <= ~layer1_out[6217];
     layer2_out[5043] <= layer1_out[4615];
     layer2_out[5044] <= layer1_out[9721] | layer1_out[9722];
     layer2_out[5045] <= ~(layer1_out[5874] & layer1_out[5875]);
     layer2_out[5046] <= ~(layer1_out[3078] | layer1_out[3079]);
     layer2_out[5047] <= ~(layer1_out[877] | layer1_out[878]);
     layer2_out[5048] <= layer1_out[2336];
     layer2_out[5049] <= layer1_out[765] | layer1_out[766];
     layer2_out[5050] <= layer1_out[2605] & ~layer1_out[2606];
     layer2_out[5051] <= layer1_out[8712] ^ layer1_out[8713];
     layer2_out[5052] <= ~layer1_out[11188];
     layer2_out[5053] <= layer1_out[3119];
     layer2_out[5054] <= ~(layer1_out[6887] ^ layer1_out[6888]);
     layer2_out[5055] <= ~(layer1_out[5854] & layer1_out[5855]);
     layer2_out[5056] <= layer1_out[10911] ^ layer1_out[10912];
     layer2_out[5057] <= layer1_out[462] & ~layer1_out[463];
     layer2_out[5058] <= layer1_out[11045];
     layer2_out[5059] <= layer1_out[6999];
     layer2_out[5060] <= layer1_out[2253];
     layer2_out[5061] <= ~layer1_out[5389];
     layer2_out[5062] <= 1'b1;
     layer2_out[5063] <= ~(layer1_out[6618] | layer1_out[6619]);
     layer2_out[5064] <= layer1_out[5150] & ~layer1_out[5151];
     layer2_out[5065] <= ~layer1_out[8106];
     layer2_out[5066] <= ~layer1_out[3894] | layer1_out[3895];
     layer2_out[5067] <= layer1_out[2284] | layer1_out[2285];
     layer2_out[5068] <= ~layer1_out[3671];
     layer2_out[5069] <= ~layer1_out[9684];
     layer2_out[5070] <= ~(layer1_out[7644] | layer1_out[7645]);
     layer2_out[5071] <= ~layer1_out[2161] | layer1_out[2160];
     layer2_out[5072] <= ~layer1_out[4280];
     layer2_out[5073] <= layer1_out[10425];
     layer2_out[5074] <= ~layer1_out[365];
     layer2_out[5075] <= layer1_out[7860];
     layer2_out[5076] <= layer1_out[4479] & layer1_out[4480];
     layer2_out[5077] <= ~(layer1_out[2838] | layer1_out[2839]);
     layer2_out[5078] <= layer1_out[3340] & layer1_out[3341];
     layer2_out[5079] <= ~(layer1_out[497] | layer1_out[498]);
     layer2_out[5080] <= layer1_out[11963] & ~layer1_out[11962];
     layer2_out[5081] <= ~layer1_out[6502];
     layer2_out[5082] <= layer1_out[10245] ^ layer1_out[10246];
     layer2_out[5083] <= layer1_out[6323] | layer1_out[6324];
     layer2_out[5084] <= ~layer1_out[6051];
     layer2_out[5085] <= ~(layer1_out[5793] | layer1_out[5794]);
     layer2_out[5086] <= ~(layer1_out[11988] ^ layer1_out[11989]);
     layer2_out[5087] <= layer1_out[8649] & layer1_out[8650];
     layer2_out[5088] <= ~layer1_out[1757];
     layer2_out[5089] <= ~layer1_out[8012] | layer1_out[8013];
     layer2_out[5090] <= ~layer1_out[5349];
     layer2_out[5091] <= layer1_out[4692];
     layer2_out[5092] <= layer1_out[3580] ^ layer1_out[3581];
     layer2_out[5093] <= ~layer1_out[4903];
     layer2_out[5094] <= layer1_out[1526];
     layer2_out[5095] <= layer1_out[10152];
     layer2_out[5096] <= ~layer1_out[4221];
     layer2_out[5097] <= ~layer1_out[5321];
     layer2_out[5098] <= layer1_out[7879];
     layer2_out[5099] <= layer1_out[822] & ~layer1_out[821];
     layer2_out[5100] <= ~(layer1_out[4299] | layer1_out[4300]);
     layer2_out[5101] <= ~(layer1_out[531] & layer1_out[532]);
     layer2_out[5102] <= layer1_out[7090] ^ layer1_out[7091];
     layer2_out[5103] <= 1'b0;
     layer2_out[5104] <= layer1_out[10500] ^ layer1_out[10501];
     layer2_out[5105] <= ~(layer1_out[1083] & layer1_out[1084]);
     layer2_out[5106] <= layer1_out[2922] & ~layer1_out[2921];
     layer2_out[5107] <= ~layer1_out[10800];
     layer2_out[5108] <= ~layer1_out[3032];
     layer2_out[5109] <= layer1_out[5932] & layer1_out[5933];
     layer2_out[5110] <= ~layer1_out[4894];
     layer2_out[5111] <= layer1_out[10549];
     layer2_out[5112] <= ~layer1_out[68] | layer1_out[69];
     layer2_out[5113] <= ~layer1_out[4212];
     layer2_out[5114] <= layer1_out[10677];
     layer2_out[5115] <= 1'b1;
     layer2_out[5116] <= ~(layer1_out[10354] & layer1_out[10355]);
     layer2_out[5117] <= 1'b0;
     layer2_out[5118] <= ~layer1_out[11439] | layer1_out[11438];
     layer2_out[5119] <= ~(layer1_out[7128] & layer1_out[7129]);
     layer2_out[5120] <= layer1_out[2659] | layer1_out[2660];
     layer2_out[5121] <= layer1_out[6994];
     layer2_out[5122] <= ~(layer1_out[9535] | layer1_out[9536]);
     layer2_out[5123] <= ~(layer1_out[6586] | layer1_out[6587]);
     layer2_out[5124] <= layer1_out[3374];
     layer2_out[5125] <= layer1_out[6850] & ~layer1_out[6849];
     layer2_out[5126] <= ~(layer1_out[5303] ^ layer1_out[5304]);
     layer2_out[5127] <= layer1_out[2699] & layer1_out[2700];
     layer2_out[5128] <= ~layer1_out[2219] | layer1_out[2220];
     layer2_out[5129] <= layer1_out[11493];
     layer2_out[5130] <= layer1_out[1651] & layer1_out[1652];
     layer2_out[5131] <= layer1_out[586] | layer1_out[587];
     layer2_out[5132] <= ~layer1_out[583];
     layer2_out[5133] <= layer1_out[4607];
     layer2_out[5134] <= ~layer1_out[9138] | layer1_out[9137];
     layer2_out[5135] <= layer1_out[6081] & ~layer1_out[6082];
     layer2_out[5136] <= ~layer1_out[7402];
     layer2_out[5137] <= layer1_out[4874] & ~layer1_out[4875];
     layer2_out[5138] <= layer1_out[179] & layer1_out[180];
     layer2_out[5139] <= layer1_out[1933];
     layer2_out[5140] <= ~(layer1_out[4038] | layer1_out[4039]);
     layer2_out[5141] <= layer1_out[9453] | layer1_out[9454];
     layer2_out[5142] <= layer1_out[10531] & ~layer1_out[10532];
     layer2_out[5143] <= ~(layer1_out[10899] & layer1_out[10900]);
     layer2_out[5144] <= ~layer1_out[7277] | layer1_out[7278];
     layer2_out[5145] <= ~(layer1_out[11682] & layer1_out[11683]);
     layer2_out[5146] <= layer1_out[1184] & ~layer1_out[1185];
     layer2_out[5147] <= ~layer1_out[1462] | layer1_out[1463];
     layer2_out[5148] <= layer1_out[8013] | layer1_out[8014];
     layer2_out[5149] <= ~(layer1_out[10956] ^ layer1_out[10957]);
     layer2_out[5150] <= layer1_out[8983] & layer1_out[8984];
     layer2_out[5151] <= layer1_out[6440] & layer1_out[6441];
     layer2_out[5152] <= layer1_out[9878] ^ layer1_out[9879];
     layer2_out[5153] <= ~(layer1_out[7569] & layer1_out[7570]);
     layer2_out[5154] <= ~layer1_out[4992];
     layer2_out[5155] <= layer1_out[1694];
     layer2_out[5156] <= ~(layer1_out[1325] ^ layer1_out[1326]);
     layer2_out[5157] <= ~(layer1_out[4262] & layer1_out[4263]);
     layer2_out[5158] <= layer1_out[5022] & ~layer1_out[5023];
     layer2_out[5159] <= layer1_out[265];
     layer2_out[5160] <= ~layer1_out[781];
     layer2_out[5161] <= layer1_out[8401];
     layer2_out[5162] <= ~(layer1_out[11202] | layer1_out[11203]);
     layer2_out[5163] <= ~(layer1_out[6854] | layer1_out[6855]);
     layer2_out[5164] <= ~layer1_out[10833] | layer1_out[10832];
     layer2_out[5165] <= ~(layer1_out[3261] & layer1_out[3262]);
     layer2_out[5166] <= layer1_out[9505];
     layer2_out[5167] <= 1'b1;
     layer2_out[5168] <= ~(layer1_out[11724] ^ layer1_out[11725]);
     layer2_out[5169] <= layer1_out[3962];
     layer2_out[5170] <= layer1_out[5114];
     layer2_out[5171] <= ~(layer1_out[322] | layer1_out[323]);
     layer2_out[5172] <= ~layer1_out[10909] | layer1_out[10908];
     layer2_out[5173] <= layer1_out[8356];
     layer2_out[5174] <= layer1_out[542];
     layer2_out[5175] <= 1'b1;
     layer2_out[5176] <= layer1_out[8490];
     layer2_out[5177] <= layer1_out[4783] & ~layer1_out[4782];
     layer2_out[5178] <= layer1_out[3811] & ~layer1_out[3810];
     layer2_out[5179] <= ~layer1_out[9574] | layer1_out[9573];
     layer2_out[5180] <= layer1_out[5238] & ~layer1_out[5237];
     layer2_out[5181] <= layer1_out[487] & layer1_out[488];
     layer2_out[5182] <= layer1_out[8514];
     layer2_out[5183] <= ~layer1_out[6820];
     layer2_out[5184] <= ~layer1_out[2498];
     layer2_out[5185] <= ~layer1_out[10808];
     layer2_out[5186] <= layer1_out[11061] | layer1_out[11062];
     layer2_out[5187] <= layer1_out[3738] & layer1_out[3739];
     layer2_out[5188] <= ~layer1_out[2645] | layer1_out[2646];
     layer2_out[5189] <= layer1_out[5501];
     layer2_out[5190] <= layer1_out[3927];
     layer2_out[5191] <= layer1_out[11225];
     layer2_out[5192] <= ~layer1_out[292];
     layer2_out[5193] <= ~layer1_out[8704] | layer1_out[8705];
     layer2_out[5194] <= layer1_out[7827] | layer1_out[7828];
     layer2_out[5195] <= ~layer1_out[4837];
     layer2_out[5196] <= layer1_out[11448] | layer1_out[11449];
     layer2_out[5197] <= ~(layer1_out[3611] & layer1_out[3612]);
     layer2_out[5198] <= layer1_out[1678] & layer1_out[1679];
     layer2_out[5199] <= layer1_out[4568] ^ layer1_out[4569];
     layer2_out[5200] <= ~layer1_out[2221] | layer1_out[2222];
     layer2_out[5201] <= ~(layer1_out[11716] & layer1_out[11717]);
     layer2_out[5202] <= ~layer1_out[6734];
     layer2_out[5203] <= layer1_out[462];
     layer2_out[5204] <= layer1_out[9927] & ~layer1_out[9928];
     layer2_out[5205] <= ~layer1_out[389];
     layer2_out[5206] <= layer1_out[10160];
     layer2_out[5207] <= ~layer1_out[2829] | layer1_out[2830];
     layer2_out[5208] <= layer1_out[9287] | layer1_out[9288];
     layer2_out[5209] <= ~layer1_out[250] | layer1_out[251];
     layer2_out[5210] <= layer1_out[2948] ^ layer1_out[2949];
     layer2_out[5211] <= 1'b1;
     layer2_out[5212] <= ~layer1_out[6404];
     layer2_out[5213] <= layer1_out[2303] & ~layer1_out[2304];
     layer2_out[5214] <= ~layer1_out[7502] | layer1_out[7501];
     layer2_out[5215] <= ~(layer1_out[8908] ^ layer1_out[8909]);
     layer2_out[5216] <= layer1_out[9483] | layer1_out[9484];
     layer2_out[5217] <= layer1_out[2550];
     layer2_out[5218] <= ~layer1_out[932] | layer1_out[933];
     layer2_out[5219] <= ~layer1_out[11552] | layer1_out[11553];
     layer2_out[5220] <= layer1_out[3656] & ~layer1_out[3657];
     layer2_out[5221] <= ~layer1_out[11991] | layer1_out[11990];
     layer2_out[5222] <= layer1_out[9642];
     layer2_out[5223] <= ~layer1_out[9039];
     layer2_out[5224] <= ~layer1_out[8910] | layer1_out[8909];
     layer2_out[5225] <= ~layer1_out[7351];
     layer2_out[5226] <= ~layer1_out[10472];
     layer2_out[5227] <= ~layer1_out[7756] | layer1_out[7757];
     layer2_out[5228] <= ~layer1_out[11727] | layer1_out[11726];
     layer2_out[5229] <= 1'b0;
     layer2_out[5230] <= ~layer1_out[2953];
     layer2_out[5231] <= layer1_out[9574] | layer1_out[9575];
     layer2_out[5232] <= ~layer1_out[7495];
     layer2_out[5233] <= ~layer1_out[4219] | layer1_out[4218];
     layer2_out[5234] <= ~layer1_out[11103];
     layer2_out[5235] <= layer1_out[2938] ^ layer1_out[2939];
     layer2_out[5236] <= layer1_out[752];
     layer2_out[5237] <= ~(layer1_out[7771] | layer1_out[7772]);
     layer2_out[5238] <= layer1_out[4859];
     layer2_out[5239] <= ~(layer1_out[11553] | layer1_out[11554]);
     layer2_out[5240] <= layer1_out[4584] & ~layer1_out[4583];
     layer2_out[5241] <= layer1_out[4722] | layer1_out[4723];
     layer2_out[5242] <= layer1_out[6587] | layer1_out[6588];
     layer2_out[5243] <= ~(layer1_out[6122] & layer1_out[6123]);
     layer2_out[5244] <= layer1_out[9576];
     layer2_out[5245] <= ~layer1_out[6077];
     layer2_out[5246] <= ~(layer1_out[2235] & layer1_out[2236]);
     layer2_out[5247] <= ~layer1_out[11555] | layer1_out[11556];
     layer2_out[5248] <= ~layer1_out[11808];
     layer2_out[5249] <= ~(layer1_out[6377] | layer1_out[6378]);
     layer2_out[5250] <= ~(layer1_out[2708] | layer1_out[2709]);
     layer2_out[5251] <= ~layer1_out[6805] | layer1_out[6806];
     layer2_out[5252] <= ~(layer1_out[6222] | layer1_out[6223]);
     layer2_out[5253] <= ~layer1_out[2590] | layer1_out[2591];
     layer2_out[5254] <= layer1_out[1414] & layer1_out[1415];
     layer2_out[5255] <= ~layer1_out[7384];
     layer2_out[5256] <= layer1_out[833] & ~layer1_out[832];
     layer2_out[5257] <= ~(layer1_out[11538] & layer1_out[11539]);
     layer2_out[5258] <= layer1_out[10421] | layer1_out[10422];
     layer2_out[5259] <= ~(layer1_out[9697] & layer1_out[9698]);
     layer2_out[5260] <= 1'b1;
     layer2_out[5261] <= layer1_out[5853];
     layer2_out[5262] <= ~layer1_out[2691];
     layer2_out[5263] <= ~layer1_out[209] | layer1_out[208];
     layer2_out[5264] <= ~layer1_out[6857] | layer1_out[6858];
     layer2_out[5265] <= ~layer1_out[3162] | layer1_out[3163];
     layer2_out[5266] <= ~layer1_out[9724];
     layer2_out[5267] <= layer1_out[1049];
     layer2_out[5268] <= ~layer1_out[3893];
     layer2_out[5269] <= layer1_out[3851];
     layer2_out[5270] <= layer1_out[9512];
     layer2_out[5271] <= layer1_out[1498] ^ layer1_out[1499];
     layer2_out[5272] <= ~(layer1_out[1456] & layer1_out[1457]);
     layer2_out[5273] <= layer1_out[471] & layer1_out[472];
     layer2_out[5274] <= layer1_out[11534];
     layer2_out[5275] <= layer1_out[2177];
     layer2_out[5276] <= ~layer1_out[8841];
     layer2_out[5277] <= layer1_out[10560] & ~layer1_out[10561];
     layer2_out[5278] <= ~layer1_out[2492] | layer1_out[2491];
     layer2_out[5279] <= ~(layer1_out[9265] ^ layer1_out[9266]);
     layer2_out[5280] <= layer1_out[8889];
     layer2_out[5281] <= ~(layer1_out[566] | layer1_out[567]);
     layer2_out[5282] <= ~layer1_out[9612];
     layer2_out[5283] <= ~layer1_out[23];
     layer2_out[5284] <= layer1_out[0];
     layer2_out[5285] <= layer1_out[3107] & ~layer1_out[3106];
     layer2_out[5286] <= ~(layer1_out[2083] | layer1_out[2084]);
     layer2_out[5287] <= ~(layer1_out[6373] | layer1_out[6374]);
     layer2_out[5288] <= layer1_out[5182];
     layer2_out[5289] <= layer1_out[4445] & ~layer1_out[4444];
     layer2_out[5290] <= ~layer1_out[2474];
     layer2_out[5291] <= layer1_out[3969] & layer1_out[3970];
     layer2_out[5292] <= ~layer1_out[848];
     layer2_out[5293] <= layer1_out[1739];
     layer2_out[5294] <= ~(layer1_out[490] ^ layer1_out[491]);
     layer2_out[5295] <= layer1_out[4124] & ~layer1_out[4123];
     layer2_out[5296] <= layer1_out[9892] & ~layer1_out[9893];
     layer2_out[5297] <= ~layer1_out[9360] | layer1_out[9359];
     layer2_out[5298] <= ~layer1_out[7668];
     layer2_out[5299] <= layer1_out[6452] | layer1_out[6453];
     layer2_out[5300] <= ~(layer1_out[3637] & layer1_out[3638]);
     layer2_out[5301] <= layer1_out[10340] | layer1_out[10341];
     layer2_out[5302] <= ~(layer1_out[879] | layer1_out[880]);
     layer2_out[5303] <= ~layer1_out[11939] | layer1_out[11938];
     layer2_out[5304] <= layer1_out[2892];
     layer2_out[5305] <= ~layer1_out[1749] | layer1_out[1750];
     layer2_out[5306] <= ~layer1_out[1745];
     layer2_out[5307] <= layer1_out[6231];
     layer2_out[5308] <= ~layer1_out[6216] | layer1_out[6215];
     layer2_out[5309] <= layer1_out[3619] | layer1_out[3620];
     layer2_out[5310] <= ~layer1_out[2957];
     layer2_out[5311] <= layer1_out[9343] | layer1_out[9344];
     layer2_out[5312] <= layer1_out[8555];
     layer2_out[5313] <= layer1_out[6672] & layer1_out[6673];
     layer2_out[5314] <= layer1_out[7462] | layer1_out[7463];
     layer2_out[5315] <= 1'b0;
     layer2_out[5316] <= ~layer1_out[5711];
     layer2_out[5317] <= layer1_out[2896] & ~layer1_out[2897];
     layer2_out[5318] <= ~layer1_out[7571] | layer1_out[7572];
     layer2_out[5319] <= layer1_out[5679] | layer1_out[5680];
     layer2_out[5320] <= layer1_out[9154] | layer1_out[9155];
     layer2_out[5321] <= layer1_out[9046] & ~layer1_out[9047];
     layer2_out[5322] <= layer1_out[7298] & ~layer1_out[7299];
     layer2_out[5323] <= ~layer1_out[2481];
     layer2_out[5324] <= layer1_out[5258] ^ layer1_out[5259];
     layer2_out[5325] <= layer1_out[7760] ^ layer1_out[7761];
     layer2_out[5326] <= layer1_out[5487];
     layer2_out[5327] <= layer1_out[6301];
     layer2_out[5328] <= layer1_out[1535] & ~layer1_out[1534];
     layer2_out[5329] <= layer1_out[4010] & layer1_out[4011];
     layer2_out[5330] <= layer1_out[7660] & ~layer1_out[7659];
     layer2_out[5331] <= layer1_out[6451];
     layer2_out[5332] <= layer1_out[6860] & layer1_out[6861];
     layer2_out[5333] <= ~(layer1_out[11656] ^ layer1_out[11657]);
     layer2_out[5334] <= ~(layer1_out[4834] & layer1_out[4835]);
     layer2_out[5335] <= ~layer1_out[10441] | layer1_out[10442];
     layer2_out[5336] <= ~layer1_out[3014] | layer1_out[3015];
     layer2_out[5337] <= layer1_out[4638] & ~layer1_out[4637];
     layer2_out[5338] <= layer1_out[6562] & ~layer1_out[6563];
     layer2_out[5339] <= layer1_out[402];
     layer2_out[5340] <= ~(layer1_out[8218] ^ layer1_out[8219]);
     layer2_out[5341] <= layer1_out[5268];
     layer2_out[5342] <= layer1_out[9523];
     layer2_out[5343] <= layer1_out[9074] ^ layer1_out[9075];
     layer2_out[5344] <= layer1_out[5205];
     layer2_out[5345] <= ~layer1_out[2126];
     layer2_out[5346] <= ~(layer1_out[9986] & layer1_out[9987]);
     layer2_out[5347] <= ~layer1_out[10436] | layer1_out[10437];
     layer2_out[5348] <= ~layer1_out[1964] | layer1_out[1963];
     layer2_out[5349] <= layer1_out[6991] & ~layer1_out[6992];
     layer2_out[5350] <= layer1_out[3242];
     layer2_out[5351] <= ~layer1_out[3533];
     layer2_out[5352] <= ~layer1_out[7428];
     layer2_out[5353] <= ~(layer1_out[5631] ^ layer1_out[5632]);
     layer2_out[5354] <= layer1_out[6672];
     layer2_out[5355] <= ~layer1_out[3063];
     layer2_out[5356] <= layer1_out[5304] ^ layer1_out[5305];
     layer2_out[5357] <= ~layer1_out[8593] | layer1_out[8594];
     layer2_out[5358] <= ~(layer1_out[10300] & layer1_out[10301]);
     layer2_out[5359] <= ~layer1_out[5721];
     layer2_out[5360] <= layer1_out[5171] ^ layer1_out[5172];
     layer2_out[5361] <= ~layer1_out[9815];
     layer2_out[5362] <= ~layer1_out[1936];
     layer2_out[5363] <= layer1_out[10717] & layer1_out[10718];
     layer2_out[5364] <= ~(layer1_out[3767] & layer1_out[3768]);
     layer2_out[5365] <= ~layer1_out[11341];
     layer2_out[5366] <= ~layer1_out[226];
     layer2_out[5367] <= ~layer1_out[5946] | layer1_out[5947];
     layer2_out[5368] <= layer1_out[662] & ~layer1_out[663];
     layer2_out[5369] <= layer1_out[1660];
     layer2_out[5370] <= ~layer1_out[829];
     layer2_out[5371] <= ~(layer1_out[5791] | layer1_out[5792]);
     layer2_out[5372] <= ~(layer1_out[1850] ^ layer1_out[1851]);
     layer2_out[5373] <= 1'b0;
     layer2_out[5374] <= ~(layer1_out[2612] ^ layer1_out[2613]);
     layer2_out[5375] <= layer1_out[6815];
     layer2_out[5376] <= layer1_out[10793] & ~layer1_out[10794];
     layer2_out[5377] <= layer1_out[1229] ^ layer1_out[1230];
     layer2_out[5378] <= layer1_out[5633] & layer1_out[5634];
     layer2_out[5379] <= layer1_out[2680] & layer1_out[2681];
     layer2_out[5380] <= layer1_out[4580] ^ layer1_out[4581];
     layer2_out[5381] <= layer1_out[4377];
     layer2_out[5382] <= ~(layer1_out[3924] & layer1_out[3925]);
     layer2_out[5383] <= ~(layer1_out[4388] & layer1_out[4389]);
     layer2_out[5384] <= layer1_out[11629] & layer1_out[11630];
     layer2_out[5385] <= layer1_out[3713];
     layer2_out[5386] <= layer1_out[4964];
     layer2_out[5387] <= layer1_out[5378] & layer1_out[5379];
     layer2_out[5388] <= layer1_out[9074];
     layer2_out[5389] <= ~layer1_out[4329];
     layer2_out[5390] <= layer1_out[6868] | layer1_out[6869];
     layer2_out[5391] <= ~layer1_out[4092];
     layer2_out[5392] <= ~layer1_out[11574] | layer1_out[11573];
     layer2_out[5393] <= 1'b0;
     layer2_out[5394] <= layer1_out[62];
     layer2_out[5395] <= ~layer1_out[3026];
     layer2_out[5396] <= ~layer1_out[11459];
     layer2_out[5397] <= layer1_out[3967] & ~layer1_out[3968];
     layer2_out[5398] <= 1'b0;
     layer2_out[5399] <= layer1_out[3920] & ~layer1_out[3921];
     layer2_out[5400] <= ~layer1_out[9717];
     layer2_out[5401] <= ~(layer1_out[6028] ^ layer1_out[6029]);
     layer2_out[5402] <= layer1_out[749];
     layer2_out[5403] <= ~layer1_out[3237];
     layer2_out[5404] <= layer1_out[9032] & ~layer1_out[9031];
     layer2_out[5405] <= ~(layer1_out[9146] | layer1_out[9147]);
     layer2_out[5406] <= ~layer1_out[1203];
     layer2_out[5407] <= ~(layer1_out[11875] | layer1_out[11876]);
     layer2_out[5408] <= layer1_out[3990] & ~layer1_out[3989];
     layer2_out[5409] <= layer1_out[11751];
     layer2_out[5410] <= layer1_out[1385];
     layer2_out[5411] <= ~layer1_out[11698];
     layer2_out[5412] <= layer1_out[7867] ^ layer1_out[7868];
     layer2_out[5413] <= layer1_out[4411];
     layer2_out[5414] <= ~(layer1_out[4241] | layer1_out[4242]);
     layer2_out[5415] <= layer1_out[9195];
     layer2_out[5416] <= ~(layer1_out[665] | layer1_out[666]);
     layer2_out[5417] <= ~layer1_out[5190];
     layer2_out[5418] <= layer1_out[5675] ^ layer1_out[5676];
     layer2_out[5419] <= ~layer1_out[5272];
     layer2_out[5420] <= layer1_out[4632] & layer1_out[4633];
     layer2_out[5421] <= layer1_out[859] & ~layer1_out[858];
     layer2_out[5422] <= ~layer1_out[3840];
     layer2_out[5423] <= layer1_out[10288] ^ layer1_out[10289];
     layer2_out[5424] <= layer1_out[8202];
     layer2_out[5425] <= layer1_out[8787];
     layer2_out[5426] <= ~layer1_out[4044] | layer1_out[4043];
     layer2_out[5427] <= layer1_out[5472];
     layer2_out[5428] <= ~layer1_out[10725] | layer1_out[10724];
     layer2_out[5429] <= ~layer1_out[9654] | layer1_out[9655];
     layer2_out[5430] <= layer1_out[5051] & ~layer1_out[5052];
     layer2_out[5431] <= layer1_out[6188] & ~layer1_out[6189];
     layer2_out[5432] <= ~layer1_out[833] | layer1_out[834];
     layer2_out[5433] <= layer1_out[4316] & ~layer1_out[4315];
     layer2_out[5434] <= ~layer1_out[6344];
     layer2_out[5435] <= 1'b0;
     layer2_out[5436] <= layer1_out[6909] & ~layer1_out[6910];
     layer2_out[5437] <= ~(layer1_out[10440] | layer1_out[10441]);
     layer2_out[5438] <= ~layer1_out[2037];
     layer2_out[5439] <= layer1_out[3410] | layer1_out[3411];
     layer2_out[5440] <= layer1_out[8447];
     layer2_out[5441] <= layer1_out[1191];
     layer2_out[5442] <= ~layer1_out[10578];
     layer2_out[5443] <= layer1_out[10216] & ~layer1_out[10215];
     layer2_out[5444] <= layer1_out[10144];
     layer2_out[5445] <= layer1_out[11731];
     layer2_out[5446] <= 1'b0;
     layer2_out[5447] <= layer1_out[3851];
     layer2_out[5448] <= layer1_out[680];
     layer2_out[5449] <= layer1_out[9237] & ~layer1_out[9238];
     layer2_out[5450] <= ~layer1_out[8847];
     layer2_out[5451] <= layer1_out[543] & ~layer1_out[542];
     layer2_out[5452] <= 1'b1;
     layer2_out[5453] <= ~layer1_out[11926] | layer1_out[11925];
     layer2_out[5454] <= layer1_out[1423] & ~layer1_out[1422];
     layer2_out[5455] <= ~layer1_out[7818] | layer1_out[7819];
     layer2_out[5456] <= layer1_out[5158];
     layer2_out[5457] <= 1'b0;
     layer2_out[5458] <= layer1_out[9926] & ~layer1_out[9927];
     layer2_out[5459] <= layer1_out[10295];
     layer2_out[5460] <= layer1_out[7798] & ~layer1_out[7797];
     layer2_out[5461] <= layer1_out[6279];
     layer2_out[5462] <= layer1_out[11901] & ~layer1_out[11900];
     layer2_out[5463] <= layer1_out[11413] | layer1_out[11414];
     layer2_out[5464] <= layer1_out[3399] | layer1_out[3400];
     layer2_out[5465] <= ~(layer1_out[4175] ^ layer1_out[4176]);
     layer2_out[5466] <= layer1_out[803];
     layer2_out[5467] <= layer1_out[9831] & layer1_out[9832];
     layer2_out[5468] <= ~(layer1_out[3019] | layer1_out[3020]);
     layer2_out[5469] <= ~layer1_out[2178];
     layer2_out[5470] <= ~(layer1_out[10202] ^ layer1_out[10203]);
     layer2_out[5471] <= layer1_out[1409] & ~layer1_out[1410];
     layer2_out[5472] <= ~(layer1_out[2794] | layer1_out[2795]);
     layer2_out[5473] <= layer1_out[1367] & ~layer1_out[1366];
     layer2_out[5474] <= 1'b1;
     layer2_out[5475] <= layer1_out[746] & ~layer1_out[745];
     layer2_out[5476] <= layer1_out[4669] & layer1_out[4670];
     layer2_out[5477] <= ~(layer1_out[912] ^ layer1_out[913]);
     layer2_out[5478] <= ~layer1_out[8266];
     layer2_out[5479] <= layer1_out[8861] ^ layer1_out[8862];
     layer2_out[5480] <= layer1_out[7003] ^ layer1_out[7004];
     layer2_out[5481] <= layer1_out[2439];
     layer2_out[5482] <= ~(layer1_out[2001] | layer1_out[2002]);
     layer2_out[5483] <= ~layer1_out[6670];
     layer2_out[5484] <= ~layer1_out[11195];
     layer2_out[5485] <= ~layer1_out[8768] | layer1_out[8769];
     layer2_out[5486] <= layer1_out[4939] & ~layer1_out[4938];
     layer2_out[5487] <= 1'b1;
     layer2_out[5488] <= layer1_out[3246] & layer1_out[3247];
     layer2_out[5489] <= layer1_out[2391] | layer1_out[2392];
     layer2_out[5490] <= ~(layer1_out[3549] & layer1_out[3550]);
     layer2_out[5491] <= ~layer1_out[5645] | layer1_out[5646];
     layer2_out[5492] <= ~layer1_out[6750] | layer1_out[6749];
     layer2_out[5493] <= ~(layer1_out[10052] ^ layer1_out[10053]);
     layer2_out[5494] <= ~layer1_out[445];
     layer2_out[5495] <= ~(layer1_out[3651] | layer1_out[3652]);
     layer2_out[5496] <= ~layer1_out[9646];
     layer2_out[5497] <= ~layer1_out[10297];
     layer2_out[5498] <= ~layer1_out[11531];
     layer2_out[5499] <= ~layer1_out[5231];
     layer2_out[5500] <= layer1_out[1925] & ~layer1_out[1926];
     layer2_out[5501] <= layer1_out[1233];
     layer2_out[5502] <= ~(layer1_out[7001] ^ layer1_out[7002]);
     layer2_out[5503] <= layer1_out[5659] & layer1_out[5660];
     layer2_out[5504] <= layer1_out[7685] & ~layer1_out[7686];
     layer2_out[5505] <= ~layer1_out[1589];
     layer2_out[5506] <= ~(layer1_out[6033] ^ layer1_out[6034]);
     layer2_out[5507] <= ~layer1_out[1348] | layer1_out[1349];
     layer2_out[5508] <= ~layer1_out[8897] | layer1_out[8896];
     layer2_out[5509] <= layer1_out[3644] ^ layer1_out[3645];
     layer2_out[5510] <= layer1_out[2202] ^ layer1_out[2203];
     layer2_out[5511] <= layer1_out[7749] ^ layer1_out[7750];
     layer2_out[5512] <= ~layer1_out[10564] | layer1_out[10563];
     layer2_out[5513] <= layer1_out[9124];
     layer2_out[5514] <= layer1_out[9234];
     layer2_out[5515] <= ~layer1_out[954] | layer1_out[953];
     layer2_out[5516] <= layer1_out[2094] | layer1_out[2095];
     layer2_out[5517] <= layer1_out[7225];
     layer2_out[5518] <= ~(layer1_out[8133] ^ layer1_out[8134]);
     layer2_out[5519] <= ~layer1_out[11678] | layer1_out[11677];
     layer2_out[5520] <= ~(layer1_out[5658] ^ layer1_out[5659]);
     layer2_out[5521] <= layer1_out[10843] ^ layer1_out[10844];
     layer2_out[5522] <= ~layer1_out[8145];
     layer2_out[5523] <= ~layer1_out[199] | layer1_out[198];
     layer2_out[5524] <= ~layer1_out[8684];
     layer2_out[5525] <= layer1_out[11975];
     layer2_out[5526] <= layer1_out[3291];
     layer2_out[5527] <= layer1_out[2111];
     layer2_out[5528] <= ~(layer1_out[5325] | layer1_out[5326]);
     layer2_out[5529] <= ~(layer1_out[11442] | layer1_out[11443]);
     layer2_out[5530] <= ~layer1_out[8520];
     layer2_out[5531] <= ~(layer1_out[2338] & layer1_out[2339]);
     layer2_out[5532] <= ~layer1_out[579] | layer1_out[578];
     layer2_out[5533] <= ~layer1_out[10640] | layer1_out[10641];
     layer2_out[5534] <= 1'b1;
     layer2_out[5535] <= layer1_out[5367] ^ layer1_out[5368];
     layer2_out[5536] <= layer1_out[3974] ^ layer1_out[3975];
     layer2_out[5537] <= ~(layer1_out[7221] ^ layer1_out[7222]);
     layer2_out[5538] <= ~layer1_out[8964];
     layer2_out[5539] <= ~(layer1_out[387] | layer1_out[388]);
     layer2_out[5540] <= ~(layer1_out[6774] & layer1_out[6775]);
     layer2_out[5541] <= ~(layer1_out[7632] | layer1_out[7633]);
     layer2_out[5542] <= layer1_out[2293];
     layer2_out[5543] <= ~layer1_out[10029];
     layer2_out[5544] <= layer1_out[4718] ^ layer1_out[4719];
     layer2_out[5545] <= layer1_out[8373];
     layer2_out[5546] <= layer1_out[11426] & ~layer1_out[11425];
     layer2_out[5547] <= layer1_out[10491] & layer1_out[10492];
     layer2_out[5548] <= layer1_out[3155];
     layer2_out[5549] <= layer1_out[2637];
     layer2_out[5550] <= layer1_out[600];
     layer2_out[5551] <= ~layer1_out[477] | layer1_out[476];
     layer2_out[5552] <= layer1_out[2367] | layer1_out[2368];
     layer2_out[5553] <= ~layer1_out[7259];
     layer2_out[5554] <= ~layer1_out[9149];
     layer2_out[5555] <= ~layer1_out[6802] | layer1_out[6803];
     layer2_out[5556] <= layer1_out[9090];
     layer2_out[5557] <= layer1_out[3461] | layer1_out[3462];
     layer2_out[5558] <= ~layer1_out[3062];
     layer2_out[5559] <= layer1_out[3307] & ~layer1_out[3306];
     layer2_out[5560] <= ~(layer1_out[1765] | layer1_out[1766]);
     layer2_out[5561] <= ~layer1_out[64] | layer1_out[63];
     layer2_out[5562] <= ~layer1_out[4606] | layer1_out[4607];
     layer2_out[5563] <= layer1_out[10726] & ~layer1_out[10727];
     layer2_out[5564] <= ~layer1_out[11413];
     layer2_out[5565] <= layer1_out[6495];
     layer2_out[5566] <= ~layer1_out[9413] | layer1_out[9414];
     layer2_out[5567] <= layer1_out[6492];
     layer2_out[5568] <= layer1_out[11500];
     layer2_out[5569] <= layer1_out[2263] & layer1_out[2264];
     layer2_out[5570] <= layer1_out[10303];
     layer2_out[5571] <= ~(layer1_out[3829] & layer1_out[3830]);
     layer2_out[5572] <= layer1_out[809];
     layer2_out[5573] <= layer1_out[527];
     layer2_out[5574] <= ~(layer1_out[9125] ^ layer1_out[9126]);
     layer2_out[5575] <= ~layer1_out[5470] | layer1_out[5471];
     layer2_out[5576] <= layer1_out[4302];
     layer2_out[5577] <= layer1_out[6313] ^ layer1_out[6314];
     layer2_out[5578] <= ~layer1_out[10241];
     layer2_out[5579] <= ~(layer1_out[4935] & layer1_out[4936]);
     layer2_out[5580] <= ~layer1_out[4417] | layer1_out[4416];
     layer2_out[5581] <= ~layer1_out[8834];
     layer2_out[5582] <= layer1_out[374] & ~layer1_out[373];
     layer2_out[5583] <= layer1_out[5507];
     layer2_out[5584] <= layer1_out[7039] ^ layer1_out[7040];
     layer2_out[5585] <= layer1_out[321];
     layer2_out[5586] <= ~layer1_out[3071];
     layer2_out[5587] <= layer1_out[7283] & layer1_out[7284];
     layer2_out[5588] <= layer1_out[656] | layer1_out[657];
     layer2_out[5589] <= layer1_out[6966] | layer1_out[6967];
     layer2_out[5590] <= ~layer1_out[11279];
     layer2_out[5591] <= ~layer1_out[6724];
     layer2_out[5592] <= ~layer1_out[4995] | layer1_out[4996];
     layer2_out[5593] <= ~layer1_out[9750];
     layer2_out[5594] <= layer1_out[5964];
     layer2_out[5595] <= ~layer1_out[11308] | layer1_out[11307];
     layer2_out[5596] <= ~layer1_out[8677] | layer1_out[8678];
     layer2_out[5597] <= layer1_out[4620];
     layer2_out[5598] <= layer1_out[3208] & ~layer1_out[3207];
     layer2_out[5599] <= ~layer1_out[8628] | layer1_out[8627];
     layer2_out[5600] <= layer1_out[3195];
     layer2_out[5601] <= ~(layer1_out[5009] & layer1_out[5010]);
     layer2_out[5602] <= layer1_out[9649] | layer1_out[9650];
     layer2_out[5603] <= ~(layer1_out[1814] & layer1_out[1815]);
     layer2_out[5604] <= ~(layer1_out[8948] ^ layer1_out[8949]);
     layer2_out[5605] <= ~layer1_out[11906];
     layer2_out[5606] <= ~layer1_out[3791];
     layer2_out[5607] <= layer1_out[11262];
     layer2_out[5608] <= layer1_out[10442] & ~layer1_out[10443];
     layer2_out[5609] <= ~(layer1_out[6772] | layer1_out[6773]);
     layer2_out[5610] <= layer1_out[153] ^ layer1_out[154];
     layer2_out[5611] <= ~(layer1_out[4733] & layer1_out[4734]);
     layer2_out[5612] <= layer1_out[3396] & ~layer1_out[3397];
     layer2_out[5613] <= ~(layer1_out[8290] & layer1_out[8291]);
     layer2_out[5614] <= layer1_out[10970];
     layer2_out[5615] <= layer1_out[10584] & layer1_out[10585];
     layer2_out[5616] <= ~layer1_out[4355];
     layer2_out[5617] <= ~(layer1_out[10931] | layer1_out[10932]);
     layer2_out[5618] <= layer1_out[11243] ^ layer1_out[11244];
     layer2_out[5619] <= layer1_out[9398];
     layer2_out[5620] <= ~layer1_out[3986] | layer1_out[3987];
     layer2_out[5621] <= layer1_out[4817];
     layer2_out[5622] <= ~layer1_out[9542] | layer1_out[9541];
     layer2_out[5623] <= layer1_out[10857];
     layer2_out[5624] <= ~(layer1_out[666] & layer1_out[667]);
     layer2_out[5625] <= layer1_out[8553] & layer1_out[8554];
     layer2_out[5626] <= ~layer1_out[9952] | layer1_out[9953];
     layer2_out[5627] <= layer1_out[3729] & ~layer1_out[3728];
     layer2_out[5628] <= layer1_out[1860];
     layer2_out[5629] <= ~layer1_out[5310] | layer1_out[5311];
     layer2_out[5630] <= ~(layer1_out[2596] ^ layer1_out[2597]);
     layer2_out[5631] <= ~layer1_out[11605];
     layer2_out[5632] <= ~layer1_out[1468];
     layer2_out[5633] <= layer1_out[8680];
     layer2_out[5634] <= ~layer1_out[5849];
     layer2_out[5635] <= layer1_out[2209] & ~layer1_out[2208];
     layer2_out[5636] <= layer1_out[8637] & ~layer1_out[8638];
     layer2_out[5637] <= layer1_out[5429] | layer1_out[5430];
     layer2_out[5638] <= ~(layer1_out[7467] & layer1_out[7468]);
     layer2_out[5639] <= layer1_out[11838] | layer1_out[11839];
     layer2_out[5640] <= ~(layer1_out[11093] ^ layer1_out[11094]);
     layer2_out[5641] <= layer1_out[9221];
     layer2_out[5642] <= ~layer1_out[10633];
     layer2_out[5643] <= ~layer1_out[10484] | layer1_out[10483];
     layer2_out[5644] <= ~layer1_out[11465];
     layer2_out[5645] <= ~(layer1_out[4581] ^ layer1_out[4582]);
     layer2_out[5646] <= ~(layer1_out[4535] & layer1_out[4536]);
     layer2_out[5647] <= layer1_out[3664];
     layer2_out[5648] <= layer1_out[10566] & layer1_out[10567];
     layer2_out[5649] <= layer1_out[7440];
     layer2_out[5650] <= layer1_out[113];
     layer2_out[5651] <= ~(layer1_out[8498] ^ layer1_out[8499]);
     layer2_out[5652] <= ~layer1_out[3680];
     layer2_out[5653] <= layer1_out[6718] | layer1_out[6719];
     layer2_out[5654] <= 1'b1;
     layer2_out[5655] <= layer1_out[1855] | layer1_out[1856];
     layer2_out[5656] <= layer1_out[8746] & ~layer1_out[8747];
     layer2_out[5657] <= layer1_out[9654];
     layer2_out[5658] <= layer1_out[3488] ^ layer1_out[3489];
     layer2_out[5659] <= layer1_out[9065];
     layer2_out[5660] <= ~layer1_out[1704];
     layer2_out[5661] <= ~(layer1_out[5228] | layer1_out[5229]);
     layer2_out[5662] <= ~layer1_out[3989] | layer1_out[3988];
     layer2_out[5663] <= ~layer1_out[10986];
     layer2_out[5664] <= 1'b0;
     layer2_out[5665] <= layer1_out[7741] & layer1_out[7742];
     layer2_out[5666] <= ~layer1_out[11463] | layer1_out[11462];
     layer2_out[5667] <= layer1_out[8510];
     layer2_out[5668] <= layer1_out[4834];
     layer2_out[5669] <= layer1_out[4477] & ~layer1_out[4478];
     layer2_out[5670] <= ~layer1_out[5867] | layer1_out[5868];
     layer2_out[5671] <= layer1_out[8603];
     layer2_out[5672] <= ~(layer1_out[1061] & layer1_out[1062]);
     layer2_out[5673] <= layer1_out[11312] & ~layer1_out[11311];
     layer2_out[5674] <= layer1_out[5255];
     layer2_out[5675] <= layer1_out[8256];
     layer2_out[5676] <= layer1_out[7460];
     layer2_out[5677] <= layer1_out[30];
     layer2_out[5678] <= ~(layer1_out[972] & layer1_out[973]);
     layer2_out[5679] <= ~layer1_out[9693];
     layer2_out[5680] <= ~layer1_out[3740];
     layer2_out[5681] <= ~layer1_out[7405];
     layer2_out[5682] <= layer1_out[11359];
     layer2_out[5683] <= ~(layer1_out[5993] | layer1_out[5994]);
     layer2_out[5684] <= ~layer1_out[7848];
     layer2_out[5685] <= ~(layer1_out[3193] | layer1_out[3194]);
     layer2_out[5686] <= ~layer1_out[4722];
     layer2_out[5687] <= layer1_out[1108] ^ layer1_out[1109];
     layer2_out[5688] <= ~layer1_out[1624] | layer1_out[1623];
     layer2_out[5689] <= ~layer1_out[5893];
     layer2_out[5690] <= layer1_out[11161] & ~layer1_out[11162];
     layer2_out[5691] <= layer1_out[6019] & ~layer1_out[6018];
     layer2_out[5692] <= ~layer1_out[7755] | layer1_out[7756];
     layer2_out[5693] <= layer1_out[3576];
     layer2_out[5694] <= ~layer1_out[11600];
     layer2_out[5695] <= ~(layer1_out[2676] & layer1_out[2677]);
     layer2_out[5696] <= layer1_out[11299];
     layer2_out[5697] <= layer1_out[3689];
     layer2_out[5698] <= layer1_out[5265] & ~layer1_out[5266];
     layer2_out[5699] <= layer1_out[4948] & ~layer1_out[4947];
     layer2_out[5700] <= layer1_out[4948] ^ layer1_out[4949];
     layer2_out[5701] <= layer1_out[8118];
     layer2_out[5702] <= ~(layer1_out[6682] ^ layer1_out[6683]);
     layer2_out[5703] <= layer1_out[4044];
     layer2_out[5704] <= layer1_out[9648] ^ layer1_out[9649];
     layer2_out[5705] <= layer1_out[267] | layer1_out[268];
     layer2_out[5706] <= ~layer1_out[8965];
     layer2_out[5707] <= ~layer1_out[8806];
     layer2_out[5708] <= ~layer1_out[7551] | layer1_out[7550];
     layer2_out[5709] <= ~(layer1_out[266] | layer1_out[267]);
     layer2_out[5710] <= layer1_out[464] | layer1_out[465];
     layer2_out[5711] <= ~layer1_out[3255];
     layer2_out[5712] <= layer1_out[10855] | layer1_out[10856];
     layer2_out[5713] <= layer1_out[6302] & ~layer1_out[6303];
     layer2_out[5714] <= layer1_out[4641];
     layer2_out[5715] <= ~(layer1_out[6559] | layer1_out[6560]);
     layer2_out[5716] <= ~(layer1_out[886] | layer1_out[887]);
     layer2_out[5717] <= ~(layer1_out[4742] ^ layer1_out[4743]);
     layer2_out[5718] <= ~layer1_out[8025];
     layer2_out[5719] <= layer1_out[8067] & ~layer1_out[8066];
     layer2_out[5720] <= layer1_out[10585];
     layer2_out[5721] <= ~layer1_out[7056] | layer1_out[7057];
     layer2_out[5722] <= ~(layer1_out[5110] ^ layer1_out[5111]);
     layer2_out[5723] <= ~layer1_out[5348] | layer1_out[5347];
     layer2_out[5724] <= layer1_out[4400];
     layer2_out[5725] <= ~(layer1_out[7602] | layer1_out[7603]);
     layer2_out[5726] <= layer1_out[6008];
     layer2_out[5727] <= layer1_out[1459];
     layer2_out[5728] <= layer1_out[8965];
     layer2_out[5729] <= layer1_out[2154] & ~layer1_out[2153];
     layer2_out[5730] <= ~(layer1_out[6428] | layer1_out[6429]);
     layer2_out[5731] <= ~(layer1_out[4113] & layer1_out[4114]);
     layer2_out[5732] <= ~layer1_out[453];
     layer2_out[5733] <= ~layer1_out[3956] | layer1_out[3957];
     layer2_out[5734] <= 1'b1;
     layer2_out[5735] <= layer1_out[2729] ^ layer1_out[2730];
     layer2_out[5736] <= layer1_out[3123] & layer1_out[3124];
     layer2_out[5737] <= ~layer1_out[8843] | layer1_out[8842];
     layer2_out[5738] <= ~layer1_out[5066];
     layer2_out[5739] <= ~layer1_out[9253] | layer1_out[9254];
     layer2_out[5740] <= layer1_out[8121];
     layer2_out[5741] <= layer1_out[8991] ^ layer1_out[8992];
     layer2_out[5742] <= ~layer1_out[8450] | layer1_out[8451];
     layer2_out[5743] <= ~layer1_out[4921];
     layer2_out[5744] <= layer1_out[1372];
     layer2_out[5745] <= ~layer1_out[1670] | layer1_out[1671];
     layer2_out[5746] <= ~layer1_out[4272];
     layer2_out[5747] <= ~(layer1_out[7163] | layer1_out[7164]);
     layer2_out[5748] <= layer1_out[10189] & layer1_out[10190];
     layer2_out[5749] <= ~layer1_out[7185];
     layer2_out[5750] <= ~layer1_out[2751] | layer1_out[2752];
     layer2_out[5751] <= ~layer1_out[1817];
     layer2_out[5752] <= layer1_out[7570];
     layer2_out[5753] <= 1'b0;
     layer2_out[5754] <= ~layer1_out[5517];
     layer2_out[5755] <= layer1_out[51] | layer1_out[52];
     layer2_out[5756] <= layer1_out[5697] & ~layer1_out[5696];
     layer2_out[5757] <= ~(layer1_out[9028] | layer1_out[9029]);
     layer2_out[5758] <= layer1_out[10133];
     layer2_out[5759] <= ~layer1_out[9055];
     layer2_out[5760] <= layer1_out[902] | layer1_out[903];
     layer2_out[5761] <= ~layer1_out[6755] | layer1_out[6756];
     layer2_out[5762] <= layer1_out[7205] & layer1_out[7206];
     layer2_out[5763] <= ~layer1_out[11224] | layer1_out[11223];
     layer2_out[5764] <= ~layer1_out[5464];
     layer2_out[5765] <= layer1_out[9307] | layer1_out[9308];
     layer2_out[5766] <= ~(layer1_out[5212] ^ layer1_out[5213]);
     layer2_out[5767] <= ~(layer1_out[5748] ^ layer1_out[5749]);
     layer2_out[5768] <= ~layer1_out[6770] | layer1_out[6769];
     layer2_out[5769] <= ~layer1_out[1455] | layer1_out[1456];
     layer2_out[5770] <= ~(layer1_out[11191] | layer1_out[11192]);
     layer2_out[5771] <= layer1_out[4983] & ~layer1_out[4984];
     layer2_out[5772] <= layer1_out[9376];
     layer2_out[5773] <= layer1_out[8939];
     layer2_out[5774] <= ~layer1_out[6030];
     layer2_out[5775] <= layer1_out[835];
     layer2_out[5776] <= ~(layer1_out[10508] & layer1_out[10509]);
     layer2_out[5777] <= ~layer1_out[4588];
     layer2_out[5778] <= 1'b1;
     layer2_out[5779] <= ~(layer1_out[9543] ^ layer1_out[9544]);
     layer2_out[5780] <= layer1_out[241] & layer1_out[242];
     layer2_out[5781] <= layer1_out[782] & ~layer1_out[783];
     layer2_out[5782] <= ~layer1_out[1987] | layer1_out[1986];
     layer2_out[5783] <= layer1_out[6919];
     layer2_out[5784] <= ~layer1_out[9182];
     layer2_out[5785] <= ~layer1_out[10529];
     layer2_out[5786] <= layer1_out[5728];
     layer2_out[5787] <= layer1_out[3139] & layer1_out[3140];
     layer2_out[5788] <= ~(layer1_out[5071] | layer1_out[5072]);
     layer2_out[5789] <= layer1_out[1918] & ~layer1_out[1919];
     layer2_out[5790] <= ~layer1_out[3166];
     layer2_out[5791] <= ~layer1_out[6797] | layer1_out[6796];
     layer2_out[5792] <= layer1_out[3888];
     layer2_out[5793] <= ~(layer1_out[9779] ^ layer1_out[9780]);
     layer2_out[5794] <= layer1_out[6632];
     layer2_out[5795] <= ~layer1_out[10976] | layer1_out[10975];
     layer2_out[5796] <= ~(layer1_out[591] & layer1_out[592]);
     layer2_out[5797] <= layer1_out[3545] | layer1_out[3546];
     layer2_out[5798] <= ~(layer1_out[5807] ^ layer1_out[5808]);
     layer2_out[5799] <= layer1_out[11346];
     layer2_out[5800] <= layer1_out[9445] & layer1_out[9446];
     layer2_out[5801] <= layer1_out[4348] ^ layer1_out[4349];
     layer2_out[5802] <= layer1_out[4378] & layer1_out[4379];
     layer2_out[5803] <= ~layer1_out[9500];
     layer2_out[5804] <= ~(layer1_out[5092] & layer1_out[5093]);
     layer2_out[5805] <= layer1_out[4061] ^ layer1_out[4062];
     layer2_out[5806] <= layer1_out[8319] & ~layer1_out[8320];
     layer2_out[5807] <= layer1_out[6352];
     layer2_out[5808] <= ~layer1_out[4244];
     layer2_out[5809] <= layer1_out[11053];
     layer2_out[5810] <= layer1_out[11355] & ~layer1_out[11356];
     layer2_out[5811] <= 1'b0;
     layer2_out[5812] <= ~layer1_out[9864];
     layer2_out[5813] <= layer1_out[425] & ~layer1_out[424];
     layer2_out[5814] <= layer1_out[9751];
     layer2_out[5815] <= ~layer1_out[6177] | layer1_out[6176];
     layer2_out[5816] <= layer1_out[9982] & ~layer1_out[9983];
     layer2_out[5817] <= layer1_out[42] & ~layer1_out[41];
     layer2_out[5818] <= ~layer1_out[5089] | layer1_out[5090];
     layer2_out[5819] <= layer1_out[10410];
     layer2_out[5820] <= layer1_out[6146] | layer1_out[6147];
     layer2_out[5821] <= layer1_out[8904] & ~layer1_out[8903];
     layer2_out[5822] <= layer1_out[10734] & ~layer1_out[10733];
     layer2_out[5823] <= ~(layer1_out[3895] ^ layer1_out[3896]);
     layer2_out[5824] <= ~(layer1_out[4975] & layer1_out[4976]);
     layer2_out[5825] <= layer1_out[11506] | layer1_out[11507];
     layer2_out[5826] <= ~layer1_out[3724];
     layer2_out[5827] <= ~layer1_out[8154] | layer1_out[8153];
     layer2_out[5828] <= ~(layer1_out[7261] | layer1_out[7262]);
     layer2_out[5829] <= layer1_out[11266] | layer1_out[11267];
     layer2_out[5830] <= ~layer1_out[8717];
     layer2_out[5831] <= layer1_out[3309] & ~layer1_out[3308];
     layer2_out[5832] <= layer1_out[7112] & ~layer1_out[7111];
     layer2_out[5833] <= layer1_out[9912] & layer1_out[9913];
     layer2_out[5834] <= ~layer1_out[6393] | layer1_out[6394];
     layer2_out[5835] <= ~layer1_out[1723];
     layer2_out[5836] <= ~layer1_out[10316] | layer1_out[10317];
     layer2_out[5837] <= ~layer1_out[10029];
     layer2_out[5838] <= ~layer1_out[3383] | layer1_out[3382];
     layer2_out[5839] <= layer1_out[8817] & layer1_out[8818];
     layer2_out[5840] <= 1'b0;
     layer2_out[5841] <= ~(layer1_out[1004] | layer1_out[1005]);
     layer2_out[5842] <= layer1_out[7980] & layer1_out[7981];
     layer2_out[5843] <= layer1_out[7625] & layer1_out[7626];
     layer2_out[5844] <= layer1_out[429] & ~layer1_out[428];
     layer2_out[5845] <= ~layer1_out[9287];
     layer2_out[5846] <= layer1_out[3190];
     layer2_out[5847] <= layer1_out[6905] ^ layer1_out[6906];
     layer2_out[5848] <= layer1_out[11963];
     layer2_out[5849] <= ~(layer1_out[8960] | layer1_out[8961]);
     layer2_out[5850] <= ~layer1_out[10901];
     layer2_out[5851] <= ~(layer1_out[9620] ^ layer1_out[9621]);
     layer2_out[5852] <= layer1_out[10116];
     layer2_out[5853] <= layer1_out[5654] & ~layer1_out[5653];
     layer2_out[5854] <= ~layer1_out[9156];
     layer2_out[5855] <= ~layer1_out[6785];
     layer2_out[5856] <= ~layer1_out[6390];
     layer2_out[5857] <= ~layer1_out[4703];
     layer2_out[5858] <= ~layer1_out[3801];
     layer2_out[5859] <= layer1_out[5973] ^ layer1_out[5974];
     layer2_out[5860] <= ~layer1_out[6841];
     layer2_out[5861] <= layer1_out[1972];
     layer2_out[5862] <= ~layer1_out[2390] | layer1_out[2391];
     layer2_out[5863] <= layer1_out[3934] ^ layer1_out[3935];
     layer2_out[5864] <= layer1_out[85] & ~layer1_out[86];
     layer2_out[5865] <= layer1_out[10127] & layer1_out[10128];
     layer2_out[5866] <= layer1_out[4133];
     layer2_out[5867] <= layer1_out[6903];
     layer2_out[5868] <= layer1_out[9885];
     layer2_out[5869] <= ~layer1_out[5308];
     layer2_out[5870] <= ~layer1_out[6564] | layer1_out[6563];
     layer2_out[5871] <= ~(layer1_out[10631] | layer1_out[10632]);
     layer2_out[5872] <= ~(layer1_out[6489] | layer1_out[6490]);
     layer2_out[5873] <= layer1_out[5828] & ~layer1_out[5829];
     layer2_out[5874] <= layer1_out[6898];
     layer2_out[5875] <= ~(layer1_out[3993] & layer1_out[3994]);
     layer2_out[5876] <= ~(layer1_out[10723] | layer1_out[10724]);
     layer2_out[5877] <= ~layer1_out[3425] | layer1_out[3424];
     layer2_out[5878] <= layer1_out[7864] | layer1_out[7865];
     layer2_out[5879] <= layer1_out[9743] & ~layer1_out[9744];
     layer2_out[5880] <= ~layer1_out[413] | layer1_out[414];
     layer2_out[5881] <= ~(layer1_out[5996] | layer1_out[5997]);
     layer2_out[5882] <= layer1_out[3033] & layer1_out[3034];
     layer2_out[5883] <= layer1_out[4383];
     layer2_out[5884] <= ~(layer1_out[5118] & layer1_out[5119]);
     layer2_out[5885] <= ~layer1_out[2676];
     layer2_out[5886] <= layer1_out[10180] | layer1_out[10181];
     layer2_out[5887] <= layer1_out[2123];
     layer2_out[5888] <= layer1_out[915] & ~layer1_out[916];
     layer2_out[5889] <= ~layer1_out[3460];
     layer2_out[5890] <= ~(layer1_out[1552] & layer1_out[1553]);
     layer2_out[5891] <= layer1_out[6205] | layer1_out[6206];
     layer2_out[5892] <= layer1_out[10059];
     layer2_out[5893] <= ~(layer1_out[2479] & layer1_out[2480]);
     layer2_out[5894] <= layer1_out[5872] & ~layer1_out[5871];
     layer2_out[5895] <= layer1_out[7572];
     layer2_out[5896] <= layer1_out[3045];
     layer2_out[5897] <= layer1_out[9705] & ~layer1_out[9704];
     layer2_out[5898] <= ~layer1_out[7467];
     layer2_out[5899] <= ~layer1_out[3540];
     layer2_out[5900] <= layer1_out[3875];
     layer2_out[5901] <= layer1_out[3086];
     layer2_out[5902] <= layer1_out[4111] & ~layer1_out[4110];
     layer2_out[5903] <= layer1_out[7125] & ~layer1_out[7124];
     layer2_out[5904] <= ~layer1_out[1324];
     layer2_out[5905] <= layer1_out[186];
     layer2_out[5906] <= ~(layer1_out[7792] & layer1_out[7793]);
     layer2_out[5907] <= layer1_out[735];
     layer2_out[5908] <= ~layer1_out[5856];
     layer2_out[5909] <= ~(layer1_out[5245] ^ layer1_out[5246]);
     layer2_out[5910] <= layer1_out[7865] | layer1_out[7866];
     layer2_out[5911] <= layer1_out[6935];
     layer2_out[5912] <= ~(layer1_out[7720] | layer1_out[7721]);
     layer2_out[5913] <= layer1_out[3403] & ~layer1_out[3402];
     layer2_out[5914] <= ~(layer1_out[2329] ^ layer1_out[2330]);
     layer2_out[5915] <= layer1_out[3606] ^ layer1_out[3607];
     layer2_out[5916] <= layer1_out[10103] & ~layer1_out[10104];
     layer2_out[5917] <= layer1_out[5385] & ~layer1_out[5386];
     layer2_out[5918] <= ~layer1_out[2725];
     layer2_out[5919] <= ~layer1_out[3487];
     layer2_out[5920] <= layer1_out[1403];
     layer2_out[5921] <= layer1_out[5644] ^ layer1_out[5645];
     layer2_out[5922] <= ~layer1_out[7780];
     layer2_out[5923] <= ~(layer1_out[11802] ^ layer1_out[11803]);
     layer2_out[5924] <= layer1_out[6648] & layer1_out[6649];
     layer2_out[5925] <= ~layer1_out[131];
     layer2_out[5926] <= ~layer1_out[4712];
     layer2_out[5927] <= layer1_out[3021] | layer1_out[3022];
     layer2_out[5928] <= layer1_out[5838];
     layer2_out[5929] <= ~(layer1_out[5273] ^ layer1_out[5274]);
     layer2_out[5930] <= layer1_out[11380] ^ layer1_out[11381];
     layer2_out[5931] <= layer1_out[9681];
     layer2_out[5932] <= layer1_out[5515];
     layer2_out[5933] <= layer1_out[2937] | layer1_out[2938];
     layer2_out[5934] <= layer1_out[11023];
     layer2_out[5935] <= layer1_out[1697];
     layer2_out[5936] <= ~(layer1_out[9994] & layer1_out[9995]);
     layer2_out[5937] <= ~layer1_out[9200] | layer1_out[9199];
     layer2_out[5938] <= layer1_out[8109];
     layer2_out[5939] <= ~(layer1_out[6990] & layer1_out[6991]);
     layer2_out[5940] <= ~layer1_out[2115] | layer1_out[2116];
     layer2_out[5941] <= layer1_out[1124] & layer1_out[1125];
     layer2_out[5942] <= layer1_out[4159] & layer1_out[4160];
     layer2_out[5943] <= layer1_out[7366];
     layer2_out[5944] <= ~layer1_out[4785];
     layer2_out[5945] <= layer1_out[10486] ^ layer1_out[10487];
     layer2_out[5946] <= ~layer1_out[6658];
     layer2_out[5947] <= ~layer1_out[3090] | layer1_out[3091];
     layer2_out[5948] <= ~(layer1_out[5123] | layer1_out[5124]);
     layer2_out[5949] <= ~layer1_out[8446];
     layer2_out[5950] <= ~(layer1_out[5005] & layer1_out[5006]);
     layer2_out[5951] <= layer1_out[9563] & ~layer1_out[9564];
     layer2_out[5952] <= layer1_out[9450];
     layer2_out[5953] <= layer1_out[9547] & ~layer1_out[9548];
     layer2_out[5954] <= layer1_out[796] ^ layer1_out[797];
     layer2_out[5955] <= ~(layer1_out[5519] & layer1_out[5520]);
     layer2_out[5956] <= layer1_out[11280];
     layer2_out[5957] <= ~layer1_out[4397] | layer1_out[4396];
     layer2_out[5958] <= ~(layer1_out[6894] | layer1_out[6895]);
     layer2_out[5959] <= ~layer1_out[8866];
     layer2_out[5960] <= ~layer1_out[9467];
     layer2_out[5961] <= layer1_out[5376] & ~layer1_out[5375];
     layer2_out[5962] <= ~layer1_out[1745];
     layer2_out[5963] <= ~(layer1_out[4992] | layer1_out[4993]);
     layer2_out[5964] <= layer1_out[4143] ^ layer1_out[4144];
     layer2_out[5965] <= ~layer1_out[10452];
     layer2_out[5966] <= layer1_out[9857];
     layer2_out[5967] <= ~(layer1_out[4690] ^ layer1_out[4691]);
     layer2_out[5968] <= layer1_out[10737] & ~layer1_out[10738];
     layer2_out[5969] <= ~layer1_out[2023] | layer1_out[2024];
     layer2_out[5970] <= ~(layer1_out[7608] | layer1_out[7609]);
     layer2_out[5971] <= layer1_out[2989] ^ layer1_out[2990];
     layer2_out[5972] <= layer1_out[655] & ~layer1_out[654];
     layer2_out[5973] <= ~(layer1_out[6615] ^ layer1_out[6616]);
     layer2_out[5974] <= ~(layer1_out[3770] | layer1_out[3771]);
     layer2_out[5975] <= ~(layer1_out[6506] & layer1_out[6507]);
     layer2_out[5976] <= ~(layer1_out[7896] | layer1_out[7897]);
     layer2_out[5977] <= layer1_out[8723] & ~layer1_out[8722];
     layer2_out[5978] <= ~(layer1_out[9469] | layer1_out[9470]);
     layer2_out[5979] <= layer1_out[7708] & layer1_out[7709];
     layer2_out[5980] <= ~layer1_out[3169];
     layer2_out[5981] <= ~layer1_out[5147];
     layer2_out[5982] <= ~(layer1_out[4338] & layer1_out[4339]);
     layer2_out[5983] <= layer1_out[3643] & layer1_out[3644];
     layer2_out[5984] <= ~(layer1_out[817] | layer1_out[818]);
     layer2_out[5985] <= layer1_out[6226] ^ layer1_out[6227];
     layer2_out[5986] <= layer1_out[4466] & ~layer1_out[4467];
     layer2_out[5987] <= ~layer1_out[1031] | layer1_out[1030];
     layer2_out[5988] <= ~layer1_out[3948];
     layer2_out[5989] <= layer1_out[3448] ^ layer1_out[3449];
     layer2_out[5990] <= layer1_out[1529] & ~layer1_out[1528];
     layer2_out[5991] <= ~layer1_out[11228];
     layer2_out[5992] <= layer1_out[11501];
     layer2_out[5993] <= layer1_out[11050] & ~layer1_out[11051];
     layer2_out[5994] <= ~(layer1_out[9738] & layer1_out[9739]);
     layer2_out[5995] <= ~layer1_out[4544];
     layer2_out[5996] <= layer1_out[9209] | layer1_out[9210];
     layer2_out[5997] <= layer1_out[7489] & ~layer1_out[7490];
     layer2_out[5998] <= layer1_out[4538] & ~layer1_out[4537];
     layer2_out[5999] <= ~(layer1_out[10672] | layer1_out[10673]);
     layer2_out[6000] <= layer1_out[9935] & ~layer1_out[9936];
     layer2_out[6001] <= layer1_out[3114] | layer1_out[3115];
     layer2_out[6002] <= ~layer1_out[10003];
     layer2_out[6003] <= ~layer1_out[9714];
     layer2_out[6004] <= ~layer1_out[11586];
     layer2_out[6005] <= layer1_out[2607] | layer1_out[2608];
     layer2_out[6006] <= ~(layer1_out[7889] & layer1_out[7890]);
     layer2_out[6007] <= ~(layer1_out[5689] | layer1_out[5690]);
     layer2_out[6008] <= layer1_out[10075];
     layer2_out[6009] <= ~(layer1_out[949] & layer1_out[950]);
     layer2_out[6010] <= layer1_out[7399] ^ layer1_out[7400];
     layer2_out[6011] <= ~layer1_out[7994] | layer1_out[7993];
     layer2_out[6012] <= layer1_out[1085] & ~layer1_out[1084];
     layer2_out[6013] <= ~(layer1_out[10038] & layer1_out[10039]);
     layer2_out[6014] <= ~layer1_out[1284];
     layer2_out[6015] <= layer1_out[1158] & ~layer1_out[1157];
     layer2_out[6016] <= layer1_out[11457] & layer1_out[11458];
     layer2_out[6017] <= layer1_out[10502] & ~layer1_out[10501];
     layer2_out[6018] <= layer1_out[2032];
     layer2_out[6019] <= layer1_out[7876];
     layer2_out[6020] <= ~layer1_out[3520];
     layer2_out[6021] <= layer1_out[579];
     layer2_out[6022] <= layer1_out[5636] | layer1_out[5637];
     layer2_out[6023] <= ~layer1_out[8825];
     layer2_out[6024] <= layer1_out[66];
     layer2_out[6025] <= layer1_out[11106] | layer1_out[11107];
     layer2_out[6026] <= ~layer1_out[5334];
     layer2_out[6027] <= layer1_out[3479] & ~layer1_out[3478];
     layer2_out[6028] <= layer1_out[7531];
     layer2_out[6029] <= layer1_out[8802] & ~layer1_out[8801];
     layer2_out[6030] <= ~layer1_out[3088];
     layer2_out[6031] <= layer1_out[6423] ^ layer1_out[6424];
     layer2_out[6032] <= ~layer1_out[10305];
     layer2_out[6033] <= ~(layer1_out[10919] ^ layer1_out[10920]);
     layer2_out[6034] <= layer1_out[5072] | layer1_out[5073];
     layer2_out[6035] <= ~(layer1_out[4795] ^ layer1_out[4796]);
     layer2_out[6036] <= layer1_out[7358];
     layer2_out[6037] <= layer1_out[9420];
     layer2_out[6038] <= layer1_out[1181] & ~layer1_out[1180];
     layer2_out[6039] <= ~layer1_out[11269] | layer1_out[11268];
     layer2_out[6040] <= layer1_out[6754];
     layer2_out[6041] <= ~(layer1_out[4174] & layer1_out[4175]);
     layer2_out[6042] <= layer1_out[1913];
     layer2_out[6043] <= ~layer1_out[7353];
     layer2_out[6044] <= layer1_out[827] ^ layer1_out[828];
     layer2_out[6045] <= ~(layer1_out[10984] ^ layer1_out[10985]);
     layer2_out[6046] <= layer1_out[8217] | layer1_out[8218];
     layer2_out[6047] <= ~layer1_out[10551];
     layer2_out[6048] <= ~(layer1_out[9053] & layer1_out[9054]);
     layer2_out[6049] <= ~layer1_out[10767];
     layer2_out[6050] <= ~layer1_out[3712];
     layer2_out[6051] <= layer1_out[6124];
     layer2_out[6052] <= ~layer1_out[9753] | layer1_out[9754];
     layer2_out[6053] <= 1'b0;
     layer2_out[6054] <= ~layer1_out[2119];
     layer2_out[6055] <= layer1_out[3619];
     layer2_out[6056] <= layer1_out[7208] & layer1_out[7209];
     layer2_out[6057] <= layer1_out[6417] | layer1_out[6418];
     layer2_out[6058] <= ~(layer1_out[8003] ^ layer1_out[8004]);
     layer2_out[6059] <= ~(layer1_out[7390] ^ layer1_out[7391]);
     layer2_out[6060] <= layer1_out[11856];
     layer2_out[6061] <= layer1_out[9466];
     layer2_out[6062] <= ~(layer1_out[10262] & layer1_out[10263]);
     layer2_out[6063] <= 1'b1;
     layer2_out[6064] <= layer1_out[11338];
     layer2_out[6065] <= layer1_out[11830];
     layer2_out[6066] <= ~(layer1_out[11407] | layer1_out[11408]);
     layer2_out[6067] <= ~layer1_out[2479] | layer1_out[2478];
     layer2_out[6068] <= layer1_out[22];
     layer2_out[6069] <= layer1_out[5068] & ~layer1_out[5067];
     layer2_out[6070] <= ~layer1_out[4087] | layer1_out[4088];
     layer2_out[6071] <= layer1_out[5];
     layer2_out[6072] <= ~layer1_out[1226];
     layer2_out[6073] <= layer1_out[11731];
     layer2_out[6074] <= layer1_out[4267] & ~layer1_out[4266];
     layer2_out[6075] <= ~layer1_out[1563];
     layer2_out[6076] <= ~(layer1_out[4507] & layer1_out[4508]);
     layer2_out[6077] <= ~layer1_out[6397];
     layer2_out[6078] <= ~(layer1_out[6765] ^ layer1_out[6766]);
     layer2_out[6079] <= ~(layer1_out[2518] & layer1_out[2519]);
     layer2_out[6080] <= layer1_out[8368];
     layer2_out[6081] <= ~layer1_out[6460];
     layer2_out[6082] <= ~layer1_out[7124];
     layer2_out[6083] <= ~(layer1_out[10775] & layer1_out[10776]);
     layer2_out[6084] <= layer1_out[11791];
     layer2_out[6085] <= ~layer1_out[4470];
     layer2_out[6086] <= ~(layer1_out[10402] ^ layer1_out[10403]);
     layer2_out[6087] <= layer1_out[9826];
     layer2_out[6088] <= ~layer1_out[7762];
     layer2_out[6089] <= layer1_out[6351] & ~layer1_out[6352];
     layer2_out[6090] <= ~layer1_out[6464];
     layer2_out[6091] <= ~layer1_out[6085];
     layer2_out[6092] <= ~layer1_out[47] | layer1_out[46];
     layer2_out[6093] <= layer1_out[9823];
     layer2_out[6094] <= ~(layer1_out[7823] & layer1_out[7824]);
     layer2_out[6095] <= ~layer1_out[4968];
     layer2_out[6096] <= ~(layer1_out[228] ^ layer1_out[229]);
     layer2_out[6097] <= layer1_out[7254];
     layer2_out[6098] <= layer1_out[5913] & ~layer1_out[5912];
     layer2_out[6099] <= ~layer1_out[287];
     layer2_out[6100] <= ~layer1_out[3066];
     layer2_out[6101] <= layer1_out[11732] & ~layer1_out[11733];
     layer2_out[6102] <= ~(layer1_out[11994] & layer1_out[11995]);
     layer2_out[6103] <= ~(layer1_out[4667] & layer1_out[4668]);
     layer2_out[6104] <= ~layer1_out[11716] | layer1_out[11715];
     layer2_out[6105] <= layer1_out[10705];
     layer2_out[6106] <= ~layer1_out[8081];
     layer2_out[6107] <= layer1_out[11324];
     layer2_out[6108] <= ~layer1_out[5973];
     layer2_out[6109] <= layer1_out[911] & layer1_out[912];
     layer2_out[6110] <= layer1_out[4223] ^ layer1_out[4224];
     layer2_out[6111] <= ~layer1_out[1859] | layer1_out[1860];
     layer2_out[6112] <= 1'b1;
     layer2_out[6113] <= ~(layer1_out[1277] ^ layer1_out[1278]);
     layer2_out[6114] <= layer1_out[3898];
     layer2_out[6115] <= ~layer1_out[11112] | layer1_out[11111];
     layer2_out[6116] <= layer1_out[3770] & ~layer1_out[3769];
     layer2_out[6117] <= layer1_out[10362];
     layer2_out[6118] <= ~layer1_out[7834] | layer1_out[7835];
     layer2_out[6119] <= layer1_out[7853] | layer1_out[7854];
     layer2_out[6120] <= layer1_out[11992];
     layer2_out[6121] <= layer1_out[4311] ^ layer1_out[4312];
     layer2_out[6122] <= ~layer1_out[8613];
     layer2_out[6123] <= layer1_out[11562] & layer1_out[11563];
     layer2_out[6124] <= layer1_out[8393] & ~layer1_out[8392];
     layer2_out[6125] <= ~layer1_out[3325];
     layer2_out[6126] <= ~(layer1_out[6327] & layer1_out[6328]);
     layer2_out[6127] <= layer1_out[5968];
     layer2_out[6128] <= ~(layer1_out[2758] & layer1_out[2759]);
     layer2_out[6129] <= ~(layer1_out[3456] ^ layer1_out[3457]);
     layer2_out[6130] <= ~(layer1_out[5665] | layer1_out[5666]);
     layer2_out[6131] <= layer1_out[6079];
     layer2_out[6132] <= layer1_out[4066] & ~layer1_out[4067];
     layer2_out[6133] <= layer1_out[11052] & layer1_out[11053];
     layer2_out[6134] <= layer1_out[10983] | layer1_out[10984];
     layer2_out[6135] <= layer1_out[10747] | layer1_out[10748];
     layer2_out[6136] <= layer1_out[1258] | layer1_out[1259];
     layer2_out[6137] <= ~layer1_out[7126];
     layer2_out[6138] <= layer1_out[11650];
     layer2_out[6139] <= ~layer1_out[9500];
     layer2_out[6140] <= ~layer1_out[271] | layer1_out[272];
     layer2_out[6141] <= layer1_out[6974] | layer1_out[6975];
     layer2_out[6142] <= ~layer1_out[6985];
     layer2_out[6143] <= layer1_out[5489] & ~layer1_out[5490];
     layer2_out[6144] <= ~(layer1_out[3750] | layer1_out[3751]);
     layer2_out[6145] <= layer1_out[1250] & ~layer1_out[1249];
     layer2_out[6146] <= layer1_out[8954] & ~layer1_out[8955];
     layer2_out[6147] <= ~layer1_out[2404];
     layer2_out[6148] <= ~layer1_out[8876] | layer1_out[8877];
     layer2_out[6149] <= ~layer1_out[623] | layer1_out[624];
     layer2_out[6150] <= ~layer1_out[3871] | layer1_out[3872];
     layer2_out[6151] <= ~layer1_out[5650];
     layer2_out[6152] <= layer1_out[9374] & ~layer1_out[9373];
     layer2_out[6153] <= ~(layer1_out[8336] ^ layer1_out[8337]);
     layer2_out[6154] <= layer1_out[6022] & ~layer1_out[6023];
     layer2_out[6155] <= layer1_out[11646] & layer1_out[11647];
     layer2_out[6156] <= layer1_out[5701] & ~layer1_out[5702];
     layer2_out[6157] <= ~layer1_out[7927];
     layer2_out[6158] <= layer1_out[3034];
     layer2_out[6159] <= ~(layer1_out[7301] ^ layer1_out[7302]);
     layer2_out[6160] <= layer1_out[8658] ^ layer1_out[8659];
     layer2_out[6161] <= layer1_out[3165] & layer1_out[3166];
     layer2_out[6162] <= ~(layer1_out[8629] & layer1_out[8630]);
     layer2_out[6163] <= layer1_out[3005];
     layer2_out[6164] <= ~layer1_out[11868] | layer1_out[11867];
     layer2_out[6165] <= ~(layer1_out[8289] ^ layer1_out[8290]);
     layer2_out[6166] <= layer1_out[9890];
     layer2_out[6167] <= ~layer1_out[4726] | layer1_out[4725];
     layer2_out[6168] <= ~layer1_out[4240] | layer1_out[4239];
     layer2_out[6169] <= ~layer1_out[1987];
     layer2_out[6170] <= layer1_out[5043] | layer1_out[5044];
     layer2_out[6171] <= ~layer1_out[9887];
     layer2_out[6172] <= layer1_out[10740] & layer1_out[10741];
     layer2_out[6173] <= ~(layer1_out[9403] | layer1_out[9404]);
     layer2_out[6174] <= layer1_out[7214] | layer1_out[7215];
     layer2_out[6175] <= layer1_out[876] | layer1_out[877];
     layer2_out[6176] <= layer1_out[4390] | layer1_out[4391];
     layer2_out[6177] <= ~layer1_out[2919];
     layer2_out[6178] <= ~layer1_out[7363] | layer1_out[7364];
     layer2_out[6179] <= ~layer1_out[9465];
     layer2_out[6180] <= layer1_out[8949];
     layer2_out[6181] <= ~layer1_out[5238] | layer1_out[5239];
     layer2_out[6182] <= ~layer1_out[7961];
     layer2_out[6183] <= ~(layer1_out[5453] & layer1_out[5454]);
     layer2_out[6184] <= ~layer1_out[3955];
     layer2_out[6185] <= layer1_out[1628];
     layer2_out[6186] <= layer1_out[3413] | layer1_out[3414];
     layer2_out[6187] <= layer1_out[47];
     layer2_out[6188] <= layer1_out[9893];
     layer2_out[6189] <= layer1_out[10012] & layer1_out[10013];
     layer2_out[6190] <= layer1_out[10909] & layer1_out[10910];
     layer2_out[6191] <= layer1_out[977] ^ layer1_out[978];
     layer2_out[6192] <= layer1_out[398];
     layer2_out[6193] <= layer1_out[5198] & layer1_out[5199];
     layer2_out[6194] <= ~(layer1_out[816] ^ layer1_out[817]);
     layer2_out[6195] <= ~layer1_out[10765];
     layer2_out[6196] <= ~(layer1_out[2279] ^ layer1_out[2280]);
     layer2_out[6197] <= layer1_out[5149] ^ layer1_out[5150];
     layer2_out[6198] <= layer1_out[2276] ^ layer1_out[2277];
     layer2_out[6199] <= layer1_out[8736] ^ layer1_out[8737];
     layer2_out[6200] <= ~layer1_out[885] | layer1_out[884];
     layer2_out[6201] <= layer1_out[1572] ^ layer1_out[1573];
     layer2_out[6202] <= 1'b0;
     layer2_out[6203] <= layer1_out[55];
     layer2_out[6204] <= ~layer1_out[3431] | layer1_out[3432];
     layer2_out[6205] <= ~layer1_out[8082] | layer1_out[8083];
     layer2_out[6206] <= ~layer1_out[11014] | layer1_out[11015];
     layer2_out[6207] <= layer1_out[10314];
     layer2_out[6208] <= ~(layer1_out[1074] | layer1_out[1075]);
     layer2_out[6209] <= layer1_out[6707];
     layer2_out[6210] <= ~(layer1_out[7925] & layer1_out[7926]);
     layer2_out[6211] <= ~(layer1_out[11727] & layer1_out[11728]);
     layer2_out[6212] <= ~layer1_out[1291];
     layer2_out[6213] <= ~layer1_out[4972];
     layer2_out[6214] <= ~layer1_out[9992] | layer1_out[9991];
     layer2_out[6215] <= ~(layer1_out[3588] | layer1_out[3589]);
     layer2_out[6216] <= layer1_out[9510];
     layer2_out[6217] <= ~layer1_out[9181] | layer1_out[9180];
     layer2_out[6218] <= layer1_out[3047];
     layer2_out[6219] <= layer1_out[1650];
     layer2_out[6220] <= layer1_out[11426] & layer1_out[11427];
     layer2_out[6221] <= ~layer1_out[763] | layer1_out[762];
     layer2_out[6222] <= ~layer1_out[7442] | layer1_out[7441];
     layer2_out[6223] <= ~layer1_out[4801];
     layer2_out[6224] <= ~layer1_out[1150];
     layer2_out[6225] <= ~(layer1_out[2236] ^ layer1_out[2237]);
     layer2_out[6226] <= layer1_out[4129] & layer1_out[4130];
     layer2_out[6227] <= 1'b1;
     layer2_out[6228] <= layer1_out[8061] | layer1_out[8062];
     layer2_out[6229] <= layer1_out[2554] | layer1_out[2555];
     layer2_out[6230] <= layer1_out[8090] & ~layer1_out[8089];
     layer2_out[6231] <= ~layer1_out[9659] | layer1_out[9660];
     layer2_out[6232] <= ~layer1_out[9972] | layer1_out[9973];
     layer2_out[6233] <= ~layer1_out[1471];
     layer2_out[6234] <= ~layer1_out[4037] | layer1_out[4038];
     layer2_out[6235] <= ~layer1_out[11872];
     layer2_out[6236] <= ~layer1_out[4173];
     layer2_out[6237] <= layer1_out[9066] & layer1_out[9067];
     layer2_out[6238] <= ~(layer1_out[11230] & layer1_out[11231]);
     layer2_out[6239] <= layer1_out[5221];
     layer2_out[6240] <= ~(layer1_out[2376] ^ layer1_out[2377]);
     layer2_out[6241] <= layer1_out[10476] & layer1_out[10477];
     layer2_out[6242] <= ~layer1_out[8264] | layer1_out[8265];
     layer2_out[6243] <= ~(layer1_out[8171] & layer1_out[8172]);
     layer2_out[6244] <= ~(layer1_out[8638] ^ layer1_out[8639]);
     layer2_out[6245] <= ~layer1_out[2477] | layer1_out[2476];
     layer2_out[6246] <= ~layer1_out[5914];
     layer2_out[6247] <= layer1_out[11233] ^ layer1_out[11234];
     layer2_out[6248] <= layer1_out[4004];
     layer2_out[6249] <= layer1_out[5290] & ~layer1_out[5289];
     layer2_out[6250] <= layer1_out[5888];
     layer2_out[6251] <= ~(layer1_out[2823] ^ layer1_out[2824]);
     layer2_out[6252] <= ~layer1_out[10843];
     layer2_out[6253] <= ~layer1_out[6254];
     layer2_out[6254] <= ~layer1_out[7469];
     layer2_out[6255] <= ~layer1_out[9949] | layer1_out[9950];
     layer2_out[6256] <= layer1_out[1923];
     layer2_out[6257] <= ~layer1_out[2324] | layer1_out[2325];
     layer2_out[6258] <= ~layer1_out[11022];
     layer2_out[6259] <= ~(layer1_out[997] & layer1_out[998]);
     layer2_out[6260] <= layer1_out[7200] & layer1_out[7201];
     layer2_out[6261] <= 1'b1;
     layer2_out[6262] <= ~layer1_out[6790];
     layer2_out[6263] <= ~layer1_out[6926];
     layer2_out[6264] <= layer1_out[10636];
     layer2_out[6265] <= ~layer1_out[9970];
     layer2_out[6266] <= layer1_out[1903];
     layer2_out[6267] <= ~layer1_out[3623] | layer1_out[3622];
     layer2_out[6268] <= ~(layer1_out[5188] & layer1_out[5189]);
     layer2_out[6269] <= layer1_out[2227] & ~layer1_out[2226];
     layer2_out[6270] <= ~layer1_out[4495];
     layer2_out[6271] <= ~layer1_out[5449] | layer1_out[5448];
     layer2_out[6272] <= ~layer1_out[4045] | layer1_out[4046];
     layer2_out[6273] <= layer1_out[7916] | layer1_out[7917];
     layer2_out[6274] <= ~layer1_out[9121];
     layer2_out[6275] <= layer1_out[7820];
     layer2_out[6276] <= ~layer1_out[5865] | layer1_out[5864];
     layer2_out[6277] <= ~(layer1_out[10221] | layer1_out[10222]);
     layer2_out[6278] <= layer1_out[4993];
     layer2_out[6279] <= ~layer1_out[8508];
     layer2_out[6280] <= ~layer1_out[474];
     layer2_out[6281] <= layer1_out[3860] & ~layer1_out[3861];
     layer2_out[6282] <= layer1_out[7588];
     layer2_out[6283] <= layer1_out[7714];
     layer2_out[6284] <= ~layer1_out[2390];
     layer2_out[6285] <= ~layer1_out[2697];
     layer2_out[6286] <= 1'b0;
     layer2_out[6287] <= layer1_out[6178];
     layer2_out[6288] <= layer1_out[384] & layer1_out[385];
     layer2_out[6289] <= layer1_out[3501] & ~layer1_out[3500];
     layer2_out[6290] <= ~(layer1_out[1579] ^ layer1_out[1580]);
     layer2_out[6291] <= layer1_out[2632];
     layer2_out[6292] <= layer1_out[9851];
     layer2_out[6293] <= layer1_out[4549] & ~layer1_out[4550];
     layer2_out[6294] <= ~layer1_out[4363] | layer1_out[4364];
     layer2_out[6295] <= layer1_out[1864] & ~layer1_out[1863];
     layer2_out[6296] <= ~layer1_out[9726];
     layer2_out[6297] <= ~(layer1_out[3571] ^ layer1_out[3572]);
     layer2_out[6298] <= ~(layer1_out[7237] & layer1_out[7238]);
     layer2_out[6299] <= ~layer1_out[9607] | layer1_out[9606];
     layer2_out[6300] <= layer1_out[6794] & ~layer1_out[6793];
     layer2_out[6301] <= ~layer1_out[8857];
     layer2_out[6302] <= ~layer1_out[3160];
     layer2_out[6303] <= layer1_out[10904] & layer1_out[10905];
     layer2_out[6304] <= layer1_out[4201] | layer1_out[4202];
     layer2_out[6305] <= ~layer1_out[443] | layer1_out[444];
     layer2_out[6306] <= ~layer1_out[1636];
     layer2_out[6307] <= layer1_out[742];
     layer2_out[6308] <= 1'b1;
     layer2_out[6309] <= ~(layer1_out[8165] | layer1_out[8166]);
     layer2_out[6310] <= layer1_out[1138];
     layer2_out[6311] <= layer1_out[2706] & ~layer1_out[2707];
     layer2_out[6312] <= ~layer1_out[10179];
     layer2_out[6313] <= 1'b0;
     layer2_out[6314] <= ~layer1_out[1862];
     layer2_out[6315] <= layer1_out[1153];
     layer2_out[6316] <= ~(layer1_out[4421] | layer1_out[4422]);
     layer2_out[6317] <= ~(layer1_out[10790] | layer1_out[10791]);
     layer2_out[6318] <= ~(layer1_out[5326] & layer1_out[5327]);
     layer2_out[6319] <= layer1_out[1917];
     layer2_out[6320] <= ~layer1_out[9827];
     layer2_out[6321] <= layer1_out[2833];
     layer2_out[6322] <= layer1_out[3688];
     layer2_out[6323] <= layer1_out[5969] | layer1_out[5970];
     layer2_out[6324] <= layer1_out[3185] & ~layer1_out[3186];
     layer2_out[6325] <= ~layer1_out[11305] | layer1_out[11306];
     layer2_out[6326] <= layer1_out[11955] & ~layer1_out[11956];
     layer2_out[6327] <= ~layer1_out[7625] | layer1_out[7624];
     layer2_out[6328] <= layer1_out[6798] ^ layer1_out[6799];
     layer2_out[6329] <= layer1_out[3342];
     layer2_out[6330] <= layer1_out[8645] & layer1_out[8646];
     layer2_out[6331] <= ~(layer1_out[640] & layer1_out[641]);
     layer2_out[6332] <= layer1_out[11095] ^ layer1_out[11096];
     layer2_out[6333] <= ~layer1_out[4168];
     layer2_out[6334] <= ~(layer1_out[3526] ^ layer1_out[3527]);
     layer2_out[6335] <= layer1_out[10906] | layer1_out[10907];
     layer2_out[6336] <= ~layer1_out[5539];
     layer2_out[6337] <= ~layer1_out[3498] | layer1_out[3497];
     layer2_out[6338] <= ~(layer1_out[275] | layer1_out[276]);
     layer2_out[6339] <= layer1_out[632] & ~layer1_out[633];
     layer2_out[6340] <= ~(layer1_out[6311] & layer1_out[6312]);
     layer2_out[6341] <= layer1_out[321];
     layer2_out[6342] <= 1'b0;
     layer2_out[6343] <= ~(layer1_out[6023] | layer1_out[6024]);
     layer2_out[6344] <= ~layer1_out[3201] | layer1_out[3202];
     layer2_out[6345] <= ~layer1_out[6402];
     layer2_out[6346] <= layer1_out[5506];
     layer2_out[6347] <= layer1_out[3996] & ~layer1_out[3997];
     layer2_out[6348] <= layer1_out[7611] & layer1_out[7612];
     layer2_out[6349] <= layer1_out[7143] & ~layer1_out[7142];
     layer2_out[6350] <= layer1_out[5591] ^ layer1_out[5592];
     layer2_out[6351] <= layer1_out[375];
     layer2_out[6352] <= ~(layer1_out[8203] & layer1_out[8204]);
     layer2_out[6353] <= ~layer1_out[6667] | layer1_out[6666];
     layer2_out[6354] <= 1'b1;
     layer2_out[6355] <= layer1_out[8338];
     layer2_out[6356] <= ~layer1_out[3410];
     layer2_out[6357] <= layer1_out[7787];
     layer2_out[6358] <= ~(layer1_out[7079] | layer1_out[7080]);
     layer2_out[6359] <= ~layer1_out[3907];
     layer2_out[6360] <= ~(layer1_out[11597] ^ layer1_out[11598]);
     layer2_out[6361] <= layer1_out[236];
     layer2_out[6362] <= layer1_out[8400];
     layer2_out[6363] <= layer1_out[3237];
     layer2_out[6364] <= ~(layer1_out[11190] | layer1_out[11191]);
     layer2_out[6365] <= ~layer1_out[1063];
     layer2_out[6366] <= ~layer1_out[9251];
     layer2_out[6367] <= ~(layer1_out[11142] ^ layer1_out[11143]);
     layer2_out[6368] <= layer1_out[11418] & ~layer1_out[11417];
     layer2_out[6369] <= layer1_out[6301];
     layer2_out[6370] <= ~(layer1_out[8499] ^ layer1_out[8500]);
     layer2_out[6371] <= ~layer1_out[5440];
     layer2_out[6372] <= layer1_out[6902];
     layer2_out[6373] <= layer1_out[6907];
     layer2_out[6374] <= layer1_out[4758] & layer1_out[4759];
     layer2_out[6375] <= ~layer1_out[5227];
     layer2_out[6376] <= layer1_out[9077] ^ layer1_out[9078];
     layer2_out[6377] <= ~(layer1_out[2741] & layer1_out[2742]);
     layer2_out[6378] <= ~layer1_out[8980];
     layer2_out[6379] <= ~(layer1_out[4979] & layer1_out[4980]);
     layer2_out[6380] <= 1'b0;
     layer2_out[6381] <= ~(layer1_out[7594] & layer1_out[7595]);
     layer2_out[6382] <= layer1_out[1005];
     layer2_out[6383] <= ~layer1_out[8698];
     layer2_out[6384] <= ~layer1_out[8415];
     layer2_out[6385] <= ~layer1_out[5704];
     layer2_out[6386] <= layer1_out[2342] & ~layer1_out[2341];
     layer2_out[6387] <= layer1_out[5831] & ~layer1_out[5830];
     layer2_out[6388] <= ~(layer1_out[2627] ^ layer1_out[2628]);
     layer2_out[6389] <= ~layer1_out[7271];
     layer2_out[6390] <= layer1_out[7382];
     layer2_out[6391] <= layer1_out[3345] | layer1_out[3346];
     layer2_out[6392] <= layer1_out[11618] ^ layer1_out[11619];
     layer2_out[6393] <= layer1_out[7817] & ~layer1_out[7816];
     layer2_out[6394] <= layer1_out[8273];
     layer2_out[6395] <= layer1_out[1710];
     layer2_out[6396] <= layer1_out[5098] & ~layer1_out[5097];
     layer2_out[6397] <= ~layer1_out[6823];
     layer2_out[6398] <= layer1_out[4156];
     layer2_out[6399] <= layer1_out[7221] & ~layer1_out[7220];
     layer2_out[6400] <= ~(layer1_out[2722] ^ layer1_out[2723]);
     layer2_out[6401] <= ~layer1_out[9132];
     layer2_out[6402] <= ~(layer1_out[3621] ^ layer1_out[3622]);
     layer2_out[6403] <= ~(layer1_out[290] | layer1_out[291]);
     layer2_out[6404] <= layer1_out[11194] & ~layer1_out[11193];
     layer2_out[6405] <= ~layer1_out[4928];
     layer2_out[6406] <= ~layer1_out[2610];
     layer2_out[6407] <= ~layer1_out[11627] | layer1_out[11626];
     layer2_out[6408] <= ~layer1_out[5567] | layer1_out[5566];
     layer2_out[6409] <= layer1_out[4952];
     layer2_out[6410] <= ~(layer1_out[11344] & layer1_out[11345]);
     layer2_out[6411] <= layer1_out[4344] ^ layer1_out[4345];
     layer2_out[6412] <= layer1_out[9639];
     layer2_out[6413] <= layer1_out[2622];
     layer2_out[6414] <= layer1_out[5253] | layer1_out[5254];
     layer2_out[6415] <= ~(layer1_out[800] | layer1_out[801]);
     layer2_out[6416] <= layer1_out[818] ^ layer1_out[819];
     layer2_out[6417] <= ~layer1_out[6473];
     layer2_out[6418] <= layer1_out[2092] | layer1_out[2093];
     layer2_out[6419] <= layer1_out[9310] & ~layer1_out[9311];
     layer2_out[6420] <= layer1_out[946] & ~layer1_out[947];
     layer2_out[6421] <= layer1_out[11032] ^ layer1_out[11033];
     layer2_out[6422] <= ~(layer1_out[7700] ^ layer1_out[7701]);
     layer2_out[6423] <= layer1_out[11085];
     layer2_out[6424] <= ~(layer1_out[4508] ^ layer1_out[4509]);
     layer2_out[6425] <= layer1_out[5288] & ~layer1_out[5289];
     layer2_out[6426] <= layer1_out[4293];
     layer2_out[6427] <= ~layer1_out[10438];
     layer2_out[6428] <= ~layer1_out[11247];
     layer2_out[6429] <= ~(layer1_out[4865] | layer1_out[4866]);
     layer2_out[6430] <= ~(layer1_out[7847] & layer1_out[7848]);
     layer2_out[6431] <= layer1_out[1807];
     layer2_out[6432] <= ~layer1_out[10142] | layer1_out[10141];
     layer2_out[6433] <= ~layer1_out[5184] | layer1_out[5185];
     layer2_out[6434] <= layer1_out[2260];
     layer2_out[6435] <= ~layer1_out[2688] | layer1_out[2689];
     layer2_out[6436] <= ~layer1_out[8578];
     layer2_out[6437] <= layer1_out[7513];
     layer2_out[6438] <= layer1_out[11653] & layer1_out[11654];
     layer2_out[6439] <= layer1_out[10865] & layer1_out[10866];
     layer2_out[6440] <= layer1_out[3234];
     layer2_out[6441] <= ~(layer1_out[681] ^ layer1_out[682]);
     layer2_out[6442] <= layer1_out[9916];
     layer2_out[6443] <= layer1_out[6702];
     layer2_out[6444] <= layer1_out[1106];
     layer2_out[6445] <= layer1_out[4900] | layer1_out[4901];
     layer2_out[6446] <= ~(layer1_out[8932] & layer1_out[8933]);
     layer2_out[6447] <= ~layer1_out[8325];
     layer2_out[6448] <= layer1_out[6922] | layer1_out[6923];
     layer2_out[6449] <= 1'b1;
     layer2_out[6450] <= layer1_out[3112];
     layer2_out[6451] <= layer1_out[5577];
     layer2_out[6452] <= ~layer1_out[1925];
     layer2_out[6453] <= ~layer1_out[4579];
     layer2_out[6454] <= ~(layer1_out[3828] & layer1_out[3829]);
     layer2_out[6455] <= ~layer1_out[7843];
     layer2_out[6456] <= ~layer1_out[8354];
     layer2_out[6457] <= ~layer1_out[8099];
     layer2_out[6458] <= layer1_out[7045];
     layer2_out[6459] <= ~layer1_out[6839] | layer1_out[6838];
     layer2_out[6460] <= ~layer1_out[11151];
     layer2_out[6461] <= layer1_out[11557];
     layer2_out[6462] <= layer1_out[1779] | layer1_out[1780];
     layer2_out[6463] <= ~layer1_out[7036];
     layer2_out[6464] <= layer1_out[6279] & layer1_out[6280];
     layer2_out[6465] <= ~layer1_out[10222] | layer1_out[10223];
     layer2_out[6466] <= layer1_out[8654];
     layer2_out[6467] <= ~(layer1_out[587] | layer1_out[588]);
     layer2_out[6468] <= layer1_out[2943];
     layer2_out[6469] <= layer1_out[6627] ^ layer1_out[6628];
     layer2_out[6470] <= ~layer1_out[4105];
     layer2_out[6471] <= ~(layer1_out[8545] ^ layer1_out[8546]);
     layer2_out[6472] <= ~layer1_out[10231] | layer1_out[10230];
     layer2_out[6473] <= ~layer1_out[9805] | layer1_out[9804];
     layer2_out[6474] <= ~layer1_out[715];
     layer2_out[6475] <= layer1_out[2081] & ~layer1_out[2080];
     layer2_out[6476] <= ~(layer1_out[8583] & layer1_out[8584]);
     layer2_out[6477] <= layer1_out[720] ^ layer1_out[721];
     layer2_out[6478] <= layer1_out[11700] & ~layer1_out[11699];
     layer2_out[6479] <= layer1_out[10451] & ~layer1_out[10450];
     layer2_out[6480] <= ~(layer1_out[7986] | layer1_out[7987]);
     layer2_out[6481] <= layer1_out[8444] & layer1_out[8445];
     layer2_out[6482] <= layer1_out[1894];
     layer2_out[6483] <= layer1_out[5692] & layer1_out[5693];
     layer2_out[6484] <= ~(layer1_out[11578] ^ layer1_out[11579]);
     layer2_out[6485] <= layer1_out[530] & layer1_out[531];
     layer2_out[6486] <= ~(layer1_out[9544] & layer1_out[9545]);
     layer2_out[6487] <= layer1_out[2279] & ~layer1_out[2278];
     layer2_out[6488] <= layer1_out[8023] & ~layer1_out[8022];
     layer2_out[6489] <= ~layer1_out[6754];
     layer2_out[6490] <= layer1_out[11790] & layer1_out[11791];
     layer2_out[6491] <= layer1_out[11981] & layer1_out[11982];
     layer2_out[6492] <= ~layer1_out[753];
     layer2_out[6493] <= ~layer1_out[1675] | layer1_out[1674];
     layer2_out[6494] <= layer1_out[5047];
     layer2_out[6495] <= layer1_out[8718] & ~layer1_out[8717];
     layer2_out[6496] <= ~(layer1_out[3291] & layer1_out[3292]);
     layer2_out[6497] <= layer1_out[10315] & layer1_out[10316];
     layer2_out[6498] <= ~layer1_out[4238];
     layer2_out[6499] <= ~layer1_out[11072];
     layer2_out[6500] <= ~(layer1_out[7509] & layer1_out[7510]);
     layer2_out[6501] <= ~layer1_out[8128] | layer1_out[8129];
     layer2_out[6502] <= ~layer1_out[2205] | layer1_out[2204];
     layer2_out[6503] <= ~layer1_out[7323] | layer1_out[7322];
     layer2_out[6504] <= layer1_out[4577] | layer1_out[4578];
     layer2_out[6505] <= layer1_out[5850];
     layer2_out[6506] <= ~(layer1_out[1466] | layer1_out[1467]);
     layer2_out[6507] <= layer1_out[7901] | layer1_out[7902];
     layer2_out[6508] <= layer1_out[10739];
     layer2_out[6509] <= layer1_out[9604] | layer1_out[9605];
     layer2_out[6510] <= layer1_out[7867];
     layer2_out[6511] <= layer1_out[11000] & ~layer1_out[11001];
     layer2_out[6512] <= layer1_out[4449];
     layer2_out[6513] <= ~(layer1_out[10679] & layer1_out[10680]);
     layer2_out[6514] <= ~layer1_out[1242];
     layer2_out[6515] <= layer1_out[10802];
     layer2_out[6516] <= 1'b0;
     layer2_out[6517] <= layer1_out[1296] | layer1_out[1297];
     layer2_out[6518] <= ~(layer1_out[3321] | layer1_out[3322]);
     layer2_out[6519] <= ~layer1_out[8020];
     layer2_out[6520] <= layer1_out[6962] & ~layer1_out[6961];
     layer2_out[6521] <= layer1_out[7514] & ~layer1_out[7515];
     layer2_out[6522] <= layer1_out[8706];
     layer2_out[6523] <= layer1_out[5130] & layer1_out[5131];
     layer2_out[6524] <= layer1_out[8869] ^ layer1_out[8870];
     layer2_out[6525] <= ~layer1_out[1527] | layer1_out[1526];
     layer2_out[6526] <= layer1_out[10224];
     layer2_out[6527] <= layer1_out[7265] | layer1_out[7266];
     layer2_out[6528] <= layer1_out[5217] & ~layer1_out[5216];
     layer2_out[6529] <= layer1_out[7012];
     layer2_out[6530] <= layer1_out[7650];
     layer2_out[6531] <= layer1_out[529];
     layer2_out[6532] <= ~(layer1_out[6219] ^ layer1_out[6220]);
     layer2_out[6533] <= ~layer1_out[9532] | layer1_out[9531];
     layer2_out[6534] <= layer1_out[11444] & ~layer1_out[11445];
     layer2_out[6535] <= layer1_out[3560] ^ layer1_out[3561];
     layer2_out[6536] <= ~layer1_out[8282] | layer1_out[8281];
     layer2_out[6537] <= layer1_out[300] & layer1_out[301];
     layer2_out[6538] <= ~layer1_out[11007];
     layer2_out[6539] <= ~(layer1_out[1438] & layer1_out[1439]);
     layer2_out[6540] <= layer1_out[1637];
     layer2_out[6541] <= ~(layer1_out[7526] | layer1_out[7527]);
     layer2_out[6542] <= ~layer1_out[5458];
     layer2_out[6543] <= layer1_out[135] ^ layer1_out[136];
     layer2_out[6544] <= layer1_out[466];
     layer2_out[6545] <= ~layer1_out[11542];
     layer2_out[6546] <= layer1_out[8076] & ~layer1_out[8077];
     layer2_out[6547] <= ~(layer1_out[1934] | layer1_out[1935]);
     layer2_out[6548] <= layer1_out[3763] & ~layer1_out[3764];
     layer2_out[6549] <= layer1_out[3426] & ~layer1_out[3425];
     layer2_out[6550] <= layer1_out[2971] | layer1_out[2972];
     layer2_out[6551] <= ~(layer1_out[5028] & layer1_out[5029]);
     layer2_out[6552] <= ~(layer1_out[9858] & layer1_out[9859]);
     layer2_out[6553] <= ~layer1_out[6235];
     layer2_out[6554] <= ~layer1_out[7043];
     layer2_out[6555] <= layer1_out[9351] & ~layer1_out[9352];
     layer2_out[6556] <= layer1_out[10095] | layer1_out[10096];
     layer2_out[6557] <= ~layer1_out[10946];
     layer2_out[6558] <= layer1_out[4754];
     layer2_out[6559] <= ~(layer1_out[11090] | layer1_out[11091]);
     layer2_out[6560] <= ~layer1_out[6951] | layer1_out[6952];
     layer2_out[6561] <= layer1_out[1491] ^ layer1_out[1492];
     layer2_out[6562] <= ~layer1_out[6096];
     layer2_out[6563] <= layer1_out[873];
     layer2_out[6564] <= layer1_out[11622];
     layer2_out[6565] <= ~layer1_out[9015];
     layer2_out[6566] <= layer1_out[11643] & ~layer1_out[11644];
     layer2_out[6567] <= layer1_out[10996];
     layer2_out[6568] <= ~layer1_out[9479] | layer1_out[9478];
     layer2_out[6569] <= ~layer1_out[6277];
     layer2_out[6570] <= ~(layer1_out[11082] | layer1_out[11083]);
     layer2_out[6571] <= layer1_out[10434];
     layer2_out[6572] <= layer1_out[11406];
     layer2_out[6573] <= ~layer1_out[5210];
     layer2_out[6574] <= ~layer1_out[6596];
     layer2_out[6575] <= layer1_out[9731];
     layer2_out[6576] <= ~layer1_out[8176];
     layer2_out[6577] <= layer1_out[11287] & layer1_out[11288];
     layer2_out[6578] <= ~layer1_out[10519];
     layer2_out[6579] <= ~layer1_out[7968] | layer1_out[7969];
     layer2_out[6580] <= layer1_out[3427] ^ layer1_out[3428];
     layer2_out[6581] <= layer1_out[4733];
     layer2_out[6582] <= ~layer1_out[8600] | layer1_out[8599];
     layer2_out[6583] <= ~layer1_out[10998];
     layer2_out[6584] <= ~layer1_out[3044] | layer1_out[3043];
     layer2_out[6585] <= ~layer1_out[74];
     layer2_out[6586] <= ~(layer1_out[4381] ^ layer1_out[4382]);
     layer2_out[6587] <= layer1_out[7454] ^ layer1_out[7455];
     layer2_out[6588] <= layer1_out[3935] & layer1_out[3936];
     layer2_out[6589] <= ~(layer1_out[4186] & layer1_out[4187]);
     layer2_out[6590] <= ~layer1_out[8054];
     layer2_out[6591] <= ~layer1_out[129];
     layer2_out[6592] <= layer1_out[9865] | layer1_out[9866];
     layer2_out[6593] <= ~layer1_out[10161];
     layer2_out[6594] <= layer1_out[8921] & ~layer1_out[8920];
     layer2_out[6595] <= layer1_out[7392] & ~layer1_out[7393];
     layer2_out[6596] <= layer1_out[3925];
     layer2_out[6597] <= ~layer1_out[3301];
     layer2_out[6598] <= layer1_out[11365] & ~layer1_out[11364];
     layer2_out[6599] <= ~layer1_out[9001] | layer1_out[9002];
     layer2_out[6600] <= layer1_out[10250];
     layer2_out[6601] <= layer1_out[4314];
     layer2_out[6602] <= layer1_out[9316] & ~layer1_out[9317];
     layer2_out[6603] <= layer1_out[7293];
     layer2_out[6604] <= ~layer1_out[4561];
     layer2_out[6605] <= layer1_out[7886] | layer1_out[7887];
     layer2_out[6606] <= ~(layer1_out[2240] & layer1_out[2241]);
     layer2_out[6607] <= layer1_out[6456] ^ layer1_out[6457];
     layer2_out[6608] <= ~(layer1_out[1632] ^ layer1_out[1633]);
     layer2_out[6609] <= ~(layer1_out[11858] | layer1_out[11859]);
     layer2_out[6610] <= ~(layer1_out[3294] | layer1_out[3295]);
     layer2_out[6611] <= ~(layer1_out[9042] & layer1_out[9043]);
     layer2_out[6612] <= ~layer1_out[1852];
     layer2_out[6613] <= layer1_out[9958] ^ layer1_out[9959];
     layer2_out[6614] <= layer1_out[8691] & layer1_out[8692];
     layer2_out[6615] <= ~layer1_out[11708] | layer1_out[11707];
     layer2_out[6616] <= layer1_out[103] & ~layer1_out[102];
     layer2_out[6617] <= ~layer1_out[5286];
     layer2_out[6618] <= layer1_out[5954];
     layer2_out[6619] <= ~layer1_out[3453] | layer1_out[3452];
     layer2_out[6620] <= layer1_out[8974] & ~layer1_out[8975];
     layer2_out[6621] <= layer1_out[4060];
     layer2_out[6622] <= layer1_out[1090] ^ layer1_out[1091];
     layer2_out[6623] <= layer1_out[4316] | layer1_out[4317];
     layer2_out[6624] <= layer1_out[8387];
     layer2_out[6625] <= layer1_out[3589] & ~layer1_out[3590];
     layer2_out[6626] <= layer1_out[10205];
     layer2_out[6627] <= layer1_out[4671] & ~layer1_out[4672];
     layer2_out[6628] <= layer1_out[2774] & ~layer1_out[2773];
     layer2_out[6629] <= layer1_out[5461];
     layer2_out[6630] <= layer1_out[78] | layer1_out[79];
     layer2_out[6631] <= ~layer1_out[8289] | layer1_out[8288];
     layer2_out[6632] <= layer1_out[9150] | layer1_out[9151];
     layer2_out[6633] <= ~layer1_out[6208];
     layer2_out[6634] <= ~layer1_out[9503];
     layer2_out[6635] <= ~layer1_out[8212] | layer1_out[8211];
     layer2_out[6636] <= layer1_out[8246] & ~layer1_out[8247];
     layer2_out[6637] <= layer1_out[6048] & ~layer1_out[6049];
     layer2_out[6638] <= ~(layer1_out[4847] & layer1_out[4848]);
     layer2_out[6639] <= layer1_out[10532] & layer1_out[10533];
     layer2_out[6640] <= ~(layer1_out[9298] | layer1_out[9299]);
     layer2_out[6641] <= ~layer1_out[8502];
     layer2_out[6642] <= layer1_out[2034] & ~layer1_out[2033];
     layer2_out[6643] <= ~layer1_out[2988];
     layer2_out[6644] <= 1'b0;
     layer2_out[6645] <= ~layer1_out[3336];
     layer2_out[6646] <= ~(layer1_out[9564] | layer1_out[9565]);
     layer2_out[6647] <= ~(layer1_out[2293] | layer1_out[2294]);
     layer2_out[6648] <= layer1_out[11218] | layer1_out[11219];
     layer2_out[6649] <= ~(layer1_out[6801] & layer1_out[6802]);
     layer2_out[6650] <= ~layer1_out[2591] | layer1_out[2592];
     layer2_out[6651] <= layer1_out[5600] | layer1_out[5601];
     layer2_out[6652] <= ~(layer1_out[4007] ^ layer1_out[4008]);
     layer2_out[6653] <= ~layer1_out[10293] | layer1_out[10292];
     layer2_out[6654] <= ~layer1_out[5050];
     layer2_out[6655] <= ~layer1_out[8216];
     layer2_out[6656] <= ~layer1_out[2328];
     layer2_out[6657] <= layer1_out[1452] & ~layer1_out[1453];
     layer2_out[6658] <= layer1_out[9677] | layer1_out[9678];
     layer2_out[6659] <= ~layer1_out[8798];
     layer2_out[6660] <= ~layer1_out[4452] | layer1_out[4451];
     layer2_out[6661] <= layer1_out[5698] & ~layer1_out[5699];
     layer2_out[6662] <= ~(layer1_out[6070] ^ layer1_out[6071]);
     layer2_out[6663] <= layer1_out[1434] & layer1_out[1435];
     layer2_out[6664] <= ~(layer1_out[11849] | layer1_out[11850]);
     layer2_out[6665] <= ~(layer1_out[10993] | layer1_out[10994]);
     layer2_out[6666] <= layer1_out[5628] ^ layer1_out[5629];
     layer2_out[6667] <= layer1_out[4191] & ~layer1_out[4192];
     layer2_out[6668] <= layer1_out[5549] & ~layer1_out[5548];
     layer2_out[6669] <= ~(layer1_out[524] & layer1_out[525]);
     layer2_out[6670] <= ~(layer1_out[4234] & layer1_out[4235]);
     layer2_out[6671] <= ~(layer1_out[9981] ^ layer1_out[9982]);
     layer2_out[6672] <= ~layer1_out[2561] | layer1_out[2560];
     layer2_out[6673] <= ~(layer1_out[791] ^ layer1_out[792]);
     layer2_out[6674] <= layer1_out[7776] & ~layer1_out[7775];
     layer2_out[6675] <= ~layer1_out[5798];
     layer2_out[6676] <= ~layer1_out[10393];
     layer2_out[6677] <= layer1_out[6372];
     layer2_out[6678] <= layer1_out[93] & layer1_out[94];
     layer2_out[6679] <= ~layer1_out[2586];
     layer2_out[6680] <= ~(layer1_out[11821] | layer1_out[11822]);
     layer2_out[6681] <= layer1_out[11836];
     layer2_out[6682] <= ~layer1_out[8551] | layer1_out[8550];
     layer2_out[6683] <= ~layer1_out[10924];
     layer2_out[6684] <= layer1_out[5035] & ~layer1_out[5036];
     layer2_out[6685] <= layer1_out[3742];
     layer2_out[6686] <= ~layer1_out[10323];
     layer2_out[6687] <= ~layer1_out[8719];
     layer2_out[6688] <= layer1_out[2639] & ~layer1_out[2640];
     layer2_out[6689] <= ~layer1_out[280];
     layer2_out[6690] <= ~layer1_out[2104];
     layer2_out[6691] <= layer1_out[7233] & ~layer1_out[7232];
     layer2_out[6692] <= ~(layer1_out[2595] | layer1_out[2596]);
     layer2_out[6693] <= ~layer1_out[5213];
     layer2_out[6694] <= ~layer1_out[10465];
     layer2_out[6695] <= ~layer1_out[3325];
     layer2_out[6696] <= 1'b1;
     layer2_out[6697] <= ~(layer1_out[440] | layer1_out[441]);
     layer2_out[6698] <= ~layer1_out[11958];
     layer2_out[6699] <= ~(layer1_out[4942] & layer1_out[4943]);
     layer2_out[6700] <= ~layer1_out[11207] | layer1_out[11208];
     layer2_out[6701] <= ~layer1_out[3979];
     layer2_out[6702] <= ~(layer1_out[5197] ^ layer1_out[5198]);
     layer2_out[6703] <= layer1_out[6783];
     layer2_out[6704] <= ~layer1_out[6948];
     layer2_out[6705] <= layer1_out[2970] | layer1_out[2971];
     layer2_out[6706] <= layer1_out[4783];
     layer2_out[6707] <= ~(layer1_out[10607] | layer1_out[10608]);
     layer2_out[6708] <= layer1_out[8872] & layer1_out[8873];
     layer2_out[6709] <= layer1_out[9269];
     layer2_out[6710] <= ~layer1_out[1170];
     layer2_out[6711] <= layer1_out[5837];
     layer2_out[6712] <= layer1_out[5283] & ~layer1_out[5284];
     layer2_out[6713] <= layer1_out[1187] & layer1_out[1188];
     layer2_out[6714] <= ~(layer1_out[8941] | layer1_out[8942]);
     layer2_out[6715] <= layer1_out[7735] & ~layer1_out[7736];
     layer2_out[6716] <= ~layer1_out[969] | layer1_out[970];
     layer2_out[6717] <= layer1_out[683];
     layer2_out[6718] <= ~(layer1_out[6024] ^ layer1_out[6025]);
     layer2_out[6719] <= layer1_out[9832];
     layer2_out[6720] <= ~(layer1_out[4196] | layer1_out[4197]);
     layer2_out[6721] <= 1'b0;
     layer2_out[6722] <= ~layer1_out[10342];
     layer2_out[6723] <= ~layer1_out[6938] | layer1_out[6937];
     layer2_out[6724] <= ~layer1_out[10516];
     layer2_out[6725] <= ~layer1_out[4422];
     layer2_out[6726] <= layer1_out[296];
     layer2_out[6727] <= ~(layer1_out[10171] & layer1_out[10172]);
     layer2_out[6728] <= layer1_out[6130] & layer1_out[6131];
     layer2_out[6729] <= layer1_out[1318];
     layer2_out[6730] <= ~layer1_out[5290];
     layer2_out[6731] <= ~layer1_out[6521];
     layer2_out[6732] <= ~layer1_out[2522] | layer1_out[2521];
     layer2_out[6733] <= ~layer1_out[10344] | layer1_out[10343];
     layer2_out[6734] <= ~layer1_out[1878] | layer1_out[1879];
     layer2_out[6735] <= ~layer1_out[7303];
     layer2_out[6736] <= ~layer1_out[7526];
     layer2_out[6737] <= layer1_out[9936] | layer1_out[9937];
     layer2_out[6738] <= ~layer1_out[2771];
     layer2_out[6739] <= ~layer1_out[7595];
     layer2_out[6740] <= ~layer1_out[4906];
     layer2_out[6741] <= ~layer1_out[5604];
     layer2_out[6742] <= ~layer1_out[6074] | layer1_out[6073];
     layer2_out[6743] <= layer1_out[6344] & ~layer1_out[6345];
     layer2_out[6744] <= layer1_out[7005] & ~layer1_out[7004];
     layer2_out[6745] <= layer1_out[2113];
     layer2_out[6746] <= layer1_out[1239];
     layer2_out[6747] <= ~layer1_out[6570];
     layer2_out[6748] <= layer1_out[1094];
     layer2_out[6749] <= ~(layer1_out[2817] | layer1_out[2818]);
     layer2_out[6750] <= ~layer1_out[6094];
     layer2_out[6751] <= ~layer1_out[11922];
     layer2_out[6752] <= layer1_out[1336] & layer1_out[1337];
     layer2_out[6753] <= ~layer1_out[11097];
     layer2_out[6754] <= ~(layer1_out[7707] | layer1_out[7708]);
     layer2_out[6755] <= ~layer1_out[5512] | layer1_out[5511];
     layer2_out[6756] <= ~layer1_out[840];
     layer2_out[6757] <= ~layer1_out[6026];
     layer2_out[6758] <= ~layer1_out[11736];
     layer2_out[6759] <= layer1_out[8186];
     layer2_out[6760] <= ~(layer1_out[11420] & layer1_out[11421]);
     layer2_out[6761] <= ~(layer1_out[11119] | layer1_out[11120]);
     layer2_out[6762] <= layer1_out[10239];
     layer2_out[6763] <= ~(layer1_out[3392] ^ layer1_out[3393]);
     layer2_out[6764] <= ~layer1_out[2578];
     layer2_out[6765] <= ~(layer1_out[8048] & layer1_out[8049]);
     layer2_out[6766] <= ~layer1_out[11080] | layer1_out[11081];
     layer2_out[6767] <= layer1_out[3943] | layer1_out[3944];
     layer2_out[6768] <= layer1_out[2092];
     layer2_out[6769] <= layer1_out[7734] & ~layer1_out[7733];
     layer2_out[6770] <= layer1_out[4230] & layer1_out[4231];
     layer2_out[6771] <= ~(layer1_out[11182] ^ layer1_out[11183]);
     layer2_out[6772] <= layer1_out[2031] & ~layer1_out[2032];
     layer2_out[6773] <= layer1_out[4138];
     layer2_out[6774] <= layer1_out[11371] & ~layer1_out[11372];
     layer2_out[6775] <= ~layer1_out[4025];
     layer2_out[6776] <= layer1_out[11155];
     layer2_out[6777] <= ~layer1_out[10855];
     layer2_out[6778] <= layer1_out[5736];
     layer2_out[6779] <= layer1_out[5881] & layer1_out[5882];
     layer2_out[6780] <= ~layer1_out[3950];
     layer2_out[6781] <= layer1_out[1444] & layer1_out[1445];
     layer2_out[6782] <= layer1_out[517] & ~layer1_out[516];
     layer2_out[6783] <= layer1_out[3203] & ~layer1_out[3204];
     layer2_out[6784] <= 1'b1;
     layer2_out[6785] <= layer1_out[11381];
     layer2_out[6786] <= ~layer1_out[7349] | layer1_out[7348];
     layer2_out[6787] <= ~layer1_out[9881];
     layer2_out[6788] <= layer1_out[3298];
     layer2_out[6789] <= ~(layer1_out[3415] ^ layer1_out[3416]);
     layer2_out[6790] <= ~layer1_out[226] | layer1_out[225];
     layer2_out[6791] <= ~layer1_out[6215] | layer1_out[6214];
     layer2_out[6792] <= layer1_out[722] & ~layer1_out[721];
     layer2_out[6793] <= layer1_out[5820] & ~layer1_out[5819];
     layer2_out[6794] <= ~layer1_out[9881];
     layer2_out[6795] <= layer1_out[3847];
     layer2_out[6796] <= ~layer1_out[5647];
     layer2_out[6797] <= layer1_out[1927] & layer1_out[1928];
     layer2_out[6798] <= ~(layer1_out[11177] & layer1_out[11178]);
     layer2_out[6799] <= layer1_out[8984];
     layer2_out[6800] <= layer1_out[9722];
     layer2_out[6801] <= ~(layer1_out[11385] ^ layer1_out[11386]);
     layer2_out[6802] <= layer1_out[1316] & ~layer1_out[1317];
     layer2_out[6803] <= layer1_out[11303] & ~layer1_out[11304];
     layer2_out[6804] <= layer1_out[4022];
     layer2_out[6805] <= ~layer1_out[8621] | layer1_out[8620];
     layer2_out[6806] <= 1'b0;
     layer2_out[6807] <= ~(layer1_out[9914] & layer1_out[9915]);
     layer2_out[6808] <= layer1_out[1524] & ~layer1_out[1523];
     layer2_out[6809] <= layer1_out[3016];
     layer2_out[6810] <= ~layer1_out[3666] | layer1_out[3667];
     layer2_out[6811] <= layer1_out[1996] & layer1_out[1997];
     layer2_out[6812] <= layer1_out[10599] & ~layer1_out[10598];
     layer2_out[6813] <= ~(layer1_out[11290] ^ layer1_out[11291]);
     layer2_out[6814] <= layer1_out[8458] & layer1_out[8459];
     layer2_out[6815] <= ~(layer1_out[10336] | layer1_out[10337]);
     layer2_out[6816] <= layer1_out[7856];
     layer2_out[6817] <= layer1_out[6240];
     layer2_out[6818] <= layer1_out[508];
     layer2_out[6819] <= layer1_out[8022] & ~layer1_out[8021];
     layer2_out[6820] <= layer1_out[8960];
     layer2_out[6821] <= ~layer1_out[7276];
     layer2_out[6822] <= ~(layer1_out[10786] ^ layer1_out[10787]);
     layer2_out[6823] <= ~layer1_out[4084] | layer1_out[4085];
     layer2_out[6824] <= ~layer1_out[4913];
     layer2_out[6825] <= ~layer1_out[733];
     layer2_out[6826] <= layer1_out[160] | layer1_out[161];
     layer2_out[6827] <= ~layer1_out[3259];
     layer2_out[6828] <= layer1_out[8155];
     layer2_out[6829] <= ~layer1_out[2571];
     layer2_out[6830] <= ~(layer1_out[9374] & layer1_out[9375]);
     layer2_out[6831] <= 1'b1;
     layer2_out[6832] <= layer1_out[11972] | layer1_out[11973];
     layer2_out[6833] <= layer1_out[11446];
     layer2_out[6834] <= ~layer1_out[6312] | layer1_out[6313];
     layer2_out[6835] <= ~(layer1_out[10952] | layer1_out[10953]);
     layer2_out[6836] <= layer1_out[7937] & ~layer1_out[7938];
     layer2_out[6837] <= layer1_out[8364];
     layer2_out[6838] <= ~layer1_out[11042];
     layer2_out[6839] <= ~layer1_out[7813];
     layer2_out[6840] <= layer1_out[7216] ^ layer1_out[7217];
     layer2_out[6841] <= layer1_out[4644];
     layer2_out[6842] <= layer1_out[3167] ^ layer1_out[3168];
     layer2_out[6843] <= layer1_out[5186];
     layer2_out[6844] <= ~layer1_out[2364];
     layer2_out[6845] <= layer1_out[3466];
     layer2_out[6846] <= ~layer1_out[2443];
     layer2_out[6847] <= ~(layer1_out[3705] ^ layer1_out[3706]);
     layer2_out[6848] <= ~layer1_out[1017];
     layer2_out[6849] <= ~layer1_out[5143] | layer1_out[5142];
     layer2_out[6850] <= ~layer1_out[7066];
     layer2_out[6851] <= 1'b0;
     layer2_out[6852] <= layer1_out[11819];
     layer2_out[6853] <= ~layer1_out[5924];
     layer2_out[6854] <= ~layer1_out[10167];
     layer2_out[6855] <= ~layer1_out[10280] | layer1_out[10281];
     layer2_out[6856] <= ~(layer1_out[1144] & layer1_out[1145]);
     layer2_out[6857] <= layer1_out[8888] & layer1_out[8889];
     layer2_out[6858] <= ~layer1_out[9041];
     layer2_out[6859] <= layer1_out[2104];
     layer2_out[6860] <= ~(layer1_out[9383] & layer1_out[9384]);
     layer2_out[6861] <= ~layer1_out[6447] | layer1_out[6446];
     layer2_out[6862] <= layer1_out[372] & ~layer1_out[373];
     layer2_out[6863] <= layer1_out[10122] ^ layer1_out[10123];
     layer2_out[6864] <= ~(layer1_out[3546] | layer1_out[3547]);
     layer2_out[6865] <= ~(layer1_out[11206] | layer1_out[11207]);
     layer2_out[6866] <= layer1_out[1056] ^ layer1_out[1057];
     layer2_out[6867] <= ~(layer1_out[333] | layer1_out[334]);
     layer2_out[6868] <= layer1_out[5683] & ~layer1_out[5682];
     layer2_out[6869] <= layer1_out[10010];
     layer2_out[6870] <= layer1_out[1921];
     layer2_out[6871] <= ~layer1_out[1938];
     layer2_out[6872] <= layer1_out[5136];
     layer2_out[6873] <= layer1_out[2533] & ~layer1_out[2534];
     layer2_out[6874] <= ~layer1_out[8158];
     layer2_out[6875] <= ~(layer1_out[9345] ^ layer1_out[9346]);
     layer2_out[6876] <= ~layer1_out[5892];
     layer2_out[6877] <= ~(layer1_out[4426] & layer1_out[4427]);
     layer2_out[6878] <= ~layer1_out[8822] | layer1_out[8823];
     layer2_out[6879] <= ~layer1_out[7767];
     layer2_out[6880] <= ~(layer1_out[8006] | layer1_out[8007]);
     layer2_out[6881] <= ~(layer1_out[2028] ^ layer1_out[2029]);
     layer2_out[6882] <= layer1_out[11902];
     layer2_out[6883] <= layer1_out[3793] | layer1_out[3794];
     layer2_out[6884] <= ~(layer1_out[154] ^ layer1_out[155]);
     layer2_out[6885] <= layer1_out[823] & ~layer1_out[824];
     layer2_out[6886] <= layer1_out[7891] | layer1_out[7892];
     layer2_out[6887] <= layer1_out[11088] & ~layer1_out[11087];
     layer2_out[6888] <= ~layer1_out[8742];
     layer2_out[6889] <= layer1_out[1996];
     layer2_out[6890] <= layer1_out[7964] | layer1_out[7965];
     layer2_out[6891] <= layer1_out[11035] | layer1_out[11036];
     layer2_out[6892] <= layer1_out[7033] & ~layer1_out[7034];
     layer2_out[6893] <= layer1_out[5896];
     layer2_out[6894] <= layer1_out[6885];
     layer2_out[6895] <= layer1_out[2296];
     layer2_out[6896] <= layer1_out[96];
     layer2_out[6897] <= layer1_out[4236];
     layer2_out[6898] <= ~(layer1_out[10994] & layer1_out[10995]);
     layer2_out[6899] <= layer1_out[109];
     layer2_out[6900] <= ~(layer1_out[1288] & layer1_out[1289]);
     layer2_out[6901] <= ~(layer1_out[6847] & layer1_out[6848]);
     layer2_out[6902] <= layer1_out[8148] & ~layer1_out[8149];
     layer2_out[6903] <= ~layer1_out[7311];
     layer2_out[6904] <= layer1_out[9795] | layer1_out[9796];
     layer2_out[6905] <= layer1_out[11680];
     layer2_out[6906] <= layer1_out[5796];
     layer2_out[6907] <= ~layer1_out[6290] | layer1_out[6289];
     layer2_out[6908] <= layer1_out[6576] | layer1_out[6577];
     layer2_out[6909] <= layer1_out[6919] & ~layer1_out[6918];
     layer2_out[6910] <= ~layer1_out[655];
     layer2_out[6911] <= ~(layer1_out[3159] | layer1_out[3160]);
     layer2_out[6912] <= ~layer1_out[7822] | layer1_out[7823];
     layer2_out[6913] <= layer1_out[4498] & ~layer1_out[4497];
     layer2_out[6914] <= ~layer1_out[11146] | layer1_out[11147];
     layer2_out[6915] <= layer1_out[3333];
     layer2_out[6916] <= ~layer1_out[8748];
     layer2_out[6917] <= layer1_out[10884] & ~layer1_out[10883];
     layer2_out[6918] <= layer1_out[9002] | layer1_out[9003];
     layer2_out[6919] <= layer1_out[8552];
     layer2_out[6920] <= layer1_out[11471] & ~layer1_out[11470];
     layer2_out[6921] <= layer1_out[855];
     layer2_out[6922] <= ~layer1_out[4023] | layer1_out[4024];
     layer2_out[6923] <= layer1_out[1208];
     layer2_out[6924] <= layer1_out[2805];
     layer2_out[6925] <= ~layer1_out[356];
     layer2_out[6926] <= ~layer1_out[7341];
     layer2_out[6927] <= ~layer1_out[4597];
     layer2_out[6928] <= ~layer1_out[11780] | layer1_out[11781];
     layer2_out[6929] <= layer1_out[512];
     layer2_out[6930] <= layer1_out[1530];
     layer2_out[6931] <= ~layer1_out[2722];
     layer2_out[6932] <= layer1_out[10681] & layer1_out[10682];
     layer2_out[6933] <= ~layer1_out[2745];
     layer2_out[6934] <= ~layer1_out[8182] | layer1_out[8181];
     layer2_out[6935] <= layer1_out[9957] ^ layer1_out[9958];
     layer2_out[6936] <= layer1_out[1134] ^ layer1_out[1135];
     layer2_out[6937] <= layer1_out[9763];
     layer2_out[6938] <= layer1_out[3976];
     layer2_out[6939] <= layer1_out[3344] & ~layer1_out[3343];
     layer2_out[6940] <= layer1_out[10342];
     layer2_out[6941] <= ~layer1_out[8108] | layer1_out[8109];
     layer2_out[6942] <= layer1_out[7911] | layer1_out[7912];
     layer2_out[6943] <= layer1_out[11755];
     layer2_out[6944] <= ~layer1_out[2653];
     layer2_out[6945] <= ~layer1_out[5877] | layer1_out[5876];
     layer2_out[6946] <= layer1_out[3449] ^ layer1_out[3450];
     layer2_out[6947] <= 1'b0;
     layer2_out[6948] <= ~layer1_out[3443];
     layer2_out[6949] <= ~layer1_out[5527];
     layer2_out[6950] <= layer1_out[9940] & ~layer1_out[9941];
     layer2_out[6951] <= ~(layer1_out[2359] & layer1_out[2360]);
     layer2_out[6952] <= layer1_out[7531];
     layer2_out[6953] <= ~(layer1_out[3135] ^ layer1_out[3136]);
     layer2_out[6954] <= ~layer1_out[9738] | layer1_out[9737];
     layer2_out[6955] <= ~layer1_out[8890];
     layer2_out[6956] <= layer1_out[6900] ^ layer1_out[6901];
     layer2_out[6957] <= ~(layer1_out[457] ^ layer1_out[458]);
     layer2_out[6958] <= ~(layer1_out[7680] ^ layer1_out[7681]);
     layer2_out[6959] <= ~(layer1_out[8885] & layer1_out[8886]);
     layer2_out[6960] <= layer1_out[4709] ^ layer1_out[4710];
     layer2_out[6961] <= layer1_out[5805] | layer1_out[5806];
     layer2_out[6962] <= ~layer1_out[10398];
     layer2_out[6963] <= ~layer1_out[8651] | layer1_out[8652];
     layer2_out[6964] <= layer1_out[758] & ~layer1_out[757];
     layer2_out[6965] <= ~(layer1_out[9844] | layer1_out[9845]);
     layer2_out[6966] <= ~(layer1_out[6780] & layer1_out[6781]);
     layer2_out[6967] <= ~(layer1_out[10146] & layer1_out[10147]);
     layer2_out[6968] <= ~layer1_out[4387] | layer1_out[4386];
     layer2_out[6969] <= ~(layer1_out[3939] & layer1_out[3940]);
     layer2_out[6970] <= layer1_out[3210];
     layer2_out[6971] <= layer1_out[10537] & layer1_out[10538];
     layer2_out[6972] <= layer1_out[8251] & layer1_out[8252];
     layer2_out[6973] <= ~layer1_out[2333] | layer1_out[2332];
     layer2_out[6974] <= ~layer1_out[9408];
     layer2_out[6975] <= ~layer1_out[1442];
     layer2_out[6976] <= ~layer1_out[8383];
     layer2_out[6977] <= layer1_out[165];
     layer2_out[6978] <= layer1_out[5910] | layer1_out[5911];
     layer2_out[6979] <= layer1_out[9717] ^ layer1_out[9718];
     layer2_out[6980] <= layer1_out[5178] | layer1_out[5179];
     layer2_out[6981] <= layer1_out[2098] | layer1_out[2099];
     layer2_out[6982] <= layer1_out[11515];
     layer2_out[6983] <= ~layer1_out[10933];
     layer2_out[6984] <= ~layer1_out[7657] | layer1_out[7656];
     layer2_out[6985] <= ~(layer1_out[10841] | layer1_out[10842]);
     layer2_out[6986] <= layer1_out[8369];
     layer2_out[6987] <= layer1_out[8554];
     layer2_out[6988] <= layer1_out[1381] & ~layer1_out[1380];
     layer2_out[6989] <= layer1_out[5993];
     layer2_out[6990] <= layer1_out[2934] | layer1_out[2935];
     layer2_out[6991] <= layer1_out[7424] & ~layer1_out[7425];
     layer2_out[6992] <= ~(layer1_out[5423] | layer1_out[5424]);
     layer2_out[6993] <= ~(layer1_out[1172] & layer1_out[1173]);
     layer2_out[6994] <= ~layer1_out[3022];
     layer2_out[6995] <= layer1_out[6019];
     layer2_out[6996] <= layer1_out[1810] ^ layer1_out[1811];
     layer2_out[6997] <= layer1_out[5961];
     layer2_out[6998] <= layer1_out[296] & ~layer1_out[297];
     layer2_out[6999] <= layer1_out[5901];
     layer2_out[7000] <= layer1_out[3613];
     layer2_out[7001] <= ~layer1_out[6107];
     layer2_out[7002] <= ~layer1_out[6303] | layer1_out[6304];
     layer2_out[7003] <= layer1_out[2841];
     layer2_out[7004] <= ~(layer1_out[725] | layer1_out[726]);
     layer2_out[7005] <= ~layer1_out[236] | layer1_out[235];
     layer2_out[7006] <= layer1_out[4727];
     layer2_out[7007] <= layer1_out[6338] & ~layer1_out[6337];
     layer2_out[7008] <= layer1_out[2828] & layer1_out[2829];
     layer2_out[7009] <= layer1_out[8459] & layer1_out[8460];
     layer2_out[7010] <= ~(layer1_out[10392] & layer1_out[10393]);
     layer2_out[7011] <= layer1_out[3505] | layer1_out[3506];
     layer2_out[7012] <= layer1_out[11144] & ~layer1_out[11143];
     layer2_out[7013] <= ~layer1_out[5417] | layer1_out[5418];
     layer2_out[7014] <= layer1_out[7607];
     layer2_out[7015] <= layer1_out[7178] & layer1_out[7179];
     layer2_out[7016] <= layer1_out[11281] | layer1_out[11282];
     layer2_out[7017] <= layer1_out[2815];
     layer2_out[7018] <= layer1_out[9384] & ~layer1_out[9385];
     layer2_out[7019] <= layer1_out[4226] & layer1_out[4227];
     layer2_out[7020] <= layer1_out[17] & layer1_out[18];
     layer2_out[7021] <= ~layer1_out[3897] | layer1_out[3898];
     layer2_out[7022] <= ~layer1_out[6342];
     layer2_out[7023] <= layer1_out[9382];
     layer2_out[7024] <= layer1_out[6771];
     layer2_out[7025] <= layer1_out[1802];
     layer2_out[7026] <= layer1_out[3876] | layer1_out[3877];
     layer2_out[7027] <= layer1_out[329] & ~layer1_out[328];
     layer2_out[7028] <= ~(layer1_out[2203] ^ layer1_out[2204]);
     layer2_out[7029] <= ~(layer1_out[9852] | layer1_out[9853]);
     layer2_out[7030] <= 1'b0;
     layer2_out[7031] <= layer1_out[10258];
     layer2_out[7032] <= ~layer1_out[7929];
     layer2_out[7033] <= ~(layer1_out[10745] & layer1_out[10746]);
     layer2_out[7034] <= layer1_out[10963] | layer1_out[10964];
     layer2_out[7035] <= ~layer1_out[7801] | layer1_out[7800];
     layer2_out[7036] <= layer1_out[11204];
     layer2_out[7037] <= ~layer1_out[439] | layer1_out[440];
     layer2_out[7038] <= layer1_out[1872] & layer1_out[1873];
     layer2_out[7039] <= ~layer1_out[9255] | layer1_out[9254];
     layer2_out[7040] <= layer1_out[6959] & ~layer1_out[6960];
     layer2_out[7041] <= ~layer1_out[4896] | layer1_out[4895];
     layer2_out[7042] <= ~layer1_out[2145];
     layer2_out[7043] <= layer1_out[7528] & layer1_out[7529];
     layer2_out[7044] <= layer1_out[7948];
     layer2_out[7045] <= ~(layer1_out[1720] ^ layer1_out[1721]);
     layer2_out[7046] <= ~layer1_out[4862];
     layer2_out[7047] <= layer1_out[4937] & ~layer1_out[4936];
     layer2_out[7048] <= ~layer1_out[9481];
     layer2_out[7049] <= layer1_out[11325];
     layer2_out[7050] <= layer1_out[7188] | layer1_out[7189];
     layer2_out[7051] <= ~layer1_out[7613];
     layer2_out[7052] <= layer1_out[2660];
     layer2_out[7053] <= layer1_out[1766];
     layer2_out[7054] <= ~layer1_out[11828] | layer1_out[11829];
     layer2_out[7055] <= layer1_out[11347] ^ layer1_out[11348];
     layer2_out[7056] <= ~(layer1_out[8000] & layer1_out[8001]);
     layer2_out[7057] <= layer1_out[7369] | layer1_out[7370];
     layer2_out[7058] <= ~layer1_out[2488];
     layer2_out[7059] <= layer1_out[9040] & ~layer1_out[9041];
     layer2_out[7060] <= layer1_out[217];
     layer2_out[7061] <= ~(layer1_out[11036] | layer1_out[11037]);
     layer2_out[7062] <= ~layer1_out[5056] | layer1_out[5057];
     layer2_out[7063] <= layer1_out[11314];
     layer2_out[7064] <= ~layer1_out[11471] | layer1_out[11472];
     layer2_out[7065] <= layer1_out[661];
     layer2_out[7066] <= ~layer1_out[1977];
     layer2_out[7067] <= ~layer1_out[6140];
     layer2_out[7068] <= layer1_out[8884] ^ layer1_out[8885];
     layer2_out[7069] <= ~layer1_out[942];
     layer2_out[7070] <= layer1_out[9147];
     layer2_out[7071] <= layer1_out[8198];
     layer2_out[7072] <= 1'b1;
     layer2_out[7073] <= ~layer1_out[3455];
     layer2_out[7074] <= ~(layer1_out[8248] & layer1_out[8249]);
     layer2_out[7075] <= ~(layer1_out[2996] ^ layer1_out[2997]);
     layer2_out[7076] <= layer1_out[724] ^ layer1_out[725];
     layer2_out[7077] <= layer1_out[6401] ^ layer1_out[6402];
     layer2_out[7078] <= ~(layer1_out[8699] | layer1_out[8700]);
     layer2_out[7079] <= layer1_out[8789] ^ layer1_out[8790];
     layer2_out[7080] <= ~(layer1_out[6572] | layer1_out[6573]);
     layer2_out[7081] <= layer1_out[8342] ^ layer1_out[8343];
     layer2_out[7082] <= ~(layer1_out[5377] & layer1_out[5378]);
     layer2_out[7083] <= layer1_out[591] & ~layer1_out[590];
     layer2_out[7084] <= layer1_out[3694] & ~layer1_out[3695];
     layer2_out[7085] <= ~(layer1_out[9559] ^ layer1_out[9560]);
     layer2_out[7086] <= layer1_out[1136];
     layer2_out[7087] <= ~layer1_out[1993];
     layer2_out[7088] <= layer1_out[6509];
     layer2_out[7089] <= layer1_out[7409] ^ layer1_out[7410];
     layer2_out[7090] <= layer1_out[11798];
     layer2_out[7091] <= ~layer1_out[7064] | layer1_out[7063];
     layer2_out[7092] <= layer1_out[1945];
     layer2_out[7093] <= ~layer1_out[6099] | layer1_out[6098];
     layer2_out[7094] <= layer1_out[2865];
     layer2_out[7095] <= ~(layer1_out[6924] & layer1_out[6925]);
     layer2_out[7096] <= layer1_out[2] & layer1_out[3];
     layer2_out[7097] <= layer1_out[2977];
     layer2_out[7098] <= ~layer1_out[1816];
     layer2_out[7099] <= layer1_out[7374] & ~layer1_out[7375];
     layer2_out[7100] <= ~(layer1_out[945] & layer1_out[946]);
     layer2_out[7101] <= layer1_out[6591] | layer1_out[6592];
     layer2_out[7102] <= layer1_out[9243] | layer1_out[9244];
     layer2_out[7103] <= layer1_out[9341];
     layer2_out[7104] <= layer1_out[4551];
     layer2_out[7105] <= layer1_out[10811] & layer1_out[10812];
     layer2_out[7106] <= ~layer1_out[11787] | layer1_out[11786];
     layer2_out[7107] <= ~(layer1_out[3841] & layer1_out[3842]);
     layer2_out[7108] <= ~layer1_out[1789];
     layer2_out[7109] <= ~(layer1_out[310] & layer1_out[311]);
     layer2_out[7110] <= ~layer1_out[7604];
     layer2_out[7111] <= layer1_out[1535] & ~layer1_out[1536];
     layer2_out[7112] <= layer1_out[2496] & ~layer1_out[2495];
     layer2_out[7113] <= layer1_out[5583];
     layer2_out[7114] <= layer1_out[9787];
     layer2_out[7115] <= layer1_out[7351] | layer1_out[7352];
     layer2_out[7116] <= layer1_out[11361] & ~layer1_out[11362];
     layer2_out[7117] <= layer1_out[5556] | layer1_out[5557];
     layer2_out[7118] <= layer1_out[8488] | layer1_out[8489];
     layer2_out[7119] <= layer1_out[4029] & layer1_out[4030];
     layer2_out[7120] <= layer1_out[9034] & ~layer1_out[9033];
     layer2_out[7121] <= ~(layer1_out[7318] & layer1_out[7319]);
     layer2_out[7122] <= layer1_out[8058];
     layer2_out[7123] <= layer1_out[11483];
     layer2_out[7124] <= layer1_out[9389] ^ layer1_out[9390];
     layer2_out[7125] <= ~layer1_out[9077];
     layer2_out[7126] <= layer1_out[5311];
     layer2_out[7127] <= ~layer1_out[9206];
     layer2_out[7128] <= ~(layer1_out[5835] & layer1_out[5836]);
     layer2_out[7129] <= ~layer1_out[357] | layer1_out[358];
     layer2_out[7130] <= ~(layer1_out[5424] | layer1_out[5425]);
     layer2_out[7131] <= layer1_out[9038];
     layer2_out[7132] <= ~(layer1_out[5041] | layer1_out[5042]);
     layer2_out[7133] <= ~(layer1_out[9592] ^ layer1_out[9593]);
     layer2_out[7134] <= ~layer1_out[962] | layer1_out[963];
     layer2_out[7135] <= 1'b0;
     layer2_out[7136] <= layer1_out[4603];
     layer2_out[7137] <= ~layer1_out[10927];
     layer2_out[7138] <= layer1_out[3465] & ~layer1_out[3464];
     layer2_out[7139] <= layer1_out[5802] ^ layer1_out[5803];
     layer2_out[7140] <= layer1_out[10927];
     layer2_out[7141] <= layer1_out[3245] & ~layer1_out[3246];
     layer2_out[7142] <= layer1_out[7638] & ~layer1_out[7637];
     layer2_out[7143] <= layer1_out[10257] ^ layer1_out[10258];
     layer2_out[7144] <= ~layer1_out[8096];
     layer2_out[7145] <= ~(layer1_out[3405] | layer1_out[3406]);
     layer2_out[7146] <= ~(layer1_out[4594] & layer1_out[4595]);
     layer2_out[7147] <= layer1_out[2246] & ~layer1_out[2245];
     layer2_out[7148] <= ~layer1_out[10236] | layer1_out[10235];
     layer2_out[7149] <= ~layer1_out[7627] | layer1_out[7626];
     layer2_out[7150] <= ~layer1_out[10829];
     layer2_out[7151] <= ~layer1_out[9691];
     layer2_out[7152] <= 1'b0;
     layer2_out[7153] <= ~(layer1_out[6111] & layer1_out[6112]);
     layer2_out[7154] <= ~layer1_out[1886];
     layer2_out[7155] <= layer1_out[3579];
     layer2_out[7156] <= ~(layer1_out[2901] ^ layer1_out[2902]);
     layer2_out[7157] <= layer1_out[9334] & ~layer1_out[9335];
     layer2_out[7158] <= layer1_out[7549] | layer1_out[7550];
     layer2_out[7159] <= ~(layer1_out[1486] | layer1_out[1487]);
     layer2_out[7160] <= ~layer1_out[9424];
     layer2_out[7161] <= layer1_out[7804];
     layer2_out[7162] <= layer1_out[1139];
     layer2_out[7163] <= layer1_out[2809];
     layer2_out[7164] <= layer1_out[1783];
     layer2_out[7165] <= layer1_out[10091] & ~layer1_out[10090];
     layer2_out[7166] <= layer1_out[7238] | layer1_out[7239];
     layer2_out[7167] <= ~layer1_out[2762] | layer1_out[2763];
     layer2_out[7168] <= ~layer1_out[3318] | layer1_out[3319];
     layer2_out[7169] <= layer1_out[1607] & ~layer1_out[1606];
     layer2_out[7170] <= ~(layer1_out[10475] & layer1_out[10476]);
     layer2_out[7171] <= layer1_out[11492] | layer1_out[11493];
     layer2_out[7172] <= layer1_out[6599] | layer1_out[6600];
     layer2_out[7173] <= layer1_out[1161] | layer1_out[1162];
     layer2_out[7174] <= layer1_out[10786] & ~layer1_out[10785];
     layer2_out[7175] <= layer1_out[3067];
     layer2_out[7176] <= layer1_out[4014];
     layer2_out[7177] <= layer1_out[9269] & ~layer1_out[9268];
     layer2_out[7178] <= ~layer1_out[0];
     layer2_out[7179] <= ~layer1_out[7360];
     layer2_out[7180] <= ~layer1_out[9640];
     layer2_out[7181] <= ~layer1_out[5510];
     layer2_out[7182] <= ~layer1_out[8462];
     layer2_out[7183] <= layer1_out[10791] & ~layer1_out[10792];
     layer2_out[7184] <= ~(layer1_out[2962] ^ layer1_out[2963]);
     layer2_out[7185] <= layer1_out[2719];
     layer2_out[7186] <= ~layer1_out[5358];
     layer2_out[7187] <= layer1_out[1047];
     layer2_out[7188] <= layer1_out[3853] & layer1_out[3854];
     layer2_out[7189] <= ~(layer1_out[4436] & layer1_out[4437]);
     layer2_out[7190] <= ~layer1_out[2863] | layer1_out[2862];
     layer2_out[7191] <= layer1_out[1700] ^ layer1_out[1701];
     layer2_out[7192] <= ~layer1_out[6810] | layer1_out[6811];
     layer2_out[7193] <= ~layer1_out[10589];
     layer2_out[7194] <= layer1_out[4625];
     layer2_out[7195] <= ~(layer1_out[1433] ^ layer1_out[1434]);
     layer2_out[7196] <= layer1_out[11401];
     layer2_out[7197] <= layer1_out[6046] | layer1_out[6047];
     layer2_out[7198] <= layer1_out[4342];
     layer2_out[7199] <= ~(layer1_out[7926] & layer1_out[7927]);
     layer2_out[7200] <= layer1_out[5039];
     layer2_out[7201] <= layer1_out[1077];
     layer2_out[7202] <= ~layer1_out[4206];
     layer2_out[7203] <= ~layer1_out[9891] | layer1_out[9890];
     layer2_out[7204] <= ~layer1_out[11136];
     layer2_out[7205] <= ~layer1_out[9295];
     layer2_out[7206] <= layer1_out[2815] & ~layer1_out[2816];
     layer2_out[7207] <= ~layer1_out[10520] | layer1_out[10521];
     layer2_out[7208] <= layer1_out[10047];
     layer2_out[7209] <= ~layer1_out[6837];
     layer2_out[7210] <= layer1_out[6395] & layer1_out[6396];
     layer2_out[7211] <= ~layer1_out[8506];
     layer2_out[7212] <= ~layer1_out[4427] | layer1_out[4428];
     layer2_out[7213] <= layer1_out[4905] | layer1_out[4906];
     layer2_out[7214] <= ~(layer1_out[2540] ^ layer1_out[2541]);
     layer2_out[7215] <= layer1_out[10151];
     layer2_out[7216] <= layer1_out[644] & layer1_out[645];
     layer2_out[7217] <= layer1_out[9790] & ~layer1_out[9789];
     layer2_out[7218] <= layer1_out[8280] | layer1_out[8281];
     layer2_out[7219] <= ~layer1_out[6420] | layer1_out[6419];
     layer2_out[7220] <= ~(layer1_out[2178] | layer1_out[2179]);
     layer2_out[7221] <= layer1_out[3530] & ~layer1_out[3531];
     layer2_out[7222] <= layer1_out[8977] & ~layer1_out[8978];
     layer2_out[7223] <= layer1_out[6800];
     layer2_out[7224] <= ~layer1_out[7182];
     layer2_out[7225] <= ~(layer1_out[9768] & layer1_out[9769]);
     layer2_out[7226] <= layer1_out[6073] & ~layer1_out[6072];
     layer2_out[7227] <= layer1_out[10113] & ~layer1_out[10112];
     layer2_out[7228] <= layer1_out[4836];
     layer2_out[7229] <= ~(layer1_out[3111] | layer1_out[3112]);
     layer2_out[7230] <= ~(layer1_out[4464] & layer1_out[4465]);
     layer2_out[7231] <= ~(layer1_out[7389] ^ layer1_out[7390]);
     layer2_out[7232] <= ~layer1_out[10571];
     layer2_out[7233] <= ~layer1_out[6509];
     layer2_out[7234] <= ~layer1_out[3402];
     layer2_out[7235] <= 1'b1;
     layer2_out[7236] <= layer1_out[7895];
     layer2_out[7237] <= layer1_out[9968];
     layer2_out[7238] <= layer1_out[285];
     layer2_out[7239] <= layer1_out[3240] & ~layer1_out[3241];
     layer2_out[7240] <= ~layer1_out[10863] | layer1_out[10862];
     layer2_out[7241] <= ~layer1_out[1287] | layer1_out[1288];
     layer2_out[7242] <= layer1_out[11020];
     layer2_out[7243] <= ~layer1_out[8181];
     layer2_out[7244] <= layer1_out[794];
     layer2_out[7245] <= layer1_out[1396] ^ layer1_out[1397];
     layer2_out[7246] <= ~layer1_out[6002];
     layer2_out[7247] <= layer1_out[9560] & ~layer1_out[9561];
     layer2_out[7248] <= ~layer1_out[3287];
     layer2_out[7249] <= layer1_out[6047] | layer1_out[6048];
     layer2_out[7250] <= layer1_out[10033];
     layer2_out[7251] <= layer1_out[6712];
     layer2_out[7252] <= ~layer1_out[3362] | layer1_out[3363];
     layer2_out[7253] <= layer1_out[8896];
     layer2_out[7254] <= ~layer1_out[1052];
     layer2_out[7255] <= ~layer1_out[4211] | layer1_out[4210];
     layer2_out[7256] <= layer1_out[5114];
     layer2_out[7257] <= layer1_out[10907] | layer1_out[10908];
     layer2_out[7258] <= layer1_out[6541];
     layer2_out[7259] <= layer1_out[8349];
     layer2_out[7260] <= layer1_out[5691];
     layer2_out[7261] <= ~(layer1_out[11833] | layer1_out[11834]);
     layer2_out[7262] <= layer1_out[477] | layer1_out[478];
     layer2_out[7263] <= layer1_out[4774] ^ layer1_out[4775];
     layer2_out[7264] <= layer1_out[8260];
     layer2_out[7265] <= ~layer1_out[1370];
     layer2_out[7266] <= ~layer1_out[2347];
     layer2_out[7267] <= layer1_out[10516] & ~layer1_out[10515];
     layer2_out[7268] <= ~layer1_out[9705] | layer1_out[9706];
     layer2_out[7269] <= ~layer1_out[10751] | layer1_out[10750];
     layer2_out[7270] <= ~layer1_out[6556];
     layer2_out[7271] <= ~(layer1_out[3252] | layer1_out[3253]);
     layer2_out[7272] <= ~(layer1_out[10618] & layer1_out[10619]);
     layer2_out[7273] <= ~(layer1_out[10175] | layer1_out[10176]);
     layer2_out[7274] <= ~(layer1_out[8347] ^ layer1_out[8348]);
     layer2_out[7275] <= layer1_out[10296] & ~layer1_out[10295];
     layer2_out[7276] <= ~(layer1_out[8317] | layer1_out[8318]);
     layer2_out[7277] <= ~layer1_out[9174] | layer1_out[9173];
     layer2_out[7278] <= layer1_out[5008] ^ layer1_out[5009];
     layer2_out[7279] <= layer1_out[8200] & ~layer1_out[8201];
     layer2_out[7280] <= ~layer1_out[9861];
     layer2_out[7281] <= ~(layer1_out[3103] & layer1_out[3104]);
     layer2_out[7282] <= 1'b1;
     layer2_out[7283] <= layer1_out[851];
     layer2_out[7284] <= layer1_out[11648] ^ layer1_out[11649];
     layer2_out[7285] <= ~(layer1_out[172] & layer1_out[173]);
     layer2_out[7286] <= ~layer1_out[922] | layer1_out[921];
     layer2_out[7287] <= ~layer1_out[1285] | layer1_out[1286];
     layer2_out[7288] <= ~(layer1_out[10054] | layer1_out[10055]);
     layer2_out[7289] <= ~layer1_out[10387];
     layer2_out[7290] <= ~layer1_out[7942];
     layer2_out[7291] <= ~layer1_out[7041] | layer1_out[7040];
     layer2_out[7292] <= layer1_out[6966];
     layer2_out[7293] <= ~(layer1_out[4181] & layer1_out[4182]);
     layer2_out[7294] <= layer1_out[10660] & ~layer1_out[10661];
     layer2_out[7295] <= layer1_out[6144] & ~layer1_out[6143];
     layer2_out[7296] <= layer1_out[11160] ^ layer1_out[11161];
     layer2_out[7297] <= layer1_out[7963] ^ layer1_out[7964];
     layer2_out[7298] <= layer1_out[2061];
     layer2_out[7299] <= layer1_out[7223];
     layer2_out[7300] <= layer1_out[481] | layer1_out[482];
     layer2_out[7301] <= layer1_out[6084] & ~layer1_out[6083];
     layer2_out[7302] <= layer1_out[6117] & layer1_out[6118];
     layer2_out[7303] <= layer1_out[1359];
     layer2_out[7304] <= ~layer1_out[3818];
     layer2_out[7305] <= layer1_out[1608] & ~layer1_out[1609];
     layer2_out[7306] <= ~layer1_out[5682];
     layer2_out[7307] <= ~layer1_out[3179] | layer1_out[3178];
     layer2_out[7308] <= ~layer1_out[6840] | layer1_out[6839];
     layer2_out[7309] <= ~layer1_out[6732];
     layer2_out[7310] <= layer1_out[8814];
     layer2_out[7311] <= ~layer1_out[11770] | layer1_out[11769];
     layer2_out[7312] <= layer1_out[5975] | layer1_out[5976];
     layer2_out[7313] <= ~(layer1_out[4498] ^ layer1_out[4499]);
     layer2_out[7314] <= ~layer1_out[1014] | layer1_out[1013];
     layer2_out[7315] <= ~(layer1_out[10869] & layer1_out[10870]);
     layer2_out[7316] <= ~(layer1_out[5608] & layer1_out[5609]);
     layer2_out[7317] <= ~(layer1_out[2364] | layer1_out[2365]);
     layer2_out[7318] <= layer1_out[1170] | layer1_out[1171];
     layer2_out[7319] <= ~layer1_out[4162];
     layer2_out[7320] <= layer1_out[429];
     layer2_out[7321] <= layer1_out[3762] & ~layer1_out[3761];
     layer2_out[7322] <= layer1_out[11792] | layer1_out[11793];
     layer2_out[7323] <= ~(layer1_out[11067] & layer1_out[11068]);
     layer2_out[7324] <= layer1_out[11617] & ~layer1_out[11616];
     layer2_out[7325] <= layer1_out[11880] & layer1_out[11881];
     layer2_out[7326] <= 1'b1;
     layer2_out[7327] <= layer1_out[191];
     layer2_out[7328] <= ~layer1_out[11636];
     layer2_out[7329] <= ~layer1_out[3131];
     layer2_out[7330] <= ~layer1_out[5710];
     layer2_out[7331] <= layer1_out[5294];
     layer2_out[7332] <= ~layer1_out[8085] | layer1_out[8086];
     layer2_out[7333] <= ~(layer1_out[6475] ^ layer1_out[6476]);
     layer2_out[7334] <= ~(layer1_out[3532] ^ layer1_out[3533]);
     layer2_out[7335] <= layer1_out[10878] & layer1_out[10879];
     layer2_out[7336] <= layer1_out[9685];
     layer2_out[7337] <= layer1_out[1370] & ~layer1_out[1371];
     layer2_out[7338] <= ~layer1_out[5126];
     layer2_out[7339] <= layer1_out[552] | layer1_out[553];
     layer2_out[7340] <= layer1_out[2434];
     layer2_out[7341] <= layer1_out[7450] | layer1_out[7451];
     layer2_out[7342] <= layer1_out[394] & ~layer1_out[395];
     layer2_out[7343] <= layer1_out[3146] & layer1_out[3147];
     layer2_out[7344] <= layer1_out[9114];
     layer2_out[7345] <= ~layer1_out[5635];
     layer2_out[7346] <= ~layer1_out[10915];
     layer2_out[7347] <= ~layer1_out[1914] | layer1_out[1913];
     layer2_out[7348] <= layer1_out[1615];
     layer2_out[7349] <= 1'b0;
     layer2_out[7350] <= ~layer1_out[8369];
     layer2_out[7351] <= layer1_out[10232];
     layer2_out[7352] <= layer1_out[6333] & ~layer1_out[6334];
     layer2_out[7353] <= layer1_out[7068] | layer1_out[7069];
     layer2_out[7354] <= layer1_out[2042];
     layer2_out[7355] <= layer1_out[9203] ^ layer1_out[9204];
     layer2_out[7356] <= ~(layer1_out[8568] ^ layer1_out[8569]);
     layer2_out[7357] <= layer1_out[8734] & ~layer1_out[8735];
     layer2_out[7358] <= ~layer1_out[11554];
     layer2_out[7359] <= layer1_out[11300] | layer1_out[11301];
     layer2_out[7360] <= layer1_out[8264] & ~layer1_out[8263];
     layer2_out[7361] <= ~layer1_out[7870];
     layer2_out[7362] <= ~(layer1_out[11639] | layer1_out[11640]);
     layer2_out[7363] <= ~layer1_out[5887] | layer1_out[5886];
     layer2_out[7364] <= ~layer1_out[6153];
     layer2_out[7365] <= layer1_out[991] & layer1_out[992];
     layer2_out[7366] <= ~layer1_out[5128];
     layer2_out[7367] <= ~layer1_out[6238];
     layer2_out[7368] <= layer1_out[7922];
     layer2_out[7369] <= ~layer1_out[9435];
     layer2_out[7370] <= ~layer1_out[5765];
     layer2_out[7371] <= layer1_out[3508] ^ layer1_out[3509];
     layer2_out[7372] <= 1'b0;
     layer2_out[7373] <= ~layer1_out[2652] | layer1_out[2651];
     layer2_out[7374] <= layer1_out[7396] | layer1_out[7397];
     layer2_out[7375] <= ~layer1_out[2360] | layer1_out[2361];
     layer2_out[7376] <= layer1_out[11135] & ~layer1_out[11136];
     layer2_out[7377] <= layer1_out[11147] & ~layer1_out[11148];
     layer2_out[7378] <= ~layer1_out[9871];
     layer2_out[7379] <= layer1_out[2946] ^ layer1_out[2947];
     layer2_out[7380] <= ~layer1_out[3731] | layer1_out[3732];
     layer2_out[7381] <= ~(layer1_out[7054] & layer1_out[7055]);
     layer2_out[7382] <= layer1_out[8693] ^ layer1_out[8694];
     layer2_out[7383] <= layer1_out[9699] | layer1_out[9700];
     layer2_out[7384] <= layer1_out[6620] & ~layer1_out[6619];
     layer2_out[7385] <= 1'b1;
     layer2_out[7386] <= ~layer1_out[4627] | layer1_out[4626];
     layer2_out[7387] <= layer1_out[8123] & ~layer1_out[8124];
     layer2_out[7388] <= ~layer1_out[11310];
     layer2_out[7389] <= layer1_out[7240] | layer1_out[7241];
     layer2_out[7390] <= layer1_out[5839] & layer1_out[5840];
     layer2_out[7391] <= ~layer1_out[961];
     layer2_out[7392] <= layer1_out[3054] & layer1_out[3055];
     layer2_out[7393] <= layer1_out[405] & layer1_out[406];
     layer2_out[7394] <= layer1_out[11462];
     layer2_out[7395] <= layer1_out[5570] ^ layer1_out[5571];
     layer2_out[7396] <= ~layer1_out[5313] | layer1_out[5314];
     layer2_out[7397] <= layer1_out[7186] & ~layer1_out[7187];
     layer2_out[7398] <= ~(layer1_out[1037] | layer1_out[1038]);
     layer2_out[7399] <= ~layer1_out[9476] | layer1_out[9477];
     layer2_out[7400] <= ~layer1_out[7892];
     layer2_out[7401] <= layer1_out[2443];
     layer2_out[7402] <= ~layer1_out[7676] | layer1_out[7677];
     layer2_out[7403] <= ~layer1_out[7486];
     layer2_out[7404] <= layer1_out[2207];
     layer2_out[7405] <= ~(layer1_out[869] ^ layer1_out[870]);
     layer2_out[7406] <= layer1_out[7774];
     layer2_out[7407] <= ~layer1_out[5480] | layer1_out[5479];
     layer2_out[7408] <= ~layer1_out[8553] | layer1_out[8552];
     layer2_out[7409] <= 1'b0;
     layer2_out[7410] <= ~(layer1_out[2082] | layer1_out[2083]);
     layer2_out[7411] <= ~(layer1_out[9436] | layer1_out[9437]);
     layer2_out[7412] <= ~layer1_out[11625];
     layer2_out[7413] <= ~(layer1_out[7762] | layer1_out[7763]);
     layer2_out[7414] <= ~layer1_out[2577];
     layer2_out[7415] <= layer1_out[11724] & ~layer1_out[11723];
     layer2_out[7416] <= ~layer1_out[4066] | layer1_out[4065];
     layer2_out[7417] <= ~(layer1_out[9913] & layer1_out[9914]);
     layer2_out[7418] <= ~(layer1_out[11690] | layer1_out[11691]);
     layer2_out[7419] <= ~(layer1_out[1726] & layer1_out[1727]);
     layer2_out[7420] <= layer1_out[1747];
     layer2_out[7421] <= layer1_out[3649] & ~layer1_out[3650];
     layer2_out[7422] <= layer1_out[6175];
     layer2_out[7423] <= layer1_out[3379];
     layer2_out[7424] <= layer1_out[10027];
     layer2_out[7425] <= layer1_out[9429] ^ layer1_out[9430];
     layer2_out[7426] <= layer1_out[7688] | layer1_out[7689];
     layer2_out[7427] <= ~layer1_out[10847];
     layer2_out[7428] <= ~layer1_out[5677];
     layer2_out[7429] <= ~layer1_out[1207] | layer1_out[1206];
     layer2_out[7430] <= ~(layer1_out[5000] | layer1_out[5001]);
     layer2_out[7431] <= ~layer1_out[3969];
     layer2_out[7432] <= ~layer1_out[8467];
     layer2_out[7433] <= ~layer1_out[8136] | layer1_out[8135];
     layer2_out[7434] <= layer1_out[2515] & layer1_out[2516];
     layer2_out[7435] <= ~layer1_out[4425];
     layer2_out[7436] <= layer1_out[6775] ^ layer1_out[6776];
     layer2_out[7437] <= layer1_out[11354];
     layer2_out[7438] <= layer1_out[137];
     layer2_out[7439] <= layer1_out[2403];
     layer2_out[7440] <= layer1_out[3303] | layer1_out[3304];
     layer2_out[7441] <= ~layer1_out[6363];
     layer2_out[7442] <= ~layer1_out[11277] | layer1_out[11278];
     layer2_out[7443] <= 1'b0;
     layer2_out[7444] <= layer1_out[9004] & ~layer1_out[9003];
     layer2_out[7445] <= ~(layer1_out[9458] | layer1_out[9459]);
     layer2_out[7446] <= layer1_out[11927] & layer1_out[11928];
     layer2_out[7447] <= layer1_out[617];
     layer2_out[7448] <= layer1_out[9360] | layer1_out[9361];
     layer2_out[7449] <= ~(layer1_out[5124] | layer1_out[5125]);
     layer2_out[7450] <= layer1_out[88] & ~layer1_out[87];
     layer2_out[7451] <= ~layer1_out[929] | layer1_out[928];
     layer2_out[7452] <= layer1_out[10157] & layer1_out[10158];
     layer2_out[7453] <= ~(layer1_out[6064] ^ layer1_out[6065]);
     layer2_out[7454] <= layer1_out[7592] & ~layer1_out[7593];
     layer2_out[7455] <= layer1_out[7174];
     layer2_out[7456] <= ~layer1_out[7540];
     layer2_out[7457] <= layer1_out[343] & ~layer1_out[342];
     layer2_out[7458] <= ~layer1_out[8383];
     layer2_out[7459] <= layer1_out[9546];
     layer2_out[7460] <= layer1_out[6960] & ~layer1_out[6961];
     layer2_out[7461] <= layer1_out[6014];
     layer2_out[7462] <= ~layer1_out[11180];
     layer2_out[7463] <= layer1_out[4767] ^ layer1_out[4768];
     layer2_out[7464] <= ~(layer1_out[8448] | layer1_out[8449]);
     layer2_out[7465] <= layer1_out[4806] & layer1_out[4807];
     layer2_out[7466] <= layer1_out[6207] | layer1_out[6208];
     layer2_out[7467] <= layer1_out[9511];
     layer2_out[7468] <= layer1_out[10165];
     layer2_out[7469] <= layer1_out[3358] | layer1_out[3359];
     layer2_out[7470] <= ~(layer1_out[1120] & layer1_out[1121]);
     layer2_out[7471] <= ~layer1_out[3354];
     layer2_out[7472] <= layer1_out[10011];
     layer2_out[7473] <= layer1_out[1567];
     layer2_out[7474] <= ~layer1_out[8899];
     layer2_out[7475] <= layer1_out[10415] ^ layer1_out[10416];
     layer2_out[7476] <= layer1_out[7145];
     layer2_out[7477] <= layer1_out[4205];
     layer2_out[7478] <= ~(layer1_out[6777] | layer1_out[6778]);
     layer2_out[7479] <= layer1_out[1956] | layer1_out[1957];
     layer2_out[7480] <= ~layer1_out[4899] | layer1_out[4900];
     layer2_out[7481] <= layer1_out[140] & layer1_out[141];
     layer2_out[7482] <= layer1_out[1055];
     layer2_out[7483] <= ~layer1_out[7445] | layer1_out[7444];
     layer2_out[7484] <= ~(layer1_out[11394] & layer1_out[11395]);
     layer2_out[7485] <= ~layer1_out[3047];
     layer2_out[7486] <= layer1_out[6481] ^ layer1_out[6482];
     layer2_out[7487] <= ~layer1_out[5048];
     layer2_out[7488] <= layer1_out[120];
     layer2_out[7489] <= layer1_out[3161] | layer1_out[3162];
     layer2_out[7490] <= layer1_out[6041] & layer1_out[6042];
     layer2_out[7491] <= layer1_out[10174] & ~layer1_out[10175];
     layer2_out[7492] <= layer1_out[10876] ^ layer1_out[10877];
     layer2_out[7493] <= ~layer1_out[8149];
     layer2_out[7494] <= layer1_out[6913] & layer1_out[6914];
     layer2_out[7495] <= ~layer1_out[3125];
     layer2_out[7496] <= layer1_out[4457] & ~layer1_out[4456];
     layer2_out[7497] <= layer1_out[6468] & ~layer1_out[6467];
     layer2_out[7498] <= ~layer1_out[11140];
     layer2_out[7499] <= 1'b1;
     layer2_out[7500] <= layer1_out[3914] | layer1_out[3915];
     layer2_out[7501] <= ~layer1_out[4545];
     layer2_out[7502] <= layer1_out[2700] | layer1_out[2701];
     layer2_out[7503] <= layer1_out[2078] | layer1_out[2079];
     layer2_out[7504] <= ~(layer1_out[5247] ^ layer1_out[5248]);
     layer2_out[7505] <= layer1_out[5850] | layer1_out[5851];
     layer2_out[7506] <= layer1_out[11158] ^ layer1_out[11159];
     layer2_out[7507] <= layer1_out[3122] & ~layer1_out[3121];
     layer2_out[7508] <= layer1_out[3117] & layer1_out[3118];
     layer2_out[7509] <= ~layer1_out[10617] | layer1_out[10618];
     layer2_out[7510] <= ~layer1_out[7113];
     layer2_out[7511] <= layer1_out[6641];
     layer2_out[7512] <= layer1_out[4730] | layer1_out[4731];
     layer2_out[7513] <= ~layer1_out[3099];
     layer2_out[7514] <= layer1_out[4984] | layer1_out[4985];
     layer2_out[7515] <= layer1_out[7248] & ~layer1_out[7247];
     layer2_out[7516] <= layer1_out[668];
     layer2_out[7517] <= ~(layer1_out[8214] | layer1_out[8215]);
     layer2_out[7518] <= ~layer1_out[16] | layer1_out[15];
     layer2_out[7519] <= layer1_out[10001] & ~layer1_out[10002];
     layer2_out[7520] <= layer1_out[7432] | layer1_out[7433];
     layer2_out[7521] <= ~layer1_out[11109] | layer1_out[11110];
     layer2_out[7522] <= ~layer1_out[9887];
     layer2_out[7523] <= ~layer1_out[11399];
     layer2_out[7524] <= ~(layer1_out[10816] & layer1_out[10817]);
     layer2_out[7525] <= layer1_out[3640] & ~layer1_out[3641];
     layer2_out[7526] <= layer1_out[6126] ^ layer1_out[6127];
     layer2_out[7527] <= ~(layer1_out[4882] & layer1_out[4883]);
     layer2_out[7528] <= ~layer1_out[9369];
     layer2_out[7529] <= layer1_out[2020] ^ layer1_out[2021];
     layer2_out[7530] <= layer1_out[1899] & ~layer1_out[1898];
     layer2_out[7531] <= layer1_out[3170] & layer1_out[3171];
     layer2_out[7532] <= layer1_out[4199] & ~layer1_out[4200];
     layer2_out[7533] <= ~(layer1_out[5957] ^ layer1_out[5958]);
     layer2_out[7534] <= layer1_out[767];
     layer2_out[7535] <= ~layer1_out[3564];
     layer2_out[7536] <= ~(layer1_out[754] | layer1_out[755]);
     layer2_out[7537] <= ~layer1_out[6006];
     layer2_out[7538] <= ~layer1_out[6723] | layer1_out[6724];
     layer2_out[7539] <= ~(layer1_out[634] | layer1_out[635]);
     layer2_out[7540] <= ~(layer1_out[10541] | layer1_out[10542]);
     layer2_out[7541] <= ~(layer1_out[1524] & layer1_out[1525]);
     layer2_out[7542] <= ~layer1_out[10742] | layer1_out[10741];
     layer2_out[7543] <= ~(layer1_out[5798] & layer1_out[5799]);
     layer2_out[7544] <= ~layer1_out[6963];
     layer2_out[7545] <= layer1_out[10030] | layer1_out[10031];
     layer2_out[7546] <= ~(layer1_out[1228] ^ layer1_out[1229]);
     layer2_out[7547] <= ~layer1_out[713];
     layer2_out[7548] <= ~layer1_out[2780];
     layer2_out[7549] <= layer1_out[4438];
     layer2_out[7550] <= ~layer1_out[354];
     layer2_out[7551] <= ~layer1_out[9171];
     layer2_out[7552] <= layer1_out[2123];
     layer2_out[7553] <= layer1_out[167] | layer1_out[168];
     layer2_out[7554] <= ~layer1_out[7562];
     layer2_out[7555] <= ~layer1_out[11292];
     layer2_out[7556] <= ~(layer1_out[9098] & layer1_out[9099]);
     layer2_out[7557] <= layer1_out[5174] | layer1_out[5175];
     layer2_out[7558] <= layer1_out[4440] & ~layer1_out[4439];
     layer2_out[7559] <= layer1_out[5339] & ~layer1_out[5340];
     layer2_out[7560] <= ~(layer1_out[2064] | layer1_out[2065]);
     layer2_out[7561] <= ~layer1_out[9991];
     layer2_out[7562] <= layer1_out[6538];
     layer2_out[7563] <= ~layer1_out[11556];
     layer2_out[7564] <= ~layer1_out[2256] | layer1_out[2257];
     layer2_out[7565] <= ~(layer1_out[8278] | layer1_out[8279]);
     layer2_out[7566] <= ~layer1_out[11985];
     layer2_out[7567] <= layer1_out[11701] | layer1_out[11702];
     layer2_out[7568] <= ~(layer1_out[4587] | layer1_out[4588]);
     layer2_out[7569] <= layer1_out[318] & ~layer1_out[319];
     layer2_out[7570] <= ~layer1_out[58];
     layer2_out[7571] <= ~(layer1_out[5404] ^ layer1_out[5405]);
     layer2_out[7572] <= ~(layer1_out[3076] ^ layer1_out[3077]);
     layer2_out[7573] <= layer1_out[10538] & ~layer1_out[10539];
     layer2_out[7574] <= ~layer1_out[1041] | layer1_out[1040];
     layer2_out[7575] <= layer1_out[9361];
     layer2_out[7576] <= layer1_out[4647];
     layer2_out[7577] <= layer1_out[9877];
     layer2_out[7578] <= layer1_out[1848] & ~layer1_out[1849];
     layer2_out[7579] <= ~(layer1_out[4491] ^ layer1_out[4492]);
     layer2_out[7580] <= layer1_out[10769];
     layer2_out[7581] <= ~layer1_out[2224];
     layer2_out[7582] <= layer1_out[8079];
     layer2_out[7583] <= layer1_out[671] & layer1_out[672];
     layer2_out[7584] <= ~(layer1_out[5415] & layer1_out[5416]);
     layer2_out[7585] <= ~(layer1_out[958] & layer1_out[959]);
     layer2_out[7586] <= layer1_out[1830] & layer1_out[1831];
     layer2_out[7587] <= layer1_out[4660] | layer1_out[4661];
     layer2_out[7588] <= layer1_out[4592];
     layer2_out[7589] <= ~(layer1_out[1166] ^ layer1_out[1167]);
     layer2_out[7590] <= 1'b0;
     layer2_out[7591] <= ~layer1_out[7107];
     layer2_out[7592] <= layer1_out[2798] | layer1_out[2799];
     layer2_out[7593] <= layer1_out[4085];
     layer2_out[7594] <= ~layer1_out[5888] | layer1_out[5889];
     layer2_out[7595] <= layer1_out[917] & ~layer1_out[916];
     layer2_out[7596] <= ~layer1_out[6896];
     layer2_out[7597] <= ~layer1_out[9428] | layer1_out[9427];
     layer2_out[7598] <= ~layer1_out[5620];
     layer2_out[7599] <= ~layer1_out[10355];
     layer2_out[7600] <= layer1_out[2845] ^ layer1_out[2846];
     layer2_out[7601] <= layer1_out[11031];
     layer2_out[7602] <= layer1_out[9105];
     layer2_out[7603] <= ~(layer1_out[492] & layer1_out[493]);
     layer2_out[7604] <= ~layer1_out[7989];
     layer2_out[7605] <= ~layer1_out[8405] | layer1_out[8404];
     layer2_out[7606] <= layer1_out[1301];
     layer2_out[7607] <= layer1_out[3592];
     layer2_out[7608] <= layer1_out[11853] ^ layer1_out[11854];
     layer2_out[7609] <= layer1_out[543] | layer1_out[544];
     layer2_out[7610] <= ~(layer1_out[8773] & layer1_out[8774]);
     layer2_out[7611] <= ~(layer1_out[7209] | layer1_out[7210]);
     layer2_out[7612] <= ~layer1_out[9974];
     layer2_out[7613] <= ~layer1_out[11705];
     layer2_out[7614] <= ~(layer1_out[2599] ^ layer1_out[2600]);
     layer2_out[7615] <= layer1_out[3049] | layer1_out[3050];
     layer2_out[7616] <= ~layer1_out[9749];
     layer2_out[7617] <= ~layer1_out[5241] | layer1_out[5240];
     layer2_out[7618] <= layer1_out[11593] & layer1_out[11594];
     layer2_out[7619] <= layer1_out[6877] & ~layer1_out[6876];
     layer2_out[7620] <= layer1_out[10333];
     layer2_out[7621] <= ~layer1_out[6310];
     layer2_out[7622] <= ~layer1_out[10948];
     layer2_out[7623] <= layer1_out[9089] & ~layer1_out[9088];
     layer2_out[7624] <= ~layer1_out[1012];
     layer2_out[7625] <= layer1_out[1941] & layer1_out[1942];
     layer2_out[7626] <= layer1_out[11255] ^ layer1_out[11256];
     layer2_out[7627] <= ~(layer1_out[10359] | layer1_out[10360]);
     layer2_out[7628] <= ~layer1_out[5422];
     layer2_out[7629] <= ~layer1_out[256] | layer1_out[257];
     layer2_out[7630] <= layer1_out[4978] & ~layer1_out[4979];
     layer2_out[7631] <= ~layer1_out[6618];
     layer2_out[7632] <= ~(layer1_out[3418] ^ layer1_out[3419]);
     layer2_out[7633] <= layer1_out[5761] & ~layer1_out[5760];
     layer2_out[7634] <= layer1_out[1558];
     layer2_out[7635] <= ~layer1_out[10765];
     layer2_out[7636] <= ~(layer1_out[10659] ^ layer1_out[10660]);
     layer2_out[7637] <= layer1_out[9447] | layer1_out[9448];
     layer2_out[7638] <= ~layer1_out[773];
     layer2_out[7639] <= ~layer1_out[7435];
     layer2_out[7640] <= layer1_out[6151];
     layer2_out[7641] <= ~layer1_out[7722] | layer1_out[7721];
     layer2_out[7642] <= layer1_out[9984];
     layer2_out[7643] <= layer1_out[2318] & ~layer1_out[2317];
     layer2_out[7644] <= ~(layer1_out[846] & layer1_out[847]);
     layer2_out[7645] <= layer1_out[3461];
     layer2_out[7646] <= ~(layer1_out[11204] & layer1_out[11205]);
     layer2_out[7647] <= ~layer1_out[7177];
     layer2_out[7648] <= ~layer1_out[9392];
     layer2_out[7649] <= layer1_out[8912] | layer1_out[8913];
     layer2_out[7650] <= layer1_out[6636] | layer1_out[6637];
     layer2_out[7651] <= layer1_out[9963];
     layer2_out[7652] <= ~(layer1_out[10282] & layer1_out[10283]);
     layer2_out[7653] <= layer1_out[10917] & ~layer1_out[10918];
     layer2_out[7654] <= ~(layer1_out[10779] & layer1_out[10780]);
     layer2_out[7655] <= ~(layer1_out[7620] & layer1_out[7621]);
     layer2_out[7656] <= ~(layer1_out[4214] | layer1_out[4215]);
     layer2_out[7657] <= ~layer1_out[1363];
     layer2_out[7658] <= ~layer1_out[1352];
     layer2_out[7659] <= ~(layer1_out[8678] | layer1_out[8679]);
     layer2_out[7660] <= layer1_out[5891] | layer1_out[5892];
     layer2_out[7661] <= ~layer1_out[8840] | layer1_out[8839];
     layer2_out[7662] <= layer1_out[9793] & ~layer1_out[9794];
     layer2_out[7663] <= ~layer1_out[11234];
     layer2_out[7664] <= ~layer1_out[3504] | layer1_out[3503];
     layer2_out[7665] <= ~layer1_out[9113];
     layer2_out[7666] <= layer1_out[1088] & ~layer1_out[1087];
     layer2_out[7667] <= 1'b1;
     layer2_out[7668] <= layer1_out[10665] & layer1_out[10666];
     layer2_out[7669] <= layer1_out[8412];
     layer2_out[7670] <= layer1_out[8595] & ~layer1_out[8596];
     layer2_out[7671] <= ~layer1_out[9618] | layer1_out[9617];
     layer2_out[7672] <= layer1_out[3655];
     layer2_out[7673] <= ~layer1_out[1110] | layer1_out[1109];
     layer2_out[7674] <= layer1_out[7955] ^ layer1_out[7956];
     layer2_out[7675] <= layer1_out[10973] ^ layer1_out[10974];
     layer2_out[7676] <= layer1_out[7314] ^ layer1_out[7315];
     layer2_out[7677] <= layer1_out[4981] | layer1_out[4982];
     layer2_out[7678] <= ~(layer1_out[6995] ^ layer1_out[6996]);
     layer2_out[7679] <= layer1_out[6129] & ~layer1_out[6128];
     layer2_out[7680] <= layer1_out[7914];
     layer2_out[7681] <= ~layer1_out[8517];
     layer2_out[7682] <= ~(layer1_out[4006] & layer1_out[4007]);
     layer2_out[7683] <= layer1_out[3365] & layer1_out[3366];
     layer2_out[7684] <= ~layer1_out[10109];
     layer2_out[7685] <= layer1_out[8779] & ~layer1_out[8780];
     layer2_out[7686] <= ~layer1_out[6228];
     layer2_out[7687] <= ~layer1_out[11270];
     layer2_out[7688] <= ~layer1_out[6814];
     layer2_out[7689] <= ~layer1_out[8351];
     layer2_out[7690] <= layer1_out[6603] & ~layer1_out[6604];
     layer2_out[7691] <= layer1_out[5553] & ~layer1_out[5554];
     layer2_out[7692] <= ~(layer1_out[1968] ^ layer1_out[1969]);
     layer2_out[7693] <= layer1_out[9066];
     layer2_out[7694] <= ~layer1_out[6846];
     layer2_out[7695] <= layer1_out[10374];
     layer2_out[7696] <= ~(layer1_out[7321] & layer1_out[7322]);
     layer2_out[7697] <= layer1_out[7994] ^ layer1_out[7995];
     layer2_out[7698] <= ~layer1_out[3607];
     layer2_out[7699] <= ~layer1_out[4930] | layer1_out[4931];
     layer2_out[7700] <= ~layer1_out[7298] | layer1_out[7297];
     layer2_out[7701] <= layer1_out[1892] & layer1_out[1893];
     layer2_out[7702] <= ~layer1_out[7547];
     layer2_out[7703] <= layer1_out[3006];
     layer2_out[7704] <= ~(layer1_out[450] ^ layer1_out[451]);
     layer2_out[7705] <= layer1_out[2826] | layer1_out[2827];
     layer2_out[7706] <= ~layer1_out[11760];
     layer2_out[7707] <= layer1_out[9088] & ~layer1_out[9087];
     layer2_out[7708] <= layer1_out[5384];
     layer2_out[7709] <= ~(layer1_out[1943] ^ layer1_out[1944]);
     layer2_out[7710] <= layer1_out[7509] & ~layer1_out[7508];
     layer2_out[7711] <= ~layer1_out[4555];
     layer2_out[7712] <= ~(layer1_out[2849] | layer1_out[2850]);
     layer2_out[7713] <= layer1_out[6287] | layer1_out[6288];
     layer2_out[7714] <= ~(layer1_out[8132] & layer1_out[8133]);
     layer2_out[7715] <= ~layer1_out[10758];
     layer2_out[7716] <= layer1_out[5643] & ~layer1_out[5644];
     layer2_out[7717] <= ~(layer1_out[5405] ^ layer1_out[5406]);
     layer2_out[7718] <= layer1_out[2598] | layer1_out[2599];
     layer2_out[7719] <= layer1_out[6191];
     layer2_out[7720] <= ~(layer1_out[3907] & layer1_out[3908]);
     layer2_out[7721] <= layer1_out[7750];
     layer2_out[7722] <= ~layer1_out[6610];
     layer2_out[7723] <= ~(layer1_out[9735] | layer1_out[9736]);
     layer2_out[7724] <= ~(layer1_out[5586] & layer1_out[5587]);
     layer2_out[7725] <= layer1_out[10147] & ~layer1_out[10148];
     layer2_out[7726] <= layer1_out[4302];
     layer2_out[7727] <= ~layer1_out[4974];
     layer2_out[7728] <= layer1_out[7728] & layer1_out[7729];
     layer2_out[7729] <= ~layer1_out[1203];
     layer2_out[7730] <= layer1_out[7845];
     layer2_out[7731] <= ~(layer1_out[11569] ^ layer1_out[11570]);
     layer2_out[7732] <= layer1_out[161];
     layer2_out[7733] <= layer1_out[7524];
     layer2_out[7734] <= layer1_out[2415];
     layer2_out[7735] <= layer1_out[152];
     layer2_out[7736] <= layer1_out[3745] & ~layer1_out[3746];
     layer2_out[7737] <= ~layer1_out[6481];
     layer2_out[7738] <= ~layer1_out[10081] | layer1_out[10080];
     layer2_out[7739] <= ~(layer1_out[5121] & layer1_out[5122]);
     layer2_out[7740] <= layer1_out[4960];
     layer2_out[7741] <= ~(layer1_out[5434] | layer1_out[5435]);
     layer2_out[7742] <= ~layer1_out[4865];
     layer2_out[7743] <= ~layer1_out[7645];
     layer2_out[7744] <= layer1_out[8581];
     layer2_out[7745] <= ~layer1_out[7156] | layer1_out[7157];
     layer2_out[7746] <= layer1_out[2889] & layer1_out[2890];
     layer2_out[7747] <= ~layer1_out[5225];
     layer2_out[7748] <= layer1_out[522];
     layer2_out[7749] <= ~layer1_out[1189];
     layer2_out[7750] <= layer1_out[5202] & ~layer1_out[5201];
     layer2_out[7751] <= layer1_out[10506];
     layer2_out[7752] <= layer1_out[9063];
     layer2_out[7753] <= ~(layer1_out[3267] ^ layer1_out[3268]);
     layer2_out[7754] <= layer1_out[11591];
     layer2_out[7755] <= ~layer1_out[2466];
     layer2_out[7756] <= layer1_out[3059];
     layer2_out[7757] <= ~layer1_out[11661];
     layer2_out[7758] <= ~layer1_out[589];
     layer2_out[7759] <= ~layer1_out[10771];
     layer2_out[7760] <= layer1_out[5464] & ~layer1_out[5465];
     layer2_out[7761] <= ~layer1_out[385] | layer1_out[386];
     layer2_out[7762] <= layer1_out[1822] ^ layer1_out[1823];
     layer2_out[7763] <= ~(layer1_out[493] & layer1_out[494]);
     layer2_out[7764] <= ~layer1_out[9694] | layer1_out[9695];
     layer2_out[7765] <= ~layer1_out[1336];
     layer2_out[7766] <= 1'b0;
     layer2_out[7767] <= ~layer1_out[8831] | layer1_out[8830];
     layer2_out[7768] <= ~layer1_out[2249];
     layer2_out[7769] <= layer1_out[3198] & ~layer1_out[3199];
     layer2_out[7770] <= 1'b1;
     layer2_out[7771] <= layer1_out[11805];
     layer2_out[7772] <= ~layer1_out[9767];
     layer2_out[7773] <= layer1_out[2871] & layer1_out[2872];
     layer2_out[7774] <= layer1_out[7367];
     layer2_out[7775] <= ~layer1_out[6567];
     layer2_out[7776] <= layer1_out[2865] & ~layer1_out[2864];
     layer2_out[7777] <= ~(layer1_out[10771] | layer1_out[10772]);
     layer2_out[7778] <= ~(layer1_out[10332] & layer1_out[10333]);
     layer2_out[7779] <= layer1_out[6522] & layer1_out[6523];
     layer2_out[7780] <= ~layer1_out[11589];
     layer2_out[7781] <= ~(layer1_out[1685] ^ layer1_out[1686]);
     layer2_out[7782] <= ~layer1_out[4490] | layer1_out[4491];
     layer2_out[7783] <= ~layer1_out[1015];
     layer2_out[7784] <= ~layer1_out[3354] | layer1_out[3355];
     layer2_out[7785] <= ~layer1_out[6152];
     layer2_out[7786] <= ~layer1_out[469];
     layer2_out[7787] <= ~(layer1_out[5340] ^ layer1_out[5341]);
     layer2_out[7788] <= ~layer1_out[6319] | layer1_out[6320];
     layer2_out[7789] <= ~layer1_out[10825] | layer1_out[10824];
     layer2_out[7790] <= layer1_out[8857] & ~layer1_out[8856];
     layer2_out[7791] <= layer1_out[11037];
     layer2_out[7792] <= layer1_out[10925] & layer1_out[10926];
     layer2_out[7793] <= layer1_out[3980] | layer1_out[3981];
     layer2_out[7794] <= layer1_out[3610] | layer1_out[3611];
     layer2_out[7795] <= ~layer1_out[9489];
     layer2_out[7796] <= layer1_out[6553] & ~layer1_out[6554];
     layer2_out[7797] <= ~(layer1_out[6621] ^ layer1_out[6622]);
     layer2_out[7798] <= layer1_out[7447] & ~layer1_out[7448];
     layer2_out[7799] <= layer1_out[5271] & ~layer1_out[5270];
     layer2_out[7800] <= ~layer1_out[5149] | layer1_out[5148];
     layer2_out[7801] <= layer1_out[943];
     layer2_out[7802] <= ~(layer1_out[2157] & layer1_out[2158]);
     layer2_out[7803] <= layer1_out[10142] & ~layer1_out[10143];
     layer2_out[7804] <= 1'b0;
     layer2_out[7805] <= layer1_out[6498];
     layer2_out[7806] <= ~layer1_out[6172];
     layer2_out[7807] <= layer1_out[10864];
     layer2_out[7808] <= ~layer1_out[1120] | layer1_out[1119];
     layer2_out[7809] <= ~layer1_out[1836];
     layer2_out[7810] <= ~layer1_out[7264];
     layer2_out[7811] <= 1'b0;
     layer2_out[7812] <= layer1_out[10018] & ~layer1_out[10019];
     layer2_out[7813] <= ~layer1_out[7945];
     layer2_out[7814] <= layer1_out[2558] & layer1_out[2559];
     layer2_out[7815] <= layer1_out[6091];
     layer2_out[7816] <= layer1_out[957] & layer1_out[958];
     layer2_out[7817] <= layer1_out[7376] & layer1_out[7377];
     layer2_out[7818] <= layer1_out[168] & layer1_out[169];
     layer2_out[7819] <= ~(layer1_out[9385] & layer1_out[9386]);
     layer2_out[7820] <= layer1_out[8571] | layer1_out[8572];
     layer2_out[7821] <= ~layer1_out[1620];
     layer2_out[7822] <= layer1_out[6243];
     layer2_out[7823] <= ~layer1_out[11911];
     layer2_out[7824] <= layer1_out[1155];
     layer2_out[7825] <= layer1_out[10482] | layer1_out[10483];
     layer2_out[7826] <= layer1_out[1540] ^ layer1_out[1541];
     layer2_out[7827] <= layer1_out[219];
     layer2_out[7828] <= ~(layer1_out[11351] ^ layer1_out[11352]);
     layer2_out[7829] <= layer1_out[10296];
     layer2_out[7830] <= ~layer1_out[159] | layer1_out[160];
     layer2_out[7831] <= layer1_out[1678] & ~layer1_out[1677];
     layer2_out[7832] <= ~(layer1_out[9428] ^ layer1_out[9429]);
     layer2_out[7833] <= ~layer1_out[2311];
     layer2_out[7834] <= ~(layer1_out[9215] | layer1_out[9216]);
     layer2_out[7835] <= layer1_out[7722];
     layer2_out[7836] <= ~layer1_out[11769];
     layer2_out[7837] <= layer1_out[4184] & ~layer1_out[4185];
     layer2_out[7838] <= ~layer1_out[2039];
     layer2_out[7839] <= ~layer1_out[6131] | layer1_out[6132];
     layer2_out[7840] <= layer1_out[171] & ~layer1_out[172];
     layer2_out[7841] <= ~(layer1_out[8428] ^ layer1_out[8429]);
     layer2_out[7842] <= ~layer1_out[10110] | layer1_out[10109];
     layer2_out[7843] <= layer1_out[1636] & ~layer1_out[1635];
     layer2_out[7844] <= layer1_out[11232];
     layer2_out[7845] <= layer1_out[719];
     layer2_out[7846] <= ~layer1_out[11747];
     layer2_out[7847] <= layer1_out[2138];
     layer2_out[7848] <= ~layer1_out[894] | layer1_out[893];
     layer2_out[7849] <= ~layer1_out[9598];
     layer2_out[7850] <= ~layer1_out[3292];
     layer2_out[7851] <= ~(layer1_out[1930] | layer1_out[1931]);
     layer2_out[7852] <= ~layer1_out[9576];
     layer2_out[7853] <= ~(layer1_out[10212] ^ layer1_out[10213]);
     layer2_out[7854] <= layer1_out[9999] & ~layer1_out[10000];
     layer2_out[7855] <= layer1_out[4614];
     layer2_out[7856] <= layer1_out[3816];
     layer2_out[7857] <= layer1_out[1395];
     layer2_out[7858] <= ~(layer1_out[4705] | layer1_out[4706]);
     layer2_out[7859] <= layer1_out[361];
     layer2_out[7860] <= ~layer1_out[8837];
     layer2_out[7861] <= layer1_out[2769];
     layer2_out[7862] <= ~(layer1_out[9248] | layer1_out[9249]);
     layer2_out[7863] <= layer1_out[1388];
     layer2_out[7864] <= layer1_out[7912];
     layer2_out[7865] <= layer1_out[1890];
     layer2_out[7866] <= layer1_out[2584] & layer1_out[2585];
     layer2_out[7867] <= layer1_out[5755] & ~layer1_out[5756];
     layer2_out[7868] <= ~layer1_out[2951];
     layer2_out[7869] <= ~(layer1_out[5279] & layer1_out[5280]);
     layer2_out[7870] <= layer1_out[5684] & layer1_out[5685];
     layer2_out[7871] <= layer1_out[1292] & layer1_out[1293];
     layer2_out[7872] <= layer1_out[6828];
     layer2_out[7873] <= layer1_out[1413] & ~layer1_out[1414];
     layer2_out[7874] <= layer1_out[3282] | layer1_out[3283];
     layer2_out[7875] <= ~layer1_out[2466];
     layer2_out[7876] <= layer1_out[2966];
     layer2_out[7877] <= layer1_out[1795];
     layer2_out[7878] <= layer1_out[1339] & layer1_out[1340];
     layer2_out[7879] <= ~(layer1_out[1638] ^ layer1_out[1639]);
     layer2_out[7880] <= layer1_out[7522] & ~layer1_out[7521];
     layer2_out[7881] <= ~layer1_out[8997];
     layer2_out[7882] <= ~layer1_out[2657] | layer1_out[2658];
     layer2_out[7883] <= ~layer1_out[6469];
     layer2_out[7884] <= 1'b1;
     layer2_out[7885] <= ~layer1_out[8961];
     layer2_out[7886] <= ~layer1_out[11920];
     layer2_out[7887] <= layer1_out[7500];
     layer2_out[7888] <= layer1_out[5708] ^ layer1_out[5709];
     layer2_out[7889] <= layer1_out[8530] & ~layer1_out[8531];
     layer2_out[7890] <= layer1_out[2257];
     layer2_out[7891] <= ~layer1_out[5455] | layer1_out[5456];
     layer2_out[7892] <= layer1_out[2070] & ~layer1_out[2069];
     layer2_out[7893] <= ~layer1_out[11785] | layer1_out[11786];
     layer2_out[7894] <= 1'b0;
     layer2_out[7895] <= ~layer1_out[9546];
     layer2_out[7896] <= ~layer1_out[2718];
     layer2_out[7897] <= ~(layer1_out[263] ^ layer1_out[264]);
     layer2_out[7898] <= ~(layer1_out[3013] | layer1_out[3014]);
     layer2_out[7899] <= layer1_out[3886];
     layer2_out[7900] <= layer1_out[6609] | layer1_out[6610];
     layer2_out[7901] <= ~(layer1_out[2351] ^ layer1_out[2352]);
     layer2_out[7902] <= ~layer1_out[8339];
     layer2_out[7903] <= ~layer1_out[10242];
     layer2_out[7904] <= ~(layer1_out[3276] & layer1_out[3277]);
     layer2_out[7905] <= ~(layer1_out[1959] | layer1_out[1960]);
     layer2_out[7906] <= layer1_out[1320] & ~layer1_out[1319];
     layer2_out[7907] <= ~layer1_out[4688];
     layer2_out[7908] <= layer1_out[7330] & layer1_out[7331];
     layer2_out[7909] <= ~(layer1_out[5266] & layer1_out[5267]);
     layer2_out[7910] <= ~(layer1_out[10744] ^ layer1_out[10745]);
     layer2_out[7911] <= layer1_out[4565] ^ layer1_out[4566];
     layer2_out[7912] <= layer1_out[9274] & layer1_out[9275];
     layer2_out[7913] <= layer1_out[3029] & layer1_out[3030];
     layer2_out[7914] <= ~layer1_out[7271] | layer1_out[7270];
     layer2_out[7915] <= ~layer1_out[6480];
     layer2_out[7916] <= ~layer1_out[8095] | layer1_out[8096];
     layer2_out[7917] <= layer1_out[6883];
     layer2_out[7918] <= ~layer1_out[234];
     layer2_out[7919] <= layer1_out[1782];
     layer2_out[7920] <= layer1_out[501];
     layer2_out[7921] <= layer1_out[11272] | layer1_out[11273];
     layer2_out[7922] <= layer1_out[6531] & ~layer1_out[6532];
     layer2_out[7923] <= layer1_out[11418] ^ layer1_out[11419];
     layer2_out[7924] <= ~(layer1_out[697] & layer1_out[698]);
     layer2_out[7925] <= layer1_out[9859] ^ layer1_out[9860];
     layer2_out[7926] <= layer1_out[10115];
     layer2_out[7927] <= ~layer1_out[11960];
     layer2_out[7928] <= ~layer1_out[8239];
     layer2_out[7929] <= ~layer1_out[5207] | layer1_out[5206];
     layer2_out[7930] <= layer1_out[2261];
     layer2_out[7931] <= ~(layer1_out[4212] | layer1_out[4213]);
     layer2_out[7932] <= layer1_out[830] | layer1_out[831];
     layer2_out[7933] <= layer1_out[3665];
     layer2_out[7934] <= layer1_out[9030] ^ layer1_out[9031];
     layer2_out[7935] <= ~(layer1_out[8267] & layer1_out[8268]);
     layer2_out[7936] <= ~layer1_out[7095];
     layer2_out[7937] <= layer1_out[3261];
     layer2_out[7938] <= ~(layer1_out[8854] ^ layer1_out[8855]);
     layer2_out[7939] <= layer1_out[9846] ^ layer1_out[9847];
     layer2_out[7940] <= layer1_out[11050] & ~layer1_out[11049];
     layer2_out[7941] <= layer1_out[5236];
     layer2_out[7942] <= ~layer1_out[3715];
     layer2_out[7943] <= layer1_out[10416] & ~layer1_out[10417];
     layer2_out[7944] <= ~(layer1_out[2816] | layer1_out[2817]);
     layer2_out[7945] <= ~layer1_out[393];
     layer2_out[7946] <= layer1_out[10395];
     layer2_out[7947] <= layer1_out[6493];
     layer2_out[7948] <= layer1_out[4510] & ~layer1_out[4509];
     layer2_out[7949] <= layer1_out[8978] ^ layer1_out[8979];
     layer2_out[7950] <= ~layer1_out[4522];
     layer2_out[7951] <= ~layer1_out[9405];
     layer2_out[7952] <= layer1_out[9100];
     layer2_out[7953] <= layer1_out[8185] & layer1_out[8186];
     layer2_out[7954] <= ~layer1_out[3510];
     layer2_out[7955] <= ~layer1_out[2837] | layer1_out[2838];
     layer2_out[7956] <= ~layer1_out[2159];
     layer2_out[7957] <= ~layer1_out[4479] | layer1_out[4478];
     layer2_out[7958] <= layer1_out[3332];
     layer2_out[7959] <= layer1_out[9278];
     layer2_out[7960] <= ~layer1_out[9356] | layer1_out[9357];
     layer2_out[7961] <= ~layer1_out[7345] | layer1_out[7344];
     layer2_out[7962] <= ~layer1_out[10020];
     layer2_out[7963] <= layer1_out[10104];
     layer2_out[7964] <= layer1_out[5820];
     layer2_out[7965] <= ~layer1_out[8797];
     layer2_out[7966] <= layer1_out[4352] | layer1_out[4353];
     layer2_out[7967] <= ~(layer1_out[10527] | layer1_out[10528]);
     layer2_out[7968] <= ~layer1_out[10987];
     layer2_out[7969] <= ~layer1_out[8006];
     layer2_out[7970] <= layer1_out[9595];
     layer2_out[7971] <= layer1_out[4062] & ~layer1_out[4063];
     layer2_out[7972] <= layer1_out[8167] & ~layer1_out[8168];
     layer2_out[7973] <= ~layer1_out[691];
     layer2_out[7974] <= ~layer1_out[2960] | layer1_out[2961];
     layer2_out[7975] <= ~layer1_out[1304];
     layer2_out[7976] <= layer1_out[6270] | layer1_out[6271];
     layer2_out[7977] <= layer1_out[3282];
     layer2_out[7978] <= layer1_out[2562];
     layer2_out[7979] <= ~layer1_out[10153] | layer1_out[10154];
     layer2_out[7980] <= layer1_out[6728];
     layer2_out[7981] <= layer1_out[7536] & layer1_out[7537];
     layer2_out[7982] <= ~(layer1_out[9366] & layer1_out[9367]);
     layer2_out[7983] <= ~(layer1_out[7055] ^ layer1_out[7056]);
     layer2_out[7984] <= ~layer1_out[7808];
     layer2_out[7985] <= ~(layer1_out[9569] | layer1_out[9570]);
     layer2_out[7986] <= ~layer1_out[2189];
     layer2_out[7987] <= ~layer1_out[10793];
     layer2_out[7988] <= layer1_out[5173];
     layer2_out[7989] <= ~layer1_out[2797] | layer1_out[2796];
     layer2_out[7990] <= ~(layer1_out[901] ^ layer1_out[902]);
     layer2_out[7991] <= ~layer1_out[4665];
     layer2_out[7992] <= ~(layer1_out[8252] | layer1_out[8253]);
     layer2_out[7993] <= ~(layer1_out[7841] ^ layer1_out[7842]);
     layer2_out[7994] <= layer1_out[11505] | layer1_out[11506];
     layer2_out[7995] <= ~layer1_out[1418];
     layer2_out[7996] <= layer1_out[10041] ^ layer1_out[10042];
     layer2_out[7997] <= ~layer1_out[10167];
     layer2_out[7998] <= layer1_out[1658];
     layer2_out[7999] <= layer1_out[5666] | layer1_out[5667];
     layer2_out[8000] <= layer1_out[1673];
     layer2_out[8001] <= layer1_out[1049];
     layer2_out[8002] <= ~(layer1_out[4127] & layer1_out[4128]);
     layer2_out[8003] <= ~(layer1_out[5789] ^ layer1_out[5790]);
     layer2_out[8004] <= ~layer1_out[9187];
     layer2_out[8005] <= ~layer1_out[6014] | layer1_out[6013];
     layer2_out[8006] <= layer1_out[3344] & ~layer1_out[3345];
     layer2_out[8007] <= ~(layer1_out[7566] | layer1_out[7567]);
     layer2_out[8008] <= ~layer1_out[6284];
     layer2_out[8009] <= ~(layer1_out[2704] ^ layer1_out[2705]);
     layer2_out[8010] <= ~(layer1_out[11711] | layer1_out[11712]);
     layer2_out[8011] <= ~layer1_out[4902] | layer1_out[4903];
     layer2_out[8012] <= ~layer1_out[11738];
     layer2_out[8013] <= ~(layer1_out[7778] ^ layer1_out[7779]);
     layer2_out[8014] <= layer1_out[6697] & layer1_out[6698];
     layer2_out[8015] <= layer1_out[1073] & ~layer1_out[1072];
     layer2_out[8016] <= layer1_out[10903];
     layer2_out[8017] <= layer1_out[8640] | layer1_out[8641];
     layer2_out[8018] <= ~layer1_out[2107];
     layer2_out[8019] <= ~layer1_out[4801];
     layer2_out[8020] <= layer1_out[5594] ^ layer1_out[5595];
     layer2_out[8021] <= ~layer1_out[11584];
     layer2_out[8022] <= layer1_out[5336] | layer1_out[5337];
     layer2_out[8023] <= ~(layer1_out[9242] ^ layer1_out[9243]);
     layer2_out[8024] <= layer1_out[8605];
     layer2_out[8025] <= 1'b1;
     layer2_out[8026] <= layer1_out[4554] ^ layer1_out[4555];
     layer2_out[8027] <= layer1_out[10547] | layer1_out[10548];
     layer2_out[8028] <= ~(layer1_out[8351] | layer1_out[8352]);
     layer2_out[8029] <= ~layer1_out[9527];
     layer2_out[8030] <= ~layer1_out[6859];
     layer2_out[8031] <= layer1_out[9443];
     layer2_out[8032] <= ~(layer1_out[9761] | layer1_out[9762]);
     layer2_out[8033] <= layer1_out[3386];
     layer2_out[8034] <= ~(layer1_out[8464] | layer1_out[8465]);
     layer2_out[8035] <= layer1_out[8268];
     layer2_out[8036] <= layer1_out[5309] & ~layer1_out[5310];
     layer2_out[8037] <= layer1_out[7476] & ~layer1_out[7477];
     layer2_out[8038] <= layer1_out[2950];
     layer2_out[8039] <= ~(layer1_out[10949] & layer1_out[10950]);
     layer2_out[8040] <= layer1_out[7196] | layer1_out[7197];
     layer2_out[8041] <= ~(layer1_out[8632] ^ layer1_out[8633]);
     layer2_out[8042] <= layer1_out[2539];
     layer2_out[8043] <= ~layer1_out[8324] | layer1_out[8323];
     layer2_out[8044] <= ~layer1_out[7911];
     layer2_out[8045] <= layer1_out[4343] & ~layer1_out[4344];
     layer2_out[8046] <= layer1_out[3995];
     layer2_out[8047] <= layer1_out[2982] & ~layer1_out[2983];
     layer2_out[8048] <= ~(layer1_out[9906] & layer1_out[9907]);
     layer2_out[8049] <= ~layer1_out[5027] | layer1_out[5028];
     layer2_out[8050] <= layer1_out[202];
     layer2_out[8051] <= ~(layer1_out[7881] ^ layer1_out[7882]);
     layer2_out[8052] <= ~layer1_out[5256];
     layer2_out[8053] <= layer1_out[10951];
     layer2_out[8054] <= layer1_out[3447] & layer1_out[3448];
     layer2_out[8055] <= ~(layer1_out[5334] & layer1_out[5335]);
     layer2_out[8056] <= ~layer1_out[436];
     layer2_out[8057] <= 1'b0;
     layer2_out[8058] <= layer1_out[3774] ^ layer1_out[3775];
     layer2_out[8059] <= ~(layer1_out[1347] | layer1_out[1348]);
     layer2_out[8060] <= layer1_out[11822] ^ layer1_out[11823];
     layer2_out[8061] <= layer1_out[7293] | layer1_out[7294];
     layer2_out[8062] <= ~layer1_out[4504] | layer1_out[4503];
     layer2_out[8063] <= ~layer1_out[5452];
     layer2_out[8064] <= ~layer1_out[9518] | layer1_out[9519];
     layer2_out[8065] <= layer1_out[3042] & ~layer1_out[3041];
     layer2_out[8066] <= ~(layer1_out[2168] ^ layer1_out[2169]);
     layer2_out[8067] <= ~layer1_out[1786] | layer1_out[1785];
     layer2_out[8068] <= layer1_out[3596] | layer1_out[3597];
     layer2_out[8069] <= ~layer1_out[7339];
     layer2_out[8070] <= layer1_out[2820];
     layer2_out[8071] <= layer1_out[340];
     layer2_out[8072] <= layer1_out[9778] | layer1_out[9779];
     layer2_out[8073] <= ~(layer1_out[3553] | layer1_out[3554]);
     layer2_out[8074] <= layer1_out[5891];
     layer2_out[8075] <= ~layer1_out[5063];
     layer2_out[8076] <= ~layer1_out[11173];
     layer2_out[8077] <= ~layer1_out[6272] | layer1_out[6271];
     layer2_out[8078] <= layer1_out[5036];
     layer2_out[8079] <= layer1_out[5195] ^ layer1_out[5196];
     layer2_out[8080] <= ~(layer1_out[8867] & layer1_out[8868]);
     layer2_out[8081] <= ~layer1_out[8858] | layer1_out[8859];
     layer2_out[8082] <= layer1_out[8668];
     layer2_out[8083] <= ~(layer1_out[8460] | layer1_out[8461]);
     layer2_out[8084] <= layer1_out[11087] & ~layer1_out[11086];
     layer2_out[8085] <= layer1_out[9305];
     layer2_out[8086] <= ~layer1_out[3137];
     layer2_out[8087] <= ~(layer1_out[6113] & layer1_out[6114]);
     layer2_out[8088] <= ~layer1_out[4322];
     layer2_out[8089] <= ~layer1_out[9091];
     layer2_out[8090] <= layer1_out[5480] | layer1_out[5481];
     layer2_out[8091] <= ~layer1_out[5514];
     layer2_out[8092] <= layer1_out[6292] & ~layer1_out[6293];
     layer2_out[8093] <= ~layer1_out[3481] | layer1_out[3482];
     layer2_out[8094] <= layer1_out[5964] & layer1_out[5965];
     layer2_out[8095] <= ~(layer1_out[1786] ^ layer1_out[1787]);
     layer2_out[8096] <= layer1_out[3200];
     layer2_out[8097] <= layer1_out[1183] ^ layer1_out[1184];
     layer2_out[8098] <= layer1_out[6830];
     layer2_out[8099] <= layer1_out[648] & layer1_out[649];
     layer2_out[8100] <= ~layer1_out[2398];
     layer2_out[8101] <= ~(layer1_out[48] ^ layer1_out[49]);
     layer2_out[8102] <= ~layer1_out[11912];
     layer2_out[8103] <= ~layer1_out[9216];
     layer2_out[8104] <= layer1_out[7667] & ~layer1_out[7666];
     layer2_out[8105] <= ~(layer1_out[7709] | layer1_out[7710]);
     layer2_out[8106] <= layer1_out[1764];
     layer2_out[8107] <= 1'b0;
     layer2_out[8108] <= ~layer1_out[4327];
     layer2_out[8109] <= ~(layer1_out[5527] & layer1_out[5528]);
     layer2_out[8110] <= layer1_out[6179] | layer1_out[6180];
     layer2_out[8111] <= 1'b0;
     layer2_out[8112] <= layer1_out[6999] ^ layer1_out[7000];
     layer2_out[8113] <= ~layer1_out[8859];
     layer2_out[8114] <= ~(layer1_out[9082] & layer1_out[9083]);
     layer2_out[8115] <= layer1_out[691] & layer1_out[692];
     layer2_out[8116] <= ~layer1_out[10625] | layer1_out[10626];
     layer2_out[8117] <= layer1_out[3665];
     layer2_out[8118] <= ~layer1_out[9314];
     layer2_out[8119] <= ~layer1_out[4886];
     layer2_out[8120] <= layer1_out[2494] ^ layer1_out[2495];
     layer2_out[8121] <= ~layer1_out[6798];
     layer2_out[8122] <= ~layer1_out[11349];
     layer2_out[8123] <= ~layer1_out[2185];
     layer2_out[8124] <= layer1_out[1569];
     layer2_out[8125] <= ~layer1_out[7697];
     layer2_out[8126] <= layer1_out[4000];
     layer2_out[8127] <= ~layer1_out[1702] | layer1_out[1701];
     layer2_out[8128] <= ~layer1_out[11851] | layer1_out[11852];
     layer2_out[8129] <= layer1_out[2649] & ~layer1_out[2648];
     layer2_out[8130] <= ~(layer1_out[10098] ^ layer1_out[10099]);
     layer2_out[8131] <= ~layer1_out[5869] | layer1_out[5870];
     layer2_out[8132] <= layer1_out[1038] | layer1_out[1039];
     layer2_out[8133] <= 1'b1;
     layer2_out[8134] <= ~(layer1_out[2580] ^ layer1_out[2581]);
     layer2_out[8135] <= ~(layer1_out[4989] | layer1_out[4990]);
     layer2_out[8136] <= ~layer1_out[6460];
     layer2_out[8137] <= layer1_out[6020] & ~layer1_out[6021];
     layer2_out[8138] <= ~layer1_out[278];
     layer2_out[8139] <= ~layer1_out[8000] | layer1_out[7999];
     layer2_out[8140] <= layer1_out[4693];
     layer2_out[8141] <= ~layer1_out[2165];
     layer2_out[8142] <= layer1_out[5436] & ~layer1_out[5435];
     layer2_out[8143] <= layer1_out[4911] & layer1_out[4912];
     layer2_out[8144] <= ~layer1_out[8615] | layer1_out[8616];
     layer2_out[8145] <= layer1_out[2745] & layer1_out[2746];
     layer2_out[8146] <= layer1_out[7917] & layer1_out[7918];
     layer2_out[8147] <= ~layer1_out[4468];
     layer2_out[8148] <= ~(layer1_out[3436] | layer1_out[3437]);
     layer2_out[8149] <= ~(layer1_out[2766] ^ layer1_out[2767]);
     layer2_out[8150] <= layer1_out[4054] & ~layer1_out[4055];
     layer2_out[8151] <= layer1_out[11456];
     layer2_out[8152] <= layer1_out[3816] & ~layer1_out[3817];
     layer2_out[8153] <= layer1_out[7163];
     layer2_out[8154] <= layer1_out[10900] ^ layer1_out[10901];
     layer2_out[8155] <= layer1_out[9333];
     layer2_out[8156] <= ~(layer1_out[11138] & layer1_out[11139]);
     layer2_out[8157] <= ~layer1_out[8591] | layer1_out[8590];
     layer2_out[8158] <= layer1_out[3953] & ~layer1_out[3952];
     layer2_out[8159] <= ~(layer1_out[2592] | layer1_out[2593]);
     layer2_out[8160] <= layer1_out[10751] & ~layer1_out[10752];
     layer2_out[8161] <= layer1_out[4193];
     layer2_out[8162] <= ~(layer1_out[8068] ^ layer1_out[8069]);
     layer2_out[8163] <= layer1_out[793];
     layer2_out[8164] <= ~(layer1_out[4961] ^ layer1_out[4962]);
     layer2_out[8165] <= layer1_out[3234];
     layer2_out[8166] <= layer1_out[4747];
     layer2_out[8167] <= layer1_out[10505] | layer1_out[10506];
     layer2_out[8168] <= ~layer1_out[4348];
     layer2_out[8169] <= ~layer1_out[5410] | layer1_out[5411];
     layer2_out[8170] <= ~layer1_out[11075];
     layer2_out[8171] <= ~layer1_out[1461];
     layer2_out[8172] <= ~(layer1_out[10075] & layer1_out[10076]);
     layer2_out[8173] <= ~layer1_out[2018];
     layer2_out[8174] <= layer1_out[9372] & ~layer1_out[9373];
     layer2_out[8175] <= layer1_out[6591];
     layer2_out[8176] <= ~(layer1_out[11416] ^ layer1_out[11417]);
     layer2_out[8177] <= ~layer1_out[9836] | layer1_out[9835];
     layer2_out[8178] <= ~layer1_out[5380] | layer1_out[5381];
     layer2_out[8179] <= layer1_out[5157] | layer1_out[5158];
     layer2_out[8180] <= layer1_out[5101] & ~layer1_out[5100];
     layer2_out[8181] <= layer1_out[8740];
     layer2_out[8182] <= ~layer1_out[1073] | layer1_out[1074];
     layer2_out[8183] <= ~layer1_out[3031];
     layer2_out[8184] <= layer1_out[5785];
     layer2_out[8185] <= ~(layer1_out[3390] | layer1_out[3391]);
     layer2_out[8186] <= ~(layer1_out[630] ^ layer1_out[631]);
     layer2_out[8187] <= layer1_out[1126];
     layer2_out[8188] <= layer1_out[2950] | layer1_out[2951];
     layer2_out[8189] <= ~layer1_out[9891] | layer1_out[9892];
     layer2_out[8190] <= layer1_out[1804] & ~layer1_out[1803];
     layer2_out[8191] <= layer1_out[4465] ^ layer1_out[4466];
     layer2_out[8192] <= layer1_out[700] ^ layer1_out[701];
     layer2_out[8193] <= ~layer1_out[4489];
     layer2_out[8194] <= ~(layer1_out[8101] & layer1_out[8102]);
     layer2_out[8195] <= ~layer1_out[10331] | layer1_out[10330];
     layer2_out[8196] <= layer1_out[6500] & ~layer1_out[6501];
     layer2_out[8197] <= ~layer1_out[7017];
     layer2_out[8198] <= layer1_out[142] & ~layer1_out[141];
     layer2_out[8199] <= ~layer1_out[4985];
     layer2_out[8200] <= layer1_out[4068] & layer1_out[4069];
     layer2_out[8201] <= ~layer1_out[4891];
     layer2_out[8202] <= layer1_out[11025] & layer1_out[11026];
     layer2_out[8203] <= ~layer1_out[4930] | layer1_out[4929];
     layer2_out[8204] <= layer1_out[9520];
     layer2_out[8205] <= ~layer1_out[11293];
     layer2_out[8206] <= ~(layer1_out[8385] | layer1_out[8386]);
     layer2_out[8207] <= ~layer1_out[2624];
     layer2_out[8208] <= ~(layer1_out[10325] | layer1_out[10326]);
     layer2_out[8209] <= layer1_out[11512] ^ layer1_out[11513];
     layer2_out[8210] <= layer1_out[7982] & ~layer1_out[7983];
     layer2_out[8211] <= ~layer1_out[5095] | layer1_out[5094];
     layer2_out[8212] <= ~layer1_out[10720] | layer1_out[10719];
     layer2_out[8213] <= layer1_out[7103];
     layer2_out[8214] <= ~(layer1_out[2782] & layer1_out[2783]);
     layer2_out[8215] <= layer1_out[3157] ^ layer1_out[3158];
     layer2_out[8216] <= ~(layer1_out[3899] ^ layer1_out[3900]);
     layer2_out[8217] <= layer1_out[5081];
     layer2_out[8218] <= layer1_out[2837];
     layer2_out[8219] <= layer1_out[3146];
     layer2_out[8220] <= ~(layer1_out[10736] & layer1_out[10737]);
     layer2_out[8221] <= layer1_out[8083] | layer1_out[8084];
     layer2_out[8222] <= ~layer1_out[8567] | layer1_out[8568];
     layer2_out[8223] <= ~(layer1_out[2493] & layer1_out[2494]);
     layer2_out[8224] <= ~(layer1_out[2940] & layer1_out[2941]);
     layer2_out[8225] <= layer1_out[8440];
     layer2_out[8226] <= ~layer1_out[9819] | layer1_out[9820];
     layer2_out[8227] <= layer1_out[6182];
     layer2_out[8228] <= ~layer1_out[3270];
     layer2_out[8229] <= ~layer1_out[4027];
     layer2_out[8230] <= layer1_out[8116];
     layer2_out[8231] <= 1'b1;
     layer2_out[8232] <= ~layer1_out[1362];
     layer2_out[8233] <= ~layer1_out[9895];
     layer2_out[8234] <= ~layer1_out[2611];
     layer2_out[8235] <= layer1_out[9802];
     layer2_out[8236] <= ~layer1_out[7052];
     layer2_out[8237] <= ~layer1_out[5555];
     layer2_out[8238] <= layer1_out[11461];
     layer2_out[8239] <= ~layer1_out[420] | layer1_out[421];
     layer2_out[8240] <= ~layer1_out[7119];
     layer2_out[8241] <= layer1_out[9723];
     layer2_out[8242] <= layer1_out[5691];
     layer2_out[8243] <= ~layer1_out[7412];
     layer2_out[8244] <= layer1_out[8087];
     layer2_out[8245] <= 1'b1;
     layer2_out[8246] <= layer1_out[1200] & ~layer1_out[1199];
     layer2_out[8247] <= layer1_out[10261] & layer1_out[10262];
     layer2_out[8248] <= layer1_out[9226] & ~layer1_out[9227];
     layer2_out[8249] <= ~layer1_out[4806];
     layer2_out[8250] <= ~layer1_out[7648] | layer1_out[7647];
     layer2_out[8251] <= layer1_out[1039] | layer1_out[1040];
     layer2_out[8252] <= ~(layer1_out[5988] & layer1_out[5989]);
     layer2_out[8253] <= layer1_out[1803] & ~layer1_out[1802];
     layer2_out[8254] <= layer1_out[10197] & layer1_out[10198];
     layer2_out[8255] <= ~(layer1_out[10539] & layer1_out[10540]);
     layer2_out[8256] <= layer1_out[3992] | layer1_out[3993];
     layer2_out[8257] <= layer1_out[7786];
     layer2_out[8258] <= ~layer1_out[10735];
     layer2_out[8259] <= layer1_out[9230];
     layer2_out[8260] <= layer1_out[5078];
     layer2_out[8261] <= ~layer1_out[6358] | layer1_out[6357];
     layer2_out[8262] <= layer1_out[24];
     layer2_out[8263] <= ~layer1_out[1663] | layer1_out[1662];
     layer2_out[8264] <= layer1_out[10610] & layer1_out[10611];
     layer2_out[8265] <= layer1_out[11277];
     layer2_out[8266] <= layer1_out[6265] ^ layer1_out[6266];
     layer2_out[8267] <= layer1_out[576];
     layer2_out[8268] <= ~layer1_out[10573] | layer1_out[10572];
     layer2_out[8269] <= ~layer1_out[6478] | layer1_out[6477];
     layer2_out[8270] <= layer1_out[7978] ^ layer1_out[7979];
     layer2_out[8271] <= layer1_out[10378];
     layer2_out[8272] <= layer1_out[7012];
     layer2_out[8273] <= ~layer1_out[3183];
     layer2_out[8274] <= layer1_out[4858] & ~layer1_out[4857];
     layer2_out[8275] <= ~layer1_out[11391] | layer1_out[11392];
     layer2_out[8276] <= ~layer1_out[7775];
     layer2_out[8277] <= ~layer1_out[7355];
     layer2_out[8278] <= ~layer1_out[4441];
     layer2_out[8279] <= layer1_out[3663] & ~layer1_out[3662];
     layer2_out[8280] <= ~(layer1_out[1440] & layer1_out[1441]);
     layer2_out[8281] <= layer1_out[1127] & ~layer1_out[1128];
     layer2_out[8282] <= ~layer1_out[11479] | layer1_out[11478];
     layer2_out[8283] <= layer1_out[2448];
     layer2_out[8284] <= layer1_out[9658];
     layer2_out[8285] <= ~layer1_out[1657];
     layer2_out[8286] <= ~layer1_out[10286];
     layer2_out[8287] <= ~layer1_out[11558];
     layer2_out[8288] <= ~(layer1_out[843] ^ layer1_out[844]);
     layer2_out[8289] <= ~layer1_out[2313];
     layer2_out[8290] <= layer1_out[10513] | layer1_out[10514];
     layer2_out[8291] <= ~layer1_out[11848] | layer1_out[11847];
     layer2_out[8292] <= ~layer1_out[2191] | layer1_out[2192];
     layer2_out[8293] <= layer1_out[8813] ^ layer1_out[8814];
     layer2_out[8294] <= ~layer1_out[1483] | layer1_out[1482];
     layer2_out[8295] <= layer1_out[1007];
     layer2_out[8296] <= ~layer1_out[6658];
     layer2_out[8297] <= layer1_out[8783];
     layer2_out[8298] <= ~layer1_out[5426] | layer1_out[5425];
     layer2_out[8299] <= layer1_out[7542];
     layer2_out[8300] <= ~layer1_out[3502];
     layer2_out[8301] <= ~(layer1_out[1910] & layer1_out[1911]);
     layer2_out[8302] <= layer1_out[11495] & ~layer1_out[11494];
     layer2_out[8303] <= layer1_out[11658] ^ layer1_out[11659];
     layer2_out[8304] <= ~(layer1_out[5255] | layer1_out[5256]);
     layer2_out[8305] <= layer1_out[845] & layer1_out[846];
     layer2_out[8306] <= ~(layer1_out[9961] & layer1_out[9962]);
     layer2_out[8307] <= layer1_out[7557] & ~layer1_out[7558];
     layer2_out[8308] <= ~layer1_out[11195];
     layer2_out[8309] <= ~layer1_out[1347];
     layer2_out[8310] <= ~(layer1_out[6705] | layer1_out[6706]);
     layer2_out[8311] <= layer1_out[2437];
     layer2_out[8312] <= ~layer1_out[11406];
     layer2_out[8313] <= layer1_out[6295];
     layer2_out[8314] <= ~(layer1_out[6257] & layer1_out[6258]);
     layer2_out[8315] <= ~(layer1_out[2189] | layer1_out[2190]);
     layer2_out[8316] <= layer1_out[11129] & layer1_out[11130];
     layer2_out[8317] <= ~(layer1_out[11679] | layer1_out[11680]);
     layer2_out[8318] <= ~(layer1_out[11215] ^ layer1_out[11216]);
     layer2_out[8319] <= ~(layer1_out[10497] ^ layer1_out[10498]);
     layer2_out[8320] <= ~layer1_out[6156];
     layer2_out[8321] <= ~layer1_out[1562];
     layer2_out[8322] <= layer1_out[797] | layer1_out[798];
     layer2_out[8323] <= layer1_out[4779] ^ layer1_out[4780];
     layer2_out[8324] <= ~(layer1_out[1598] & layer1_out[1599]);
     layer2_out[8325] <= ~layer1_out[896] | layer1_out[897];
     layer2_out[8326] <= ~(layer1_out[4760] ^ layer1_out[4761]);
     layer2_out[8327] <= layer1_out[10123];
     layer2_out[8328] <= layer1_out[9921];
     layer2_out[8329] <= ~layer1_out[7735] | layer1_out[7734];
     layer2_out[8330] <= ~layer1_out[7497] | layer1_out[7498];
     layer2_out[8331] <= layer1_out[1085] & ~layer1_out[1086];
     layer2_out[8332] <= layer1_out[127];
     layer2_out[8333] <= ~(layer1_out[2358] & layer1_out[2359]);
     layer2_out[8334] <= ~layer1_out[11603] | layer1_out[11604];
     layer2_out[8335] <= ~layer1_out[1537];
     layer2_out[8336] <= ~layer1_out[9256];
     layer2_out[8337] <= layer1_out[10220] | layer1_out[10221];
     layer2_out[8338] <= ~layer1_out[1450];
     layer2_out[8339] <= ~layer1_out[10805];
     layer2_out[8340] <= layer1_out[1253];
     layer2_out[8341] <= ~layer1_out[7872] | layer1_out[7873];
     layer2_out[8342] <= ~layer1_out[1468];
     layer2_out[8343] <= layer1_out[7952];
     layer2_out[8344] <= layer1_out[11859] ^ layer1_out[11860];
     layer2_out[8345] <= layer1_out[3843];
     layer2_out[8346] <= ~(layer1_out[7704] | layer1_out[7705]);
     layer2_out[8347] <= layer1_out[6634];
     layer2_out[8348] <= layer1_out[5104];
     layer2_out[8349] <= layer1_out[10858];
     layer2_out[8350] <= ~(layer1_out[7242] ^ layer1_out[7243]);
     layer2_out[8351] <= ~layer1_out[7468];
     layer2_out[8352] <= ~layer1_out[10287] | layer1_out[10288];
     layer2_out[8353] <= layer1_out[4183];
     layer2_out[8354] <= layer1_out[9049];
     layer2_out[8355] <= ~(layer1_out[10228] & layer1_out[10229]);
     layer2_out[8356] <= layer1_out[6261];
     layer2_out[8357] <= ~layer1_out[5179] | layer1_out[5180];
     layer2_out[8358] <= ~layer1_out[4548];
     layer2_out[8359] <= ~layer1_out[7521];
     layer2_out[8360] <= layer1_out[6552] & ~layer1_out[6553];
     layer2_out[8361] <= layer1_out[7084] ^ layer1_out[7085];
     layer2_out[8362] <= ~layer1_out[2103];
     layer2_out[8363] <= ~(layer1_out[5117] | layer1_out[5118]);
     layer2_out[8364] <= ~(layer1_out[7406] | layer1_out[7407]);
     layer2_out[8365] <= ~(layer1_out[7288] | layer1_out[7289]);
     layer2_out[8366] <= layer1_out[7135];
     layer2_out[8367] <= ~layer1_out[11669] | layer1_out[11670];
     layer2_out[8368] <= layer1_out[10447];
     layer2_out[8369] <= layer1_out[126] | layer1_out[127];
     layer2_out[8370] <= layer1_out[11486] | layer1_out[11487];
     layer2_out[8371] <= ~layer1_out[3250];
     layer2_out[8372] <= layer1_out[7559] | layer1_out[7560];
     layer2_out[8373] <= layer1_out[4350] | layer1_out[4351];
     layer2_out[8374] <= layer1_out[5316];
     layer2_out[8375] <= layer1_out[11419] & layer1_out[11420];
     layer2_out[8376] <= layer1_out[3733] & layer1_out[3734];
     layer2_out[8377] <= ~(layer1_out[11939] ^ layer1_out[11940]);
     layer2_out[8378] <= ~(layer1_out[6739] | layer1_out[6740]);
     layer2_out[8379] <= ~layer1_out[5857] | layer1_out[5858];
     layer2_out[8380] <= layer1_out[11504] & ~layer1_out[11505];
     layer2_out[8381] <= ~(layer1_out[8235] ^ layer1_out[8236]);
     layer2_out[8382] <= ~layer1_out[1596] | layer1_out[1597];
     layer2_out[8383] <= ~layer1_out[3346];
     layer2_out[8384] <= ~layer1_out[4642];
     layer2_out[8385] <= layer1_out[3052] | layer1_out[3053];
     layer2_out[8386] <= layer1_out[2410] | layer1_out[2411];
     layer2_out[8387] <= ~layer1_out[3027];
     layer2_out[8388] <= ~layer1_out[1778] | layer1_out[1779];
     layer2_out[8389] <= layer1_out[4921] & layer1_out[4922];
     layer2_out[8390] <= ~layer1_out[7195] | layer1_out[7196];
     layer2_out[8391] <= layer1_out[2225] | layer1_out[2226];
     layer2_out[8392] <= layer1_out[5922] | layer1_out[5923];
     layer2_out[8393] <= ~layer1_out[8356];
     layer2_out[8394] <= layer1_out[10404] & ~layer1_out[10403];
     layer2_out[8395] <= ~(layer1_out[2868] ^ layer1_out[2869]);
     layer2_out[8396] <= layer1_out[2633] & layer1_out[2634];
     layer2_out[8397] <= ~layer1_out[11672];
     layer2_out[8398] <= layer1_out[8002] | layer1_out[8003];
     layer2_out[8399] <= layer1_out[10621];
     layer2_out[8400] <= ~layer1_out[10182];
     layer2_out[8401] <= layer1_out[8343] ^ layer1_out[8344];
     layer2_out[8402] <= layer1_out[9950] & ~layer1_out[9951];
     layer2_out[8403] <= layer1_out[3179];
     layer2_out[8404] <= layer1_out[6412] & layer1_out[6413];
     layer2_out[8405] <= ~(layer1_out[9901] & layer1_out[9902]);
     layer2_out[8406] <= ~layer1_out[6954];
     layer2_out[8407] <= layer1_out[4245];
     layer2_out[8408] <= layer1_out[7897];
     layer2_out[8409] <= layer1_out[1455] & ~layer1_out[1454];
     layer2_out[8410] <= layer1_out[791];
     layer2_out[8411] <= layer1_out[7957] & layer1_out[7958];
     layer2_out[8412] <= ~(layer1_out[5200] ^ layer1_out[5201]);
     layer2_out[8413] <= ~(layer1_out[3003] & layer1_out[3004]);
     layer2_out[8414] <= layer1_out[11770] & ~layer1_out[11771];
     layer2_out[8415] <= layer1_out[10410];
     layer2_out[8416] <= ~layer1_out[1818];
     layer2_out[8417] <= ~layer1_out[979];
     layer2_out[8418] <= ~(layer1_out[8612] ^ layer1_out[8613]);
     layer2_out[8419] <= layer1_out[3372];
     layer2_out[8420] <= ~layer1_out[2990];
     layer2_out[8421] <= ~layer1_out[9396];
     layer2_out[8422] <= ~layer1_out[11713];
     layer2_out[8423] <= 1'b1;
     layer2_out[8424] <= layer1_out[1175] | layer1_out[1176];
     layer2_out[8425] <= layer1_out[6059] | layer1_out[6060];
     layer2_out[8426] <= ~(layer1_out[1708] ^ layer1_out[1709]);
     layer2_out[8427] <= layer1_out[10204];
     layer2_out[8428] <= ~layer1_out[7859] | layer1_out[7858];
     layer2_out[8429] <= ~layer1_out[11967] | layer1_out[11966];
     layer2_out[8430] <= layer1_out[7840] & ~layer1_out[7839];
     layer2_out[8431] <= layer1_out[10208];
     layer2_out[8432] <= ~layer1_out[10272] | layer1_out[10271];
     layer2_out[8433] <= layer1_out[11761] | layer1_out[11762];
     layer2_out[8434] <= layer1_out[10970] & ~layer1_out[10969];
     layer2_out[8435] <= layer1_out[10131];
     layer2_out[8436] <= ~layer1_out[7371];
     layer2_out[8437] <= ~layer1_out[9201];
     layer2_out[8438] <= layer1_out[3486];
     layer2_out[8439] <= ~layer1_out[5586] | layer1_out[5585];
     layer2_out[8440] <= ~(layer1_out[10068] | layer1_out[10069]);
     layer2_out[8441] <= layer1_out[970];
     layer2_out[8442] <= ~(layer1_out[4033] | layer1_out[4034]);
     layer2_out[8443] <= 1'b0;
     layer2_out[8444] <= layer1_out[6536] | layer1_out[6537];
     layer2_out[8445] <= layer1_out[6847] & ~layer1_out[6846];
     layer2_out[8446] <= ~layer1_out[4363];
     layer2_out[8447] <= ~layer1_out[4659] | layer1_out[4658];
     layer2_out[8448] <= layer1_out[8911] | layer1_out[8912];
     layer2_out[8449] <= layer1_out[11431] & ~layer1_out[11432];
     layer2_out[8450] <= ~layer1_out[4695] | layer1_out[4696];
     layer2_out[8451] <= layer1_out[4150];
     layer2_out[8452] <= layer1_out[1904];
     layer2_out[8453] <= layer1_out[6650];
     layer2_out[8454] <= ~layer1_out[2694] | layer1_out[2693];
     layer2_out[8455] <= ~(layer1_out[6102] ^ layer1_out[6103]);
     layer2_out[8456] <= ~(layer1_out[8080] ^ layer1_out[8081]);
     layer2_out[8457] <= ~layer1_out[258];
     layer2_out[8458] <= layer1_out[2162] | layer1_out[2163];
     layer2_out[8459] <= layer1_out[5538] ^ layer1_out[5539];
     layer2_out[8460] <= layer1_out[8435];
     layer2_out[8461] <= layer1_out[8295] | layer1_out[8296];
     layer2_out[8462] <= ~(layer1_out[9616] ^ layer1_out[9617]);
     layer2_out[8463] <= ~layer1_out[7223];
     layer2_out[8464] <= layer1_out[3792];
     layer2_out[8465] <= ~layer1_out[4357];
     layer2_out[8466] <= ~(layer1_out[4792] | layer1_out[4793]);
     layer2_out[8467] <= layer1_out[5440];
     layer2_out[8468] <= layer1_out[1345];
     layer2_out[8469] <= layer1_out[3051] & layer1_out[3052];
     layer2_out[8470] <= layer1_out[5262];
     layer2_out[8471] <= ~(layer1_out[10604] & layer1_out[10605]);
     layer2_out[8472] <= ~layer1_out[9644];
     layer2_out[8473] <= layer1_out[855];
     layer2_out[8474] <= ~(layer1_out[1008] & layer1_out[1009]);
     layer2_out[8475] <= ~layer1_out[8140] | layer1_out[8141];
     layer2_out[8476] <= ~layer1_out[6379];
     layer2_out[8477] <= ~(layer1_out[584] & layer1_out[585]);
     layer2_out[8478] <= ~layer1_out[3133] | layer1_out[3132];
     layer2_out[8479] <= layer1_out[7256] | layer1_out[7257];
     layer2_out[8480] <= ~(layer1_out[9176] & layer1_out[9177]);
     layer2_out[8481] <= ~layer1_out[4871];
     layer2_out[8482] <= ~layer1_out[1003];
     layer2_out[8483] <= layer1_out[948] & layer1_out[949];
     layer2_out[8484] <= layer1_out[6651];
     layer2_out[8485] <= layer1_out[2714] & layer1_out[2715];
     layer2_out[8486] <= layer1_out[10132];
     layer2_out[8487] <= ~layer1_out[2444];
     layer2_out[8488] <= ~layer1_out[4106];
     layer2_out[8489] <= layer1_out[9006] | layer1_out[9007];
     layer2_out[8490] <= layer1_out[39];
     layer2_out[8491] <= ~layer1_out[9350];
     layer2_out[8492] <= layer1_out[9896] ^ layer1_out[9897];
     layer2_out[8493] <= layer1_out[9259] & ~layer1_out[9258];
     layer2_out[8494] <= ~layer1_out[4587];
     layer2_out[8495] <= ~layer1_out[2571] | layer1_out[2570];
     layer2_out[8496] <= ~layer1_out[4053];
     layer2_out[8497] <= layer1_out[5632];
     layer2_out[8498] <= ~layer1_out[2537];
     layer2_out[8499] <= layer1_out[8127] & ~layer1_out[8126];
     layer2_out[8500] <= ~layer1_out[3650];
     layer2_out[8501] <= layer1_out[10025];
     layer2_out[8502] <= layer1_out[1867] & layer1_out[1868];
     layer2_out[8503] <= layer1_out[4461];
     layer2_out[8504] <= ~layer1_out[7308];
     layer2_out[8505] <= layer1_out[5917];
     layer2_out[8506] <= layer1_out[3524];
     layer2_out[8507] <= ~layer1_out[1590];
     layer2_out[8508] <= layer1_out[2923] | layer1_out[2924];
     layer2_out[8509] <= layer1_out[6665];
     layer2_out[8510] <= layer1_out[5776] | layer1_out[5777];
     layer2_out[8511] <= layer1_out[11692];
     layer2_out[8512] <= layer1_out[2531] & ~layer1_out[2530];
     layer2_out[8513] <= ~layer1_out[6342];
     layer2_out[8514] <= layer1_out[5721] | layer1_out[5722];
     layer2_out[8515] <= ~layer1_out[3933];
     layer2_out[8516] <= layer1_out[11367] ^ layer1_out[11368];
     layer2_out[8517] <= layer1_out[4916] & layer1_out[4917];
     layer2_out[8518] <= layer1_out[6546] & ~layer1_out[6547];
     layer2_out[8519] <= layer1_out[9420] & ~layer1_out[9419];
     layer2_out[8520] <= ~layer1_out[11830];
     layer2_out[8521] <= ~layer1_out[2728];
     layer2_out[8522] <= layer1_out[7597] & ~layer1_out[7596];
     layer2_out[8523] <= layer1_out[9325] & ~layer1_out[9324];
     layer2_out[8524] <= ~layer1_out[372];
     layer2_out[8525] <= ~(layer1_out[3614] ^ layer1_out[3615]);
     layer2_out[8526] <= layer1_out[5930];
     layer2_out[8527] <= ~layer1_out[1577];
     layer2_out[8528] <= layer1_out[1313];
     layer2_out[8529] <= layer1_out[11674];
     layer2_out[8530] <= layer1_out[4960] & layer1_out[4961];
     layer2_out[8531] <= layer1_out[4463];
     layer2_out[8532] <= ~layer1_out[315];
     layer2_out[8533] <= ~layer1_out[3560];
     layer2_out[8534] <= ~(layer1_out[6418] & layer1_out[6419]);
     layer2_out[8535] <= ~layer1_out[8221];
     layer2_out[8536] <= layer1_out[4764] & ~layer1_out[4763];
     layer2_out[8537] <= layer1_out[5345];
     layer2_out[8538] <= layer1_out[2115];
     layer2_out[8539] <= layer1_out[309];
     layer2_out[8540] <= layer1_out[10043];
     layer2_out[8541] <= ~(layer1_out[10651] & layer1_out[10652]);
     layer2_out[8542] <= ~layer1_out[11310] | layer1_out[11311];
     layer2_out[8543] <= ~layer1_out[7806] | layer1_out[7807];
     layer2_out[8544] <= ~layer1_out[9680];
     layer2_out[8545] <= layer1_out[9905];
     layer2_out[8546] <= ~layer1_out[2027];
     layer2_out[8547] <= 1'b1;
     layer2_out[8548] <= layer1_out[7457] & layer1_out[7458];
     layer2_out[8549] <= ~layer1_out[336];
     layer2_out[8550] <= layer1_out[10078] & ~layer1_out[10079];
     layer2_out[8551] <= ~(layer1_out[6230] & layer1_out[6231]);
     layer2_out[8552] <= layer1_out[4891] | layer1_out[4892];
     layer2_out[8553] <= ~(layer1_out[7404] ^ layer1_out[7405]);
     layer2_out[8554] <= layer1_out[10595] | layer1_out[10596];
     layer2_out[8555] <= 1'b1;
     layer2_out[8556] <= ~layer1_out[9284] | layer1_out[9285];
     layer2_out[8557] <= layer1_out[1099];
     layer2_out[8558] <= ~(layer1_out[11511] | layer1_out[11512]);
     layer2_out[8559] <= 1'b1;
     layer2_out[8560] <= layer1_out[646] & ~layer1_out[647];
     layer2_out[8561] <= ~layer1_out[7417];
     layer2_out[8562] <= layer1_out[5536] | layer1_out[5537];
     layer2_out[8563] <= layer1_out[1183];
     layer2_out[8564] <= ~layer1_out[6880] | layer1_out[6881];
     layer2_out[8565] <= layer1_out[11285] ^ layer1_out[11286];
     layer2_out[8566] <= ~(layer1_out[11362] ^ layer1_out[11363]);
     layer2_out[8567] <= ~layer1_out[10266];
     layer2_out[8568] <= ~layer1_out[194] | layer1_out[195];
     layer2_out[8569] <= layer1_out[11784] & ~layer1_out[11783];
     layer2_out[8570] <= layer1_out[1400];
     layer2_out[8571] <= layer1_out[6459];
     layer2_out[8572] <= layer1_out[11480] ^ layer1_out[11481];
     layer2_out[8573] <= ~layer1_out[1884];
     layer2_out[8574] <= layer1_out[849];
     layer2_out[8575] <= layer1_out[9924];
     layer2_out[8576] <= layer1_out[11744];
     layer2_out[8577] <= layer1_out[3128];
     layer2_out[8578] <= ~layer1_out[11549];
     layer2_out[8579] <= layer1_out[263] & ~layer1_out[262];
     layer2_out[8580] <= layer1_out[1014] & layer1_out[1015];
     layer2_out[8581] <= layer1_out[8747] & layer1_out[8748];
     layer2_out[8582] <= ~layer1_out[2088] | layer1_out[2089];
     layer2_out[8583] <= ~(layer1_out[1972] | layer1_out[1973]);
     layer2_out[8584] <= ~layer1_out[10858];
     layer2_out[8585] <= ~(layer1_out[4771] & layer1_out[4772]);
     layer2_out[8586] <= ~layer1_out[7895] | layer1_out[7896];
     layer2_out[8587] <= ~(layer1_out[4907] & layer1_out[4908]);
     layer2_out[8588] <= ~layer1_out[8692];
     layer2_out[8589] <= ~(layer1_out[9283] & layer1_out[9284]);
     layer2_out[8590] <= layer1_out[6700] & layer1_out[6701];
     layer2_out[8591] <= layer1_out[2601] | layer1_out[2602];
     layer2_out[8592] <= layer1_out[10627] ^ layer1_out[10628];
     layer2_out[8593] <= 1'b1;
     layer2_out[8594] <= layer1_out[1464];
     layer2_out[8595] <= layer1_out[44] & ~layer1_out[45];
     layer2_out[8596] <= ~layer1_out[2859] | layer1_out[2858];
     layer2_out[8597] <= layer1_out[5790] & ~layer1_out[5791];
     layer2_out[8598] <= layer1_out[4308] & ~layer1_out[4309];
     layer2_out[8599] <= layer1_out[11066] ^ layer1_out[11067];
     layer2_out[8600] <= layer1_out[10860];
     layer2_out[8601] <= layer1_out[50] & layer1_out[51];
     layer2_out[8602] <= layer1_out[9554];
     layer2_out[8603] <= ~layer1_out[1734];
     layer2_out[8604] <= ~layer1_out[918];
     layer2_out[8605] <= ~(layer1_out[10946] & layer1_out[10947]);
     layer2_out[8606] <= ~(layer1_out[4883] & layer1_out[4884]);
     layer2_out[8607] <= ~(layer1_out[8419] & layer1_out[8420]);
     layer2_out[8608] <= ~layer1_out[2566] | layer1_out[2565];
     layer2_out[8609] <= layer1_out[5694] | layer1_out[5695];
     layer2_out[8610] <= ~layer1_out[8720];
     layer2_out[8611] <= layer1_out[8146] ^ layer1_out[8147];
     layer2_out[8612] <= layer1_out[1267];
     layer2_out[8613] <= ~(layer1_out[2526] | layer1_out[2527]);
     layer2_out[8614] <= 1'b1;
     layer2_out[8615] <= layer1_out[9870];
     layer2_out[8616] <= ~layer1_out[1162];
     layer2_out[8617] <= layer1_out[4402] & ~layer1_out[4403];
     layer2_out[8618] <= ~layer1_out[11599];
     layer2_out[8619] <= layer1_out[7300];
     layer2_out[8620] <= ~(layer1_out[3534] ^ layer1_out[3535]);
     layer2_out[8621] <= ~(layer1_out[10129] | layer1_out[10130]);
     layer2_out[8622] <= ~layer1_out[139];
     layer2_out[8623] <= ~layer1_out[1809];
     layer2_out[8624] <= layer1_out[1095] & ~layer1_out[1094];
     layer2_out[8625] <= layer1_out[8429];
     layer2_out[8626] <= ~layer1_out[11189];
     layer2_out[8627] <= layer1_out[6828];
     layer2_out[8628] <= layer1_out[4756] | layer1_out[4757];
     layer2_out[8629] <= ~layer1_out[533];
     layer2_out[8630] <= ~layer1_out[4737] | layer1_out[4738];
     layer2_out[8631] <= layer1_out[5038];
     layer2_out[8632] <= layer1_out[7607];
     layer2_out[8633] <= layer1_out[9184] & ~layer1_out[9185];
     layer2_out[8634] <= layer1_out[5329];
     layer2_out[8635] <= layer1_out[274];
     layer2_out[8636] <= layer1_out[7581] & ~layer1_out[7580];
     layer2_out[8637] <= layer1_out[11127] & ~layer1_out[11128];
     layer2_out[8638] <= layer1_out[9201];
     layer2_out[8639] <= layer1_out[789];
     layer2_out[8640] <= layer1_out[1548];
     layer2_out[8641] <= ~(layer1_out[8472] ^ layer1_out[8473]);
     layer2_out[8642] <= layer1_out[11196] ^ layer1_out[11197];
     layer2_out[8643] <= layer1_out[222] & ~layer1_out[223];
     layer2_out[8644] <= layer1_out[8919] & ~layer1_out[8920];
     layer2_out[8645] <= layer1_out[11928] & layer1_out[11929];
     layer2_out[8646] <= ~layer1_out[10493];
     layer2_out[8647] <= layer1_out[4068] & ~layer1_out[4067];
     layer2_out[8648] <= layer1_out[2346] & ~layer1_out[2347];
     layer2_out[8649] <= ~layer1_out[3009];
     layer2_out[8650] <= layer1_out[4470] ^ layer1_out[4471];
     layer2_out[8651] <= ~(layer1_out[7493] | layer1_out[7494]);
     layer2_out[8652] <= ~(layer1_out[2148] & layer1_out[2149]);
     layer2_out[8653] <= layer1_out[6515];
     layer2_out[8654] <= 1'b0;
     layer2_out[8655] <= ~(layer1_out[9632] & layer1_out[9633]);
     layer2_out[8656] <= ~layer1_out[8271];
     layer2_out[8657] <= 1'b0;
     layer2_out[8658] <= layer1_out[11832];
     layer2_out[8659] <= ~layer1_out[11132];
     layer2_out[8660] <= ~layer1_out[10935] | layer1_out[10936];
     layer2_out[8661] <= ~layer1_out[2308];
     layer2_out[8662] <= ~layer1_out[11929] | layer1_out[11930];
     layer2_out[8663] <= ~(layer1_out[1252] & layer1_out[1253]);
     layer2_out[8664] <= ~(layer1_out[5537] | layer1_out[5538]);
     layer2_out[8665] <= layer1_out[3985] | layer1_out[3986];
     layer2_out[8666] <= layer1_out[4573];
     layer2_out[8667] <= ~layer1_out[6738];
     layer2_out[8668] <= layer1_out[4055] & ~layer1_out[4056];
     layer2_out[8669] <= layer1_out[10276] & layer1_out[10277];
     layer2_out[8670] <= ~layer1_out[6281];
     layer2_out[8671] <= ~layer1_out[2981];
     layer2_out[8672] <= layer1_out[4875] ^ layer1_out[4876];
     layer2_out[8673] <= ~layer1_out[6767];
     layer2_out[8674] <= layer1_out[10279];
     layer2_out[8675] <= layer1_out[313] & layer1_out[314];
     layer2_out[8676] <= layer1_out[9126] | layer1_out[9127];
     layer2_out[8677] <= ~(layer1_out[4925] | layer1_out[4926]);
     layer2_out[8678] <= ~layer1_out[7826] | layer1_out[7827];
     layer2_out[8679] <= ~layer1_out[7037];
     layer2_out[8680] <= layer1_out[5971] ^ layer1_out[5972];
     layer2_out[8681] <= layer1_out[2015] & ~layer1_out[2016];
     layer2_out[8682] <= layer1_out[9933];
     layer2_out[8683] <= layer1_out[723] & ~layer1_out[722];
     layer2_out[8684] <= layer1_out[11141];
     layer2_out[8685] <= ~layer1_out[1383] | layer1_out[1382];
     layer2_out[8686] <= layer1_out[4216];
     layer2_out[8687] <= layer1_out[6650];
     layer2_out[8688] <= ~(layer1_out[6135] | layer1_out[6136]);
     layer2_out[8689] <= ~layer1_out[6764] | layer1_out[6765];
     layer2_out[8690] <= layer1_out[11241];
     layer2_out[8691] <= layer1_out[5591] & ~layer1_out[5590];
     layer2_out[8692] <= layer1_out[989] ^ layer1_out[990];
     layer2_out[8693] <= ~layer1_out[6189];
     layer2_out[8694] <= layer1_out[8575];
     layer2_out[8695] <= layer1_out[3018];
     layer2_out[8696] <= layer1_out[679] ^ layer1_out[680];
     layer2_out[8697] <= ~(layer1_out[4627] ^ layer1_out[4628]);
     layer2_out[8698] <= layer1_out[103] & ~layer1_out[104];
     layer2_out[8699] <= layer1_out[2344];
     layer2_out[8700] <= layer1_out[5439];
     layer2_out[8701] <= layer1_out[5371] & layer1_out[5372];
     layer2_out[8702] <= layer1_out[9945];
     layer2_out[8703] <= layer1_out[8405];
     layer2_out[8704] <= ~layer1_out[741] | layer1_out[742];
     layer2_out[8705] <= ~layer1_out[5687];
     layer2_out[8706] <= ~layer1_out[9851];
     layer2_out[8707] <= layer1_out[4876] & ~layer1_out[4877];
     layer2_out[8708] <= layer1_out[4481];
     layer2_out[8709] <= ~layer1_out[7274];
     layer2_out[8710] <= layer1_out[10550] & ~layer1_out[10551];
     layer2_out[8711] <= ~layer1_out[10063];
     layer2_out[8712] <= ~layer1_out[11958];
     layer2_out[8713] <= layer1_out[8334] & layer1_out[8335];
     layer2_out[8714] <= ~(layer1_out[7311] & layer1_out[7312]);
     layer2_out[8715] <= ~layer1_out[3610] | layer1_out[3609];
     layer2_out[8716] <= ~(layer1_out[1112] ^ layer1_out[1113]);
     layer2_out[8717] <= layer1_out[3144];
     layer2_out[8718] <= layer1_out[1616] & layer1_out[1617];
     layer2_out[8719] <= layer1_out[8646] & ~layer1_out[8647];
     layer2_out[8720] <= layer1_out[2926];
     layer2_out[8721] <= layer1_out[10388];
     layer2_out[8722] <= layer1_out[2590] & ~layer1_out[2589];
     layer2_out[8723] <= ~layer1_out[5609] | layer1_out[5610];
     layer2_out[8724] <= layer1_out[9833];
     layer2_out[8725] <= ~(layer1_out[8713] ^ layer1_out[8714]);
     layer2_out[8726] <= layer1_out[7189] & layer1_out[7190];
     layer2_out[8727] <= layer1_out[5020] ^ layer1_out[5021];
     layer2_out[8728] <= ~(layer1_out[6932] | layer1_out[6933]);
     layer2_out[8729] <= layer1_out[8565] ^ layer1_out[8566];
     layer2_out[8730] <= layer1_out[5825] & ~layer1_out[5826];
     layer2_out[8731] <= layer1_out[5357];
     layer2_out[8732] <= layer1_out[4271] & ~layer1_out[4272];
     layer2_out[8733] <= ~layer1_out[2256];
     layer2_out[8734] <= ~layer1_out[3557] | layer1_out[3556];
     layer2_out[8735] <= ~(layer1_out[6818] & layer1_out[6819]);
     layer2_out[8736] <= ~layer1_out[10454];
     layer2_out[8737] <= ~layer1_out[7965] | layer1_out[7966];
     layer2_out[8738] <= layer1_out[5499] ^ layer1_out[5500];
     layer2_out[8739] <= 1'b0;
     layer2_out[8740] <= layer1_out[255];
     layer2_out[8741] <= ~layer1_out[2427];
     layer2_out[8742] <= ~layer1_out[4282];
     layer2_out[8743] <= layer1_out[11924] ^ layer1_out[11925];
     layer2_out[8744] <= ~(layer1_out[2972] | layer1_out[2973]);
     layer2_out[8745] <= layer1_out[8358] ^ layer1_out[8359];
     layer2_out[8746] <= ~layer1_out[6973];
     layer2_out[8747] <= ~layer1_out[3370] | layer1_out[3369];
     layer2_out[8748] <= ~(layer1_out[1682] | layer1_out[1683]);
     layer2_out[8749] <= layer1_out[2500] & layer1_out[2501];
     layer2_out[8750] <= layer1_out[8834];
     layer2_out[8751] <= ~layer1_out[9411] | layer1_out[9412];
     layer2_out[8752] <= ~(layer1_out[9707] | layer1_out[9708]);
     layer2_out[8753] <= layer1_out[10275];
     layer2_out[8754] <= layer1_out[11171] & ~layer1_out[11172];
     layer2_out[8755] <= layer1_out[6259] ^ layer1_out[6260];
     layer2_out[8756] <= ~layer1_out[5315] | layer1_out[5316];
     layer2_out[8757] <= ~(layer1_out[5994] | layer1_out[5995]);
     layer2_out[8758] <= ~layer1_out[4704];
     layer2_out[8759] <= ~layer1_out[3574];
     layer2_out[8760] <= layer1_out[8589] & ~layer1_out[8590];
     layer2_out[8761] <= ~layer1_out[1437];
     layer2_out[8762] <= layer1_out[5617];
     layer2_out[8763] <= ~layer1_out[9534];
     layer2_out[8764] <= ~(layer1_out[307] | layer1_out[308]);
     layer2_out[8765] <= layer1_out[608] ^ layer1_out[609];
     layer2_out[8766] <= ~layer1_out[5544] | layer1_out[5543];
     layer2_out[8767] <= layer1_out[7809];
     layer2_out[8768] <= layer1_out[11137] & layer1_out[11138];
     layer2_out[8769] <= ~layer1_out[9612] | layer1_out[9611];
     layer2_out[8770] <= ~layer1_out[4800];
     layer2_out[8771] <= ~layer1_out[10084];
     layer2_out[8772] <= layer1_out[5782] & ~layer1_out[5781];
     layer2_out[8773] <= ~(layer1_out[5392] & layer1_out[5393]);
     layer2_out[8774] <= layer1_out[9807];
     layer2_out[8775] <= ~layer1_out[4797];
     layer2_out[8776] <= ~(layer1_out[8308] & layer1_out[8309]);
     layer2_out[8777] <= layer1_out[2016] ^ layer1_out[2017];
     layer2_out[8778] <= layer1_out[116] | layer1_out[117];
     layer2_out[8779] <= layer1_out[1879];
     layer2_out[8780] <= ~layer1_out[10529] | layer1_out[10528];
     layer2_out[8781] <= layer1_out[8244] & ~layer1_out[8243];
     layer2_out[8782] <= layer1_out[4370];
     layer2_out[8783] <= layer1_out[3918] ^ layer1_out[3919];
     layer2_out[8784] <= ~layer1_out[4249] | layer1_out[4248];
     layer2_out[8785] <= layer1_out[7358] & ~layer1_out[7357];
     layer2_out[8786] <= layer1_out[9963] ^ layer1_out[9964];
     layer2_out[8787] <= ~layer1_out[2295];
     layer2_out[8788] <= layer1_out[2611];
     layer2_out[8789] <= ~(layer1_out[2009] ^ layer1_out[2010]);
     layer2_out[8790] <= layer1_out[8058] & ~layer1_out[8057];
     layer2_out[8791] <= ~(layer1_out[3949] ^ layer1_out[3950]);
     layer2_out[8792] <= layer1_out[10136];
     layer2_out[8793] <= layer1_out[11029];
     layer2_out[8794] <= layer1_out[3830] & layer1_out[3831];
     layer2_out[8795] <= ~(layer1_out[8807] | layer1_out[8808]);
     layer2_out[8796] <= layer1_out[1568];
     layer2_out[8797] <= layer1_out[6355] & ~layer1_out[6354];
     layer2_out[8798] <= ~layer1_out[9188] | layer1_out[9189];
     layer2_out[8799] <= ~layer1_out[7107];
     layer2_out[8800] <= ~layer1_out[7304];
     layer2_out[8801] <= ~(layer1_out[10569] & layer1_out[10570]);
     layer2_out[8802] <= layer1_out[3910];
     layer2_out[8803] <= ~layer1_out[11121] | layer1_out[11120];
     layer2_out[8804] <= ~layer1_out[5499];
     layer2_out[8805] <= ~layer1_out[2912];
     layer2_out[8806] <= layer1_out[8425];
     layer2_out[8807] <= layer1_out[11602];
     layer2_out[8808] <= layer1_out[11402] & layer1_out[11403];
     layer2_out[8809] <= layer1_out[5811] & ~layer1_out[5810];
     layer2_out[8810] <= ~layer1_out[8591] | layer1_out[8592];
     layer2_out[8811] <= ~(layer1_out[5985] ^ layer1_out[5986]);
     layer2_out[8812] <= layer1_out[6756] | layer1_out[6757];
     layer2_out[8813] <= ~(layer1_out[11383] | layer1_out[11384]);
     layer2_out[8814] <= layer1_out[6128];
     layer2_out[8815] <= ~(layer1_out[8407] | layer1_out[8408]);
     layer2_out[8816] <= layer1_out[2806] | layer1_out[2807];
     layer2_out[8817] <= ~layer1_out[10572];
     layer2_out[8818] <= ~layer1_out[1722];
     layer2_out[8819] <= layer1_out[2551] | layer1_out[2552];
     layer2_out[8820] <= ~(layer1_out[2300] | layer1_out[2301]);
     layer2_out[8821] <= layer1_out[10020] | layer1_out[10021];
     layer2_out[8822] <= ~layer1_out[5788];
     layer2_out[8823] <= ~layer1_out[9741];
     layer2_out[8824] <= ~(layer1_out[438] | layer1_out[439]);
     layer2_out[8825] <= layer1_out[10159] & layer1_out[10160];
     layer2_out[8826] <= ~layer1_out[5812];
     layer2_out[8827] <= layer1_out[3978] & ~layer1_out[3979];
     layer2_out[8828] <= layer1_out[967];
     layer2_out[8829] <= ~(layer1_out[9127] & layer1_out[9128]);
     layer2_out[8830] <= layer1_out[6593];
     layer2_out[8831] <= ~(layer1_out[5765] ^ layer1_out[5766]);
     layer2_out[8832] <= ~layer1_out[8944] | layer1_out[8943];
     layer2_out[8833] <= layer1_out[1211];
     layer2_out[8834] <= ~(layer1_out[11931] | layer1_out[11932]);
     layer2_out[8835] <= layer1_out[7697] & ~layer1_out[7698];
     layer2_out[8836] <= ~layer1_out[4680];
     layer2_out[8837] <= ~layer1_out[4924];
     layer2_out[8838] <= ~(layer1_out[4719] ^ layer1_out[4720]);
     layer2_out[8839] <= layer1_out[626] ^ layer1_out[627];
     layer2_out[8840] <= ~layer1_out[10658];
     layer2_out[8841] <= layer1_out[7086];
     layer2_out[8842] <= ~layer1_out[2117];
     layer2_out[8843] <= ~layer1_out[4122];
     layer2_out[8844] <= layer1_out[11133] & ~layer1_out[11134];
     layer2_out[8845] <= layer1_out[1275];
     layer2_out[8846] <= ~layer1_out[6159] | layer1_out[6158];
     layer2_out[8847] <= layer1_out[4431] | layer1_out[4432];
     layer2_out[8848] <= ~layer1_out[6997] | layer1_out[6998];
     layer2_out[8849] <= layer1_out[7651];
     layer2_out[8850] <= ~(layer1_out[2705] & layer1_out[2706]);
     layer2_out[8851] <= layer1_out[10602];
     layer2_out[8852] <= ~layer1_out[11799];
     layer2_out[8853] <= layer1_out[4262] & ~layer1_out[4261];
     layer2_out[8854] <= ~(layer1_out[730] ^ layer1_out[731]);
     layer2_out[8855] <= layer1_out[6781] & ~layer1_out[6782];
     layer2_out[8856] <= ~layer1_out[1145] | layer1_out[1146];
     layer2_out[8857] <= layer1_out[11808] & ~layer1_out[11809];
     layer2_out[8858] <= layer1_out[2528];
     layer2_out[8859] <= layer1_out[105] | layer1_out[106];
     layer2_out[8860] <= layer1_out[9188] & ~layer1_out[9187];
     layer2_out[8861] <= ~layer1_out[11952];
     layer2_out[8862] <= layer1_out[8723] ^ layer1_out[8724];
     layer2_out[8863] <= layer1_out[7048] | layer1_out[7049];
     layer2_out[8864] <= layer1_out[1148] & ~layer1_out[1149];
     layer2_out[8865] <= ~layer1_out[2412];
     layer2_out[8866] <= layer1_out[3976] | layer1_out[3977];
     layer2_out[8867] <= layer1_out[3875];
     layer2_out[8868] <= layer1_out[3074];
     layer2_out[8869] <= layer1_out[11900];
     layer2_out[8870] <= ~layer1_out[7505] | layer1_out[7504];
     layer2_out[8871] <= layer1_out[8062] & layer1_out[8063];
     layer2_out[8872] <= ~layer1_out[2751];
     layer2_out[8873] <= ~layer1_out[1510] | layer1_out[1511];
     layer2_out[8874] <= layer1_out[7880] & layer1_out[7881];
     layer2_out[8875] <= layer1_out[4376] & ~layer1_out[4375];
     layer2_out[8876] <= layer1_out[7267] ^ layer1_out[7268];
     layer2_out[8877] <= layer1_out[10504] ^ layer1_out[10505];
     layer2_out[8878] <= ~layer1_out[4269] | layer1_out[4268];
     layer2_out[8879] <= layer1_out[3953];
     layer2_out[8880] <= ~layer1_out[354];
     layer2_out[8881] <= layer1_out[572] & ~layer1_out[573];
     layer2_out[8882] <= ~(layer1_out[1110] | layer1_out[1111]);
     layer2_out[8883] <= layer1_out[11919];
     layer2_out[8884] <= ~(layer1_out[11453] ^ layer1_out[11454]);
     layer2_out[8885] <= layer1_out[3998] ^ layer1_out[3999];
     layer2_out[8886] <= ~layer1_out[499];
     layer2_out[8887] <= layer1_out[7031];
     layer2_out[8888] <= layer1_out[36] ^ layer1_out[37];
     layer2_out[8889] <= layer1_out[6647];
     layer2_out[8890] <= ~(layer1_out[8805] | layer1_out[8806]);
     layer2_out[8891] <= layer1_out[8416];
     layer2_out[8892] <= ~(layer1_out[9472] & layer1_out[9473]);
     layer2_out[8893] <= 1'b0;
     layer2_out[8894] <= ~layer1_out[1028];
     layer2_out[8895] <= ~layer1_out[11153] | layer1_out[11152];
     layer2_out[8896] <= ~(layer1_out[1410] | layer1_out[1411]);
     layer2_out[8897] <= ~(layer1_out[2726] | layer1_out[2727]);
     layer2_out[8898] <= layer1_out[10179] ^ layer1_out[10180];
     layer2_out[8899] <= layer1_out[4511] ^ layer1_out[4512];
     layer2_out[8900] <= ~layer1_out[8115] | layer1_out[8114];
     layer2_out[8901] <= layer1_out[1760];
     layer2_out[8902] <= layer1_out[7837] & ~layer1_out[7836];
     layer2_out[8903] <= layer1_out[5946] & ~layer1_out[5945];
     layer2_out[8904] <= ~layer1_out[4104];
     layer2_out[8905] <= 1'b1;
     layer2_out[8906] <= layer1_out[5420] ^ layer1_out[5421];
     layer2_out[8907] <= ~(layer1_out[8040] | layer1_out[8041]);
     layer2_out[8908] <= ~layer1_out[10383];
     layer2_out[8909] <= layer1_out[2007] & ~layer1_out[2008];
     layer2_out[8910] <= layer1_out[467] & ~layer1_out[468];
     layer2_out[8911] <= ~layer1_out[8074] | layer1_out[8073];
     layer2_out[8912] <= layer1_out[7252];
     layer2_out[8913] <= ~layer1_out[4293];
     layer2_out[8914] <= layer1_out[11496] & layer1_out[11497];
     layer2_out[8915] <= layer1_out[9152];
     layer2_out[8916] <= ~(layer1_out[1905] & layer1_out[1906]);
     layer2_out[8917] <= layer1_out[11764] | layer1_out[11765];
     layer2_out[8918] <= ~(layer1_out[9438] | layer1_out[9439]);
     layer2_out[8919] <= layer1_out[7982];
     layer2_out[8920] <= layer1_out[6449] | layer1_out[6450];
     layer2_out[8921] <= ~layer1_out[2101];
     layer2_out[8922] <= layer1_out[6112] & ~layer1_out[6113];
     layer2_out[8923] <= layer1_out[5408] & layer1_out[5409];
     layer2_out[8924] <= layer1_out[1342];
     layer2_out[8925] <= layer1_out[3991];
     layer2_out[8926] <= layer1_out[581] & layer1_out[582];
     layer2_out[8927] <= ~layer1_out[4455] | layer1_out[4456];
     layer2_out[8928] <= ~layer1_out[8751] | layer1_out[8752];
     layer2_out[8929] <= ~layer1_out[9426] | layer1_out[9427];
     layer2_out[8930] <= ~layer1_out[11238];
     layer2_out[8931] <= layer1_out[10186];
     layer2_out[8932] <= ~layer1_out[10597] | layer1_out[10596];
     layer2_out[8933] <= ~layer1_out[1602];
     layer2_out[8934] <= layer1_out[5040];
     layer2_out[8935] <= ~layer1_out[9349];
     layer2_out[8936] <= layer1_out[7889];
     layer2_out[8937] <= ~layer1_out[3109];
     layer2_out[8938] <= layer1_out[194];
     layer2_out[8939] <= layer1_out[6934] & ~layer1_out[6935];
     layer2_out[8940] <= ~(layer1_out[10957] ^ layer1_out[10958]);
     layer2_out[8941] <= ~layer1_out[10587] | layer1_out[10586];
     layer2_out[8942] <= layer1_out[8421];
     layer2_out[8943] <= ~layer1_out[2416] | layer1_out[2415];
     layer2_out[8944] <= layer1_out[8886] & ~layer1_out[8887];
     layer2_out[8945] <= layer1_out[4739] & ~layer1_out[4740];
     layer2_out[8946] <= ~layer1_out[8191] | layer1_out[8192];
     layer2_out[8947] <= layer1_out[3930] | layer1_out[3931];
     layer2_out[8948] <= layer1_out[10831];
     layer2_out[8949] <= layer1_out[8396] & ~layer1_out[8395];
     layer2_out[8950] <= ~layer1_out[10073] | layer1_out[10074];
     layer2_out[8951] <= ~layer1_out[1051];
     layer2_out[8952] <= layer1_out[2906];
     layer2_out[8953] <= layer1_out[8242] & ~layer1_out[8243];
     layer2_out[8954] <= layer1_out[4828] & ~layer1_out[4829];
     layer2_out[8955] <= layer1_out[3512];
     layer2_out[8956] <= layer1_out[11476];
     layer2_out[8957] <= layer1_out[10972];
     layer2_out[8958] <= layer1_out[10451];
     layer2_out[8959] <= layer1_out[11834];
     layer2_out[8960] <= layer1_out[10303] | layer1_out[10304];
     layer2_out[8961] <= ~layer1_out[8621] | layer1_out[8622];
     layer2_out[8962] <= layer1_out[1747] & ~layer1_out[1746];
     layer2_out[8963] <= layer1_out[7387] & layer1_out[7388];
     layer2_out[8964] <= ~(layer1_out[9816] | layer1_out[9817]);
     layer2_out[8965] <= ~(layer1_out[11045] & layer1_out[11046]);
     layer2_out[8966] <= 1'b0;
     layer2_out[8967] <= ~layer1_out[8151] | layer1_out[8152];
     layer2_out[8968] <= layer1_out[7561];
     layer2_out[8969] <= layer1_out[573] | layer1_out[574];
     layer2_out[8970] <= layer1_out[1159] | layer1_out[1160];
     layer2_out[8971] <= layer1_out[4814];
     layer2_out[8972] <= layer1_out[1514];
     layer2_out[8973] <= layer1_out[7715] & ~layer1_out[7716];
     layer2_out[8974] <= 1'b1;
     layer2_out[8975] <= layer1_out[7920] ^ layer1_out[7921];
     layer2_out[8976] <= ~layer1_out[3981] | layer1_out[3982];
     layer2_out[8977] <= ~layer1_out[4035];
     layer2_out[8978] <= layer1_out[1024] | layer1_out[1025];
     layer2_out[8979] <= ~(layer1_out[5777] | layer1_out[5778]);
     layer2_out[8980] <= layer1_out[10113] ^ layer1_out[10114];
     layer2_out[8981] <= layer1_out[11908] & ~layer1_out[11907];
     layer2_out[8982] <= ~layer1_out[10921];
     layer2_out[8983] <= layer1_out[4198] & layer1_out[4199];
     layer2_out[8984] <= layer1_out[9651] ^ layer1_out[9652];
     layer2_out[8985] <= ~(layer1_out[7021] | layer1_out[7022]);
     layer2_out[8986] <= ~layer1_out[1058];
     layer2_out[8987] <= layer1_out[10349] & layer1_out[10350];
     layer2_out[8988] <= ~layer1_out[6454];
     layer2_out[8989] <= layer1_out[10252];
     layer2_out[8990] <= ~layer1_out[7403];
     layer2_out[8991] <= ~layer1_out[10819] | layer1_out[10820];
     layer2_out[8992] <= ~layer1_out[6713] | layer1_out[6712];
     layer2_out[8993] <= ~layer1_out[8618];
     layer2_out[8994] <= layer1_out[4747] & ~layer1_out[4746];
     layer2_out[8995] <= layer1_out[2143] & layer1_out[2144];
     layer2_out[8996] <= layer1_out[2397];
     layer2_out[8997] <= ~(layer1_out[7378] ^ layer1_out[7379]);
     layer2_out[8998] <= layer1_out[4063] | layer1_out[4064];
     layer2_out[8999] <= ~(layer1_out[34] | layer1_out[35]);
     layer2_out[9000] <= ~layer1_out[11491];
     layer2_out[9001] <= ~layer1_out[11537] | layer1_out[11536];
     layer2_out[9002] <= layer1_out[1191] & layer1_out[1192];
     layer2_out[9003] <= layer1_out[3033];
     layer2_out[9004] <= ~layer1_out[10890];
     layer2_out[9005] <= layer1_out[11299] & ~layer1_out[11300];
     layer2_out[9006] <= ~(layer1_out[133] & layer1_out[134]);
     layer2_out[9007] <= layer1_out[9703];
     layer2_out[9008] <= layer1_out[6943];
     layer2_out[9009] <= layer1_out[8492] | layer1_out[8493];
     layer2_out[9010] <= ~(layer1_out[2969] | layer1_out[2970]);
     layer2_out[9011] <= layer1_out[11275] & layer1_out[11276];
     layer2_out[9012] <= layer1_out[9758];
     layer2_out[9013] <= layer1_out[7657];
     layer2_out[9014] <= layer1_out[6332] ^ layer1_out[6333];
     layer2_out[9015] <= layer1_out[8228] & ~layer1_out[8227];
     layer2_out[9016] <= ~layer1_out[6864] | layer1_out[6865];
     layer2_out[9017] <= ~(layer1_out[1735] | layer1_out[1736]);
     layer2_out[9018] <= layer1_out[8657];
     layer2_out[9019] <= 1'b0;
     layer2_out[9020] <= layer1_out[10480] & ~layer1_out[10479];
     layer2_out[9021] <= ~(layer1_out[11772] & layer1_out[11773]);
     layer2_out[9022] <= ~layer1_out[6276] | layer1_out[6275];
     layer2_out[9023] <= ~layer1_out[6289];
     layer2_out[9024] <= layer1_out[5133] | layer1_out[5134];
     layer2_out[9025] <= layer1_out[5928] ^ layer1_out[5929];
     layer2_out[9026] <= layer1_out[785] & ~layer1_out[784];
     layer2_out[9027] <= ~layer1_out[11649];
     layer2_out[9028] <= ~layer1_out[5545];
     layer2_out[9029] <= ~(layer1_out[7180] & layer1_out[7181]);
     layer2_out[9030] <= layer1_out[10227] | layer1_out[10228];
     layer2_out[9031] <= ~(layer1_out[5574] ^ layer1_out[5575]);
     layer2_out[9032] <= ~layer1_out[6183] | layer1_out[6184];
     layer2_out[9033] <= layer1_out[1937];
     layer2_out[9034] <= layer1_out[3479] & layer1_out[3480];
     layer2_out[9035] <= layer1_out[7108];
     layer2_out[9036] <= ~layer1_out[7001];
     layer2_out[9037] <= ~(layer1_out[11946] ^ layer1_out[11947]);
     layer2_out[9038] <= layer1_out[4636] ^ layer1_out[4637];
     layer2_out[9039] <= layer1_out[11723] & ~layer1_out[11722];
     layer2_out[9040] <= layer1_out[6191] & ~layer1_out[6190];
     layer2_out[9041] <= layer1_out[10344] & ~layer1_out[10345];
     layer2_out[9042] <= ~layer1_out[2629] | layer1_out[2628];
     layer2_out[9043] <= layer1_out[10318] & layer1_out[10319];
     layer2_out[9044] <= layer1_out[7375] & layer1_out[7376];
     layer2_out[9045] <= ~layer1_out[1511] | layer1_out[1512];
     layer2_out[9046] <= layer1_out[8777] & ~layer1_out[8776];
     layer2_out[9047] <= ~(layer1_out[5465] ^ layer1_out[5466]);
     layer2_out[9048] <= ~(layer1_out[11930] & layer1_out[11931]);
     layer2_out[9049] <= ~layer1_out[11579];
     layer2_out[9050] <= ~layer1_out[2023];
     layer2_out[9051] <= ~layer1_out[11979];
     layer2_out[9052] <= layer1_out[3373] | layer1_out[3374];
     layer2_out[9053] <= ~(layer1_out[6407] ^ layer1_out[6408]);
     layer2_out[9054] <= layer1_out[6968] & ~layer1_out[6969];
     layer2_out[9055] <= ~(layer1_out[3528] & layer1_out[3529]);
     layer2_out[9056] <= ~(layer1_out[8883] & layer1_out[8884]);
     layer2_out[9057] <= ~(layer1_out[9437] & layer1_out[9438]);
     layer2_out[9058] <= ~layer1_out[2425];
     layer2_out[9059] <= ~layer1_out[1176];
     layer2_out[9060] <= layer1_out[8521] & ~layer1_out[8522];
     layer2_out[9061] <= ~(layer1_out[7819] | layer1_out[7820]);
     layer2_out[9062] <= ~layer1_out[6722] | layer1_out[6721];
     layer2_out[9063] <= ~(layer1_out[10021] | layer1_out[10022]);
     layer2_out[9064] <= ~(layer1_out[4346] | layer1_out[4347]);
     layer2_out[9065] <= ~layer1_out[1327];
     layer2_out[9066] <= layer1_out[11326] | layer1_out[11327];
     layer2_out[9067] <= layer1_out[9032] & layer1_out[9033];
     layer2_out[9068] <= ~layer1_out[10178] | layer1_out[10177];
     layer2_out[9069] <= ~(layer1_out[4768] | layer1_out[4769]);
     layer2_out[9070] <= layer1_out[1617];
     layer2_out[9071] <= layer1_out[10064] | layer1_out[10065];
     layer2_out[9072] <= ~layer1_out[7408];
     layer2_out[9073] <= layer1_out[8051];
     layer2_out[9074] <= 1'b1;
     layer2_out[9075] <= ~layer1_out[4854];
     layer2_out[9076] <= layer1_out[9364] & ~layer1_out[9363];
     layer2_out[9077] <= layer1_out[10189];
     layer2_out[9078] <= layer1_out[7245];
     layer2_out[9079] <= layer1_out[4797] & ~layer1_out[4796];
     layer2_out[9080] <= layer1_out[10219] & ~layer1_out[10220];
     layer2_out[9081] <= ~layer1_out[10120] | layer1_out[10121];
     layer2_out[9082] <= ~(layer1_out[8374] | layer1_out[8375]);
     layer2_out[9083] <= layer1_out[11184];
     layer2_out[9084] <= ~layer1_out[449];
     layer2_out[9085] <= ~layer1_out[3175];
     layer2_out[9086] <= layer1_out[4601] & ~layer1_out[4602];
     layer2_out[9087] <= layer1_out[8206] & ~layer1_out[8205];
     layer2_out[9088] <= layer1_out[11092] & layer1_out[11093];
     layer2_out[9089] <= ~layer1_out[5940] | layer1_out[5939];
     layer2_out[9090] <= layer1_out[4571] ^ layer1_out[4572];
     layer2_out[9091] <= layer1_out[2999] & ~layer1_out[2998];
     layer2_out[9092] <= layer1_out[8020] | layer1_out[8021];
     layer2_out[9093] <= ~(layer1_out[3072] & layer1_out[3073]);
     layer2_out[9094] <= layer1_out[11387] & ~layer1_out[11388];
     layer2_out[9095] <= ~layer1_out[1751] | layer1_out[1752];
     layer2_out[9096] <= layer1_out[4888];
     layer2_out[9097] <= layer1_out[9063] | layer1_out[9064];
     layer2_out[9098] <= ~layer1_out[3090];
     layer2_out[9099] <= layer1_out[5462] | layer1_out[5463];
     layer2_out[9100] <= layer1_out[4832];
     layer2_out[9101] <= ~(layer1_out[3999] ^ layer1_out[4000]);
     layer2_out[9102] <= layer1_out[11450];
     layer2_out[9103] <= layer1_out[11170] ^ layer1_out[11171];
     layer2_out[9104] <= layer1_out[1631] ^ layer1_out[1632];
     layer2_out[9105] <= layer1_out[4933];
     layer2_out[9106] <= ~(layer1_out[7093] | layer1_out[7094]);
     layer2_out[9107] <= ~layer1_out[11952];
     layer2_out[9108] <= layer1_out[9624];
     layer2_out[9109] <= layer1_out[897] & layer1_out[898];
     layer2_out[9110] <= ~layer1_out[2658] | layer1_out[2659];
     layer2_out[9111] <= ~(layer1_out[10652] | layer1_out[10653]);
     layer2_out[9112] <= layer1_out[5458] & layer1_out[5459];
     layer2_out[9113] <= layer1_out[11875] & ~layer1_out[11874];
     layer2_out[9114] <= layer1_out[11760];
     layer2_out[9115] <= layer1_out[4749] & layer1_out[4750];
     layer2_out[9116] <= ~layer1_out[9223];
     layer2_out[9117] <= layer1_out[4083] ^ layer1_out[4084];
     layer2_out[9118] <= layer1_out[9306];
     layer2_out[9119] <= ~(layer1_out[10683] ^ layer1_out[10684]);
     layer2_out[9120] <= ~layer1_out[6737];
     layer2_out[9121] <= ~layer1_out[10477];
     layer2_out[9122] <= ~layer1_out[1957] | layer1_out[1958];
     layer2_out[9123] <= layer1_out[6773] ^ layer1_out[6774];
     layer2_out[9124] <= ~(layer1_out[8664] | layer1_out[8665]);
     layer2_out[9125] <= layer1_out[6052];
     layer2_out[9126] <= ~layer1_out[1708];
     layer2_out[9127] <= ~layer1_out[10252];
     layer2_out[9128] <= layer1_out[6691] ^ layer1_out[6692];
     layer2_out[9129] <= ~layer1_out[11564];
     layer2_out[9130] <= layer1_out[8637] & ~layer1_out[8636];
     layer2_out[9131] <= ~(layer1_out[8945] & layer1_out[8946]);
     layer2_out[9132] <= ~layer1_out[7555];
     layer2_out[9133] <= ~layer1_out[7212];
     layer2_out[9134] <= ~(layer1_out[4047] ^ layer1_out[4048]);
     layer2_out[9135] <= ~layer1_out[593];
     layer2_out[9136] <= layer1_out[11877];
     layer2_out[9137] <= ~layer1_out[11998];
     layer2_out[9138] <= layer1_out[6092] ^ layer1_out[6093];
     layer2_out[9139] <= ~(layer1_out[1713] & layer1_out[1714]);
     layer2_out[9140] <= layer1_out[4973] & ~layer1_out[4974];
     layer2_out[9141] <= ~(layer1_out[8173] & layer1_out[8174]);
     layer2_out[9142] <= ~layer1_out[11893];
     layer2_out[9143] <= layer1_out[7155];
     layer2_out[9144] <= layer1_out[6206] & ~layer1_out[6207];
     layer2_out[9145] <= layer1_out[2866] ^ layer1_out[2867];
     layer2_out[9146] <= ~layer1_out[7864];
     layer2_out[9147] <= ~(layer1_out[11741] & layer1_out[11742]);
     layer2_out[9148] <= ~layer1_out[9081];
     layer2_out[9149] <= layer1_out[2714] & ~layer1_out[2713];
     layer2_out[9150] <= layer1_out[3149] & layer1_out[3150];
     layer2_out[9151] <= layer1_out[9647];
     layer2_out[9152] <= layer1_out[8838] & layer1_out[8839];
     layer2_out[9153] <= ~(layer1_out[4323] | layer1_out[4324]);
     layer2_out[9154] <= layer1_out[7799];
     layer2_out[9155] <= layer1_out[1021] & ~layer1_out[1022];
     layer2_out[9156] <= layer1_out[3359] | layer1_out[3360];
     layer2_out[9157] <= ~(layer1_out[124] & layer1_out[125]);
     layer2_out[9158] <= layer1_out[7183] ^ layer1_out[7184];
     layer2_out[9159] <= ~(layer1_out[325] & layer1_out[326]);
     layer2_out[9160] <= ~layer1_out[3083] | layer1_out[3082];
     layer2_out[9161] <= ~layer1_out[3314];
     layer2_out[9162] <= layer1_out[3717] ^ layer1_out[3718];
     layer2_out[9163] <= ~layer1_out[8485];
     layer2_out[9164] <= layer1_out[5905];
     layer2_out[9165] <= layer1_out[9990];
     layer2_out[9166] <= ~(layer1_out[4441] | layer1_out[4442]);
     layer2_out[9167] <= ~layer1_out[1082] | layer1_out[1081];
     layer2_out[9168] <= ~(layer1_out[5351] & layer1_out[5352]);
     layer2_out[9169] <= 1'b0;
     layer2_out[9170] <= ~layer1_out[1570] | layer1_out[1571];
     layer2_out[9171] <= layer1_out[4291] ^ layer1_out[4292];
     layer2_out[9172] <= ~(layer1_out[5140] | layer1_out[5141]);
     layer2_out[9173] <= ~(layer1_out[2234] | layer1_out[2235]);
     layer2_out[9174] <= layer1_out[2438];
     layer2_out[9175] <= layer1_out[4253];
     layer2_out[9176] <= layer1_out[10426];
     layer2_out[9177] <= ~(layer1_out[7534] & layer1_out[7535]);
     layer2_out[9178] <= layer1_out[11033];
     layer2_out[9179] <= layer1_out[4684] & ~layer1_out[4685];
     layer2_out[9180] <= layer1_out[1856] & layer1_out[1857];
     layer2_out[9181] <= ~(layer1_out[4454] & layer1_out[4455]);
     layer2_out[9182] <= layer1_out[3213] & ~layer1_out[3212];
     layer2_out[9183] <= ~layer1_out[3600];
     layer2_out[9184] <= ~(layer1_out[1308] ^ layer1_out[1309]);
     layer2_out[9185] <= layer1_out[2375];
     layer2_out[9186] <= ~(layer1_out[4815] | layer1_out[4816]);
     layer2_out[9187] <= ~(layer1_out[10699] | layer1_out[10700]);
     layer2_out[9188] <= layer1_out[9117] & layer1_out[9118];
     layer2_out[9189] <= layer1_out[4505] & ~layer1_out[4504];
     layer2_out[9190] <= layer1_out[10929] ^ layer1_out[10930];
     layer2_out[9191] <= layer1_out[7069] ^ layer1_out[7070];
     layer2_out[9192] <= ~(layer1_out[811] & layer1_out[812]);
     layer2_out[9193] <= layer1_out[11954] & ~layer1_out[11955];
     layer2_out[9194] <= layer1_out[6760] | layer1_out[6761];
     layer2_out[9195] <= ~layer1_out[2784] | layer1_out[2785];
     layer2_out[9196] <= layer1_out[2186];
     layer2_out[9197] <= ~layer1_out[7569] | layer1_out[7568];
     layer2_out[9198] <= ~(layer1_out[4645] & layer1_out[4646]);
     layer2_out[9199] <= layer1_out[1992] & ~layer1_out[1991];
     layer2_out[9200] <= layer1_out[6445];
     layer2_out[9201] <= ~(layer1_out[5829] ^ layer1_out[5830]);
     layer2_out[9202] <= 1'b0;
     layer2_out[9203] <= ~layer1_out[327] | layer1_out[328];
     layer2_out[9204] <= layer1_out[10806] & ~layer1_out[10807];
     layer2_out[9205] <= ~layer1_out[6633];
     layer2_out[9206] <= ~layer1_out[9225] | layer1_out[9224];
     layer2_out[9207] <= ~layer1_out[9688] | layer1_out[9687];
     layer2_out[9208] <= layer1_out[2435];
     layer2_out[9209] <= layer1_out[11729];
     layer2_out[9210] <= 1'b1;
     layer2_out[9211] <= ~layer1_out[6837];
     layer2_out[9212] <= layer1_out[9330] & ~layer1_out[9329];
     layer2_out[9213] <= layer1_out[1281] & ~layer1_out[1280];
     layer2_out[9214] <= ~(layer1_out[5936] & layer1_out[5937]);
     layer2_out[9215] <= layer1_out[11316];
     layer2_out[9216] <= ~layer1_out[8711] | layer1_out[8710];
     layer2_out[9217] <= layer1_out[2968] & ~layer1_out[2967];
     layer2_out[9218] <= ~layer1_out[10190];
     layer2_out[9219] <= layer1_out[7083];
     layer2_out[9220] <= ~layer1_out[6787];
     layer2_out[9221] <= ~layer1_out[3288] | layer1_out[3289];
     layer2_out[9222] <= layer1_out[10172];
     layer2_out[9223] <= layer1_out[9673] | layer1_out[9674];
     layer2_out[9224] <= layer1_out[10201] | layer1_out[10202];
     layer2_out[9225] <= layer1_out[6518] & ~layer1_out[6519];
     layer2_out[9226] <= layer1_out[8980] & ~layer1_out[8981];
     layer2_out[9227] <= ~layer1_out[11306];
     layer2_out[9228] <= layer1_out[5280] | layer1_out[5281];
     layer2_out[9229] <= ~(layer1_out[7677] | layer1_out[7678]);
     layer2_out[9230] <= ~layer1_out[4096];
     layer2_out[9231] <= layer1_out[2739];
     layer2_out[9232] <= ~(layer1_out[4317] ^ layer1_out[4318]);
     layer2_out[9233] <= ~(layer1_out[10364] | layer1_out[10365]);
     layer2_out[9234] <= ~layer1_out[88] | layer1_out[89];
     layer2_out[9235] <= ~layer1_out[9020] | layer1_out[9019];
     layer2_out[9236] <= layer1_out[11198];
     layer2_out[9237] <= layer1_out[1313];
     layer2_out[9238] <= ~(layer1_out[7278] | layer1_out[7279]);
     layer2_out[9239] <= layer1_out[7829];
     layer2_out[9240] <= 1'b1;
     layer2_out[9241] <= ~(layer1_out[11058] ^ layer1_out[11059]);
     layer2_out[9242] <= ~layer1_out[8844];
     layer2_out[9243] <= ~layer1_out[4740];
     layer2_out[9244] <= layer1_out[786];
     layer2_out[9245] <= ~(layer1_out[8796] & layer1_out[8797]);
     layer2_out[9246] <= layer1_out[7639] ^ layer1_out[7640];
     layer2_out[9247] <= ~layer1_out[3323];
     layer2_out[9248] <= layer1_out[4005] ^ layer1_out[4006];
     layer2_out[9249] <= ~(layer1_out[8952] & layer1_out[8953]);
     layer2_out[9250] <= layer1_out[5995];
     layer2_out[9251] <= ~layer1_out[9120];
     layer2_out[9252] <= layer1_out[3409] & ~layer1_out[3408];
     layer2_out[9253] <= layer1_out[3577];
     layer2_out[9254] <= ~(layer1_out[710] | layer1_out[711]);
     layer2_out[9255] <= ~layer1_out[7497];
     layer2_out[9256] <= ~layer1_out[5420];
     layer2_out[9257] <= ~layer1_out[10673] | layer1_out[10674];
     layer2_out[9258] <= layer1_out[8027];
     layer2_out[9259] <= ~(layer1_out[507] & layer1_out[508]);
     layer2_out[9260] <= layer1_out[4442];
     layer2_out[9261] <= ~(layer1_out[5747] | layer1_out[5748]);
     layer2_out[9262] <= ~(layer1_out[8330] & layer1_out[8331]);
     layer2_out[9263] <= ~layer1_out[100] | layer1_out[99];
     layer2_out[9264] <= layer1_out[2213] & ~layer1_out[2214];
     layer2_out[9265] <= ~layer1_out[7702] | layer1_out[7701];
     layer2_out[9266] <= layer1_out[9164] & ~layer1_out[9165];
     layer2_out[9267] <= layer1_out[8210];
     layer2_out[9268] <= ~layer1_out[1653] | layer1_out[1654];
     layer2_out[9269] <= layer1_out[9154] & ~layer1_out[9153];
     layer2_out[9270] <= ~(layer1_out[3590] ^ layer1_out[3591]);
     layer2_out[9271] <= layer1_out[1009] & layer1_out[1010];
     layer2_out[9272] <= ~layer1_out[10269];
     layer2_out[9273] <= 1'b0;
     layer2_out[9274] <= layer1_out[8810] & layer1_out[8811];
     layer2_out[9275] <= layer1_out[3707] | layer1_out[3708];
     layer2_out[9276] <= ~layer1_out[5714];
     layer2_out[9277] <= layer1_out[4117];
     layer2_out[9278] <= layer1_out[7533] ^ layer1_out[7534];
     layer2_out[9279] <= ~layer1_out[9616] | layer1_out[9615];
     layer2_out[9280] <= ~layer1_out[11302] | layer1_out[11301];
     layer2_out[9281] <= layer1_out[6730];
     layer2_out[9282] <= ~layer1_out[3869] | layer1_out[3868];
     layer2_out[9283] <= ~(layer1_out[2270] & layer1_out[2271]);
     layer2_out[9284] <= layer1_out[2842];
     layer2_out[9285] <= layer1_out[6622] & ~layer1_out[6623];
     layer2_out[9286] <= ~layer1_out[8829] | layer1_out[8830];
     layer2_out[9287] <= ~layer1_out[8867] | layer1_out[8866];
     layer2_out[9288] <= layer1_out[9459] | layer1_out[9460];
     layer2_out[9289] <= layer1_out[1706] & ~layer1_out[1705];
     layer2_out[9290] <= layer1_out[8793];
     layer2_out[9291] <= ~layer1_out[214];
     layer2_out[9292] <= layer1_out[6305] & layer1_out[6306];
     layer2_out[9293] <= layer1_out[11879] & layer1_out[11880];
     layer2_out[9294] <= layer1_out[7018];
     layer2_out[9295] <= ~layer1_out[9908];
     layer2_out[9296] <= ~layer1_out[7795] | layer1_out[7796];
     layer2_out[9297] <= layer1_out[727] & layer1_out[728];
     layer2_out[9298] <= layer1_out[2740] & ~layer1_out[2741];
     layer2_out[9299] <= layer1_out[9008];
     layer2_out[9300] <= ~layer1_out[2284] | layer1_out[2283];
     layer2_out[9301] <= layer1_out[11217];
     layer2_out[9302] <= layer1_out[11585] & layer1_out[11586];
     layer2_out[9303] <= ~(layer1_out[239] ^ layer1_out[240]);
     layer2_out[9304] <= layer1_out[8418];
     layer2_out[9305] <= layer1_out[3508];
     layer2_out[9306] <= ~layer1_out[6714];
     layer2_out[9307] <= layer1_out[2635] & ~layer1_out[2634];
     layer2_out[9308] <= ~(layer1_out[5717] & layer1_out[5718]);
     layer2_out[9309] <= ~(layer1_out[8835] | layer1_out[8836]);
     layer2_out[9310] <= 1'b1;
     layer2_out[9311] <= ~(layer1_out[11561] & layer1_out[11562]);
     layer2_out[9312] <= layer1_out[6185];
     layer2_out[9313] <= ~layer1_out[11318];
     layer2_out[9314] <= ~(layer1_out[3020] & layer1_out[3021]);
     layer2_out[9315] <= ~layer1_out[10599];
     layer2_out[9316] <= ~layer1_out[5318] | layer1_out[5317];
     layer2_out[9317] <= ~layer1_out[717] | layer1_out[718];
     layer2_out[9318] <= layer1_out[10329] & ~layer1_out[10328];
     layer2_out[9319] <= ~(layer1_out[6058] & layer1_out[6059]);
     layer2_out[9320] <= layer1_out[4872] & layer1_out[4873];
     layer2_out[9321] <= ~layer1_out[3883];
     layer2_out[9322] <= ~layer1_out[10754] | layer1_out[10753];
     layer2_out[9323] <= layer1_out[11608] & ~layer1_out[11607];
     layer2_out[9324] <= ~(layer1_out[4513] | layer1_out[4514]);
     layer2_out[9325] <= ~layer1_out[5816];
     layer2_out[9326] <= layer1_out[6174] ^ layer1_out[6175];
     layer2_out[9327] <= ~layer1_out[6883] | layer1_out[6882];
     layer2_out[9328] <= ~(layer1_out[6685] | layer1_out[6686]);
     layer2_out[9329] <= layer1_out[9514] & layer1_out[9515];
     layer2_out[9330] <= ~layer1_out[2253] | layer1_out[2252];
     layer2_out[9331] <= ~layer1_out[3211];
     layer2_out[9332] <= ~(layer1_out[1807] & layer1_out[1808]);
     layer2_out[9333] <= ~layer1_out[1342] | layer1_out[1343];
     layer2_out[9334] <= ~(layer1_out[10654] ^ layer1_out[10655]);
     layer2_out[9335] <= layer1_out[5889] ^ layer1_out[5890];
     layer2_out[9336] <= layer1_out[11459] & layer1_out[11460];
     layer2_out[9337] <= ~layer1_out[2393];
     layer2_out[9338] <= ~(layer1_out[11766] ^ layer1_out[11767]);
     layer2_out[9339] <= ~(layer1_out[8581] & layer1_out[8582]);
     layer2_out[9340] <= ~layer1_out[3377];
     layer2_out[9341] <= ~layer1_out[2419];
     layer2_out[9342] <= ~(layer1_out[3068] ^ layer1_out[3069]);
     layer2_out[9343] <= layer1_out[3483] | layer1_out[3484];
     layer2_out[9344] <= layer1_out[9797] & ~layer1_out[9796];
     layer2_out[9345] <= layer1_out[6159] & ~layer1_out[6160];
     layer2_out[9346] <= ~(layer1_out[214] | layer1_out[215]);
     layer2_out[9347] <= layer1_out[8055] | layer1_out[8056];
     layer2_out[9348] <= layer1_out[2848] & ~layer1_out[2849];
     layer2_out[9349] <= layer1_out[1826] & layer1_out[1827];
     layer2_out[9350] <= ~layer1_out[6389];
     layer2_out[9351] <= ~layer1_out[11108];
     layer2_out[9352] <= ~layer1_out[9828];
     layer2_out[9353] <= ~layer1_out[10350] | layer1_out[10351];
     layer2_out[9354] <= ~layer1_out[7456];
     layer2_out[9355] <= layer1_out[10338] | layer1_out[10339];
     layer2_out[9356] <= layer1_out[868] ^ layer1_out[869];
     layer2_out[9357] <= layer1_out[11293] ^ layer1_out[11294];
     layer2_out[9358] <= ~layer1_out[8340];
     layer2_out[9359] <= layer1_out[4657] | layer1_out[4658];
     layer2_out[9360] <= ~layer1_out[5412] | layer1_out[5411];
     layer2_out[9361] <= ~(layer1_out[3422] & layer1_out[3423]);
     layer2_out[9362] <= ~layer1_out[4860];
     layer2_out[9363] <= layer1_out[6036] & ~layer1_out[6035];
     layer2_out[9364] <= ~(layer1_out[11762] & layer1_out[11763]);
     layer2_out[9365] <= layer1_out[7403];
     layer2_out[9366] <= layer1_out[5878] & ~layer1_out[5879];
     layer2_out[9367] <= layer1_out[558];
     layer2_out[9368] <= layer1_out[3962] & ~layer1_out[3961];
     layer2_out[9369] <= ~layer1_out[10553];
     layer2_out[9370] <= ~layer1_out[1950] | layer1_out[1951];
     layer2_out[9371] <= ~(layer1_out[9581] | layer1_out[9582]);
     layer2_out[9372] <= layer1_out[1212] | layer1_out[1213];
     layer2_out[9373] <= ~(layer1_out[4851] & layer1_out[4852]);
     layer2_out[9374] <= ~layer1_out[8044] | layer1_out[8045];
     layer2_out[9375] <= 1'b1;
     layer2_out[9376] <= layer1_out[2748];
     layer2_out[9377] <= ~(layer1_out[11581] ^ layer1_out[11582]);
     layer2_out[9378] <= layer1_out[2535] | layer1_out[2536];
     layer2_out[9379] <= layer1_out[8284];
     layer2_out[9380] <= layer1_out[6751];
     layer2_out[9381] <= ~(layer1_out[2099] ^ layer1_out[2100]);
     layer2_out[9382] <= ~layer1_out[6524];
     layer2_out[9383] <= layer1_out[6668];
     layer2_out[9384] <= ~(layer1_out[2126] ^ layer1_out[2127]);
     layer2_out[9385] <= layer1_out[8223] & layer1_out[8224];
     layer2_out[9386] <= ~layer1_out[6040];
     layer2_out[9387] <= ~(layer1_out[4844] ^ layer1_out[4845]);
     layer2_out[9388] <= ~(layer1_out[3912] ^ layer1_out[3913]);
     layer2_out[9389] <= ~layer1_out[3209] | layer1_out[3208];
     layer2_out[9390] <= layer1_out[5505] & ~layer1_out[5506];
     layer2_out[9391] <= ~(layer1_out[8222] | layer1_out[8223]);
     layer2_out[9392] <= layer1_out[4129];
     layer2_out[9393] <= ~layer1_out[10653];
     layer2_out[9394] <= ~(layer1_out[698] & layer1_out[699]);
     layer2_out[9395] <= layer1_out[8513] & ~layer1_out[8512];
     layer2_out[9396] <= layer1_out[1430] & ~layer1_out[1429];
     layer2_out[9397] <= layer1_out[2263];
     layer2_out[9398] <= layer1_out[2155];
     layer2_out[9399] <= layer1_out[3931];
     layer2_out[9400] <= layer1_out[2873];
     layer2_out[9401] <= layer1_out[550] | layer1_out[551];
     layer2_out[9402] <= layer1_out[7553];
     layer2_out[9403] <= ~layer1_out[460];
     layer2_out[9404] <= ~layer1_out[1571] | layer1_out[1572];
     layer2_out[9405] <= ~layer1_out[2394];
     layer2_out[9406] <= layer1_out[9572];
     layer2_out[9407] <= layer1_out[1058];
     layer2_out[9408] <= layer1_out[1768];
     layer2_out[9409] <= ~(layer1_out[7582] & layer1_out[7583]);
     layer2_out[9410] <= layer1_out[885] | layer1_out[886];
     layer2_out[9411] <= layer1_out[11267];
     layer2_out[9412] <= ~layer1_out[6827] | layer1_out[6826];
     layer2_out[9413] <= ~(layer1_out[2199] & layer1_out[2200]);
     layer2_out[9414] <= ~layer1_out[11854];
     layer2_out[9415] <= ~(layer1_out[11986] & layer1_out[11987]);
     layer2_out[9416] <= layer1_out[2386] & layer1_out[2387];
     layer2_out[9417] <= ~(layer1_out[8206] ^ layer1_out[8207]);
     layer2_out[9418] <= layer1_out[8084] | layer1_out[8085];
     layer2_out[9419] <= ~(layer1_out[9377] ^ layer1_out[9378]);
     layer2_out[9420] <= ~layer1_out[1907] | layer1_out[1906];
     layer2_out[9421] <= layer1_out[5486];
     layer2_out[9422] <= layer1_out[6376] ^ layer1_out[6377];
     layer2_out[9423] <= ~(layer1_out[3536] | layer1_out[3537]);
     layer2_out[9424] <= layer1_out[4120] | layer1_out[4121];
     layer2_out[9425] <= layer1_out[7414] & ~layer1_out[7413];
     layer2_out[9426] <= ~layer1_out[10649] | layer1_out[10650];
     layer2_out[9427] <= layer1_out[11108] & ~layer1_out[11107];
     layer2_out[9428] <= layer1_out[8543] & ~layer1_out[8544];
     layer2_out[9429] <= ~(layer1_out[2321] & layer1_out[2322]);
     layer2_out[9430] <= ~layer1_out[7907] | layer1_out[7908];
     layer2_out[9431] <= layer1_out[4112] ^ layer1_out[4113];
     layer2_out[9432] <= ~layer1_out[4701];
     layer2_out[9433] <= layer1_out[7073] ^ layer1_out[7074];
     layer2_out[9434] <= layer1_out[3926] & ~layer1_out[3927];
     layer2_out[9435] <= ~(layer1_out[5062] | layer1_out[5063]);
     layer2_out[9436] <= layer1_out[9585] & ~layer1_out[9586];
     layer2_out[9437] <= ~(layer1_out[5520] | layer1_out[5521]);
     layer2_out[9438] <= layer1_out[3414] | layer1_out[3415];
     layer2_out[9439] <= layer1_out[11251] & ~layer1_out[11252];
     layer2_out[9440] <= layer1_out[4030];
     layer2_out[9441] <= layer1_out[10851] & layer1_out[10852];
     layer2_out[9442] <= ~layer1_out[10088];
     layer2_out[9443] <= ~(layer1_out[2909] & layer1_out[2910]);
     layer2_out[9444] <= ~layer1_out[11718] | layer1_out[11719];
     layer2_out[9445] <= ~layer1_out[8507];
     layer2_out[9446] <= ~layer1_out[5775] | layer1_out[5774];
     layer2_out[9447] <= ~layer1_out[6439];
     layer2_out[9448] <= layer1_out[7885] ^ layer1_out[7886];
     layer2_out[9449] <= ~(layer1_out[3124] & layer1_out[3125]);
     layer2_out[9450] <= ~layer1_out[4542] | layer1_out[4541];
     layer2_out[9451] <= ~layer1_out[9037];
     layer2_out[9452] <= layer1_out[7532] ^ layer1_out[7533];
     layer2_out[9453] <= layer1_out[7752] & ~layer1_out[7753];
     layer2_out[9454] <= ~(layer1_out[7671] & layer1_out[7672]);
     layer2_out[9455] <= ~layer1_out[7959] | layer1_out[7958];
     layer2_out[9456] <= ~layer1_out[6404];
     layer2_out[9457] <= layer1_out[7972] & layer1_out[7973];
     layer2_out[9458] <= layer1_out[1798];
     layer2_out[9459] <= layer1_out[9847] ^ layer1_out[9848];
     layer2_out[9460] <= layer1_out[5737];
     layer2_out[9461] <= ~layer1_out[1656];
     layer2_out[9462] <= ~layer1_out[5867];
     layer2_out[9463] <= ~layer1_out[4896];
     layer2_out[9464] <= layer1_out[9387] & ~layer1_out[9386];
     layer2_out[9465] <= layer1_out[9123];
     layer2_out[9466] <= layer1_out[2888] & ~layer1_out[2889];
     layer2_out[9467] <= layer1_out[674];
     layer2_out[9468] <= layer1_out[4908] & layer1_out[4909];
     layer2_out[9469] <= layer1_out[6548] | layer1_out[6549];
     layer2_out[9470] <= ~(layer1_out[8325] ^ layer1_out[8326]);
     layer2_out[9471] <= ~layer1_out[568];
     layer2_out[9472] <= ~layer1_out[8389];
     layer2_out[9473] <= ~(layer1_out[3837] | layer1_out[3838]);
     layer2_out[9474] <= layer1_out[5868] ^ layer1_out[5869];
     layer2_out[9475] <= ~(layer1_out[5535] | layer1_out[5536]);
     layer2_out[9476] <= layer1_out[99] & ~layer1_out[98];
     layer2_out[9477] <= layer1_out[3048] ^ layer1_out[3049];
     layer2_out[9478] <= ~(layer1_out[11825] ^ layer1_out[11826]);
     layer2_out[9479] <= layer1_out[11329] ^ layer1_out[11330];
     layer2_out[9480] <= layer1_out[1178];
     layer2_out[9481] <= layer1_out[4447] & ~layer1_out[4446];
     layer2_out[9482] <= ~layer1_out[2120];
     layer2_out[9483] <= layer1_out[282] & ~layer1_out[281];
     layer2_out[9484] <= ~layer1_out[11455];
     layer2_out[9485] <= ~layer1_out[10032];
     layer2_out[9486] <= layer1_out[5033] & ~layer1_out[5034];
     layer2_out[9487] <= ~layer1_out[4839] | layer1_out[4838];
     layer2_out[9488] <= layer1_out[8642] & layer1_out[8643];
     layer2_out[9489] <= ~layer1_out[1236];
     layer2_out[9490] <= ~layer1_out[10905] | layer1_out[10906];
     layer2_out[9491] <= layer1_out[2147] | layer1_out[2148];
     layer2_out[9492] <= ~layer1_out[9472] | layer1_out[9471];
     layer2_out[9493] <= ~(layer1_out[10695] ^ layer1_out[10696]);
     layer2_out[9494] <= layer1_out[6870] ^ layer1_out[6871];
     layer2_out[9495] <= ~(layer1_out[8781] ^ layer1_out[8782]);
     layer2_out[9496] <= layer1_out[1497];
     layer2_out[9497] <= ~layer1_out[2904];
     layer2_out[9498] <= layer1_out[1555];
     layer2_out[9499] <= ~layer1_out[1019];
     layer2_out[9500] <= layer1_out[234] & ~layer1_out[233];
     layer2_out[9501] <= ~layer1_out[4802];
     layer2_out[9502] <= layer1_out[8966] & layer1_out[8967];
     layer2_out[9503] <= layer1_out[2354];
     layer2_out[9504] <= ~layer1_out[563];
     layer2_out[9505] <= layer1_out[6977] & ~layer1_out[6978];
     layer2_out[9506] <= ~layer1_out[8905];
     layer2_out[9507] <= layer1_out[10254] | layer1_out[10255];
     layer2_out[9508] <= layer1_out[10346] & ~layer1_out[10347];
     layer2_out[9509] <= ~(layer1_out[11632] & layer1_out[11633]);
     layer2_out[9510] <= layer1_out[5593];
     layer2_out[9511] <= ~(layer1_out[1769] | layer1_out[1770]);
     layer2_out[9512] <= layer1_out[9426];
     layer2_out[9513] <= layer1_out[4699] & ~layer1_out[4700];
     layer2_out[9514] <= layer1_out[7032];
     layer2_out[9515] <= ~layer1_out[6298] | layer1_out[6297];
     layer2_out[9516] <= ~layer1_out[19];
     layer2_out[9517] <= layer1_out[9930] & ~layer1_out[9929];
     layer2_out[9518] <= layer1_out[10713] & ~layer1_out[10712];
     layer2_out[9519] <= layer1_out[10162] | layer1_out[10163];
     layer2_out[9520] <= layer1_out[3897];
     layer2_out[9521] <= ~(layer1_out[7954] | layer1_out[7955]);
     layer2_out[9522] <= ~(layer1_out[7984] & layer1_out[7985]);
     layer2_out[9523] <= layer1_out[1126];
     layer2_out[9524] <= ~layer1_out[5432] | layer1_out[5433];
     layer2_out[9525] <= layer1_out[10676];
     layer2_out[9526] <= layer1_out[564] & ~layer1_out[563];
     layer2_out[9527] <= layer1_out[9247];
     layer2_out[9528] <= layer1_out[539] & ~layer1_out[540];
     layer2_out[9529] <= layer1_out[5084];
     layer2_out[9530] <= ~layer1_out[6550];
     layer2_out[9531] <= layer1_out[8828] & ~layer1_out[8829];
     layer2_out[9532] <= ~layer1_out[938] | layer1_out[937];
     layer2_out[9533] <= layer1_out[178];
     layer2_out[9534] <= ~layer1_out[11364];
     layer2_out[9535] <= ~layer1_out[10810];
     layer2_out[9536] <= layer1_out[9021] ^ layer1_out[9022];
     layer2_out[9537] <= layer1_out[8465] | layer1_out[8466];
     layer2_out[9538] <= ~layer1_out[1436] | layer1_out[1437];
     layer2_out[9539] <= ~layer1_out[7116];
     layer2_out[9540] <= layer1_out[594];
     layer2_out[9541] <= ~layer1_out[1625] | layer1_out[1624];
     layer2_out[9542] <= ~layer1_out[9820];
     layer2_out[9543] <= layer1_out[7251];
     layer2_out[9544] <= layer1_out[11040];
     layer2_out[9545] <= layer1_out[5168] & layer1_out[5169];
     layer2_out[9546] <= layer1_out[110] & layer1_out[111];
     layer2_out[9547] <= layer1_out[1847];
     layer2_out[9548] <= ~(layer1_out[10682] | layer1_out[10683]);
     layer2_out[9549] <= layer1_out[895];
     layer2_out[9550] <= layer1_out[5589] & ~layer1_out[5590];
     layer2_out[9551] <= layer1_out[4451];
     layer2_out[9552] <= layer1_out[1640] & ~layer1_out[1639];
     layer2_out[9553] <= layer1_out[10663] & ~layer1_out[10662];
     layer2_out[9554] <= ~layer1_out[5628] | layer1_out[5627];
     layer2_out[9555] <= layer1_out[7781] & ~layer1_out[7782];
     layer2_out[9556] <= ~layer1_out[9493];
     layer2_out[9557] <= layer1_out[10559] ^ layer1_out[10560];
     layer2_out[9558] <= layer1_out[5090] | layer1_out[5091];
     layer2_out[9559] <= layer1_out[6454] & ~layer1_out[6453];
     layer2_out[9560] <= layer1_out[3882] & ~layer1_out[3881];
     layer2_out[9561] <= ~(layer1_out[6910] ^ layer1_out[6911]);
     layer2_out[9562] <= layer1_out[482] ^ layer1_out[483];
     layer2_out[9563] <= layer1_out[8155] | layer1_out[8156];
     layer2_out[9564] <= layer1_out[3218] & layer1_out[3219];
     layer2_out[9565] <= layer1_out[9656];
     layer2_out[9566] <= ~layer1_out[4220] | layer1_out[4219];
     layer2_out[9567] <= ~layer1_out[11533];
     layer2_out[9568] <= layer1_out[4613] & ~layer1_out[4612];
     layer2_out[9569] <= ~layer1_out[10519];
     layer2_out[9570] <= ~layer1_out[9935] | layer1_out[9934];
     layer2_out[9571] <= ~layer1_out[6335] | layer1_out[6334];
     layer2_out[9572] <= layer1_out[5187];
     layer2_out[9573] <= ~(layer1_out[8672] ^ layer1_out[8673]);
     layer2_out[9574] <= layer1_out[1508] ^ layer1_out[1509];
     layer2_out[9575] <= ~(layer1_out[11370] ^ layer1_out[11371]);
     layer2_out[9576] <= ~(layer1_out[10429] & layer1_out[10430]);
     layer2_out[9577] <= layer1_out[1463] & ~layer1_out[1464];
     layer2_out[9578] <= layer1_out[3498];
     layer2_out[9579] <= layer1_out[7694] & ~layer1_out[7695];
     layer2_out[9580] <= ~layer1_out[7148] | layer1_out[7149];
     layer2_out[9581] <= layer1_out[702] | layer1_out[703];
     layer2_out[9582] <= ~(layer1_out[435] & layer1_out[436]);
     layer2_out[9583] <= ~layer1_out[2953];
     layer2_out[9584] <= ~layer1_out[2641];
     layer2_out[9585] <= ~(layer1_out[1501] & layer1_out[1502]);
     layer2_out[9586] <= ~layer1_out[2441] | layer1_out[2442];
     layer2_out[9587] <= ~layer1_out[9749];
     layer2_out[9588] <= ~layer1_out[1991];
     layer2_out[9589] <= ~layer1_out[1751] | layer1_out[1750];
     layer2_out[9590] <= layer1_out[1182] & ~layer1_out[1181];
     layer2_out[9591] <= ~(layer1_out[10404] & layer1_out[10405]);
     layer2_out[9592] <= layer1_out[3250] | layer1_out[3251];
     layer2_out[9593] <= ~(layer1_out[7326] & layer1_out[7327]);
     layer2_out[9594] <= ~layer1_out[7536] | layer1_out[7535];
     layer2_out[9595] <= ~layer1_out[11863] | layer1_out[11862];
     layer2_out[9596] <= ~layer1_out[2054] | layer1_out[2053];
     layer2_out[9597] <= layer1_out[8792];
     layer2_out[9598] <= layer1_out[11356] & layer1_out[11357];
     layer2_out[9599] <= ~(layer1_out[1045] ^ layer1_out[1046]);
     layer2_out[9600] <= layer1_out[8409];
     layer2_out[9601] <= ~layer1_out[3635];
     layer2_out[9602] <= ~layer1_out[951];
     layer2_out[9603] <= ~(layer1_out[1947] ^ layer1_out[1948]);
     layer2_out[9604] <= layer1_out[8772] & layer1_out[8773];
     layer2_out[9605] <= ~(layer1_out[5544] | layer1_out[5545]);
     layer2_out[9606] <= 1'b0;
     layer2_out[9607] <= layer1_out[3467] & layer1_out[3468];
     layer2_out[9608] <= layer1_out[5282];
     layer2_out[9609] <= layer1_out[6598] & ~layer1_out[6597];
     layer2_out[9610] <= layer1_out[4824] ^ layer1_out[4825];
     layer2_out[9611] <= ~(layer1_out[5877] ^ layer1_out[5878]);
     layer2_out[9612] <= ~(layer1_out[1147] & layer1_out[1148]);
     layer2_out[9613] <= layer1_out[9507] & layer1_out[9508];
     layer2_out[9614] <= layer1_out[5833];
     layer2_out[9615] <= ~layer1_out[1262] | layer1_out[1263];
     layer2_out[9616] <= ~layer1_out[4690];
     layer2_out[9617] <= ~layer1_out[6598] | layer1_out[6599];
     layer2_out[9618] <= layer1_out[8056] | layer1_out[8057];
     layer2_out[9619] <= ~layer1_out[7396];
     layer2_out[9620] <= layer1_out[9588];
     layer2_out[9621] <= layer1_out[11339];
     layer2_out[9622] <= layer1_out[6071] ^ layer1_out[6072];
     layer2_out[9623] <= ~layer1_out[9746] | layer1_out[9747];
     layer2_out[9624] <= layer1_out[5622] & layer1_out[5623];
     layer2_out[9625] <= layer1_out[5267];
     layer2_out[9626] <= layer1_out[3137] ^ layer1_out[3138];
     layer2_out[9627] <= layer1_out[1641];
     layer2_out[9628] <= layer1_out[7057];
     layer2_out[9629] <= ~layer1_out[8316] | layer1_out[8317];
     layer2_out[9630] <= layer1_out[6384] | layer1_out[6385];
     layer2_out[9631] <= layer1_out[3312];
     layer2_out[9632] <= layer1_out[11734];
     layer2_out[9633] <= layer1_out[4368] | layer1_out[4369];
     layer2_out[9634] <= ~layer1_out[9961];
     layer2_out[9635] <= ~(layer1_out[11156] & layer1_out[11157]);
     layer2_out[9636] <= layer1_out[4624] & layer1_out[4625];
     layer2_out[9637] <= ~layer1_out[5732] | layer1_out[5731];
     layer2_out[9638] <= layer1_out[11895];
     layer2_out[9639] <= ~(layer1_out[2060] | layer1_out[2061]);
     layer2_out[9640] <= layer1_out[9022];
     layer2_out[9641] <= ~(layer1_out[7630] ^ layer1_out[7631]);
     layer2_out[9642] <= ~layer1_out[5926] | layer1_out[5925];
     layer2_out[9643] <= ~(layer1_out[10951] ^ layer1_out[10952]);
     layer2_out[9644] <= layer1_out[5452];
     layer2_out[9645] <= layer1_out[11155];
     layer2_out[9646] <= ~layer1_out[5579];
     layer2_out[9647] <= layer1_out[10609];
     layer2_out[9648] <= layer1_out[657];
     layer2_out[9649] <= layer1_out[6690];
     layer2_out[9650] <= layer1_out[11740] & ~layer1_out[11739];
     layer2_out[9651] <= layer1_out[11333] & ~layer1_out[11332];
     layer2_out[9652] <= ~layer1_out[8394];
     layer2_out[9653] <= ~(layer1_out[4209] ^ layer1_out[4210]);
     layer2_out[9654] <= ~(layer1_out[3678] & layer1_out[3679]);
     layer2_out[9655] <= ~layer1_out[1554] | layer1_out[1555];
     layer2_out[9656] <= ~(layer1_out[10414] | layer1_out[10415]);
     layer2_out[9657] <= layer1_out[6194] & ~layer1_out[6195];
     layer2_out[9658] <= layer1_out[7861] & layer1_out[7862];
     layer2_out[9659] <= ~(layer1_out[2250] | layer1_out[2251]);
     layer2_out[9660] <= layer1_out[6679] | layer1_out[6680];
     layer2_out[9661] <= layer1_out[5095] & layer1_out[5096];
     layer2_out[9662] <= ~layer1_out[893];
     layer2_out[9663] <= layer1_out[4306];
     layer2_out[9664] <= layer1_out[9922];
     layer2_out[9665] <= layer1_out[10633] & ~layer1_out[10634];
     layer2_out[9666] <= ~layer1_out[11873] | layer1_out[11872];
     layer2_out[9667] <= layer1_out[938] ^ layer1_out[939];
     layer2_out[9668] <= ~layer1_out[1961];
     layer2_out[9669] <= ~layer1_out[1475];
     layer2_out[9670] <= layer1_out[4168] & ~layer1_out[4169];
     layer2_out[9671] <= ~layer1_out[9932] | layer1_out[9931];
     layer2_out[9672] <= layer1_out[11893] & ~layer1_out[11892];
     layer2_out[9673] <= layer1_out[11932];
     layer2_out[9674] <= layer1_out[2395];
     layer2_out[9675] <= ~layer1_out[3244];
     layer2_out[9676] <= layer1_out[8190] ^ layer1_out[8191];
     layer2_out[9677] <= layer1_out[2431] & ~layer1_out[2432];
     layer2_out[9678] <= layer1_out[4268] & ~layer1_out[4267];
     layer2_out[9679] <= layer1_out[4381] & ~layer1_out[4380];
     layer2_out[9680] <= layer1_out[8547];
     layer2_out[9681] <= ~layer1_out[5482] | layer1_out[5481];
     layer2_out[9682] <= layer1_out[7642] & ~layer1_out[7641];
     layer2_out[9683] <= ~(layer1_out[1473] | layer1_out[1474]);
     layer2_out[9684] <= ~(layer1_out[9578] | layer1_out[9579]);
     layer2_out[9685] <= layer1_out[9247];
     layer2_out[9686] <= layer1_out[4911];
     layer2_out[9687] <= layer1_out[4699];
     layer2_out[9688] <= ~layer1_out[6300];
     layer2_out[9689] <= layer1_out[5050] & layer1_out[5051];
     layer2_out[9690] <= ~layer1_out[9605] | layer1_out[9606];
     layer2_out[9691] <= layer1_out[2216] & ~layer1_out[2215];
     layer2_out[9692] <= layer1_out[1543] & layer1_out[1544];
     layer2_out[9693] <= ~(layer1_out[5301] | layer1_out[5302]);
     layer2_out[9694] <= ~layer1_out[2536];
     layer2_out[9695] <= layer1_out[6281] & ~layer1_out[6282];
     layer2_out[9696] <= ~(layer1_out[638] & layer1_out[639]);
     layer2_out[9697] <= 1'b1;
     layer2_out[9698] <= layer1_out[8657];
     layer2_out[9699] <= layer1_out[8601];
     layer2_out[9700] <= ~layer1_out[11646];
     layer2_out[9701] <= ~layer1_out[6487];
     layer2_out[9702] <= ~layer1_out[10657];
     layer2_out[9703] <= ~layer1_out[7768];
     layer2_out[9704] <= layer1_out[7308];
     layer2_out[9705] <= ~layer1_out[6241];
     layer2_out[9706] <= layer1_out[3141] & layer1_out[3142];
     layer2_out[9707] <= layer1_out[6139];
     layer2_out[9708] <= layer1_out[8821];
     layer2_out[9709] <= layer1_out[4675] & layer1_out[4676];
     layer2_out[9710] <= layer1_out[3039];
     layer2_out[9711] <= layer1_out[8065] & layer1_out[8066];
     layer2_out[9712] <= layer1_out[377] & layer1_out[378];
     layer2_out[9713] <= layer1_out[399];
     layer2_out[9714] <= layer1_out[10728];
     layer2_out[9715] <= ~layer1_out[9283] | layer1_out[9282];
     layer2_out[9716] <= ~layer1_out[474];
     layer2_out[9717] <= ~layer1_out[3701] | layer1_out[3700];
     layer2_out[9718] <= layer1_out[7368] & ~layer1_out[7367];
     layer2_out[9719] <= ~layer1_out[3748] | layer1_out[3749];
     layer2_out[9720] <= layer1_out[642];
     layer2_out[9721] <= layer1_out[8752] ^ layer1_out[8753];
     layer2_out[9722] <= layer1_out[4279] | layer1_out[4280];
     layer2_out[9723] <= ~layer1_out[7046];
     layer2_out[9724] <= ~(layer1_out[9011] | layer1_out[9012]);
     layer2_out[9725] <= layer1_out[4476];
     layer2_out[9726] <= layer1_out[11480] & ~layer1_out[11479];
     layer2_out[9727] <= ~layer1_out[5016] | layer1_out[5015];
     layer2_out[9728] <= ~layer1_out[2382];
     layer2_out[9729] <= layer1_out[8468] & ~layer1_out[8469];
     layer2_out[9730] <= layer1_out[8092] & ~layer1_out[8091];
     layer2_out[9731] <= ~(layer1_out[5934] & layer1_out[5935]);
     layer2_out[9732] <= ~layer1_out[6626] | layer1_out[6627];
     layer2_out[9733] <= layer1_out[7969] | layer1_out[7970];
     layer2_out[9734] <= layer1_out[1718] ^ layer1_out[1719];
     layer2_out[9735] <= ~layer1_out[8598];
     layer2_out[9736] <= ~layer1_out[4708];
     layer2_out[9737] <= layer1_out[569] & ~layer1_out[570];
     layer2_out[9738] <= layer1_out[9302];
     layer2_out[9739] <= ~(layer1_out[571] | layer1_out[572]);
     layer2_out[9740] <= layer1_out[8144] & ~layer1_out[8143];
     layer2_out[9741] <= layer1_out[1507];
     layer2_out[9742] <= layer1_out[615] | layer1_out[616];
     layer2_out[9743] <= layer1_out[3465] ^ layer1_out[3466];
     layer2_out[9744] <= ~layer1_out[2937] | layer1_out[2936];
     layer2_out[9745] <= ~layer1_out[3627] | layer1_out[3628];
     layer2_out[9746] <= layer1_out[9919];
     layer2_out[9747] <= layer1_out[11031];
     layer2_out[9748] <= ~layer1_out[10150];
     layer2_out[9749] <= layer1_out[3483] & ~layer1_out[3482];
     layer2_out[9750] <= ~layer1_out[8014];
     layer2_out[9751] <= layer1_out[7529] & ~layer1_out[7530];
     layer2_out[9752] <= layer1_out[7883];
     layer2_out[9753] <= ~(layer1_out[3598] | layer1_out[3599]);
     layer2_out[9754] <= layer1_out[3800] & layer1_out[3801];
     layer2_out[9755] <= ~layer1_out[6311] | layer1_out[6310];
     layer2_out[9756] <= layer1_out[1000] & ~layer1_out[999];
     layer2_out[9757] <= ~layer1_out[575];
     layer2_out[9758] <= layer1_out[9103];
     layer2_out[9759] <= layer1_out[8625] & layer1_out[8626];
     layer2_out[9760] <= layer1_out[5208];
     layer2_out[9761] <= layer1_out[5676] & ~layer1_out[5677];
     layer2_out[9762] <= ~(layer1_out[3679] | layer1_out[3680]);
     layer2_out[9763] <= layer1_out[6821] & layer1_out[6822];
     layer2_out[9764] <= layer1_out[9391] & ~layer1_out[9392];
     layer2_out[9765] <= ~layer1_out[7605];
     layer2_out[9766] <= layer1_out[9018] & ~layer1_out[9019];
     layer2_out[9767] <= ~(layer1_out[7929] ^ layer1_out[7930]);
     layer2_out[9768] <= layer1_out[4591] & layer1_out[4592];
     layer2_out[9769] <= layer1_out[3457] & ~layer1_out[3458];
     layer2_out[9770] <= layer1_out[3332];
     layer2_out[9771] <= ~(layer1_out[4423] & layer1_out[4424]);
     layer2_out[9772] <= layer1_out[183] & ~layer1_out[182];
     layer2_out[9773] <= ~layer1_out[6931] | layer1_out[6932];
     layer2_out[9774] <= layer1_out[10133];
     layer2_out[9775] <= layer1_out[9362] & layer1_out[9363];
     layer2_out[9776] <= layer1_out[6921];
     layer2_out[9777] <= ~(layer1_out[6799] & layer1_out[6800]);
     layer2_out[9778] <= ~layer1_out[4957] | layer1_out[4958];
     layer2_out[9779] <= layer1_out[675];
     layer2_out[9780] <= ~layer1_out[11392];
     layer2_out[9781] <= layer1_out[9802] & layer1_out[9803];
     layer2_out[9782] <= layer1_out[7804] & layer1_out[7805];
     layer2_out[9783] <= ~layer1_out[9029];
     layer2_out[9784] <= layer1_out[2320] & ~layer1_out[2319];
     layer2_out[9785] <= layer1_out[3555] ^ layer1_out[3556];
     layer2_out[9786] <= ~(layer1_out[8039] ^ layer1_out[8040]);
     layer2_out[9787] <= layer1_out[5541] & layer1_out[5542];
     layer2_out[9788] <= ~layer1_out[9826];
     layer2_out[9789] <= layer1_out[10762];
     layer2_out[9790] <= ~(layer1_out[7556] ^ layer1_out[7557]);
     layer2_out[9791] <= ~layer1_out[11631];
     layer2_out[9792] <= layer1_out[7610];
     layer2_out[9793] <= layer1_out[2314] & layer1_out[2315];
     layer2_out[9794] <= ~layer1_out[5610] | layer1_out[5611];
     layer2_out[9795] <= ~(layer1_out[5359] ^ layer1_out[5360]);
     layer2_out[9796] <= ~(layer1_out[11695] | layer1_out[11696]);
     layer2_out[9797] <= ~layer1_out[2441];
     layer2_out[9798] <= layer1_out[3673] | layer1_out[3674];
     layer2_out[9799] <= layer1_out[5928] & ~layer1_out[5927];
     layer2_out[9800] <= layer1_out[11054] & ~layer1_out[11055];
     layer2_out[9801] <= layer1_out[2870] & ~layer1_out[2869];
     layer2_out[9802] <= layer1_out[1530] | layer1_out[1531];
     layer2_out[9803] <= ~(layer1_out[3036] | layer1_out[3037]);
     layer2_out[9804] <= ~(layer1_out[555] ^ layer1_out[556]);
     layer2_out[9805] <= layer1_out[8311] & ~layer1_out[8310];
     layer2_out[9806] <= layer1_out[1933] | layer1_out[1934];
     layer2_out[9807] <= layer1_out[4813] | layer1_out[4814];
     layer2_out[9808] <= ~layer1_out[11023];
     layer2_out[9809] <= layer1_out[5821];
     layer2_out[9810] <= layer1_out[1820];
     layer2_out[9811] <= layer1_out[11845];
     layer2_out[9812] <= layer1_out[3696] & ~layer1_out[3697];
     layer2_out[9813] <= layer1_out[11591];
     layer2_out[9814] <= ~(layer1_out[6972] ^ layer1_out[6973]);
     layer2_out[9815] <= ~layer1_out[1381];
     layer2_out[9816] <= ~(layer1_out[8687] | layer1_out[8688]);
     layer2_out[9817] <= ~layer1_out[6186];
     layer2_out[9818] <= ~(layer1_out[5956] & layer1_out[5957]);
     layer2_out[9819] <= layer1_out[10872];
     layer2_out[9820] <= layer1_out[4148];
     layer2_out[9821] <= 1'b1;
     layer2_out[9822] <= ~layer1_out[11814];
     layer2_out[9823] <= ~(layer1_out[9281] ^ layer1_out[9282]);
     layer2_out[9824] <= ~layer1_out[4608] | layer1_out[4609];
     layer2_out[9825] <= ~(layer1_out[9448] & layer1_out[9449]);
     layer2_out[9826] <= ~layer1_out[6560];
     layer2_out[9827] <= layer1_out[8273] & layer1_out[8274];
     layer2_out[9828] <= layer1_out[5911];
     layer2_out[9829] <= layer1_out[3293] | layer1_out[3294];
     layer2_out[9830] <= layer1_out[10082] | layer1_out[10083];
     layer2_out[9831] <= ~layer1_out[10402] | layer1_out[10401];
     layer2_out[9832] <= ~(layer1_out[8234] & layer1_out[8235]);
     layer2_out[9833] <= layer1_out[9166];
     layer2_out[9834] <= ~layer1_out[3729];
     layer2_out[9835] <= ~layer1_out[2448];
     layer2_out[9836] <= layer1_out[4614] & ~layer1_out[4613];
     layer2_out[9837] <= layer1_out[7416];
     layer2_out[9838] <= layer1_out[5897] & layer1_out[5898];
     layer2_out[9839] <= layer1_out[11657] | layer1_out[11658];
     layer2_out[9840] <= layer1_out[7423];
     layer2_out[9841] <= ~layer1_out[908];
     layer2_out[9842] <= ~layer1_out[8242];
     layer2_out[9843] <= ~(layer1_out[5494] | layer1_out[5495]);
     layer2_out[9844] <= ~(layer1_out[10368] & layer1_out[10369]);
     layer2_out[9845] <= ~(layer1_out[11330] ^ layer1_out[11331]);
     layer2_out[9846] <= layer1_out[11941];
     layer2_out[9847] <= layer1_out[1752] & layer1_out[1753];
     layer2_out[9848] <= ~(layer1_out[11481] | layer1_out[11482]);
     layer2_out[9849] <= ~layer1_out[11263];
     layer2_out[9850] <= layer1_out[7740];
     layer2_out[9851] <= layer1_out[5859] & layer1_out[5860];
     layer2_out[9852] <= ~layer1_out[3704];
     layer2_out[9853] <= layer1_out[2581] ^ layer1_out[2582];
     layer2_out[9854] <= layer1_out[10645] & ~layer1_out[10644];
     layer2_out[9855] <= layer1_out[9580];
     layer2_out[9856] <= layer1_out[3184] & ~layer1_out[3183];
     layer2_out[9857] <= layer1_out[7041] & layer1_out[7042];
     layer2_out[9858] <= ~layer1_out[243];
     layer2_out[9859] <= ~layer1_out[1186] | layer1_out[1185];
     layer2_out[9860] <= ~layer1_out[10395] | layer1_out[10394];
     layer2_out[9861] <= ~(layer1_out[1819] ^ layer1_out[1820]);
     layer2_out[9862] <= layer1_out[10719];
     layer2_out[9863] <= ~layer1_out[10691];
     layer2_out[9864] <= ~layer1_out[8452] | layer1_out[8453];
     layer2_out[9865] <= ~(layer1_out[2801] ^ layer1_out[2802]);
     layer2_out[9866] <= ~layer1_out[3880] | layer1_out[3881];
     layer2_out[9867] <= layer1_out[8391] ^ layer1_out[8392];
     layer2_out[9868] <= ~layer1_out[2417];
     layer2_out[9869] <= layer1_out[10016] & ~layer1_out[10015];
     layer2_out[9870] <= ~layer1_out[5173];
     layer2_out[9871] <= ~layer1_out[4245];
     layer2_out[9872] <= layer1_out[10005] | layer1_out[10006];
     layer2_out[9873] <= layer1_out[6707] & ~layer1_out[6708];
     layer2_out[9874] <= ~layer1_out[4429] | layer1_out[4430];
     layer2_out[9875] <= layer1_out[11176];
     layer2_out[9876] <= layer1_out[5726] ^ layer1_out[5727];
     layer2_out[9877] <= layer1_out[614];
     layer2_out[9878] <= layer1_out[2006] & ~layer1_out[2005];
     layer2_out[9879] <= ~layer1_out[2697] | layer1_out[2696];
     layer2_out[9880] <= ~layer1_out[4412] | layer1_out[4411];
     layer2_out[9881] <= layer1_out[8906];
     layer2_out[9882] <= layer1_out[8826];
     layer2_out[9883] <= ~(layer1_out[11615] | layer1_out[11616]);
     layer2_out[9884] <= layer1_out[4337] | layer1_out[4338];
     layer2_out[9885] <= layer1_out[2488];
     layer2_out[9886] <= layer1_out[467] & ~layer1_out[466];
     layer2_out[9887] <= ~(layer1_out[5980] & layer1_out[5981]);
     layer2_out[9888] <= ~layer1_out[731];
     layer2_out[9889] <= ~layer1_out[1265];
     layer2_out[9890] <= ~layer1_out[2647] | layer1_out[2648];
     layer2_out[9891] <= layer1_out[10629] | layer1_out[10630];
     layer2_out[9892] <= layer1_out[4678] ^ layer1_out[4679];
     layer2_out[9893] <= ~layer1_out[11949];
     layer2_out[9894] <= ~(layer1_out[2807] & layer1_out[2808]);
     layer2_out[9895] <= layer1_out[8993];
     layer2_out[9896] <= layer1_out[2572] | layer1_out[2573];
     layer2_out[9897] <= ~(layer1_out[3812] | layer1_out[3813]);
     layer2_out[9898] <= layer1_out[1664] & ~layer1_out[1663];
     layer2_out[9899] <= layer1_out[6426] & layer1_out[6427];
     layer2_out[9900] <= layer1_out[2136] & ~layer1_out[2135];
     layer2_out[9901] <= layer1_out[11974] & ~layer1_out[11973];
     layer2_out[9902] <= ~layer1_out[4661] | layer1_out[4662];
     layer2_out[9903] <= ~layer1_out[3376];
     layer2_out[9904] <= ~(layer1_out[874] | layer1_out[875]);
     layer2_out[9905] <= layer1_out[9197] & ~layer1_out[9196];
     layer2_out[9906] <= layer1_out[5233];
     layer2_out[9907] <= layer1_out[12];
     layer2_out[9908] <= ~layer1_out[6660];
     layer2_out[9909] <= ~(layer1_out[5532] ^ layer1_out[5533]);
     layer2_out[9910] <= layer1_out[10035] | layer1_out[10036];
     layer2_out[9911] <= ~layer1_out[9131];
     layer2_out[9912] <= layer1_out[873];
     layer2_out[9913] <= ~(layer1_out[269] ^ layer1_out[270]);
     layer2_out[9914] <= layer1_out[2057] & ~layer1_out[2058];
     layer2_out[9915] <= ~(layer1_out[4229] | layer1_out[4230]);
     layer2_out[9916] <= layer1_out[6571] ^ layer1_out[6572];
     layer2_out[9917] <= ~(layer1_out[9813] & layer1_out[9814]);
     layer2_out[9918] <= ~layer1_out[2621] | layer1_out[2620];
     layer2_out[9919] <= ~layer1_out[5769];
     layer2_out[9920] <= ~layer1_out[9543];
     layer2_out[9921] <= layer1_out[11806] & layer1_out[11807];
     layer2_out[9922] <= ~(layer1_out[8305] ^ layer1_out[8306]);
     layer2_out[9923] <= ~layer1_out[510];
     layer2_out[9924] <= layer1_out[6212] & ~layer1_out[6211];
     layer2_out[9925] <= layer1_out[3258] & ~layer1_out[3257];
     layer2_out[9926] <= layer1_out[2260];
     layer2_out[9927] <= ~layer1_out[6947];
     layer2_out[9928] <= layer1_out[2737] & ~layer1_out[2738];
     layer2_out[9929] <= layer1_out[6168] & ~layer1_out[6169];
     layer2_out[9930] <= ~layer1_out[1007];
     layer2_out[9931] <= layer1_out[9485];
     layer2_out[9932] <= layer1_out[3150] | layer1_out[3151];
     layer2_out[9933] <= ~layer1_out[10573];
     layer2_out[9934] <= layer1_out[10455] & ~layer1_out[10454];
     layer2_out[9935] <= layer1_out[11977] & layer1_out[11978];
     layer2_out[9936] <= ~layer1_out[2383] | layer1_out[2382];
     layer2_out[9937] <= ~layer1_out[6315] | layer1_out[6316];
     layer2_out[9938] <= ~(layer1_out[7923] | layer1_out[7924]);
     layer2_out[9939] <= layer1_out[11613];
     layer2_out[9940] <= ~layer1_out[7953];
     layer2_out[9941] <= ~layer1_out[4501];
     layer2_out[9942] <= layer1_out[8982] & ~layer1_out[8981];
     layer2_out[9943] <= layer1_out[5528] & layer1_out[5529];
     layer2_out[9944] <= ~layer1_out[10414] | layer1_out[10413];
     layer2_out[9945] <= ~(layer1_out[9874] & layer1_out[9875]);
     layer2_out[9946] <= ~layer1_out[9628];
     layer2_out[9947] <= layer1_out[5605];
     layer2_out[9948] <= ~layer1_out[11410];
     layer2_out[9949] <= layer1_out[982] | layer1_out[983];
     layer2_out[9950] <= layer1_out[1071] | layer1_out[1072];
     layer2_out[9951] <= ~layer1_out[8046] | layer1_out[8045];
     layer2_out[9952] <= ~layer1_out[10253] | layer1_out[10254];
     layer2_out[9953] <= layer1_out[968] | layer1_out[969];
     layer2_out[9954] <= layer1_out[5242];
     layer2_out[9955] <= layer1_out[9095];
     layer2_out[9956] <= 1'b1;
     layer2_out[9957] <= ~layer1_out[6877];
     layer2_out[9958] <= ~layer1_out[2979];
     layer2_out[9959] <= layer1_out[7751] & ~layer1_out[7752];
     layer2_out[9960] <= ~layer1_out[8665] | layer1_out[8666];
     layer2_out[9961] <= ~(layer1_out[1827] & layer1_out[1828]);
     layer2_out[9962] <= layer1_out[5392];
     layer2_out[9963] <= layer1_out[1897];
     layer2_out[9964] <= ~(layer1_out[4473] & layer1_out[4474]);
     layer2_out[9965] <= ~(layer1_out[939] & layer1_out[940]);
     layer2_out[9966] <= ~layer1_out[3765];
     layer2_out[9967] <= layer1_out[11369];
     layer2_out[9968] <= ~layer1_out[4345];
     layer2_out[9969] <= layer1_out[1600];
     layer2_out[9970] <= ~layer1_out[10149];
     layer2_out[9971] <= ~(layer1_out[8939] | layer1_out[8940]);
     layer2_out[9972] <= layer1_out[2275];
     layer2_out[9973] <= layer1_out[6413] ^ layer1_out[6414];
     layer2_out[9974] <= ~layer1_out[5920];
     layer2_out[9975] <= ~(layer1_out[7518] & layer1_out[7519]);
     layer2_out[9976] <= layer1_out[9849];
     layer2_out[9977] <= ~layer1_out[6872];
     layer2_out[9978] <= ~(layer1_out[11915] & layer1_out[11916]);
     layer2_out[9979] <= ~(layer1_out[9538] ^ layer1_out[9539]);
     layer2_out[9980] <= layer1_out[7394] | layer1_out[7395];
     layer2_out[9981] <= layer1_out[7058];
     layer2_out[9982] <= ~(layer1_out[4776] ^ layer1_out[4777]);
     layer2_out[9983] <= ~(layer1_out[8850] & layer1_out[8851]);
     layer2_out[9984] <= ~layer1_out[8539];
     layer2_out[9985] <= ~layer1_out[7324];
     layer2_out[9986] <= ~layer1_out[5284];
     layer2_out[9987] <= ~(layer1_out[1724] & layer1_out[1725]);
     layer2_out[9988] <= ~(layer1_out[4140] & layer1_out[4141]);
     layer2_out[9989] <= ~(layer1_out[2265] | layer1_out[2266]);
     layer2_out[9990] <= layer1_out[9815] & ~layer1_out[9814];
     layer2_out[9991] <= ~(layer1_out[11640] & layer1_out[11641]);
     layer2_out[9992] <= layer1_out[9689];
     layer2_out[9993] <= ~layer1_out[5902];
     layer2_out[9994] <= layer1_out[11755];
     layer2_out[9995] <= layer1_out[1929] ^ layer1_out[1930];
     layer2_out[9996] <= ~(layer1_out[119] ^ layer1_out[120]);
     layer2_out[9997] <= ~(layer1_out[749] & layer1_out[750]);
     layer2_out[9998] <= layer1_out[6251] & layer1_out[6252];
     layer2_out[9999] <= ~layer1_out[7213] | layer1_out[7214];
     layer2_out[10000] <= ~(layer1_out[33] & layer1_out[34]);
     layer2_out[10001] <= ~layer1_out[2604];
     layer2_out[10002] <= ~(layer1_out[6225] ^ layer1_out[6226]);
     layer2_out[10003] <= layer1_out[4652] & ~layer1_out[4651];
     layer2_out[10004] <= ~(layer1_out[5088] | layer1_out[5089]);
     layer2_out[10005] <= layer1_out[2561];
     layer2_out[10006] <= ~layer1_out[3632];
     layer2_out[10007] <= ~layer1_out[1482];
     layer2_out[10008] <= ~layer1_out[8333] | layer1_out[8334];
     layer2_out[10009] <= layer1_out[7745] & ~layer1_out[7746];
     layer2_out[10010] <= ~layer1_out[6193];
     layer2_out[10011] <= ~(layer1_out[4530] & layer1_out[4531]);
     layer2_out[10012] <= layer1_out[10594];
     layer2_out[10013] <= layer1_out[10347] | layer1_out[10348];
     layer2_out[10014] <= ~layer1_out[3495] | layer1_out[3494];
     layer2_out[10015] <= ~layer1_out[3422];
     layer2_out[10016] <= ~(layer1_out[3714] | layer1_out[3715]);
     layer2_out[10017] <= ~(layer1_out[1141] & layer1_out[1142]);
     layer2_out[10018] <= ~(layer1_out[11848] | layer1_out[11849]);
     layer2_out[10019] <= layer1_out[11627] & ~layer1_out[11628];
     layer2_out[10020] <= layer1_out[6556] & layer1_out[6557];
     layer2_out[10021] <= layer1_out[4863] ^ layer1_out[4864];
     layer2_out[10022] <= ~layer1_out[9943] | layer1_out[9942];
     layer2_out[10023] <= layer1_out[8922] | layer1_out[8923];
     layer2_out[10024] <= layer1_out[4183] & ~layer1_out[4182];
     layer2_out[10025] <= ~layer1_out[11181];
     layer2_out[10026] <= ~layer1_out[4310];
     layer2_out[10027] <= 1'b0;
     layer2_out[10028] <= ~(layer1_out[3725] & layer1_out[3726]);
     layer2_out[10029] <= layer1_out[8967] ^ layer1_out[8968];
     layer2_out[10030] <= layer1_out[645] & layer1_out[646];
     layer2_out[10031] <= layer1_out[456] | layer1_out[457];
     layer2_out[10032] <= ~layer1_out[1977] | layer1_out[1976];
     layer2_out[10033] <= layer1_out[8846];
     layer2_out[10034] <= layer1_out[7791];
     layer2_out[10035] <= layer1_out[6762] & ~layer1_out[6763];
     layer2_out[10036] <= layer1_out[910] & layer1_out[911];
     layer2_out[10037] <= ~layer1_out[10385];
     layer2_out[10038] <= layer1_out[11509] & ~layer1_out[11508];
     layer2_out[10039] <= layer1_out[7227] & ~layer1_out[7226];
     layer2_out[10040] <= layer1_out[3639] | layer1_out[3640];
     layer2_out[10041] <= ~layer1_out[636];
     layer2_out[10042] <= layer1_out[10732] & ~layer1_out[10731];
     layer2_out[10043] <= ~(layer1_out[2340] | layer1_out[2341]);
     layer2_out[10044] <= ~layer1_out[9142];
     layer2_out[10045] <= ~layer1_out[7346];
     layer2_out[10046] <= layer1_out[2477] & ~layer1_out[2478];
     layer2_out[10047] <= ~layer1_out[964] | layer1_out[963];
     layer2_out[10048] <= layer1_out[3642];
     layer2_out[10049] <= ~layer1_out[2821];
     layer2_out[10050] <= layer1_out[4429] & ~layer1_out[4428];
     layer2_out[10051] <= 1'b1;
     layer2_out[10052] <= layer1_out[8624] & layer1_out[8625];
     layer2_out[10053] <= ~layer1_out[4715];
     layer2_out[10054] <= ~layer1_out[7];
     layer2_out[10055] <= layer1_out[4701] & ~layer1_out[4702];
     layer2_out[10056] <= ~(layer1_out[3262] & layer1_out[3263]);
     layer2_out[10057] <= layer1_out[9440] & ~layer1_out[9441];
     layer2_out[10058] <= layer1_out[5459] | layer1_out[5460];
     layer2_out[10059] <= ~layer1_out[6466];
     layer2_out[10060] <= layer1_out[4379] ^ layer1_out[4380];
     layer2_out[10061] <= ~layer1_out[728];
     layer2_out[10062] <= layer1_out[4967];
     layer2_out[10063] <= layer1_out[4904] & ~layer1_out[4905];
     layer2_out[10064] <= ~(layer1_out[9134] & layer1_out[9135]);
     layer2_out[10065] <= ~(layer1_out[10367] ^ layer1_out[10368]);
     layer2_out[10066] <= ~layer1_out[6891];
     layer2_out[10067] <= layer1_out[3331] & ~layer1_out[3330];
     layer2_out[10068] <= layer1_out[6052] & ~layer1_out[6053];
     layer2_out[10069] <= ~(layer1_out[7763] & layer1_out[7764]);
     layer2_out[10070] <= ~(layer1_out[9583] ^ layer1_out[9584]);
     layer2_out[10071] <= ~(layer1_out[7678] & layer1_out[7679]);
     layer2_out[10072] <= layer1_out[9304];
     layer2_out[10073] <= layer1_out[5490] & ~layer1_out[5491];
     layer2_out[10074] <= layer1_out[3485] & ~layer1_out[3484];
     layer2_out[10075] <= layer1_out[2486] & layer1_out[2487];
     layer2_out[10076] <= ~(layer1_out[4341] & layer1_out[4342]);
     layer2_out[10077] <= layer1_out[930] & layer1_out[931];
     layer2_out[10078] <= layer1_out[11169];
     layer2_out[10079] <= layer1_out[11788];
     layer2_out[10080] <= ~layer1_out[10449];
     layer2_out[10081] <= ~layer1_out[1843] | layer1_out[1842];
     layer2_out[10082] <= ~layer1_out[1398];
     layer2_out[10083] <= ~layer1_out[4634];
     layer2_out[10084] <= ~layer1_out[2744];
     layer2_out[10085] <= ~(layer1_out[9838] | layer1_out[9839]);
     layer2_out[10086] <= ~layer1_out[9434];
     layer2_out[10087] <= ~layer1_out[10674];
     layer2_out[10088] <= layer1_out[4519] & ~layer1_out[4518];
     layer2_out[10089] <= ~layer1_out[6092];
     layer2_out[10090] <= ~layer1_out[2372];
     layer2_out[10091] <= layer1_out[4374] & ~layer1_out[4375];
     layer2_out[10092] <= ~layer1_out[627] | layer1_out[628];
     layer2_out[10093] <= ~layer1_out[6218];
     layer2_out[10094] <= ~(layer1_out[3241] | layer1_out[3242]);
     layer2_out[10095] <= ~(layer1_out[5428] | layer1_out[5429]);
     layer2_out[10096] <= ~layer1_out[3172] | layer1_out[3171];
     layer2_out[10097] <= layer1_out[1131] & ~layer1_out[1130];
     layer2_out[10098] <= ~(layer1_out[2384] & layer1_out[2385]);
     layer2_out[10099] <= layer1_out[6988];
     layer2_out[10100] <= layer1_out[411] | layer1_out[412];
     layer2_out[10101] <= layer1_out[4179] & layer1_out[4180];
     layer2_out[10102] <= layer1_out[2900] & ~layer1_out[2901];
     layer2_out[10103] <= layer1_out[8901] ^ layer1_out[8902];
     layer2_out[10104] <= layer1_out[302];
     layer2_out[10105] <= ~(layer1_out[1448] | layer1_out[1449]);
     layer2_out[10106] <= ~layer1_out[7665] | layer1_out[7666];
     layer2_out[10107] <= layer1_out[8119];
     layer2_out[10108] <= layer1_out[6807] & ~layer1_out[6808];
     layer2_out[10109] <= ~layer1_out[9505] | layer1_out[9506];
     layer2_out[10110] <= ~layer1_out[5598] | layer1_out[5597];
     layer2_out[10111] <= layer1_out[3118];
     layer2_out[10112] <= ~(layer1_out[7218] & layer1_out[7219]);
     layer2_out[10113] <= layer1_out[5004] | layer1_out[5005];
     layer2_out[10114] <= layer1_out[3394] ^ layer1_out[3395];
     layer2_out[10115] <= ~layer1_out[985];
     layer2_out[10116] <= layer1_out[5906] & ~layer1_out[5907];
     layer2_out[10117] <= layer1_out[5531];
     layer2_out[10118] <= ~(layer1_out[3096] ^ layer1_out[3097]);
     layer2_out[10119] <= ~layer1_out[6221] | layer1_out[6222];
     layer2_out[10120] <= ~layer1_out[7662] | layer1_out[7661];
     layer2_out[10121] <= ~(layer1_out[11270] & layer1_out[11271]);
     layer2_out[10122] <= ~(layer1_out[4950] & layer1_out[4951]);
     layer2_out[10123] <= ~layer1_out[7052] | layer1_out[7051];
     layer2_out[10124] <= layer1_out[8803] & layer1_out[8804];
     layer2_out[10125] <= ~layer1_out[7026] | layer1_out[7027];
     layer2_out[10126] <= ~layer1_out[4955] | layer1_out[4954];
     layer2_out[10127] <= ~(layer1_out[10861] | layer1_out[10862]);
     layer2_out[10128] <= ~layer1_out[6228];
     layer2_out[10129] <= ~layer1_out[3266];
     layer2_out[10130] <= ~layer1_out[4766] | layer1_out[4765];
     layer2_out[10131] <= layer1_out[5436];
     layer2_out[10132] <= layer1_out[11771] & layer1_out[11772];
     layer2_out[10133] <= layer1_out[4657] & ~layer1_out[4656];
     layer2_out[10134] <= ~(layer1_out[9597] & layer1_out[9598]);
     layer2_out[10135] <= layer1_out[7824] & ~layer1_out[7825];
     layer2_out[10136] <= ~layer1_out[3158] | layer1_out[3159];
     layer2_out[10137] <= 1'b0;
     layer2_out[10138] <= layer1_out[1470] & layer1_out[1471];
     layer2_out[10139] <= ~layer1_out[10778] | layer1_out[10777];
     layer2_out[10140] <= ~layer1_out[7097] | layer1_out[7098];
     layer2_out[10141] <= ~layer1_out[369];
     layer2_out[10142] <= layer1_out[1684];
     layer2_out[10143] <= layer1_out[1050] & ~layer1_out[1051];
     layer2_out[10144] <= layer1_out[5312] & ~layer1_out[5313];
     layer2_out[10145] <= ~layer1_out[1903];
     layer2_out[10146] <= ~(layer1_out[2995] ^ layer1_out[2996]);
     layer2_out[10147] <= layer1_out[998] ^ layer1_out[999];
     layer2_out[10148] <= ~layer1_out[6713];
     layer2_out[10149] <= ~(layer1_out[5263] ^ layer1_out[5264]);
     layer2_out[10150] <= ~layer1_out[9023];
     layer2_out[10151] <= layer1_out[5564];
     layer2_out[10152] <= ~(layer1_out[6630] | layer1_out[6631]);
     layer2_out[10153] <= layer1_out[7117] ^ layer1_out[7118];
     layer2_out[10154] <= ~layer1_out[10845];
     layer2_out[10155] <= layer1_out[2717];
     layer2_out[10156] <= layer1_out[9024];
     layer2_out[10157] <= 1'b1;
     layer2_out[10158] <= layer1_out[3653] & ~layer1_out[3652];
     layer2_out[10159] <= ~(layer1_out[10742] & layer1_out[10743]);
     layer2_out[10160] <= ~layer1_out[8047];
     layer2_out[10161] <= ~layer1_out[5142];
     layer2_out[10162] <= ~layer1_out[3885] | layer1_out[3886];
     layer2_out[10163] <= layer1_out[6681] | layer1_out[6682];
     layer2_out[10164] <= ~layer1_out[9599];
     layer2_out[10165] <= 1'b1;
     layer2_out[10166] <= ~(layer1_out[1028] & layer1_out[1029]);
     layer2_out[10167] <= layer1_out[9017];
     layer2_out[10168] <= layer1_out[4787] & ~layer1_out[4786];
     layer2_out[10169] <= layer1_out[9517];
     layer2_out[10170] <= ~layer1_out[8812] | layer1_out[8813];
     layer2_out[10171] <= ~layer1_out[6179];
     layer2_out[10172] <= ~layer1_out[2772] | layer1_out[2773];
     layer2_out[10173] <= ~layer1_out[7682];
     layer2_out[10174] <= layer1_out[5292] & layer1_out[5293];
     layer2_out[10175] <= layer1_out[6292];
     layer2_out[10176] <= layer1_out[1129];
     layer2_out[10177] <= layer1_out[144] & ~layer1_out[143];
     layer2_out[10178] <= ~layer1_out[1940];
     layer2_out[10179] <= ~layer1_out[1044];
     layer2_out[10180] <= ~layer1_out[5224];
     layer2_out[10181] <= layer1_out[6487];
     layer2_out[10182] <= ~layer1_out[10609];
     layer2_out[10183] <= ~layer1_out[4810];
     layer2_out[10184] <= layer1_out[6203] & ~layer1_out[6204];
     layer2_out[10185] <= 1'b1;
     layer2_out[10186] <= ~layer1_out[54];
     layer2_out[10187] <= ~(layer1_out[7481] & layer1_out[7482]);
     layer2_out[10188] <= ~layer1_out[5521] | layer1_out[5522];
     layer2_out[10189] <= ~(layer1_out[9013] ^ layer1_out[9014]);
     layer2_out[10190] <= ~(layer1_out[964] & layer1_out[965]);
     layer2_out[10191] <= ~layer1_out[10668] | layer1_out[10669];
     layer2_out[10192] <= layer1_out[217];
     layer2_out[10193] <= ~layer1_out[2283] | layer1_out[2282];
     layer2_out[10194] <= layer1_out[1521] & ~layer1_out[1520];
     layer2_out[10195] <= layer1_out[3683] & ~layer1_out[3682];
     layer2_out[10196] <= ~layer1_out[6142];
     layer2_out[10197] <= layer1_out[5983] ^ layer1_out[5984];
     layer2_out[10198] <= ~layer1_out[9090] | layer1_out[9091];
     layer2_out[10199] <= 1'b1;
     layer2_out[10200] <= ~layer1_out[5838];
     layer2_out[10201] <= ~layer1_out[7801] | layer1_out[7802];
     layer2_out[10202] <= ~layer1_out[1953];
     layer2_out[10203] <= layer1_out[11470] & ~layer1_out[11469];
     layer2_out[10204] <= layer1_out[4060];
     layer2_out[10205] <= layer1_out[1784] & ~layer1_out[1785];
     layer2_out[10206] <= ~(layer1_out[6710] & layer1_out[6711]);
     layer2_out[10207] <= layer1_out[7377] | layer1_out[7378];
     layer2_out[10208] <= layer1_out[4972];
     layer2_out[10209] <= layer1_out[9593] ^ layer1_out[9594];
     layer2_out[10210] <= ~(layer1_out[3757] | layer1_out[3758]);
     layer2_out[10211] <= layer1_out[8138];
     layer2_out[10212] <= ~layer1_out[11251] | layer1_out[11250];
     layer2_out[10213] <= ~layer1_out[605];
     layer2_out[10214] <= layer1_out[11628] | layer1_out[11629];
     layer2_out[10215] <= ~(layer1_out[1450] & layer1_out[1451]);
     layer2_out[10216] <= ~(layer1_out[1665] & layer1_out[1666]);
     layer2_out[10217] <= ~layer1_out[10140] | layer1_out[10141];
     layer2_out[10218] <= ~layer1_out[6832];
     layer2_out[10219] <= ~layer1_out[10836];
     layer2_out[10220] <= ~layer1_out[11061];
     layer2_out[10221] <= ~layer1_out[256];
     layer2_out[10222] <= layer1_out[704];
     layer2_out[10223] <= layer1_out[8304] & ~layer1_out[8305];
     layer2_out[10224] <= layer1_out[1546];
     layer2_out[10225] <= ~(layer1_out[6752] ^ layer1_out[6753]);
     layer2_out[10226] <= ~layer1_out[10943];
     layer2_out[10227] <= layer1_out[10735];
     layer2_out[10228] <= ~layer1_out[2597];
     layer2_out[10229] <= layer1_out[4247] | layer1_out[4248];
     layer2_out[10230] <= layer1_out[6568] ^ layer1_out[6569];
     layer2_out[10231] <= ~layer1_out[664] | layer1_out[663];
     layer2_out[10232] <= ~layer1_out[4757];
     layer2_out[10233] <= ~(layer1_out[3941] & layer1_out[3942]);
     layer2_out[10234] <= layer1_out[4401] | layer1_out[4402];
     layer2_out[10235] <= layer1_out[11914] & ~layer1_out[11915];
     layer2_out[10236] <= layer1_out[8032];
     layer2_out[10237] <= ~layer1_out[10867] | layer1_out[10866];
     layer2_out[10238] <= ~(layer1_out[8946] | layer1_out[8947]);
     layer2_out[10239] <= layer1_out[11970] & layer1_out[11971];
     layer2_out[10240] <= layer1_out[1121] | layer1_out[1122];
     layer2_out[10241] <= layer1_out[8291] | layer1_out[8292];
     layer2_out[10242] <= ~layer1_out[9737];
     layer2_out[10243] <= layer1_out[1798];
     layer2_out[10244] <= layer1_out[10874] & ~layer1_out[10875];
     layer2_out[10245] <= layer1_out[527] & ~layer1_out[528];
     layer2_out[10246] <= layer1_out[7623] & ~layer1_out[7622];
     layer2_out[10247] <= layer1_out[8260] & ~layer1_out[8261];
     layer2_out[10248] <= layer1_out[6009] | layer1_out[6010];
     layer2_out[10249] <= ~layer1_out[1163] | layer1_out[1164];
     layer2_out[10250] <= ~(layer1_out[2254] | layer1_out[2255]);
     layer2_out[10251] <= ~(layer1_out[11100] ^ layer1_out[11101]);
     layer2_out[10252] <= layer1_out[8431] & ~layer1_out[8430];
     layer2_out[10253] <= ~layer1_out[11713] | layer1_out[11714];
     layer2_out[10254] <= ~(layer1_out[2931] ^ layer1_out[2932]);
     layer2_out[10255] <= layer1_out[1217] ^ layer1_out[1218];
     layer2_out[10256] <= ~layer1_out[2291] | layer1_out[2290];
     layer2_out[10257] <= layer1_out[807] & layer1_out[808];
     layer2_out[10258] <= ~(layer1_out[6461] ^ layer1_out[6462]);
     layer2_out[10259] <= ~layer1_out[4251];
     layer2_out[10260] <= layer1_out[7333] & layer1_out[7334];
     layer2_out[10261] <= ~layer1_out[8345];
     layer2_out[10262] <= ~layer1_out[7436];
     layer2_out[10263] <= layer1_out[11167] & ~layer1_out[11168];
     layer2_out[10264] <= layer1_out[4443] & ~layer1_out[4444];
     layer2_out[10265] <= layer1_out[6793];
     layer2_out[10266] <= ~(layer1_out[2201] ^ layer1_out[2202]);
     layer2_out[10267] <= ~layer1_out[3079] | layer1_out[3080];
     layer2_out[10268] <= layer1_out[2709];
     layer2_out[10269] <= layer1_out[10225] & layer1_out[10226];
     layer2_out[10270] <= ~layer1_out[5783] | layer1_out[5782];
     layer2_out[10271] <= ~layer1_out[866];
     layer2_out[10272] <= layer1_out[7654] & ~layer1_out[7655];
     layer2_out[10273] <= layer1_out[7599] & layer1_out[7600];
     layer2_out[10274] <= ~(layer1_out[3239] & layer1_out[3240]);
     layer2_out[10275] <= ~(layer1_out[8934] ^ layer1_out[8935]);
     layer2_out[10276] <= layer1_out[3304] | layer1_out[3305];
     layer2_out[10277] <= ~layer1_out[8483] | layer1_out[8482];
     layer2_out[10278] <= ~layer1_out[324] | layer1_out[325];
     layer2_out[10279] <= layer1_out[2280] & ~layer1_out[2281];
     layer2_out[10280] <= ~(layer1_out[6134] | layer1_out[6135]);
     layer2_out[10281] <= layer1_out[2306] | layer1_out[2307];
     layer2_out[10282] <= ~layer1_out[1140];
     layer2_out[10283] <= ~layer1_out[734];
     layer2_out[10284] <= ~layer1_out[5626] | layer1_out[5627];
     layer2_out[10285] <= layer1_out[2430];
     layer2_out[10286] <= layer1_out[5343] & layer1_out[5344];
     layer2_out[10287] <= layer1_out[2362] | layer1_out[2363];
     layer2_out[10288] <= 1'b0;
     layer2_out[10289] <= layer1_out[1690];
     layer2_out[10290] <= ~(layer1_out[5883] ^ layer1_out[5884]);
     layer2_out[10291] <= layer1_out[7667] & layer1_out[7668];
     layer2_out[10292] <= ~(layer1_out[2778] ^ layer1_out[2779]);
     layer2_out[10293] <= layer1_out[7604] | layer1_out[7605];
     layer2_out[10294] <= layer1_out[2968];
     layer2_out[10295] <= ~(layer1_out[10285] | layer1_out[10286]);
     layer2_out[10296] <= ~layer1_out[10];
     layer2_out[10297] <= layer1_out[520] ^ layer1_out[521];
     layer2_out[10298] <= layer1_out[159];
     layer2_out[10299] <= layer1_out[8276] | layer1_out[8277];
     layer2_out[10300] <= layer1_out[4687] & ~layer1_out[4688];
     layer2_out[10301] <= ~layer1_out[1353] | layer1_out[1352];
     layer2_out[10302] <= ~layer1_out[9966];
     layer2_out[10303] <= layer1_out[3130] | layer1_out[3131];
     layer2_out[10304] <= ~(layer1_out[5467] | layer1_out[5468]);
     layer2_out[10305] <= ~layer1_out[5673];
     layer2_out[10306] <= layer1_out[7475] & ~layer1_out[7474];
     layer2_out[10307] <= ~(layer1_out[9939] ^ layer1_out[9940]);
     layer2_out[10308] <= ~layer1_out[8088] | layer1_out[8087];
     layer2_out[10309] <= layer1_out[11302];
     layer2_out[10310] <= layer1_out[7831] | layer1_out[7832];
     layer2_out[10311] <= layer1_out[9300] | layer1_out[9301];
     layer2_out[10312] <= layer1_out[10367] & ~layer1_out[10366];
     layer2_out[10313] <= layer1_out[10915] & layer1_out[10916];
     layer2_out[10314] <= ~(layer1_out[8121] ^ layer1_out[8122]);
     layer2_out[10315] <= layer1_out[5903] ^ layer1_out[5904];
     layer2_out[10316] <= ~layer1_out[8433];
     layer2_out[10317] <= layer1_out[6623];
     layer2_out[10318] <= ~layer1_out[860];
     layer2_out[10319] <= ~layer1_out[7560];
     layer2_out[10320] <= layer1_out[10938] & layer1_out[10939];
     layer2_out[10321] <= layer1_out[5291];
     layer2_out[10322] <= layer1_out[4826];
     layer2_out[10323] <= ~(layer1_out[1479] & layer1_out[1480]);
     layer2_out[10324] <= layer1_out[913] ^ layer1_out[914];
     layer2_out[10325] <= ~(layer1_out[2051] | layer1_out[2052]);
     layer2_out[10326] <= layer1_out[7005];
     layer2_out[10327] <= layer1_out[10930];
     layer2_out[10328] <= layer1_out[15];
     layer2_out[10329] <= ~(layer1_out[10356] & layer1_out[10357]);
     layer2_out[10330] <= ~(layer1_out[11572] | layer1_out[11573]);
     layer2_out[10331] <= ~layer1_out[2735];
     layer2_out[10332] <= layer1_out[2958] | layer1_out[2959];
     layer2_out[10333] <= layer1_out[5944];
     layer2_out[10334] <= layer1_out[2681] & ~layer1_out[2682];
     layer2_out[10335] <= ~(layer1_out[5846] | layer1_out[5847]);
     layer2_out[10336] <= layer1_out[5625] & ~layer1_out[5624];
     layer2_out[10337] <= ~layer1_out[903] | layer1_out[904];
     layer2_out[10338] <= ~layer1_out[10944] | layer1_out[10943];
     layer2_out[10339] <= layer1_out[8192] | layer1_out[8193];
     layer2_out[10340] <= ~(layer1_out[1451] & layer1_out[1452]);
     layer2_out[10341] <= layer1_out[4672];
     layer2_out[10342] <= ~layer1_out[11750];
     layer2_out[10343] <= ~layer1_out[8307];
     layer2_out[10344] <= layer1_out[3903] & layer1_out[3904];
     layer2_out[10345] <= ~layer1_out[11235] | layer1_out[11236];
     layer2_out[10346] <= layer1_out[5200];
     layer2_out[10347] <= ~layer1_out[3563];
     layer2_out[10348] <= layer1_out[8475] & ~layer1_out[8476];
     layer2_out[10349] <= layer1_out[6105] ^ layer1_out[6106];
     layer2_out[10350] <= ~layer1_out[1261] | layer1_out[1262];
     layer2_out[10351] <= ~layer1_out[9984] | layer1_out[9985];
     layer2_out[10352] <= ~layer1_out[4629];
     layer2_out[10353] <= ~(layer1_out[10072] & layer1_out[10073]);
     layer2_out[10354] <= ~(layer1_out[3845] & layer1_out[3846]);
     layer2_out[10355] <= layer1_out[5643];
     layer2_out[10356] <= layer1_out[664];
     layer2_out[10357] <= ~layer1_out[10527];
     layer2_out[10358] <= ~(layer1_out[8557] ^ layer1_out[8558]);
     layer2_out[10359] <= ~(layer1_out[11888] | layer1_out[11889]);
     layer2_out[10360] <= ~(layer1_out[7153] | layer1_out[7154]);
     layer2_out[10361] <= layer1_out[5024];
     layer2_out[10362] <= ~(layer1_out[4318] ^ layer1_out[4319]);
     layer2_out[10363] <= layer1_out[4253];
     layer2_out[10364] <= ~layer1_out[3329];
     layer2_out[10365] <= layer1_out[1097] & layer1_out[1098];
     layer2_out[10366] <= ~layer1_out[1841];
     layer2_out[10367] <= ~(layer1_out[1503] & layer1_out[1504]);
     layer2_out[10368] <= ~layer1_out[10819] | layer1_out[10818];
     layer2_out[10369] <= layer1_out[1731];
     layer2_out[10370] <= layer1_out[6407] & ~layer1_out[6406];
     layer2_out[10371] <= ~layer1_out[379];
     layer2_out[10372] <= layer1_out[2188];
     layer2_out[10373] <= layer1_out[11937] ^ layer1_out[11938];
     layer2_out[10374] <= ~layer1_out[3544];
     layer2_out[10375] <= layer1_out[10205];
     layer2_out[10376] <= layer1_out[10962];
     layer2_out[10377] <= ~layer1_out[8030];
     layer2_out[10378] <= layer1_out[9480];
     layer2_out[10379] <= layer1_out[1340] & layer1_out[1341];
     layer2_out[10380] <= ~(layer1_out[3683] ^ layer1_out[3684]);
     layer2_out[10381] <= layer1_out[853] ^ layer1_out[854];
     layer2_out[10382] <= ~layer1_out[5563];
     layer2_out[10383] <= layer1_out[8238] & ~layer1_out[8237];
     layer2_out[10384] <= layer1_out[6562] & ~layer1_out[6561];
     layer2_out[10385] <= ~(layer1_out[205] | layer1_out[206]);
     layer2_out[10386] <= layer1_out[10191] & layer1_out[10192];
     layer2_out[10387] <= ~layer1_out[648];
     layer2_out[10388] <= layer1_out[5550] ^ layer1_out[5551];
     layer2_out[10389] <= layer1_out[10725] & layer1_out[10726];
     layer2_out[10390] <= ~layer1_out[1927];
     layer2_out[10391] <= ~layer1_out[9441];
     layer2_out[10392] <= layer1_out[1390];
     layer2_out[10393] <= layer1_out[5942] & layer1_out[5943];
     layer2_out[10394] <= layer1_out[8420];
     layer2_out[10395] <= layer1_out[10039];
     layer2_out[10396] <= layer1_out[1541] & ~layer1_out[1542];
     layer2_out[10397] <= ~layer1_out[6558];
     layer2_out[10398] <= ~layer1_out[2233] | layer1_out[2234];
     layer2_out[10399] <= layer1_out[5350];
     layer2_out[10400] <= ~layer1_out[1157] | layer1_out[1156];
     layer2_out[10401] <= layer1_out[2146];
     layer2_out[10402] <= layer1_out[1888];
     layer2_out[10403] <= ~layer1_out[9558] | layer1_out[9559];
     layer2_out[10404] <= ~layer1_out[10912];
     layer2_out[10405] <= layer1_out[8387] & layer1_out[8388];
     layer2_out[10406] <= layer1_out[3213] ^ layer1_out[3214];
     layer2_out[10407] <= ~layer1_out[2090];
     layer2_out[10408] <= ~layer1_out[2867];
     layer2_out[10409] <= layer1_out[783] | layer1_out[784];
     layer2_out[10410] <= layer1_out[11162] & ~layer1_out[11163];
     layer2_out[10411] <= layer1_out[2964];
     layer2_out[10412] <= ~(layer1_out[11885] | layer1_out[11886]);
     layer2_out[10413] <= ~layer1_out[9326] | layer1_out[9327];
     layer2_out[10414] <= ~layer1_out[323] | layer1_out[324];
     layer2_out[10415] <= ~layer1_out[4407];
     layer2_out[10416] <= ~layer1_out[7825];
     layer2_out[10417] <= ~layer1_out[1928];
     layer2_out[10418] <= layer1_out[10865] & ~layer1_out[10864];
     layer2_out[10419] <= layer1_out[1955] | layer1_out[1956];
     layer2_out[10420] <= ~(layer1_out[376] & layer1_out[377]);
     layer2_out[10421] <= ~(layer1_out[2723] ^ layer1_out[2724]);
     layer2_out[10422] <= layer1_out[7834] & ~layer1_out[7833];
     layer2_out[10423] <= ~layer1_out[2490] | layer1_out[2489];
     layer2_out[10424] <= layer1_out[5647];
     layer2_out[10425] <= ~layer1_out[5086];
     layer2_out[10426] <= layer1_out[3746] ^ layer1_out[3747];
     layer2_out[10427] <= layer1_out[5192];
     layer2_out[10428] <= ~layer1_out[3620];
     layer2_out[10429] <= ~(layer1_out[5496] | layer1_out[5497]);
     layer2_out[10430] <= ~(layer1_out[5567] & layer1_out[5568]);
     layer2_out[10431] <= ~layer1_out[9342] | layer1_out[9343];
     layer2_out[10432] <= ~(layer1_out[1001] & layer1_out[1002]);
     layer2_out[10433] <= ~(layer1_out[2779] ^ layer1_out[2780]);
     layer2_out[10434] <= layer1_out[6879] & layer1_out[6880];
     layer2_out[10435] <= layer1_out[2407];
     layer2_out[10436] <= ~(layer1_out[9636] | layer1_out[9637]);
     layer2_out[10437] <= layer1_out[6435];
     layer2_out[10438] <= ~(layer1_out[7019] & layer1_out[7020]);
     layer2_out[10439] <= layer1_out[5981] & ~layer1_out[5982];
     layer2_out[10440] <= layer1_out[8702];
     layer2_out[10441] <= layer1_out[3181] | layer1_out[3182];
     layer2_out[10442] <= ~(layer1_out[10575] & layer1_out[10576]);
     layer2_out[10443] <= ~layer1_out[8116] | layer1_out[8115];
     layer2_out[10444] <= layer1_out[6696] ^ layer1_out[6697];
     layer2_out[10445] <= layer1_out[6331];
     layer2_out[10446] <= ~layer1_out[1248];
     layer2_out[10447] <= ~(layer1_out[6011] | layer1_out[6012]);
     layer2_out[10448] <= ~(layer1_out[1692] & layer1_out[1693]);
     layer2_out[10449] <= layer1_out[10837];
     layer2_out[10450] <= ~layer1_out[7812];
     layer2_out[10451] <= ~(layer1_out[9508] ^ layer1_out[9509]);
     layer2_out[10452] <= ~layer1_out[10582] | layer1_out[10583];
     layer2_out[10453] <= layer1_out[2944];
     layer2_out[10454] <= layer1_out[1737] & layer1_out[1738];
     layer2_out[10455] <= layer1_out[2835];
     layer2_out[10456] <= 1'b0;
     layer2_out[10457] <= ~layer1_out[6399] | layer1_out[6398];
     layer2_out[10458] <= layer1_out[10592] & ~layer1_out[10591];
     layer2_out[10459] <= ~layer1_out[9346] | layer1_out[9347];
     layer2_out[10460] <= layer1_out[9530];
     layer2_out[10461] <= layer1_out[4680] & layer1_out[4681];
     layer2_out[10462] <= layer1_out[2588] | layer1_out[2589];
     layer2_out[10463] <= layer1_out[7700];
     layer2_out[10464] <= ~layer1_out[4551];
     layer2_out[10465] <= ~(layer1_out[5450] ^ layer1_out[5451]);
     layer2_out[10466] <= ~(layer1_out[5974] & layer1_out[5975]);
     layer2_out[10467] <= layer1_out[2749] ^ layer1_out[2750];
     layer2_out[10468] <= ~layer1_out[3561];
     layer2_out[10469] <= layer1_out[5338] & layer1_out[5339];
     layer2_out[10470] <= layer1_out[6893] ^ layer1_out[6894];
     layer2_out[10471] <= 1'b1;
     layer2_out[10472] <= ~layer1_out[7043] | layer1_out[7044];
     layer2_out[10473] <= ~(layer1_out[7013] | layer1_out[7014]);
     layer2_out[10474] <= ~(layer1_out[5697] & layer1_out[5698]);
     layer2_out[10475] <= layer1_out[9728] & ~layer1_out[9729];
     layer2_out[10476] <= ~(layer1_out[2887] ^ layer1_out[2888]);
     layer2_out[10477] <= layer1_out[486];
     layer2_out[10478] <= layer1_out[4927];
     layer2_out[10479] <= ~layer1_out[5059];
     layer2_out[10480] <= ~layer1_out[11686] | layer1_out[11685];
     layer2_out[10481] <= ~layer1_out[7492];
     layer2_out[10482] <= layer1_out[3113] | layer1_out[3114];
     layer2_out[10483] <= ~layer1_out[6364];
     layer2_out[10484] <= layer1_out[11811] | layer1_out[11812];
     layer2_out[10485] <= ~(layer1_out[3520] | layer1_out[3521]);
     layer2_out[10486] <= ~layer1_out[2756];
     layer2_out[10487] <= layer1_out[1515] | layer1_out[1516];
     layer2_out[10488] <= layer1_out[6813] & ~layer1_out[6812];
     layer2_out[10489] <= ~(layer1_out[8816] & layer1_out[8817]);
     layer2_out[10490] <= ~layer1_out[8671];
     layer2_out[10491] <= ~layer1_out[8207] | layer1_out[8208];
     layer2_out[10492] <= 1'b1;
     layer2_out[10493] <= ~layer1_out[5247] | layer1_out[5246];
     layer2_out[10494] <= layer1_out[7846] ^ layer1_out[7847];
     layer2_out[10495] <= layer1_out[1244] & ~layer1_out[1243];
     layer2_out[10496] <= ~(layer1_out[138] & layer1_out[139]);
     layer2_out[10497] <= layer1_out[10459] & layer1_out[10460];
     layer2_out[10498] <= ~(layer1_out[2665] & layer1_out[2666]);
     layer2_out[10499] <= ~layer1_out[677];
     layer2_out[10500] <= layer1_out[2505] & ~layer1_out[2506];
     layer2_out[10501] <= layer1_out[5103] & ~layer1_out[5102];
     layer2_out[10502] <= ~layer1_out[2508] | layer1_out[2509];
     layer2_out[10503] <= layer1_out[1283];
     layer2_out[10504] <= layer1_out[3676] & ~layer1_out[3677];
     layer2_out[10505] <= layer1_out[4475];
     layer2_out[10506] <= ~layer1_out[10498];
     layer2_out[10507] <= layer1_out[4527] ^ layer1_out[4528];
     layer2_out[10508] <= ~layer1_out[1851];
     layer2_out[10509] <= layer1_out[5759] ^ layer1_out[5760];
     layer2_out[10510] <= layer1_out[8363] & ~layer1_out[8362];
     layer2_out[10511] <= layer1_out[1200] & ~layer1_out[1201];
     layer2_out[10512] <= ~layer1_out[6862];
     layer2_out[10513] <= ~layer1_out[428] | layer1_out[427];
     layer2_out[10514] <= layer1_out[2197];
     layer2_out[10515] <= ~(layer1_out[5002] ^ layer1_out[5003]);
     layer2_out[10516] <= ~layer1_out[10170] | layer1_out[10169];
     layer2_out[10517] <= ~layer1_out[10678];
     layer2_out[10518] <= layer1_out[4177];
     layer2_out[10519] <= ~(layer1_out[7703] ^ layer1_out[7704]);
     layer2_out[10520] <= ~(layer1_out[10106] & layer1_out[10107]);
     layer2_out[10521] <= ~(layer1_out[6466] | layer1_out[6467]);
     layer2_out[10522] <= layer1_out[4377] | layer1_out[4378];
     layer2_out[10523] <= ~(layer1_out[6447] & layer1_out[6448]);
     layer2_out[10524] <= layer1_out[10870] | layer1_out[10871];
     layer2_out[10525] <= layer1_out[3156] & layer1_out[3157];
     layer2_out[10526] <= ~layer1_out[7096];
     layer2_out[10527] <= layer1_out[4736] & ~layer1_out[4735];
     layer2_out[10528] <= layer1_out[10645] | layer1_out[10646];
     layer2_out[10529] <= ~layer1_out[9315] | layer1_out[9316];
     layer2_out[10530] <= ~layer1_out[2066];
     layer2_out[10531] <= ~(layer1_out[366] ^ layer1_out[367]);
     layer2_out[10532] <= layer1_out[1035] & layer1_out[1036];
     layer2_out[10533] <= ~layer1_out[10177];
     layer2_out[10534] <= layer1_out[9296] & layer1_out[9297];
     layer2_out[10535] <= ~(layer1_out[10077] & layer1_out[10078]);
     layer2_out[10536] <= layer1_out[7702] & layer1_out[7703];
     layer2_out[10537] <= layer1_out[3961];
     layer2_out[10538] <= layer1_out[6692] & ~layer1_out[6693];
     layer2_out[10539] <= ~(layer1_out[260] | layer1_out[261]);
     layer2_out[10540] <= ~(layer1_out[8262] | layer1_out[8263]);
     layer2_out[10541] <= ~layer1_out[6345] | layer1_out[6346];
     layer2_out[10542] <= layer1_out[7769];
     layer2_out[10543] <= layer1_out[11589] & layer1_out[11590];
     layer2_out[10544] <= layer1_out[883];
     layer2_out[10545] <= layer1_out[5234];
     layer2_out[10546] <= ~layer1_out[10758];
     layer2_out[10547] <= ~(layer1_out[9785] | layer1_out[9786]);
     layer2_out[10548] <= layer1_out[8354];
     layer2_out[10549] <= layer1_out[4752] & layer1_out[4753];
     layer2_out[10550] <= ~layer1_out[10361];
     layer2_out[10551] <= layer1_out[7050];
     layer2_out[10552] <= layer1_out[10329];
     layer2_out[10553] <= layer1_out[7230];
     layer2_out[10554] <= ~layer1_out[8725];
     layer2_out[10555] <= layer1_out[1622] & layer1_out[1623];
     layer2_out[10556] <= layer1_out[9782] & ~layer1_out[9783];
     layer2_out[10557] <= layer1_out[11904] | layer1_out[11905];
     layer2_out[10558] <= ~(layer1_out[2355] & layer1_out[2356]);
     layer2_out[10559] <= ~layer1_out[837];
     layer2_out[10560] <= ~layer1_out[2927] | layer1_out[2928];
     layer2_out[10561] <= ~(layer1_out[8849] ^ layer1_out[8850]);
     layer2_out[10562] <= ~layer1_out[9557];
     layer2_out[10563] <= ~layer1_out[3709] | layer1_out[3708];
     layer2_out[10564] <= ~(layer1_out[7975] | layer1_out[7976]);
     layer2_out[10565] <= ~(layer1_out[11580] & layer1_out[11581]);
     layer2_out[10566] <= ~(layer1_out[1256] & layer1_out[1257]);
     layer2_out[10567] <= ~layer1_out[3780];
     layer2_out[10568] <= ~layer1_out[1261] | layer1_out[1260];
     layer2_out[10569] <= layer1_out[611] | layer1_out[612];
     layer2_out[10570] <= layer1_out[8992] ^ layer1_out[8993];
     layer2_out[10571] <= layer1_out[8331] | layer1_out[8332];
     layer2_out[10572] <= ~layer1_out[1595];
     layer2_out[10573] <= layer1_out[6804];
     layer2_out[10574] <= layer1_out[10323] & ~layer1_out[10322];
     layer2_out[10575] <= ~(layer1_out[8921] & layer1_out[8922]);
     layer2_out[10576] <= layer1_out[10340];
     layer2_out[10577] <= layer1_out[9900];
     layer2_out[10578] <= layer1_out[7586] & ~layer1_out[7585];
     layer2_out[10579] <= ~layer1_out[4510];
     layer2_out[10580] <= layer1_out[937];
     layer2_out[10581] <= ~layer1_out[8893] | layer1_out[8894];
     layer2_out[10582] <= ~layer1_out[4884];
     layer2_out[10583] <= ~layer1_out[5074];
     layer2_out[10584] <= ~layer1_out[3476];
     layer2_out[10585] <= ~layer1_out[1584];
     layer2_out[10586] <= layer1_out[6225] & ~layer1_out[6224];
     layer2_out[10587] <= layer1_out[3566];
     layer2_out[10588] <= ~layer1_out[7249] | layer1_out[7250];
     layer2_out[10589] <= ~layer1_out[2106];
     layer2_out[10590] <= ~layer1_out[603] | layer1_out[602];
     layer2_out[10591] <= ~layer1_out[5623];
     layer2_out[10592] <= ~layer1_out[9523] | layer1_out[9522];
     layer2_out[10593] <= layer1_out[7630] & ~layer1_out[7629];
     layer2_out[10594] <= ~layer1_out[5875];
     layer2_out[10595] <= ~layer1_out[10165];
     layer2_out[10596] <= layer1_out[2062] & ~layer1_out[2063];
     layer2_out[10597] <= layer1_out[7683] & layer1_out[7684];
     layer2_out[10598] <= ~layer1_out[7110];
     layer2_out[10599] <= layer1_out[6000];
     layer2_out[10600] <= layer1_out[9480];
     layer2_out[10601] <= ~layer1_out[7575] | layer1_out[7576];
     layer2_out[10602] <= layer1_out[1997] & ~layer1_out[1998];
     layer2_out[10603] <= layer1_out[8371];
     layer2_out[10604] <= ~(layer1_out[6078] & layer1_out[6079]);
     layer2_out[10605] <= ~(layer1_out[7950] | layer1_out[7951]);
     layer2_out[10606] <= ~(layer1_out[4958] & layer1_out[4959]);
     layer2_out[10607] <= layer1_out[9405];
     layer2_out[10608] <= ~layer1_out[4899];
     layer2_out[10609] <= layer1_out[6416];
     layer2_out[10610] <= layer1_out[5550] & ~layer1_out[5549];
     layer2_out[10611] <= layer1_out[973];
     layer2_out[10612] <= ~(layer1_out[1600] | layer1_out[1601]);
     layer2_out[10613] <= ~layer1_out[3224];
     layer2_out[10614] <= ~(layer1_out[5564] & layer1_out[5565]);
     layer2_out[10615] <= layer1_out[5415];
     layer2_out[10616] <= ~layer1_out[11240] | layer1_out[11239];
     layer2_out[10617] <= ~layer1_out[5705];
     layer2_out[10618] <= ~layer1_out[6654];
     layer2_out[10619] <= ~(layer1_out[2365] ^ layer1_out[2366]);
     layer2_out[10620] <= ~layer1_out[9383] | layer1_out[9382];
     layer2_out[10621] <= ~layer1_out[11200];
     layer2_out[10622] <= layer1_out[9213];
     layer2_out[10623] <= ~layer1_out[5119];
     layer2_out[10624] <= layer1_out[5771];
     layer2_out[10625] <= layer1_out[9440];
     layer2_out[10626] <= ~(layer1_out[3734] & layer1_out[3735]);
     layer2_out[10627] <= layer1_out[80] ^ layer1_out[81];
     layer2_out[10628] <= layer1_out[9732] & ~layer1_out[9733];
     layer2_out[10629] <= layer1_out[11991];
     layer2_out[10630] <= ~(layer1_out[4879] | layer1_out[4880]);
     layer2_out[10631] <= ~layer1_out[6812] | layer1_out[6811];
     layer2_out[10632] <= 1'b0;
     layer2_out[10633] <= layer1_out[668] ^ layer1_out[669];
     layer2_out[10634] <= ~(layer1_out[2446] ^ layer1_out[2447]);
     layer2_out[10635] <= ~layer1_out[2059] | layer1_out[2058];
     layer2_out[10636] <= ~layer1_out[988];
     layer2_out[10637] <= ~(layer1_out[4035] | layer1_out[4036]);
     layer2_out[10638] <= ~layer1_out[11240];
     layer2_out[10639] <= ~(layer1_out[6933] | layer1_out[6934]);
     layer2_out[10640] <= ~layer1_out[9912];
     layer2_out[10641] <= ~layer1_out[8771];
     layer2_out[10642] <= layer1_out[5938] & layer1_out[5939];
     layer2_out[10643] <= ~(layer1_out[10885] & layer1_out[10886]);
     layer2_out[10644] <= ~(layer1_out[5418] ^ layer1_out[5419]);
     layer2_out[10645] <= ~(layer1_out[352] & layer1_out[353]);
     layer2_out[10646] <= ~layer1_out[7507];
     layer2_out[10647] <= layer1_out[3701] | layer1_out[3702];
     layer2_out[10648] <= layer1_out[1278];
     layer2_out[10649] <= layer1_out[10196];
     layer2_out[10650] <= ~(layer1_out[8424] & layer1_out[8425]);
     layer2_out[10651] <= layer1_out[4047];
     layer2_out[10652] <= ~layer1_out[1310];
     layer2_out[10653] <= ~layer1_out[1770] | layer1_out[1771];
     layer2_out[10654] <= ~layer1_out[2529] | layer1_out[2528];
     layer2_out[10655] <= layer1_out[629];
     layer2_out[10656] <= layer1_out[7740] & layer1_out[7741];
     layer2_out[10657] <= layer1_out[4384] | layer1_out[4385];
     layer2_out[10658] <= ~layer1_out[11652];
     layer2_out[10659] <= ~layer1_out[11611] | layer1_out[11612];
     layer2_out[10660] <= ~(layer1_out[219] | layer1_out[220]);
     layer2_out[10661] <= ~(layer1_out[8297] & layer1_out[8298]);
     layer2_out[10662] <= layer1_out[9357] & ~layer1_out[9358];
     layer2_out[10663] <= ~layer1_out[8754];
     layer2_out[10664] <= ~layer1_out[3217] | layer1_out[3218];
     layer2_out[10665] <= ~layer1_out[1645];
     layer2_out[10666] <= ~layer1_out[7028];
     layer2_out[10667] <= ~layer1_out[11870] | layer1_out[11869];
     layer2_out[10668] <= layer1_out[2212] ^ layer1_out[2213];
     layer2_out[10669] <= layer1_out[11421];
     layer2_out[10670] <= layer1_out[7354];
     layer2_out[10671] <= ~layer1_out[3647] | layer1_out[3646];
     layer2_out[10672] <= layer1_out[10312] & ~layer1_out[10311];
     layer2_out[10673] <= ~(layer1_out[6100] ^ layer1_out[6101]);
     layer2_out[10674] <= ~(layer1_out[11134] ^ layer1_out[11135]);
     layer2_out[10675] <= layer1_out[4567] & ~layer1_out[4568];
     layer2_out[10676] <= layer1_out[9461] & ~layer1_out[9460];
     layer2_out[10677] <= ~layer1_out[3805];
     layer2_out[10678] <= layer1_out[6484] & ~layer1_out[6483];
     layer2_out[10679] <= ~(layer1_out[9625] | layer1_out[9626]);
     layer2_out[10680] <= layer1_out[3752];
     layer2_out[10681] <= layer1_out[6779] & layer1_out[6780];
     layer2_out[10682] <= ~layer1_out[7748];
     layer2_out[10683] <= ~layer1_out[945] | layer1_out[944];
     layer2_out[10684] <= ~layer1_out[10081];
     layer2_out[10685] <= layer1_out[4151];
     layer2_out[10686] <= ~(layer1_out[804] ^ layer1_out[805]);
     layer2_out[10687] <= layer1_out[11532];
     layer2_out[10688] <= ~layer1_out[9720] | layer1_out[9721];
     layer2_out[10689] <= ~layer1_out[9572] | layer1_out[9571];
     layer2_out[10690] <= layer1_out[8365];
     layer2_out[10691] <= layer1_out[11257];
     layer2_out[10692] <= ~layer1_out[795];
     layer2_out[10693] <= layer1_out[4487];
     layer2_out[10694] <= ~layer1_out[9262] | layer1_out[9261];
     layer2_out[10695] <= layer1_out[10922];
     layer2_out[10696] <= ~layer1_out[9496];
     layer2_out[10697] <= layer1_out[11285] & ~layer1_out[11284];
     layer2_out[10698] <= ~layer1_out[7258];
     layer2_out[10699] <= ~(layer1_out[1088] | layer1_out[1089]);
     layer2_out[10700] <= ~layer1_out[8940];
     layer2_out[10701] <= ~layer1_out[6647];
     layer2_out[10702] <= ~layer1_out[8958];
     layer2_out[10703] <= ~(layer1_out[11208] & layer1_out[11209]);
     layer2_out[10704] <= ~layer1_out[10233];
     layer2_out[10705] <= ~layer1_out[7989];
     layer2_out[10706] <= layer1_out[5358];
     layer2_out[10707] <= layer1_out[5191];
     layer2_out[10708] <= layer1_out[6319] & ~layer1_out[6318];
     layer2_out[10709] <= layer1_out[11072] & ~layer1_out[11071];
     layer2_out[10710] <= ~(layer1_out[10814] ^ layer1_out[10815]);
     layer2_out[10711] <= ~(layer1_out[1667] | layer1_out[1668]);
     layer2_out[10712] <= layer1_out[8262] & ~layer1_out[8261];
     layer2_out[10713] <= layer1_out[10939] & ~layer1_out[10940];
     layer2_out[10714] <= layer1_out[6387] ^ layer1_out[6388];
     layer2_out[10715] <= ~(layer1_out[5620] ^ layer1_out[5621]);
     layer2_out[10716] <= layer1_out[11373];
     layer2_out[10717] <= ~layer1_out[4792] | layer1_out[4791];
     layer2_out[10718] <= ~layer1_out[11451];
     layer2_out[10719] <= layer1_out[181] | layer1_out[182];
     layer2_out[10720] <= layer1_out[10050] & ~layer1_out[10049];
     layer2_out[10721] <= ~(layer1_out[8239] ^ layer1_out[8240]);
     layer2_out[10722] <= layer1_out[9315] & ~layer1_out[9314];
     layer2_out[10723] <= ~(layer1_out[10509] ^ layer1_out[10510]);
     layer2_out[10724] <= layer1_out[1699] & ~layer1_out[1700];
     layer2_out[10725] <= ~layer1_out[3754] | layer1_out[3755];
     layer2_out[10726] <= layer1_out[9206];
     layer2_out[10727] <= ~(layer1_out[8018] ^ layer1_out[8019]);
     layer2_out[10728] <= layer1_out[7120] ^ layer1_out[7121];
     layer2_out[10729] <= layer1_out[3942];
     layer2_out[10730] <= layer1_out[5511] & ~layer1_out[5510];
     layer2_out[10731] <= ~(layer1_out[10849] | layer1_out[10850]);
     layer2_out[10732] <= ~(layer1_out[4276] | layer1_out[4277]);
     layer2_out[10733] <= ~layer1_out[4409] | layer1_out[4410];
     layer2_out[10734] <= layer1_out[9528] & ~layer1_out[9529];
     layer2_out[10735] <= ~layer1_out[5934];
     layer2_out[10736] <= ~(layer1_out[1487] & layer1_out[1488]);
     layer2_out[10737] <= layer1_out[5305] & ~layer1_out[5306];
     layer2_out[10738] <= layer1_out[8178];
     layer2_out[10739] <= ~layer1_out[1384];
     layer2_out[10740] <= ~layer1_out[180];
     layer2_out[10741] <= 1'b0;
     layer2_out[10742] <= ~(layer1_out[2539] ^ layer1_out[2540]);
     layer2_out[10743] <= layer1_out[11148];
     layer2_out[10744] <= layer1_out[5523] & ~layer1_out[5524];
     layer2_out[10745] <= 1'b0;
     layer2_out[10746] <= ~layer1_out[2248] | layer1_out[2247];
     layer2_out[10747] <= layer1_out[1026] & ~layer1_out[1027];
     layer2_out[10748] <= layer1_out[8102] ^ layer1_out[8103];
     layer2_out[10749] <= layer1_out[9135];
     layer2_out[10750] <= 1'b0;
     layer2_out[10751] <= layer1_out[7978] & ~layer1_out[7977];
     layer2_out[10752] <= ~(layer1_out[4584] & layer1_out[4585]);
     layer2_out[10753] <= layer1_out[2929];
     layer2_out[10754] <= layer1_out[3675] & layer1_out[3676];
     layer2_out[10755] <= ~layer1_out[70];
     layer2_out[10756] <= ~layer1_out[6267];
     layer2_out[10757] <= layer1_out[3360] ^ layer1_out[3361];
     layer2_out[10758] <= ~(layer1_out[2371] ^ layer1_out[2372]);
     layer2_out[10759] <= layer1_out[2227] & layer1_out[2228];
     layer2_out[10760] <= layer1_out[6291] & ~layer1_out[6290];
     layer2_out[10761] <= layer1_out[9389] & ~layer1_out[9388];
     layer2_out[10762] <= layer1_out[8359] & layer1_out[8360];
     layer2_out[10763] <= layer1_out[7179] | layer1_out[7180];
     layer2_out[10764] <= ~layer1_out[9408];
     layer2_out[10765] <= ~(layer1_out[11065] ^ layer1_out[11066]);
     layer2_out[10766] <= ~layer1_out[8093];
     layer2_out[10767] <= ~(layer1_out[3623] | layer1_out[3624]);
     layer2_out[10768] <= layer1_out[9747];
     layer2_out[10769] <= layer1_out[11474];
     layer2_out[10770] <= ~layer1_out[934];
     layer2_out[10771] <= ~layer1_out[7795];
     layer2_out[10772] <= layer1_out[7345];
     layer2_out[10773] <= layer1_out[4649] | layer1_out[4650];
     layer2_out[10774] <= layer1_out[8827];
     layer2_out[10775] <= ~layer1_out[7663];
     layer2_out[10776] <= ~(layer1_out[5014] & layer1_out[5015]);
     layer2_out[10777] <= layer1_out[1315];
     layer2_out[10778] <= ~(layer1_out[5075] | layer1_out[5076]);
     layer2_out[10779] <= layer1_out[4075] & layer1_out[4076];
     layer2_out[10780] <= layer1_out[11965] | layer1_out[11966];
     layer2_out[10781] <= ~layer1_out[4360] | layer1_out[4359];
     layer2_out[10782] <= ~layer1_out[318];
     layer2_out[10783] <= ~(layer1_out[1122] ^ layer1_out[1123]);
     layer2_out[10784] <= layer1_out[1994] & layer1_out[1995];
     layer2_out[10785] <= ~layer1_out[4808];
     layer2_out[10786] <= layer1_out[4982];
     layer2_out[10787] <= ~layer1_out[8851];
     layer2_out[10788] <= layer1_out[8942] | layer1_out[8943];
     layer2_out[10789] <= ~(layer1_out[4621] | layer1_out[4622]);
     layer2_out[10790] <= layer1_out[9695] & layer1_out[9696];
     layer2_out[10791] <= ~layer1_out[6022] | layer1_out[6021];
     layer2_out[10792] <= ~layer1_out[5362];
     layer2_out[10793] <= ~layer1_out[2627];
     layer2_out[10794] <= ~layer1_out[4195];
     layer2_out[10795] <= layer1_out[11665] & ~layer1_out[11666];
     layer2_out[10796] <= ~(layer1_out[2352] & layer1_out[2353]);
     layer2_out[10797] <= layer1_out[5668] & ~layer1_out[5667];
     layer2_out[10798] <= ~layer1_out[4372] | layer1_out[4373];
     layer2_out[10799] <= layer1_out[8469] | layer1_out[8470];
     layer2_out[10800] <= ~layer1_out[3799];
     layer2_out[10801] <= ~layer1_out[3019];
     layer2_out[10802] <= ~(layer1_out[8754] & layer1_out[8755]);
     layer2_out[10803] <= ~(layer1_out[7122] | layer1_out[7123]);
     layer2_out[10804] <= ~layer1_out[3445];
     layer2_out[10805] <= ~(layer1_out[1502] & layer1_out[1503]);
     layer2_out[10806] <= ~layer1_out[470];
     layer2_out[10807] <= layer1_out[1495];
     layer2_out[10808] <= layer1_out[2959] & layer1_out[2960];
     layer2_out[10809] <= ~layer1_out[11681];
     layer2_out[10810] <= ~layer1_out[2992];
     layer2_out[10811] <= ~layer1_out[10137];
     layer2_out[10812] <= ~(layer1_out[5571] ^ layer1_out[5572]);
     layer2_out[10813] <= layer1_out[706] & ~layer1_out[707];
     layer2_out[10814] <= ~layer1_out[7482];
     layer2_out[10815] <= layer1_out[5678] | layer1_out[5679];
     layer2_out[10816] <= layer1_out[9402] & layer1_out[9403];
     layer2_out[10817] <= layer1_out[2769] | layer1_out[2770];
     layer2_out[10818] <= ~(layer1_out[9336] | layer1_out[9337]);
     layer2_out[10819] <= ~layer1_out[741];
     layer2_out[10820] <= layer1_out[7672] & ~layer1_out[7673];
     layer2_out[10821] <= layer1_out[4650] & layer1_out[4651];
     layer2_out[10822] <= ~(layer1_out[9657] & layer1_out[9658]);
     layer2_out[10823] <= ~layer1_out[7441];
     layer2_out[10824] <= layer1_out[6887];
     layer2_out[10825] <= layer1_out[3356];
     layer2_out[10826] <= layer1_out[538];
     layer2_out[10827] <= ~(layer1_out[3669] & layer1_out[3670]);
     layer2_out[10828] <= layer1_out[1041] & ~layer1_out[1042];
     layer2_out[10829] <= layer1_out[5794];
     layer2_out[10830] <= ~layer1_out[1306];
     layer2_out[10831] <= ~(layer1_out[9964] & layer1_out[9965]);
     layer2_out[10832] <= ~layer1_out[8225] | layer1_out[8226];
     layer2_out[10833] <= ~(layer1_out[2105] ^ layer1_out[2106]);
     layer2_out[10834] <= ~layer1_out[10305];
     layer2_out[10835] <= ~layer1_out[425] | layer1_out[426];
     layer2_out[10836] <= layer1_out[1295];
     layer2_out[10837] <= ~(layer1_out[11898] | layer1_out[11899]);
     layer2_out[10838] <= layer1_out[7438] | layer1_out[7439];
     layer2_out[10839] <= ~layer1_out[5576] | layer1_out[5575];
     layer2_out[10840] <= ~layer1_out[2193];
     layer2_out[10841] <= ~layer1_out[8002];
     layer2_out[10842] <= ~(layer1_out[2685] | layer1_out[2686]);
     layer2_out[10843] <= ~layer1_out[2624];
     layer2_out[10844] <= layer1_out[1723] | layer1_out[1724];
     layer2_out[10845] <= ~(layer1_out[2012] ^ layer1_out[2013]);
     layer2_out[10846] <= layer1_out[653] ^ layer1_out[654];
     layer2_out[10847] <= ~(layer1_out[4970] ^ layer1_out[4971]);
     layer2_out[10848] <= ~(layer1_out[622] ^ layer1_out[623]);
     layer2_out[10849] <= layer1_out[501] | layer1_out[502];
     layer2_out[10850] <= layer1_out[11575] & layer1_out[11576];
     layer2_out[10851] <= ~layer1_out[4327];
     layer2_out[10852] <= ~(layer1_out[7060] & layer1_out[7061]);
     layer2_out[10853] <= ~layer1_out[11785] | layer1_out[11784];
     layer2_out[10854] <= layer1_out[419];
     layer2_out[10855] <= ~layer1_out[8074];
     layer2_out[10856] <= ~(layer1_out[11667] | layer1_out[11668]);
     layer2_out[10857] <= layer1_out[8503] & ~layer1_out[8502];
     layer2_out[10858] <= layer1_out[1983] | layer1_out[1984];
     layer2_out[10859] <= layer1_out[9944];
     layer2_out[10860] <= layer1_out[10270];
     layer2_out[10861] <= ~layer1_out[3699];
     layer2_out[10862] <= ~layer1_out[108];
     layer2_out[10863] <= ~layer1_out[3866] | layer1_out[3865];
     layer2_out[10864] <= ~layer1_out[7166] | layer1_out[7167];
     layer2_out[10865] <= ~layer1_out[11509] | layer1_out[11510];
     layer2_out[10866] <= ~layer1_out[2334] | layer1_out[2335];
     layer2_out[10867] <= ~layer1_out[5741];
     layer2_out[10868] <= layer1_out[8298] & ~layer1_out[8299];
     layer2_out[10869] <= layer1_out[650] & ~layer1_out[649];
     layer2_out[10870] <= layer1_out[7745] & ~layer1_out[7744];
     layer2_out[10871] <= ~layer1_out[5655];
     layer2_out[10872] <= layer1_out[1754] & ~layer1_out[1753];
     layer2_out[10873] <= ~layer1_out[142] | layer1_out[143];
     layer2_out[10874] <= layer1_out[1083];
     layer2_out[10875] <= ~layer1_out[3748] | layer1_out[3747];
     layer2_out[10876] <= ~layer1_out[1403];
     layer2_out[10877] <= ~layer1_out[981] | layer1_out[982];
     layer2_out[10878] <= layer1_out[1453];
     layer2_out[10879] <= ~(layer1_out[6763] & layer1_out[6764]);
     layer2_out[10880] <= ~layer1_out[1032];
     layer2_out[10881] <= layer1_out[9782] & ~layer1_out[9781];
     layer2_out[10882] <= ~layer1_out[1384];
     layer2_out[10883] <= layer1_out[485] & ~layer1_out[484];
     layer2_out[10884] <= layer1_out[5817] | layer1_out[5818];
     layer2_out[10885] <= ~(layer1_out[3411] ^ layer1_out[3412]);
     layer2_out[10886] <= ~(layer1_out[4665] & layer1_out[4666]);
     layer2_out[10887] <= layer1_out[6666];
     layer2_out[10888] <= ~(layer1_out[7876] | layer1_out[7877]);
     layer2_out[10889] <= layer1_out[6740] ^ layer1_out[6741];
     layer2_out[10890] <= ~layer1_out[6963];
     layer2_out[10891] <= layer1_out[6678];
     layer2_out[10892] <= layer1_out[5823];
     layer2_out[10893] <= ~(layer1_out[2920] ^ layer1_out[2921]);
     layer2_out[10894] <= layer1_out[5786];
     layer2_out[10895] <= ~(layer1_out[1604] ^ layer1_out[1605]);
     layer2_out[10896] <= ~layer1_out[6395];
     layer2_out[10897] <= ~(layer1_out[5413] ^ layer1_out[5414]);
     layer2_out[10898] <= layer1_out[9515];
     layer2_out[10899] <= ~(layer1_out[11357] | layer1_out[11358]);
     layer2_out[10900] <= ~(layer1_out[11843] & layer1_out[11844]);
     layer2_out[10901] <= ~(layer1_out[4589] & layer1_out[4590]);
     layer2_out[10902] <= ~layer1_out[6097];
     layer2_out[10903] <= ~layer1_out[3297];
     layer2_out[10904] <= ~layer1_out[4820] | layer1_out[4819];
     layer2_out[10905] <= layer1_out[10004] & ~layer1_out[10003];
     layer2_out[10906] <= ~(layer1_out[11799] | layer1_out[11800]);
     layer2_out[10907] <= ~(layer1_out[7227] | layer1_out[7228]);
     layer2_out[10908] <= ~(layer1_out[10087] | layer1_out[10088]);
     layer2_out[10909] <= layer1_out[8319] & ~layer1_out[8318];
     layer2_out[10910] <= ~(layer1_out[8811] | layer1_out[8812]);
     layer2_out[10911] <= layer1_out[5558] | layer1_out[5559];
     layer2_out[10912] <= layer1_out[11495] ^ layer1_out[11496];
     layer2_out[10913] <= layer1_out[11401] & ~layer1_out[11402];
     layer2_out[10914] <= ~(layer1_out[7426] | layer1_out[7427]);
     layer2_out[10915] <= ~(layer1_out[9050] | layer1_out[9051]);
     layer2_out[10916] <= layer1_out[6889] | layer1_out[6890];
     layer2_out[10917] <= ~layer1_out[326];
     layer2_out[10918] <= layer1_out[7863] & ~layer1_out[7862];
     layer2_out[10919] <= ~(layer1_out[101] & layer1_out[102]);
     layer2_out[10920] <= ~(layer1_out[5083] ^ layer1_out[5084]);
     layer2_out[10921] <= ~layer1_out[1676];
     layer2_out[10922] <= ~layer1_out[8764];
     layer2_out[10923] <= ~layer1_out[9586] | layer1_out[9587];
     layer2_out[10924] <= layer1_out[9455];
     layer2_out[10925] <= layer1_out[9489] & layer1_out[9490];
     layer2_out[10926] <= ~(layer1_out[6881] | layer1_out[6882]);
     layer2_out[10927] <= layer1_out[10886] | layer1_out[10887];
     layer2_out[10928] <= layer1_out[6321] & ~layer1_out[6322];
     layer2_out[10929] <= ~layer1_out[6915];
     layer2_out[10930] <= ~layer1_out[2001];
     layer2_out[10931] <= layer1_out[4393];
     layer2_out[10932] <= 1'b1;
     layer2_out[10933] <= ~layer1_out[9000];
     layer2_out[10934] <= layer1_out[10643];
     layer2_out[10935] <= layer1_out[898] ^ layer1_out[899];
     layer2_out[10936] <= layer1_out[7916];
     layer2_out[10937] <= layer1_out[11057] ^ layer1_out[11058];
     layer2_out[10938] <= ~(layer1_out[1611] & layer1_out[1612]);
     layer2_out[10939] <= ~layer1_out[1086];
     layer2_out[10940] <= layer1_out[6470] & layer1_out[6471];
     layer2_out[10941] <= layer1_out[5144];
     layer2_out[10942] <= ~(layer1_out[7463] ^ layer1_out[7464]);
     layer2_out[10943] <= ~layer1_out[6635];
     layer2_out[10944] <= layer1_out[9760] & layer1_out[9761];
     layer2_out[10945] <= layer1_out[9824] & ~layer1_out[9823];
     layer2_out[10946] <= ~(layer1_out[849] & layer1_out[850]);
     layer2_out[10947] <= layer1_out[5354] & ~layer1_out[5355];
     layer2_out[10948] <= layer1_out[3602];
     layer2_out[10949] <= layer1_out[5664];
     layer2_out[10950] <= layer1_out[9461];
     layer2_out[10951] <= ~layer1_out[7724];
     layer2_out[10952] <= layer1_out[1800];
     layer2_out[10953] <= layer1_out[3855] & ~layer1_out[3854];
     layer2_out[10954] <= ~layer1_out[8927];
     layer2_out[10955] <= ~(layer1_out[8164] | layer1_out[8165]);
     layer2_out[10956] <= ~(layer1_out[4335] | layer1_out[4336]);
     layer2_out[10957] <= layer1_out[11518];
     layer2_out[10958] <= ~layer1_out[8346] | layer1_out[8347];
     layer2_out[10959] <= ~(layer1_out[11507] ^ layer1_out[11508]);
     layer2_out[10960] <= layer1_out[2919] ^ layer1_out[2920];
     layer2_out[10961] <= ~layer1_out[669] | layer1_out[670];
     layer2_out[10962] <= layer1_out[11984] & ~layer1_out[11983];
     layer2_out[10963] <= ~layer1_out[1034];
     layer2_out[10964] <= layer1_out[5834] ^ layer1_out[5835];
     layer2_out[10965] <= layer1_out[2504] & ~layer1_out[2503];
     layer2_out[10966] <= ~layer1_out[10491];
     layer2_out[10967] <= layer1_out[9289] & ~layer1_out[9290];
     layer2_out[10968] <= ~layer1_out[10391];
     layer2_out[10969] <= ~(layer1_out[4553] & layer1_out[4554]);
     layer2_out[10970] <= ~layer1_out[4352];
     layer2_out[10971] <= layer1_out[3772] & ~layer1_out[3771];
     layer2_out[10972] <= ~layer1_out[7766];
     layer2_out[10973] <= layer1_out[7018];
     layer2_out[10974] <= layer1_out[5329] & ~layer1_out[5328];
     layer2_out[10975] <= ~layer1_out[11858];
     layer2_out[10976] <= ~(layer1_out[3835] ^ layer1_out[3836]);
     layer2_out[10977] <= ~layer1_out[11946];
     layer2_out[10978] <= ~layer1_out[2025];
     layer2_out[10979] <= ~layer1_out[6864] | layer1_out[6863];
     layer2_out[10980] <= layer1_out[11910];
     layer2_out[10981] <= ~(layer1_out[8846] | layer1_out[8847]);
     layer2_out[10982] <= ~layer1_out[2878] | layer1_out[2879];
     layer2_out[10983] <= ~(layer1_out[7030] | layer1_out[7031]);
     layer2_out[10984] <= ~(layer1_out[6068] & layer1_out[6069]);
     layer2_out[10985] <= ~layer1_out[2047] | layer1_out[2048];
     layer2_out[10986] <= ~layer1_out[9020] | layer1_out[9021];
     layer2_out[10987] <= ~layer1_out[7636] | layer1_out[7637];
     layer2_out[10988] <= layer1_out[151];
     layer2_out[10989] <= layer1_out[10685] & ~layer1_out[10686];
     layer2_out[10990] <= ~layer1_out[1358] | layer1_out[1359];
     layer2_out[10991] <= ~layer1_out[2556] | layer1_out[2557];
     layer2_out[10992] <= ~(layer1_out[2239] | layer1_out[2240]);
     layer2_out[10993] <= ~layer1_out[1421];
     layer2_out[10994] <= ~layer1_out[3490] | layer1_out[3489];
     layer2_out[10995] <= layer1_out[612];
     layer2_out[10996] <= ~layer1_out[7062];
     layer2_out[10997] <= ~layer1_out[5445];
     layer2_out[10998] <= layer1_out[4736];
     layer2_out[10999] <= layer1_out[11779] & layer1_out[11780];
     layer2_out[11000] <= layer1_out[1882] ^ layer1_out[1883];
     layer2_out[11001] <= ~layer1_out[3054];
     layer2_out[11002] <= ~(layer1_out[10118] ^ layer1_out[10119]);
     layer2_out[11003] <= layer1_out[4395];
     layer2_out[11004] <= layer1_out[518];
     layer2_out[11005] <= layer1_out[2783] & layer1_out[2784];
     layer2_out[11006] <= layer1_out[8247] & layer1_out[8248];
     layer2_out[11007] <= ~layer1_out[11351] | layer1_out[11350];
     layer2_out[11008] <= layer1_out[7201] | layer1_out[7202];
     layer2_out[11009] <= layer1_out[1255] & ~layer1_out[1254];
     layer2_out[11010] <= ~(layer1_out[9765] & layer1_out[9766]);
     layer2_out[11011] <= ~(layer1_out[10206] | layer1_out[10207]);
     layer2_out[11012] <= ~(layer1_out[8696] ^ layer1_out[8697]);
     layer2_out[11013] <= layer1_out[5712] & layer1_out[5713];
     layer2_out[11014] <= layer1_out[5045] ^ layer1_out[5046];
     layer2_out[11015] <= layer1_out[8489] & layer1_out[8490];
     layer2_out[11016] <= layer1_out[5908] | layer1_out[5909];
     layer2_out[11017] <= layer1_out[7944] & ~layer1_out[7945];
     layer2_out[11018] <= layer1_out[6164];
     layer2_out[11019] <= ~layer1_out[10214] | layer1_out[10215];
     layer2_out[11020] <= layer1_out[9602] ^ layer1_out[9603];
     layer2_out[11021] <= layer1_out[2726];
     layer2_out[11022] <= ~layer1_out[3841] | layer1_out[3840];
     layer2_out[11023] <= ~layer1_out[11117];
     layer2_out[11024] <= layer1_out[3429] ^ layer1_out[3430];
     layer2_out[11025] <= layer1_out[9549] & ~layer1_out[9550];
     layer2_out[11026] <= ~(layer1_out[7652] & layer1_out[7653]);
     layer2_out[11027] <= layer1_out[9084];
     layer2_out[11028] <= layer1_out[11748] | layer1_out[11749];
     layer2_out[11029] <= layer1_out[4101];
     layer2_out[11030] <= layer1_out[3711];
     layer2_out[11031] <= layer1_out[5479] & ~layer1_out[5478];
     layer2_out[11032] <= layer1_out[5672] | layer1_out[5673];
     layer2_out[11033] <= layer1_out[4265] | layer1_out[4266];
     layer2_out[11034] <= layer1_out[6116] & ~layer1_out[6115];
     layer2_out[11035] <= layer1_out[809] & ~layer1_out[810];
     layer2_out[11036] <= ~layer1_out[9740];
     layer2_out[11037] <= ~layer1_out[2688] | layer1_out[2687];
     layer2_out[11038] <= layer1_out[9651] & ~layer1_out[9650];
     layer2_out[11039] <= layer1_out[7813] & ~layer1_out[7812];
     layer2_out[11040] <= ~layer1_out[8933];
     layer2_out[11041] <= 1'b1;
     layer2_out[11042] <= layer1_out[7192] & ~layer1_out[7191];
     layer2_out[11043] <= layer1_out[5604] | layer1_out[5605];
     layer2_out[11044] <= layer1_out[5296] & ~layer1_out[5295];
     layer2_out[11045] <= layer1_out[11490];
     layer2_out[11046] <= ~layer1_out[11373] | layer1_out[11372];
     layer2_out[11047] <= layer1_out[8728] ^ layer1_out[8729];
     layer2_out[11048] <= ~(layer1_out[1873] & layer1_out[1874]);
     layer2_out[11049] <= layer1_out[1459] & ~layer1_out[1458];
     layer2_out[11050] <= ~layer1_out[8167];
     layer2_out[11051] <= ~layer1_out[1198];
     layer2_out[11052] <= layer1_out[1603] & layer1_out[1604];
     layer2_out[11053] <= 1'b0;
     layer2_out[11054] <= 1'b1;
     layer2_out[11055] <= ~(layer1_out[2717] | layer1_out[2718]);
     layer2_out[11056] <= layer1_out[3934];
     layer2_out[11057] <= layer1_out[10154];
     layer2_out[11058] <= layer1_out[9267] & ~layer1_out[9266];
     layer2_out[11059] <= layer1_out[1965] & ~layer1_out[1966];
     layer2_out[11060] <= ~layer1_out[11839];
     layer2_out[11061] <= ~layer1_out[6835];
     layer2_out[11062] <= ~layer1_out[4620];
     layer2_out[11063] <= layer1_out[9293] | layer1_out[9294];
     layer2_out[11064] <= ~layer1_out[7434] | layer1_out[7433];
     layer2_out[11065] <= layer1_out[4901] & layer1_out[4902];
     layer2_out[11066] <= ~layer1_out[6371] | layer1_out[6370];
     layer2_out[11067] <= layer1_out[1648] & layer1_out[1649];
     layer2_out[11068] <= layer1_out[4684] & ~layer1_out[4683];
     layer2_out[11069] <= layer1_out[1970] & ~layer1_out[1969];
     layer2_out[11070] <= layer1_out[5323] ^ layer1_out[5324];
     layer2_out[11071] <= layer1_out[9771] | layer1_out[9772];
     layer2_out[11072] <= layer1_out[11587] | layer1_out[11588];
     layer2_out[11073] <= layer1_out[9093] | layer1_out[9094];
     layer2_out[11074] <= ~(layer1_out[10605] | layer1_out[10606]);
     layer2_out[11075] <= layer1_out[11005];
     layer2_out[11076] <= layer1_out[2330] | layer1_out[2331];
     layer2_out[11077] <= ~layer1_out[2695] | layer1_out[2696];
     layer2_out[11078] <= layer1_out[2230] & layer1_out[2231];
     layer2_out[11079] <= layer1_out[9225] & layer1_out[9226];
     layer2_out[11080] <= layer1_out[5895] | layer1_out[5896];
     layer2_out[11081] <= ~(layer1_out[8449] & layer1_out[8450]);
     layer2_out[11082] <= ~layer1_out[11024] | layer1_out[11025];
     layer2_out[11083] <= ~(layer1_out[10988] | layer1_out[10989]);
     layer2_out[11084] <= ~(layer1_out[7793] & layer1_out[7794]);
     layer2_out[11085] <= layer1_out[11374];
     layer2_out[11086] <= layer1_out[2294] ^ layer1_out[2295];
     layer2_out[11087] <= ~(layer1_out[9191] ^ layer1_out[9192]);
     layer2_out[11088] <= ~layer1_out[3148];
     layer2_out[11089] <= layer1_out[6463];
     layer2_out[11090] <= layer1_out[8944] & layer1_out[8945];
     layer2_out[11091] <= layer1_out[3515];
     layer2_out[11092] <= ~layer1_out[7934];
     layer2_out[11093] <= ~layer1_out[5885];
     layer2_out[11094] <= ~layer1_out[713];
     layer2_out[11095] <= layer1_out[7527] & layer1_out[7528];
     layer2_out[11096] <= layer1_out[549];
     layer2_out[11097] <= layer1_out[3104];
     layer2_out[11098] <= ~layer1_out[7830] | layer1_out[7831];
     layer2_out[11099] <= layer1_out[4049] | layer1_out[4050];
     layer2_out[11100] <= layer1_out[1730];
     layer2_out[11101] <= 1'b0;
     layer2_out[11102] <= layer1_out[7459];
     layer2_out[11103] <= layer1_out[7215] | layer1_out[7216];
     layer2_out[11104] <= layer1_out[2776] & layer1_out[2777];
     layer2_out[11105] <= ~(layer1_out[6202] & layer1_out[6203]);
     layer2_out[11106] <= layer1_out[11663] | layer1_out[11664];
     layer2_out[11107] <= layer1_out[9487];
     layer2_out[11108] <= layer1_out[9450] | layer1_out[9451];
     layer2_out[11109] <= layer1_out[6027];
     layer2_out[11110] <= ~layer1_out[5235];
     layer2_out[11111] <= layer1_out[3539] & ~layer1_out[3538];
     layer2_out[11112] <= layer1_out[1669];
     layer2_out[11113] <= layer1_out[9264] ^ layer1_out[9265];
     layer2_out[11114] <= layer1_out[9690] & layer1_out[9691];
     layer2_out[11115] <= layer1_out[11547] ^ layer1_out[11548];
     layer2_out[11116] <= layer1_out[2515];
     layer2_out[11117] <= ~layer1_out[8722] | layer1_out[8721];
     layer2_out[11118] <= ~layer1_out[4331];
     layer2_out[11119] <= layer1_out[2486];
     layer2_out[11120] <= layer1_out[11552] & ~layer1_out[11551];
     layer2_out[11121] <= ~(layer1_out[3535] ^ layer1_out[3536]);
     layer2_out[11122] <= ~layer1_out[3399];
     layer2_out[11123] <= layer1_out[49] & layer1_out[50];
     layer2_out[11124] <= ~(layer1_out[7615] ^ layer1_out[7616]);
     layer2_out[11125] <= layer1_out[1424];
     layer2_out[11126] <= layer1_out[9798] ^ layer1_out[9799];
     layer2_out[11127] <= layer1_out[9800] ^ layer1_out[9801];
     layer2_out[11128] <= layer1_out[9978] | layer1_out[9979];
     layer2_out[11129] <= ~layer1_out[882];
     layer2_out[11130] <= ~(layer1_out[4710] ^ layer1_out[4711]);
     layer2_out[11131] <= layer1_out[8745] | layer1_out[8746];
     layer2_out[11132] <= layer1_out[8576] & ~layer1_out[8575];
     layer2_out[11133] <= layer1_out[2947] & ~layer1_out[2948];
     layer2_out[11134] <= layer1_out[3861] & layer1_out[3862];
     layer2_out[11135] <= ~layer1_out[10880] | layer1_out[10879];
     layer2_out[11136] <= ~layer1_out[653] | layer1_out[652];
     layer2_out[11137] <= layer1_out[4529];
     layer2_out[11138] <= layer1_out[6430];
     layer2_out[11139] <= layer1_out[3270];
     layer2_out[11140] <= layer1_out[1358] & ~layer1_out[1357];
     layer2_out[11141] <= ~(layer1_out[1741] ^ layer1_out[1742]);
     layer2_out[11142] <= ~layer1_out[1488] | layer1_out[1489];
     layer2_out[11143] <= ~layer1_out[6785] | layer1_out[6784];
     layer2_out[11144] <= layer1_out[547];
     layer2_out[11145] <= layer1_out[1560];
     layer2_out[11146] <= layer1_out[7685] & ~layer1_out[7684];
     layer2_out[11147] <= layer1_out[5940] | layer1_out[5941];
     layer2_out[11148] <= layer1_out[2575] ^ layer1_out[2576];
     layer2_out[11149] <= ~layer1_out[7953];
     layer2_out[11150] <= layer1_out[6359];
     layer2_out[11151] <= ~layer1_out[6249];
     layer2_out[11152] <= ~layer1_out[862];
     layer2_out[11153] <= layer1_out[4421];
     layer2_out[11154] <= layer1_out[8123];
     layer2_out[11155] <= layer1_out[7021] & ~layer1_out[7020];
     layer2_out[11156] <= layer1_out[2];
     layer2_out[11157] <= ~layer1_out[1586];
     layer2_out[11158] <= layer1_out[4432];
     layer2_out[11159] <= layer1_out[3470];
     layer2_out[11160] <= ~layer1_out[4686];
     layer2_out[11161] <= layer1_out[10626] | layer1_out[10627];
     layer2_out[11162] <= ~layer1_out[3594] | layer1_out[3593];
     layer2_out[11163] <= layer1_out[3794] & ~layer1_out[3795];
     layer2_out[11164] <= layer1_out[7100];
     layer2_out[11165] <= 1'b0;
     layer2_out[11166] <= ~layer1_out[4502] | layer1_out[4501];
     layer2_out[11167] <= layer1_out[8309] & layer1_out[8310];
     layer2_out[11168] <= ~layer1_out[11624] | layer1_out[11623];
     layer2_out[11169] <= layer1_out[2199] & ~layer1_out[2198];
     layer2_out[11170] <= ~(layer1_out[6148] & layer1_out[6149]);
     layer2_out[11171] <= layer1_out[6852];
     layer2_out[11172] <= ~layer1_out[4842];
     layer2_out[11173] <= ~layer1_out[4611];
     layer2_out[11174] <= layer1_out[8064] | layer1_out[8065];
     layer2_out[11175] <= layer1_out[9235] | layer1_out[9236];
     layer2_out[11176] <= layer1_out[400] & layer1_out[401];
     layer2_out[11177] <= layer1_out[8535] | layer1_out[8536];
     layer2_out[11178] <= ~layer1_out[10755] | layer1_out[10754];
     layer2_out[11179] <= layer1_out[4197];
     layer2_out[11180] <= layer1_out[6368] & ~layer1_out[6367];
     layer2_out[11181] <= ~layer1_out[2618];
     layer2_out[11182] <= layer1_out[4158] & ~layer1_out[4157];
     layer2_out[11183] <= ~layer1_out[9257] | layer1_out[9258];
     layer2_out[11184] <= ~layer1_out[4867];
     layer2_out[11185] <= ~(layer1_out[2071] & layer1_out[2072]);
     layer2_out[11186] <= layer1_out[8524] | layer1_out[8525];
     layer2_out[11187] <= ~(layer1_out[10772] & layer1_out[10773]);
     layer2_out[11188] <= ~layer1_out[7744];
     layer2_out[11189] <= layer1_out[3407] | layer1_out[3408];
     layer2_out[11190] <= ~layer1_out[2308];
     layer2_out[11191] <= layer1_out[4641] | layer1_out[4642];
     layer2_out[11192] <= layer1_out[805] ^ layer1_out[806];
     layer2_out[11193] <= ~(layer1_out[3972] & layer1_out[3973]);
     layer2_out[11194] <= layer1_out[3787];
     layer2_out[11195] <= layer1_out[10377] & ~layer1_out[10376];
     layer2_out[11196] <= ~layer1_out[1854];
     layer2_out[11197] <= layer1_out[11153] & ~layer1_out[11154];
     layer2_out[11198] <= ~layer1_out[3737];
     layer2_out[11199] <= ~(layer1_out[4731] ^ layer1_out[4732]);
     layer2_out[11200] <= ~layer1_out[3595];
     layer2_out[11201] <= layer1_out[9634] ^ layer1_out[9635];
     layer2_out[11202] <= ~layer1_out[1682];
     layer2_out[11203] <= layer1_out[2054] | layer1_out[2055];
     layer2_out[11204] <= layer1_out[4843];
     layer2_out[11205] <= ~layer1_out[3554];
     layer2_out[11206] <= layer1_out[3551] & ~layer1_out[3552];
     layer2_out[11207] <= ~(layer1_out[1496] ^ layer1_out[1497]);
     layer2_out[11208] <= layer1_out[3523];
     layer2_out[11209] <= layer1_out[4172];
     layer2_out[11210] <= ~(layer1_out[8634] & layer1_out[8635]);
     layer2_out[11211] <= layer1_out[547] & layer1_out[548];
     layer2_out[11212] <= layer1_out[6791] & layer1_out[6792];
     layer2_out[11213] <= ~(layer1_out[11944] ^ layer1_out[11945]);
     layer2_out[11214] <= ~layer1_out[3692];
     layer2_out[11215] <= ~(layer1_out[11850] | layer1_out[11851]);
     layer2_out[11216] <= ~layer1_out[871];
     layer2_out[11217] <= layer1_out[7961] & ~layer1_out[7962];
     layer2_out[11218] <= layer1_out[4264] & ~layer1_out[4263];
     layer2_out[11219] <= layer1_out[4919];
     layer2_out[11220] <= layer1_out[3860] & ~layer1_out[3859];
     layer2_out[11221] <= layer1_out[2089] | layer1_out[2090];
     layer2_out[11222] <= ~(layer1_out[10877] & layer1_out[10878]);
     layer2_out[11223] <= layer1_out[2546];
     layer2_out[11224] <= layer1_out[11002] | layer1_out[11003];
     layer2_out[11225] <= 1'b0;
     layer2_out[11226] <= ~layer1_out[7299] | layer1_out[7300];
     layer2_out[11227] <= layer1_out[3550];
     layer2_out[11228] <= layer1_out[1151];
     layer2_out[11229] <= ~(layer1_out[2603] & layer1_out[2604]);
     layer2_out[11230] <= layer1_out[27] & layer1_out[28];
     layer2_out[11231] <= ~layer1_out[8929] | layer1_out[8928];
     layer2_out[11232] <= ~(layer1_out[9358] | layer1_out[9359]);
     layer2_out[11233] <= layer1_out[5395];
     layer2_out[11234] <= layer1_out[3822];
     layer2_out[11235] <= ~(layer1_out[2552] | layer1_out[2553]);
     layer2_out[11236] <= layer1_out[5783] | layer1_out[5784];
     layer2_out[11237] <= layer1_out[2238] & ~layer1_out[2237];
     layer2_out[11238] <= ~layer1_out[9745];
     layer2_out[11239] <= ~layer1_out[756] | layer1_out[755];
     layer2_out[11240] <= layer1_out[5824] & layer1_out[5825];
     layer2_out[11241] <= layer1_out[756] & ~layer1_out[757];
     layer2_out[11242] <= layer1_out[5935] ^ layer1_out[5936];
     layer2_out[11243] <= 1'b1;
     layer2_out[11244] <= layer1_out[9178] & layer1_out[9179];
     layer2_out[11245] <= ~layer1_out[9742];
     layer2_out[11246] <= layer1_out[1984] | layer1_out[1985];
     layer2_out[11247] <= layer1_out[3887] & layer1_out[3888];
     layer2_out[11248] <= layer1_out[2008];
     layer2_out[11249] <= ~(layer1_out[2269] | layer1_out[2270]);
     layer2_out[11250] <= ~layer1_out[8593] | layer1_out[8592];
     layer2_out[11251] <= layer1_out[2885] & layer1_out[2886];
     layer2_out[11252] <= layer1_out[4285];
     layer2_out[11253] <= layer1_out[5863];
     layer2_out[11254] <= layer1_out[9369];
     layer2_out[11255] <= layer1_out[1388];
     layer2_out[11256] <= layer1_out[2454];
     layer2_out[11257] <= ~layer1_out[4388] | layer1_out[4387];
     layer2_out[11258] <= ~layer1_out[1577];
     layer2_out[11259] <= layer1_out[3945];
     layer2_out[11260] <= layer1_out[7254];
     layer2_out[11261] <= ~(layer1_out[9075] | layer1_out[9076]);
     layer2_out[11262] <= ~layer1_out[8306];
     layer2_out[11263] <= ~layer1_out[677];
     layer2_out[11264] <= ~layer1_out[10119];
     layer2_out[11265] <= layer1_out[1876] ^ layer1_out[1877];
     layer2_out[11266] <= ~(layer1_out[7472] ^ layer1_out[7473]);
     layer2_out[11267] <= ~layer1_out[7517] | layer1_out[7518];
     layer2_out[11268] <= ~(layer1_out[2690] | layer1_out[2691]);
     layer2_out[11269] <= layer1_out[9988] & ~layer1_out[9987];
     layer2_out[11270] <= ~(layer1_out[994] & layer1_out[995]);
     layer2_out[11271] <= ~layer1_out[5725];
     layer2_out[11272] <= layer1_out[10822] & ~layer1_out[10821];
     layer2_out[11273] <= layer1_out[3871] & ~layer1_out[3870];
     layer2_out[11274] <= ~layer1_out[7330] | layer1_out[7329];
     layer2_out[11275] <= layer1_out[5274] ^ layer1_out[5275];
     layer2_out[11276] <= ~(layer1_out[10746] & layer1_out[10747]);
     layer2_out[11277] <= layer1_out[761];
     layer2_out[11278] <= layer1_out[2143] & ~layer1_out[2142];
     layer2_out[11279] <= layer1_out[5854] & ~layer1_out[5853];
     layer2_out[11280] <= layer1_out[8715];
     layer2_out[11281] <= ~layer1_out[6743];
     layer2_out[11282] <= layer1_out[10910] | layer1_out[10911];
     layer2_out[11283] <= ~(layer1_out[10383] | layer1_out[10384]);
     layer2_out[11284] <= layer1_out[1275] | layer1_out[1276];
     layer2_out[11285] <= layer1_out[112];
     layer2_out[11286] <= ~(layer1_out[9354] | layer1_out[9355]);
     layer2_out[11287] <= layer1_out[1093];
     layer2_out[11288] <= layer1_out[3074];
     layer2_out[11289] <= ~layer1_out[687];
     layer2_out[11290] <= layer1_out[9704];
     layer2_out[11291] <= ~(layer1_out[8453] | layer1_out[8454]);
     layer2_out[11292] <= ~layer1_out[7963];
     layer2_out[11293] <= layer1_out[5069] & ~layer1_out[5068];
     layer2_out[11294] <= 1'b1;
     layer2_out[11295] <= ~layer1_out[10698];
     layer2_out[11296] <= ~layer1_out[4597];
     layer2_out[11297] <= layer1_out[3911] & ~layer1_out[3910];
     layer2_out[11298] <= layer1_out[9379];
     layer2_out[11299] <= layer1_out[9971];
     layer2_out[11300] <= layer1_out[2374];
     layer2_out[11301] <= ~layer1_out[4172] | layer1_out[4173];
     layer2_out[11302] <= ~(layer1_out[10466] & layer1_out[10467]);
     layer2_out[11303] <= ~layer1_out[7364];
     layer2_out[11304] <= layer1_out[5583] & layer1_out[5584];
     layer2_out[11305] <= ~layer1_out[9986];
     layer2_out[11306] <= layer1_out[3563] & ~layer1_out[3562];
     layer2_out[11307] <= ~layer1_out[952];
     layer2_out[11308] <= layer1_out[10110] | layer1_out[10111];
     layer2_out[11309] <= ~layer1_out[8655] | layer1_out[8656];
     layer2_out[11310] <= ~layer1_out[185];
     layer2_out[11311] <= layer1_out[3341] ^ layer1_out[3342];
     layer2_out[11312] <= ~layer1_out[10024];
     layer2_out[11313] <= layer1_out[7158] & ~layer1_out[7159];
     layer2_out[11314] <= ~(layer1_out[9897] ^ layer1_out[9898]);
     layer2_out[11315] <= ~layer1_out[6615];
     layer2_out[11316] <= layer1_out[6489];
     layer2_out[11317] <= layer1_out[8935];
     layer2_out[11318] <= ~(layer1_out[3010] | layer1_out[3011]);
     layer2_out[11319] <= layer1_out[11884];
     layer2_out[11320] <= ~(layer1_out[2566] & layer1_out[2567]);
     layer2_out[11321] <= layer1_out[3431];
     layer2_out[11322] <= layer1_out[3721];
     layer2_out[11323] <= layer1_out[444];
     layer2_out[11324] <= layer1_out[9683] & ~layer1_out[9682];
     layer2_out[11325] <= layer1_out[5672];
     layer2_out[11326] <= layer1_out[3631];
     layer2_out[11327] <= ~(layer1_out[2357] | layer1_out[2358]);
     layer2_out[11328] <= ~(layer1_out[3327] | layer1_out[3328]);
     layer2_out[11329] <= ~layer1_out[5671];
     layer2_out[11330] <= ~layer1_out[126];
     layer2_out[11331] <= layer1_out[4153];
     layer2_out[11332] <= ~layer1_out[7806];
     layer2_out[11333] <= layer1_out[8588] & layer1_out[8589];
     layer2_out[11334] <= ~(layer1_out[6320] | layer1_out[6321]);
     layer2_out[11335] <= layer1_out[2388] & ~layer1_out[2387];
     layer2_out[11336] <= layer1_out[3504] & ~layer1_out[3505];
     layer2_out[11337] <= layer1_out[11116] & layer1_out[11117];
     layer2_out[11338] <= layer1_out[9635] | layer1_out[9636];
     layer2_out[11339] <= layer1_out[2424];
     layer2_out[11340] <= layer1_out[10432] | layer1_out[10433];
     layer2_out[11341] <= ~(layer1_out[6566] | layer1_out[6567]);
     layer2_out[11342] <= ~(layer1_out[4094] & layer1_out[4095]);
     layer2_out[11343] <= ~(layer1_out[415] ^ layer1_out[416]);
     layer2_out[11344] <= ~layer1_out[3154] | layer1_out[3155];
     layer2_out[11345] <= layer1_out[8053];
     layer2_out[11346] <= layer1_out[58] & ~layer1_out[57];
     layer2_out[11347] <= layer1_out[8423] ^ layer1_out[8424];
     layer2_out[11348] <= ~layer1_out[8536];
     layer2_out[11349] <= ~layer1_out[8089];
     layer2_out[11350] <= ~layer1_out[614];
     layer2_out[11351] <= ~layer1_out[5989];
     layer2_out[11352] <= layer1_out[6929] & layer1_out[6930];
     layer2_out[11353] <= layer1_out[1323];
     layer2_out[11354] <= layer1_out[6770] ^ layer1_out[6771];
     layer2_out[11355] <= layer1_out[75] | layer1_out[76];
     layer2_out[11356] <= ~(layer1_out[8113] ^ layer1_out[8114]);
     layer2_out[11357] <= layer1_out[11560] | layer1_out[11561];
     layer2_out[11358] <= ~layer1_out[347];
     layer2_out[11359] <= layer1_out[5446];
     layer2_out[11360] <= layer1_out[862];
     layer2_out[11361] <= ~layer1_out[10363];
     layer2_out[11362] <= ~layer1_out[7170];
     layer2_out[11363] <= layer1_out[2623] & ~layer1_out[2622];
     layer2_out[11364] <= layer1_out[2507];
     layer2_out[11365] <= ~(layer1_out[5923] & layer1_out[5924]);
     layer2_out[11366] <= ~(layer1_out[9101] | layer1_out[9102]);
     layer2_out[11367] <= ~layer1_out[7252];
     layer2_out[11368] <= layer1_out[3076];
     layer2_out[11369] <= ~layer1_out[9876];
     layer2_out[11370] <= ~layer1_out[5619];
     layer2_out[11371] <= layer1_out[8055];
     layer2_out[11372] <= layer1_out[5803];
     layer2_out[11373] <= ~layer1_out[7623] | layer1_out[7624];
     layer2_out[11374] <= layer1_out[10730] & ~layer1_out[10731];
     layer2_out[11375] <= ~layer1_out[9421];
     layer2_out[11376] <= layer1_out[4531] & layer1_out[4532];
     layer2_out[11377] <= ~layer1_out[3496];
     layer2_out[11378] <= ~layer1_out[3573];
     layer2_out[11379] <= ~(layer1_out[585] ^ layer1_out[586]);
     layer2_out[11380] <= layer1_out[739] & ~layer1_out[738];
     layer2_out[11381] <= ~layer1_out[8633];
     layer2_out[11382] <= layer1_out[5856] & ~layer1_out[5857];
     layer2_out[11383] <= ~layer1_out[10464] | layer1_out[10463];
     layer2_out[11384] <= ~layer1_out[7339];
     layer2_out[11385] <= ~layer1_out[6947] | layer1_out[6948];
     layer2_out[11386] <= layer1_out[935] | layer1_out[936];
     layer2_out[11387] <= ~layer1_out[2096];
     layer2_out[11388] <= ~layer1_out[986];
     layer2_out[11389] <= ~layer1_out[215] | layer1_out[216];
     layer2_out[11390] <= layer1_out[6956] | layer1_out[6957];
     layer2_out[11391] <= ~layer1_out[3978] | layer1_out[3977];
     layer2_out[11392] <= layer1_out[11096] ^ layer1_out[11097];
     layer2_out[11393] <= layer1_out[5128];
     layer2_out[11394] <= ~(layer1_out[4329] ^ layer1_out[4330]);
     layer2_out[11395] <= layer1_out[5505];
     layer2_out[11396] <= ~layer1_out[4846];
     layer2_out[11397] <= layer1_out[8659] & layer1_out[8660];
     layer2_out[11398] <= layer1_out[204] & ~layer1_out[205];
     layer2_out[11399] <= ~(layer1_out[11693] & layer1_out[11694]);
     layer2_out[11400] <= layer1_out[2323];
     layer2_out[11401] <= ~layer1_out[5587];
     layer2_out[11402] <= ~layer1_out[11887];
     layer2_out[11403] <= ~layer1_out[2031] | layer1_out[2030];
     layer2_out[11404] <= ~(layer1_out[8042] | layer1_out[8043]);
     layer2_out[11405] <= ~layer1_out[11043];
     layer2_out[11406] <= ~layer1_out[10665] | layer1_out[10664];
     layer2_out[11407] <= layer1_out[9474];
     layer2_out[11408] <= ~layer1_out[145] | layer1_out[146];
     layer2_out[11409] <= ~layer1_out[1062];
     layer2_out[11410] <= layer1_out[9671] & layer1_out[9672];
     layer2_out[11411] <= ~layer1_out[9568];
     layer2_out[11412] <= layer1_out[5508];
     layer2_out[11413] <= ~layer1_out[10100];
     layer2_out[11414] <= layer1_out[2802];
     layer2_out[11415] <= ~layer1_out[4468];
     layer2_out[11416] <= ~layer1_out[10854];
     layer2_out[11417] <= ~(layer1_out[11316] | layer1_out[11317]);
     layer2_out[11418] <= ~layer1_out[8433];
     layer2_out[11419] <= ~layer1_out[8947];
     layer2_out[11420] <= ~layer1_out[5070] | layer1_out[5071];
     layer2_out[11421] <= layer1_out[5327] & ~layer1_out[5328];
     layer2_out[11422] <= ~layer1_out[4097] | layer1_out[4096];
     layer2_out[11423] <= ~layer1_out[11332];
     layer2_out[11424] <= layer1_out[10232] | layer1_out[10233];
     layer2_out[11425] <= ~layer1_out[6142];
     layer2_out[11426] <= layer1_out[2941] & layer1_out[2942];
     layer2_out[11427] <= ~(layer1_out[6581] & layer1_out[6582]);
     layer2_out[11428] <= ~layer1_out[4678];
     layer2_out[11429] <= layer1_out[4162] & ~layer1_out[4163];
     layer2_out[11430] <= ~(layer1_out[7565] | layer1_out[7566]);
     layer2_out[11431] <= ~layer1_out[7420];
     layer2_out[11432] <= layer1_out[3205] ^ layer1_out[3206];
     layer2_out[11433] <= layer1_out[3517] & layer1_out[3518];
     layer2_out[11434] <= ~layer1_out[10422];
     layer2_out[11435] <= ~(layer1_out[67] | layer1_out[68]);
     layer2_out[11436] <= ~layer1_out[7161];
     layer2_out[11437] <= ~layer1_out[2172] | layer1_out[2171];
     layer2_out[11438] <= layer1_out[3001] ^ layer1_out[3002];
     layer2_out[11439] <= ~layer1_out[8153];
     layer2_out[11440] <= 1'b0;
     layer2_out[11441] <= ~(layer1_out[9562] | layer1_out[9563]);
     layer2_out[11442] <= layer1_out[1173] ^ layer1_out[1174];
     layer2_out[11443] <= ~layer1_out[6001] | layer1_out[6002];
     layer2_out[11444] <= layer1_out[9601] ^ layer1_out[9602];
     layer2_out[11445] <= ~layer1_out[1139];
     layer2_out[11446] <= layer1_out[2821];
     layer2_out[11447] <= ~layer1_out[9487];
     layer2_out[11448] <= layer1_out[3361] & layer1_out[3362];
     layer2_out[11449] <= layer1_out[11440];
     layer2_out[11450] <= layer1_out[890] ^ layer1_out[891];
     layer2_out[11451] <= ~(layer1_out[5858] | layer1_out[5859]);
     layer2_out[11452] <= ~(layer1_out[7008] ^ layer1_out[7009]);
     layer2_out[11453] <= layer1_out[10541];
     layer2_out[11454] <= layer1_out[1421] ^ layer1_out[1422];
     layer2_out[11455] <= layer1_out[3739] & layer1_out[3740];
     layer2_out[11456] <= ~(layer1_out[10647] | layer1_out[10648]);
     layer2_out[11457] <= ~layer1_out[8380] | layer1_out[8381];
     layer2_out[11458] <= layer1_out[4919] & ~layer1_out[4920];
     layer2_out[11459] <= ~layer1_out[8448] | layer1_out[8447];
     layer2_out[11460] <= ~layer1_out[9642];
     layer2_out[11461] <= layer1_out[7674];
     layer2_out[11462] <= layer1_out[10495] & ~layer1_out[10494];
     layer2_out[11463] <= layer1_out[9498] & ~layer1_out[9497];
     layer2_out[11464] <= layer1_out[7718] | layer1_out[7719];
     layer2_out[11465] <= ~(layer1_out[7779] | layer1_out[7780]);
     layer2_out[11466] <= ~(layer1_out[4391] & layer1_out[4392]);
     layer2_out[11467] <= layer1_out[10624];
     layer2_out[11468] <= layer1_out[4350] & ~layer1_out[4349];
     layer2_out[11469] <= layer1_out[6286] & ~layer1_out[6285];
     layer2_out[11470] <= layer1_out[1561] & ~layer1_out[1560];
     layer2_out[11471] <= ~layer1_out[781];
     layer2_out[11472] <= ~(layer1_out[3608] ^ layer1_out[3609]);
     layer2_out[11473] <= ~layer1_out[9330] | layer1_out[9331];
     layer2_out[11474] <= ~layer1_out[2331];
     layer2_out[11475] <= ~layer1_out[5541];
     layer2_out[11476] <= layer1_out[2342];
     layer2_out[11477] <= ~(layer1_out[10721] | layer1_out[10722]);
     layer2_out[11478] <= ~layer1_out[5907] | layer1_out[5908];
     layer2_out[11479] <= ~layer1_out[5412];
     layer2_out[11480] <= layer1_out[8925] & layer1_out[8926];
     layer2_out[11481] <= ~layer1_out[10928] | layer1_out[10929];
     layer2_out[11482] <= ~layer1_out[1309] | layer1_out[1310];
     layer2_out[11483] <= ~layer1_out[5399];
     layer2_out[11484] <= ~layer1_out[9286] | layer1_out[9285];
     layer2_out[11485] <= layer1_out[3327];
     layer2_out[11486] <= layer1_out[158] & ~layer1_out[157];
     layer2_out[11487] <= ~(layer1_out[2583] ^ layer1_out[2584]);
     layer2_out[11488] <= ~layer1_out[9570];
     layer2_out[11489] <= layer1_out[6184] ^ layer1_out[6185];
     layer2_out[11490] <= ~layer1_out[3173];
     layer2_out[11491] <= ~layer1_out[919] | layer1_out[920];
     layer2_out[11492] <= layer1_out[5203];
     layer2_out[11493] <= ~(layer1_out[2961] ^ layer1_out[2962]);
     layer2_out[11494] <= layer1_out[887];
     layer2_out[11495] <= layer1_out[2041] & layer1_out[2042];
     layer2_out[11496] <= layer1_out[8952] & ~layer1_out[8951];
     layer2_out[11497] <= layer1_out[3190] & layer1_out[3191];
     layer2_out[11498] <= layer1_out[1238];
     layer2_out[11499] <= ~layer1_out[955];
     layer2_out[11500] <= ~(layer1_out[5754] ^ layer1_out[5755]);
     layer2_out[11501] <= layer1_out[5366];
     layer2_out[11502] <= ~layer1_out[2019];
     layer2_out[11503] <= ~(layer1_out[793] ^ layer1_out[794]);
     layer2_out[11504] <= ~(layer1_out[4114] | layer1_out[4115]);
     layer2_out[11505] <= ~layer1_out[10796] | layer1_out[10795];
     layer2_out[11506] <= ~layer1_out[2313];
     layer2_out[11507] <= layer1_out[4602];
     layer2_out[11508] <= ~layer1_out[994] | layer1_out[993];
     layer2_out[11509] <= layer1_out[2860];
     layer2_out[11510] <= layer1_out[4562] & layer1_out[4563];
     layer2_out[11511] <= ~layer1_out[2554] | layer1_out[2553];
     layer2_out[11512] <= layer1_out[10127];
     layer2_out[11513] <= ~(layer1_out[1194] ^ layer1_out[1195]);
     layer2_out[11514] <= layer1_out[536] & ~layer1_out[535];
     layer2_out[11515] <= layer1_out[431] & layer1_out[432];
     layer2_out[11516] <= layer1_out[8295] & ~layer1_out[8294];
     layer2_out[11517] <= ~(layer1_out[5386] | layer1_out[5387]);
     layer2_out[11518] <= layer1_out[2422] & ~layer1_out[2421];
     layer2_out[11519] <= ~(layer1_out[1657] | layer1_out[1658]);
     layer2_out[11520] <= ~layer1_out[1592];
     layer2_out[11521] <= ~layer1_out[1754] | layer1_out[1755];
     layer2_out[11522] <= layer1_out[202] & layer1_out[203];
     layer2_out[11523] <= layer1_out[7499];
     layer2_out[11524] <= layer1_out[4131] & ~layer1_out[4132];
     layer2_out[11525] <= layer1_out[3878];
     layer2_out[11526] <= ~layer1_out[554] | layer1_out[555];
     layer2_out[11527] <= layer1_out[10769] | layer1_out[10770];
     layer2_out[11528] <= ~layer1_out[4074];
     layer2_out[11529] <= layer1_out[9327] & layer1_out[9328];
     layer2_out[11530] <= layer1_out[5661];
     layer2_out[11531] <= layer1_out[8112] & ~layer1_out[8111];
     layer2_out[11532] <= ~layer1_out[5244];
     layer2_out[11533] <= layer1_out[4767];
     layer2_out[11534] <= layer1_out[10803] | layer1_out[10804];
     layer2_out[11535] <= layer1_out[3287] & layer1_out[3288];
     layer2_out[11536] <= layer1_out[5880] ^ layer1_out[5881];
     layer2_out[11537] <= ~layer1_out[11514];
     layer2_out[11538] <= layer1_out[11015];
     layer2_out[11539] <= layer1_out[3042] ^ layer1_out[3043];
     layer2_out[11540] <= ~(layer1_out[10976] | layer1_out[10977]);
     layer2_out[11541] <= layer1_out[5154] | layer1_out[5155];
     layer2_out[11542] <= 1'b1;
     layer2_out[11543] <= ~layer1_out[1112] | layer1_out[1111];
     layer2_out[11544] <= layer1_out[1004];
     layer2_out[11545] <= layer1_out[10887];
     layer2_out[11546] <= ~(layer1_out[4414] & layer1_out[4415]);
     layer2_out[11547] <= layer1_out[11313];
     layer2_out[11548] <= layer1_out[4255] & ~layer1_out[4256];
     layer2_out[11549] <= layer1_out[4273] & ~layer1_out[4274];
     layer2_out[11550] <= ~(layer1_out[8566] & layer1_out[8567]);
     layer2_out[11551] <= layer1_out[9882] ^ layer1_out[9883];
     layer2_out[11552] <= layer1_out[11794] & ~layer1_out[11793];
     layer2_out[11553] <= ~(layer1_out[9633] | layer1_out[9634]);
     layer2_out[11554] <= layer1_out[8619] | layer1_out[8620];
     layer2_out[11555] <= ~layer1_out[3749];
     layer2_out[11556] <= layer1_out[8823];
     layer2_out[11557] <= ~layer1_out[7416];
     layer2_out[11558] <= layer1_out[311];
     layer2_out[11559] <= layer1_out[1954];
     layer2_out[11560] <= ~layer1_out[8404];
     layer2_out[11561] <= ~layer1_out[6855] | layer1_out[6856];
     layer2_out[11562] <= ~(layer1_out[10579] ^ layer1_out[10580]);
     layer2_out[11563] <= ~layer1_out[5599];
     layer2_out[11564] <= ~layer1_out[80];
     layer2_out[11565] <= ~(layer1_out[6822] | layer1_out[6823]);
     layer2_out[11566] <= ~(layer1_out[8887] ^ layer1_out[8888]);
     layer2_out[11567] <= ~layer1_out[6979] | layer1_out[6980];
     layer2_out[11568] <= ~layer1_out[7009];
     layer2_out[11569] <= ~layer1_out[7991];
     layer2_out[11570] <= ~layer1_out[403];
     layer2_out[11571] <= layer1_out[11797];
     layer2_out[11572] <= layer1_out[306] ^ layer1_out[307];
     layer2_out[11573] <= ~layer1_out[5641];
     layer2_out[11574] <= ~layer1_out[9548];
     layer2_out[11575] <= layer1_out[10512] | layer1_out[10513];
     layer2_out[11576] <= ~layer1_out[6261];
     layer2_out[11577] <= layer1_out[11752] & ~layer1_out[11751];
     layer2_out[11578] <= layer1_out[2416] | layer1_out[2417];
     layer2_out[11579] <= layer1_out[4546] | layer1_out[4547];
     layer2_out[11580] <= layer1_out[10537];
     layer2_out[11581] <= layer1_out[7371];
     layer2_out[11582] <= ~(layer1_out[3857] & layer1_out[3858]);
     layer2_out[11583] <= layer1_out[4852] | layer1_out[4853];
     layer2_out[11584] <= ~(layer1_out[619] | layer1_out[620]);
     layer2_out[11585] <= layer1_out[6671] & ~layer1_out[6670];
     layer2_out[11586] <= ~layer1_out[10043];
     layer2_out[11587] <= layer1_out[2711] | layer1_out[2712];
     layer2_out[11588] <= ~layer1_out[7448];
     layer2_out[11589] <= layer1_out[2640] & layer1_out[2641];
     layer2_out[11590] <= layer1_out[11651];
     layer2_out[11591] <= ~(layer1_out[4018] & layer1_out[4019]);
     layer2_out[11592] <= ~layer1_out[5941];
     layer2_out[11593] <= layer1_out[9252];
     layer2_out[11594] <= layer1_out[6604] ^ layer1_out[6605];
     layer2_out[11595] <= ~layer1_out[4310] | layer1_out[4311];
     layer2_out[11596] <= ~layer1_out[915];
     layer2_out[11597] <= ~layer1_out[1691];
     layer2_out[11598] <= layer1_out[9059];
     layer2_out[11599] <= layer1_out[2349] & layer1_out[2350];
     layer2_out[11600] <= layer1_out[10470] & ~layer1_out[10471];
     layer2_out[11601] <= ~layer1_out[565];
     layer2_out[11602] <= layer1_out[1306];
     layer2_out[11603] <= ~layer1_out[4540];
     layer2_out[11604] <= ~layer1_out[6200];
     layer2_out[11605] <= ~(layer1_out[7007] | layer1_out[7008]);
     layer2_out[11606] <= ~layer1_out[11193] | layer1_out[11192];
     layer2_out[11607] <= ~layer1_out[7122] | layer1_out[7121];
     layer2_out[11608] <= layer1_out[7538] & layer1_out[7539];
     layer2_out[11609] <= ~layer1_out[10389] | layer1_out[10390];
     layer2_out[11610] <= layer1_out[9686];
     layer2_out[11611] <= layer1_out[6500] & ~layer1_out[6499];
     layer2_out[11612] <= layer1_out[3067] & ~layer1_out[3066];
     layer2_out[11613] <= ~layer1_out[7646];
     layer2_out[11614] <= ~layer1_out[5144] | layer1_out[5143];
     layer2_out[11615] <= ~layer1_out[6356] | layer1_out[6355];
     layer2_out[11616] <= layer1_out[3587] & ~layer1_out[3588];
     layer2_out[11617] <= layer1_out[6336] & layer1_out[6337];
     layer2_out[11618] <= ~layer1_out[2793];
     layer2_out[11619] <= 1'b1;
     layer2_out[11620] <= ~layer1_out[10006];
     layer2_out[11621] <= layer1_out[11429] & layer1_out[11430];
     layer2_out[11622] <= 1'b0;
     layer2_out[11623] <= layer1_out[8507];
     layer2_out[11624] <= ~layer1_out[7191];
     layer2_out[11625] <= layer1_out[1223];
     layer2_out[11626] <= ~(layer1_out[8236] ^ layer1_out[8237]);
     layer2_out[11627] <= ~(layer1_out[4177] & layer1_out[4178]);
     layer2_out[11628] <= layer1_out[561];
     layer2_out[11629] <= ~layer1_out[7275];
     layer2_out[11630] <= ~layer1_out[8608] | layer1_out[8609];
     layer2_out[11631] <= layer1_out[2908] ^ layer1_out[2909];
     layer2_out[11632] <= ~(layer1_out[6383] | layer1_out[6384]);
     layer2_out[11633] <= ~layer1_out[920] | layer1_out[921];
     layer2_out[11634] <= ~(layer1_out[7967] ^ layer1_out[7968]);
     layer2_out[11635] <= ~layer1_out[9025] | layer1_out[9026];
     layer2_out[11636] <= layer1_out[4695];
     layer2_out[11637] <= ~layer1_out[3558];
     layer2_out[11638] <= ~layer1_out[224];
     layer2_out[11639] <= ~layer1_out[1958];
     layer2_out[11640] <= ~layer1_out[6449] | layer1_out[6448];
     layer2_out[11641] <= ~layer1_out[6986] | layer1_out[6985];
     layer2_out[11642] <= layer1_out[2999] ^ layer1_out[3000];
     layer2_out[11643] <= layer1_out[10229];
     layer2_out[11644] <= ~(layer1_out[289] ^ layer1_out[290]);
     layer2_out[11645] <= ~(layer1_out[1884] & layer1_out[1885]);
     layer2_out[11646] <= ~layer1_out[7513] | layer1_out[7512];
     layer2_out[11647] <= layer1_out[9244];
     layer2_out[11648] <= layer1_out[990];
     layer2_out[11649] <= layer1_out[4336] | layer1_out[4337];
     layer2_out[11650] <= layer1_out[10761] & ~layer1_out[10760];
     layer2_out[11651] <= layer1_out[2542] & layer1_out[2543];
     layer2_out[11652] <= layer1_out[11668];
     layer2_out[11653] <= ~layer1_out[10574];
     layer2_out[11654] <= layer1_out[6945] & ~layer1_out[6944];
     layer2_out[11655] <= layer1_out[4823] ^ layer1_out[4824];
     layer2_out[11656] <= ~(layer1_out[513] & layer1_out[514]);
     layer2_out[11657] <= layer1_out[9947];
     layer2_out[11658] <= layer1_out[9630];
     layer2_out[11659] <= ~layer1_out[9967];
     layer2_out[11660] <= layer1_out[7577] & ~layer1_out[7578];
     layer2_out[11661] <= ~layer1_out[348];
     layer2_out[11662] <= layer1_out[11721];
     layer2_out[11663] <= ~layer1_out[9551];
     layer2_out[11664] <= layer1_out[5615];
     layer2_out[11665] <= layer1_out[4118] | layer1_out[4119];
     layer2_out[11666] <= layer1_out[8998] & ~layer1_out[8997];
     layer2_out[11667] <= ~(layer1_out[11089] | layer1_out[11090]);
     layer2_out[11668] <= 1'b1;
     layer2_out[11669] <= layer1_out[11121];
     layer2_out[11670] <= layer1_out[5087];
     layer2_out[11671] <= layer1_out[11817] & layer1_out[11818];
     layer2_out[11672] <= layer1_out[5741];
     layer2_out[11673] <= ~(layer1_out[10614] | layer1_out[10615]);
     layer2_out[11674] <= ~layer1_out[2765] | layer1_out[2764];
     layer2_out[11675] <= layer1_out[7326];
     layer2_out[11676] <= layer1_out[9609] & layer1_out[9610];
     layer2_out[11677] <= ~layer1_out[2302];
     layer2_out[11678] <= ~layer1_out[6452] | layer1_out[6451];
     layer2_out[11679] <= layer1_out[6170];
     layer2_out[11680] <= layer1_out[10244] & ~layer1_out[10243];
     layer2_out[11681] <= ~(layer1_out[6520] & layer1_out[6521]);
     layer2_out[11682] <= ~layer1_out[6397];
     layer2_out[11683] <= ~layer1_out[3284] | layer1_out[3283];
     layer2_out[11684] <= ~layer1_out[4493] | layer1_out[4494];
     layer2_out[11685] <= ~layer1_out[6720];
     layer2_out[11686] <= ~layer1_out[9899] | layer1_out[9898];
     layer2_out[11687] <= ~(layer1_out[6817] ^ layer1_out[6818]);
     layer2_out[11688] <= ~(layer1_out[7248] & layer1_out[7249]);
     layer2_out[11689] <= ~layer1_out[7462];
     layer2_out[11690] <= ~layer1_out[8322] | layer1_out[8321];
     layer2_out[11691] <= layer1_out[1042] ^ layer1_out[1043];
     layer2_out[11692] <= ~layer1_out[1688];
     layer2_out[11693] <= ~(layer1_out[956] & layer1_out[957]);
     layer2_out[11694] <= layer1_out[5915];
     layer2_out[11695] <= ~layer1_out[532];
     layer2_out[11696] <= ~layer1_out[2733] | layer1_out[2732];
     layer2_out[11697] <= ~layer1_out[3220];
     layer2_out[11698] <= layer1_out[580];
     layer2_out[11699] <= ~(layer1_out[9338] | layer1_out[9339]);
     layer2_out[11700] <= ~(layer1_out[4134] & layer1_out[4135]);
     layer2_out[11701] <= layer1_out[11079];
     layer2_out[11702] <= layer1_out[1949] & layer1_out[1950];
     layer2_out[11703] <= layer1_out[4040];
     layer2_out[11704] <= layer1_out[6016];
     layer2_out[11705] <= layer1_out[1166];
     layer2_out[11706] <= ~(layer1_out[11228] | layer1_out[11229]);
     layer2_out[11707] <= ~(layer1_out[3307] & layer1_out[3308]);
     layer2_out[11708] <= layer1_out[11378];
     layer2_out[11709] <= layer1_out[6643] | layer1_out[6644];
     layer2_out[11710] <= ~(layer1_out[4019] ^ layer1_out[4020]);
     layer2_out[11711] <= layer1_out[6595];
     layer2_out[11712] <= layer1_out[8624];
     layer2_out[11713] <= ~layer1_out[7852];
     layer2_out[11714] <= ~(layer1_out[2954] | layer1_out[2955]);
     layer2_out[11715] <= ~layer1_out[5833] | layer1_out[5832];
     layer2_out[11716] <= layer1_out[10584];
     layer2_out[11717] <= 1'b0;
     layer2_out[11718] <= ~(layer1_out[8201] | layer1_out[8202]);
     layer2_out[11719] <= ~layer1_out[523];
     layer2_out[11720] <= ~layer1_out[5060];
     layer2_out[11721] <= ~layer1_out[6479];
     layer2_out[11722] <= layer1_out[932] & ~layer1_out[931];
     layer2_out[11723] <= ~layer1_out[6603];
     layer2_out[11724] <= layer1_out[5302] | layer1_out[5303];
     layer2_out[11725] <= ~layer1_out[3438];
     layer2_out[11726] <= ~(layer1_out[10371] & layer1_out[10372]);
     layer2_out[11727] <= ~(layer1_out[10139] ^ layer1_out[10140]);
     layer2_out[11728] <= ~layer1_out[9260] | layer1_out[9261];
     layer2_out[11729] <= ~layer1_out[5204] | layer1_out[5203];
     layer2_out[11730] <= ~layer1_out[6504] | layer1_out[6505];
     layer2_out[11731] <= 1'b0;
     layer2_out[11732] <= layer1_out[2491] & ~layer1_out[2490];
     layer2_out[11733] <= layer1_out[3582] & ~layer1_out[3583];
     layer2_out[11734] <= layer1_out[5006];
     layer2_out[11735] <= layer1_out[447] & layer1_out[448];
     layer2_out[11736] <= layer1_out[7061];
     layer2_out[11737] <= ~(layer1_out[2652] & layer1_out[2653]);
     layer2_out[11738] <= layer1_out[7165] | layer1_out[7166];
     layer2_out[11739] <= ~layer1_out[3937];
     layer2_out[11740] <= layer1_out[62] & ~layer1_out[61];
     layer2_out[11741] <= layer1_out[11211];
     layer2_out[11742] <= layer1_out[9780] & layer1_out[9781];
     layer2_out[11743] <= ~layer1_out[208];
     layer2_out[11744] <= ~(layer1_out[10211] | layer1_out[10212]);
     layer2_out[11745] <= layer1_out[14] & ~layer1_out[13];
     layer2_out[11746] <= ~(layer1_out[6243] | layer1_out[6244]);
     layer2_out[11747] <= layer1_out[7241] | layer1_out[7242];
     layer2_out[11748] <= ~(layer1_out[9270] | layer1_out[9271]);
     layer2_out[11749] <= layer1_out[10641];
     layer2_out[11750] <= layer1_out[1907];
     layer2_out[11751] <= ~(layer1_out[3819] | layer1_out[3820]);
     layer2_out[11752] <= ~layer1_out[5847];
     layer2_out[11753] <= layer1_out[1025] | layer1_out[1026];
     layer2_out[11754] <= layer1_out[2739] & layer1_out[2740];
     layer2_out[11755] <= ~layer1_out[10144] | layer1_out[10143];
     layer2_out[11756] <= layer1_out[699] & layer1_out[700];
     layer2_out[11757] <= ~layer1_out[2458];
     layer2_out[11758] <= layer1_out[9111] & ~layer1_out[9110];
     layer2_out[11759] <= ~layer1_out[11542];
     layer2_out[11760] <= ~(layer1_out[9809] | layer1_out[9810]);
     layer2_out[11761] <= layer1_out[2451] & ~layer1_out[2450];
     layer2_out[11762] <= layer1_out[7160];
     layer2_out[11763] <= layer1_out[10354] & ~layer1_out[10353];
     layer2_out[11764] <= ~(layer1_out[11598] & layer1_out[11599]);
     layer2_out[11765] <= layer1_out[10903];
     layer2_out[11766] <= ~layer1_out[2119];
     layer2_out[11767] <= layer1_out[1099];
     layer2_out[11768] <= ~(layer1_out[1091] & layer1_out[1092]);
     layer2_out[11769] <= layer1_out[4015] ^ layer1_out[4016];
     layer2_out[11770] <= layer1_out[8438] ^ layer1_out[8439];
     layer2_out[11771] <= layer1_out[11468];
     layer2_out[11772] <= layer1_out[8038] & layer1_out[8039];
     layer2_out[11773] <= ~layer1_out[1533];
     layer2_out[11774] <= layer1_out[821] & ~layer1_out[820];
     layer2_out[11775] <= layer1_out[6729] & layer1_out[6730];
     layer2_out[11776] <= ~layer1_out[3570];
     layer2_out[11777] <= ~(layer1_out[5482] ^ layer1_out[5483]);
     layer2_out[11778] <= layer1_out[7239];
     layer2_out[11779] <= layer1_out[5113];
     layer2_out[11780] <= layer1_out[11996];
     layer2_out[11781] <= ~(layer1_out[9495] | layer1_out[9496]);
     layer2_out[11782] <= 1'b1;
     layer2_out[11783] <= ~layer1_out[5843];
     layer2_out[11784] <= ~layer1_out[1346];
     layer2_out[11785] <= layer1_out[4116] & ~layer1_out[4117];
     layer2_out[11786] <= ~layer1_out[3567] | layer1_out[3568];
     layer2_out[11787] <= ~layer1_out[10789];
     layer2_out[11788] <= layer1_out[7681] & layer1_out[7682];
     layer2_out[11789] <= ~(layer1_out[9387] & layer1_out[9388]);
     layer2_out[11790] <= ~layer1_out[3832];
     layer2_out[11791] <= ~layer1_out[9664] | layer1_out[9665];
     layer2_out[11792] <= layer1_out[2881] & ~layer1_out[2880];
     layer2_out[11793] <= layer1_out[10827];
     layer2_out[11794] <= layer1_out[5717];
     layer2_out[11795] <= layer1_out[5517];
     layer2_out[11796] <= layer1_out[148];
     layer2_out[11797] <= layer1_out[8188] ^ layer1_out[8189];
     layer2_out[11798] <= ~layer1_out[6625];
     layer2_out[11799] <= layer1_out[5707] | layer1_out[5708];
     layer2_out[11800] <= ~(layer1_out[2323] ^ layer1_out[2324]);
     layer2_out[11801] <= layer1_out[4071] & ~layer1_out[4072];
     layer2_out[11802] <= layer1_out[7464] ^ layer1_out[7465];
     layer2_out[11803] <= ~(layer1_out[5093] | layer1_out[5094]);
     layer2_out[11804] <= ~layer1_out[7350];
     layer2_out[11805] <= ~(layer1_out[6110] & layer1_out[6111]);
     layer2_out[11806] <= layer1_out[7296] & ~layer1_out[7297];
     layer2_out[11807] <= ~(layer1_out[8510] & layer1_out[8511]);
     layer2_out[11808] <= layer1_out[7788] & layer1_out[7789];
     layer2_out[11809] <= ~layer1_out[7920];
     layer2_out[11810] <= layer1_out[3462];
     layer2_out[11811] <= layer1_out[3957];
     layer2_out[11812] <= ~layer1_out[8515];
     layer2_out[11813] <= ~layer1_out[381];
     layer2_out[11814] <= layer1_out[1946] ^ layer1_out[1947];
     layer2_out[11815] <= layer1_out[1886];
     layer2_out[11816] <= ~layer1_out[4571];
     layer2_out[11817] <= layer1_out[4360] & layer1_out[4361];
     layer2_out[11818] <= ~layer1_out[4435] | layer1_out[4436];
     layer2_out[11819] <= layer1_out[895] & layer1_out[896];
     layer2_out[11820] <= 1'b1;
     layer2_out[11821] <= layer1_out[6720] & ~layer1_out[6719];
     layer2_out[11822] <= layer1_out[3890] & layer1_out[3891];
     layer2_out[11823] <= layer1_out[11118] & layer1_out[11119];
     layer2_out[11824] <= layer1_out[10525] | layer1_out[10526];
     layer2_out[11825] <= 1'b0;
     layer2_out[11826] <= layer1_out[9241] | layer1_out[9242];
     layer2_out[11827] <= layer1_out[629] & ~layer1_out[628];
     layer2_out[11828] <= ~layer1_out[3490] | layer1_out[3491];
     layer2_out[11829] <= ~layer1_out[11676] | layer1_out[11677];
     layer2_out[11830] <= layer1_out[1874] ^ layer1_out[1875];
     layer2_out[11831] <= layer1_out[3594];
     layer2_out[11832] <= layer1_out[7642] & ~layer1_out[7643];
     layer2_out[11833] <= ~(layer1_out[8230] | layer1_out[8231]);
     layer2_out[11834] <= layer1_out[11840];
     layer2_out[11835] <= layer1_out[7006] & layer1_out[7007];
     layer2_out[11836] <= layer1_out[4107] | layer1_out[4108];
     layer2_out[11837] <= layer1_out[8049] & layer1_out[8050];
     layer2_out[11838] <= layer1_out[1870];
     layer2_out[11839] <= layer1_out[8048];
     layer2_out[11840] <= layer1_out[1773] & ~layer1_out[1774];
     layer2_out[11841] <= 1'b0;
     layer2_out[11842] <= ~layer1_out[489];
     layer2_out[11843] <= ~(layer1_out[3420] ^ layer1_out[3421]);
     layer2_out[11844] <= layer1_out[10546] | layer1_out[10547];
     layer2_out[11845] <= layer1_out[3727];
     layer2_out[11846] <= ~layer1_out[866] | layer1_out[867];
     layer2_out[11847] <= ~(layer1_out[7649] & layer1_out[7650]);
     layer2_out[11848] <= layer1_out[270] & layer1_out[271];
     layer2_out[11849] <= layer1_out[221] & ~layer1_out[222];
     layer2_out[11850] <= layer1_out[10263] & ~layer1_out[10264];
     layer2_out[11851] <= layer1_out[10290] & ~layer1_out[10291];
     layer2_out[11852] <= layer1_out[95] & ~layer1_out[96];
     layer2_out[11853] <= ~layer1_out[9656] | layer1_out[9655];
     layer2_out[11854] <= layer1_out[11610];
     layer2_out[11855] <= layer1_out[4486];
     layer2_out[11856] <= ~(layer1_out[10944] & layer1_out[10945]);
     layer2_out[11857] <= layer1_out[574] & layer1_out[575];
     layer2_out[11858] <= layer1_out[678] ^ layer1_out[679];
     layer2_out[11859] <= layer1_out[7336] & ~layer1_out[7337];
     layer2_out[11860] <= layer1_out[1811];
     layer2_out[11861] <= ~layer1_out[2842] | layer1_out[2843];
     layer2_out[11862] <= ~(layer1_out[3786] ^ layer1_out[3787]);
     layer2_out[11863] <= ~(layer1_out[2774] & layer1_out[2775]);
     layer2_out[11864] <= ~(layer1_out[8910] & layer1_out[8911]);
     layer2_out[11865] <= ~layer1_out[10622];
     layer2_out[11866] <= ~(layer1_out[2366] & layer1_out[2367]);
     layer2_out[11867] <= ~layer1_out[11020] | layer1_out[11021];
     layer2_out[11868] <= layer1_out[8676] & ~layer1_out[8675];
     layer2_out[11869] <= layer1_out[3690] & layer1_out[3691];
     layer2_out[11870] <= ~layer1_out[4154];
     layer2_out[11871] <= layer1_out[9394];
     layer2_out[11872] <= layer1_out[907];
     layer2_out[11873] <= ~layer1_out[3256];
     layer2_out[11874] <= layer1_out[6743] & layer1_out[6744];
     layer2_out[11875] <= layer1_out[4793] | layer1_out[4794];
     layer2_out[11876] <= ~layer1_out[2663] | layer1_out[2662];
     layer2_out[11877] <= ~(layer1_out[7732] & layer1_out[7733]);
     layer2_out[11878] <= layer1_out[4552] & layer1_out[4553];
     layer2_out[11879] <= ~(layer1_out[661] & layer1_out[662]);
     layer2_out[11880] <= ~(layer1_out[5431] ^ layer1_out[5432]);
     layer2_out[11881] <= ~(layer1_out[10079] & layer1_out[10080]);
     layer2_out[11882] <= layer1_out[8737] & ~layer1_out[8738];
     layer2_out[11883] <= ~(layer1_out[6420] ^ layer1_out[6421]);
     layer2_out[11884] <= layer1_out[5156] & ~layer1_out[5157];
     layer2_out[11885] <= ~(layer1_out[11451] & layer1_out[11452]);
     layer2_out[11886] <= ~layer1_out[8686];
     layer2_out[11887] <= layer1_out[8762];
     layer2_out[11888] <= ~layer1_out[1406];
     layer2_out[11889] <= layer1_out[7619];
     layer2_out[11890] <= layer1_out[7814] | layer1_out[7815];
     layer2_out[11891] <= ~layer1_out[8955];
     layer2_out[11892] <= layer1_out[7314] & ~layer1_out[7313];
     layer2_out[11893] <= layer1_out[6085] & ~layer1_out[6084];
     layer2_out[11894] <= layer1_out[2882] & layer1_out[2883];
     layer2_out[11895] <= layer1_out[7065];
     layer2_out[11896] <= layer1_out[4940] & ~layer1_out[4939];
     layer2_out[11897] <= ~layer1_out[7676];
     layer2_out[11898] <= layer1_out[4640];
     layer2_out[11899] <= layer1_out[1980] ^ layer1_out[1981];
     layer2_out[11900] <= ~layer1_out[9401] | layer1_out[9402];
     layer2_out[11901] <= layer1_out[11922];
     layer2_out[11902] <= ~(layer1_out[1343] ^ layer1_out[1344]);
     layer2_out[11903] <= 1'b1;
     layer2_out[11904] <= ~layer1_out[1655];
     layer2_out[11905] <= ~(layer1_out[3667] ^ layer1_out[3668]);
     layer2_out[11906] <= layer1_out[392];
     layer2_out[11907] <= ~layer1_out[2439];
     layer2_out[11908] <= ~(layer1_out[2734] | layer1_out[2735]);
     layer2_out[11909] <= ~(layer1_out[3846] & layer1_out[3847]);
     layer2_out[11910] <= layer1_out[4713];
     layer2_out[11911] <= ~layer1_out[4774];
     layer2_out[11912] <= ~(layer1_out[7274] ^ layer1_out[7275]);
     layer2_out[11913] <= ~layer1_out[11502] | layer1_out[11503];
     layer2_out[11914] <= ~layer1_out[3587];
     layer2_out[11915] <= layer1_out[1553] & layer1_out[1554];
     layer2_out[11916] <= ~(layer1_out[3716] | layer1_out[3717]);
     layer2_out[11917] <= ~(layer1_out[2939] ^ layer1_out[2940]);
     layer2_out[11918] <= ~(layer1_out[2361] & layer1_out[2362]);
     layer2_out[11919] <= ~layer1_out[4840];
     layer2_out[11920] <= ~layer1_out[2517];
     layer2_out[11921] <= layer1_out[7609];
     layer2_out[11922] <= layer1_out[3404] & ~layer1_out[3405];
     layer2_out[11923] <= ~layer1_out[7511] | layer1_out[7512];
     layer2_out[11924] <= ~layer1_out[3626];
     layer2_out[11925] <= ~layer1_out[253];
     layer2_out[11926] <= layer1_out[6391] ^ layer1_out[6392];
     layer2_out[11927] <= ~layer1_out[4234];
     layer2_out[11928] <= layer1_out[11969] & layer1_out[11970];
     layer2_out[11929] <= ~layer1_out[8570] | layer1_out[8571];
     layer2_out[11930] <= layer1_out[9181] ^ layer1_out[9182];
     layer2_out[11931] <= ~(layer1_out[8051] | layer1_out[8052]);
     layer2_out[11932] <= layer1_out[2682];
     layer2_out[11933] <= layer1_out[3525] & ~layer1_out[3524];
     layer2_out[11934] <= 1'b1;
     layer2_out[11935] <= ~layer1_out[11437];
     layer2_out[11936] <= ~layer1_out[6035];
     layer2_out[11937] <= ~layer1_out[3278] | layer1_out[3279];
     layer2_out[11938] <= layer1_out[8332];
     layer2_out[11939] <= ~(layer1_out[10289] & layer1_out[10290]);
     layer2_out[11940] <= layer1_out[1136] & ~layer1_out[1137];
     layer2_out[11941] <= ~(layer1_out[1107] | layer1_out[1108]);
     layer2_out[11942] <= ~layer1_out[3017];
     layer2_out[11943] <= ~(layer1_out[6082] | layer1_out[6083]);
     layer2_out[11944] <= ~(layer1_out[7711] & layer1_out[7712]);
     layer2_out[11945] <= layer1_out[6411];
     layer2_out[11946] <= layer1_out[10794] | layer1_out[10795];
     layer2_out[11947] <= layer1_out[3743] ^ layer1_out[3744];
     layer2_out[11948] <= layer1_out[819] & ~layer1_out[820];
     layer2_out[11949] <= ~layer1_out[10473];
     layer2_out[11950] <= ~layer1_out[3286] | layer1_out[3285];
     layer2_out[11951] <= ~(layer1_out[9715] | layer1_out[9716]);
     layer2_out[11952] <= ~layer1_out[7083] | layer1_out[7082];
     layer2_out[11953] <= ~layer1_out[170];
     layer2_out[11954] <= ~layer1_out[9150] | layer1_out[9149];
     layer2_out[11955] <= layer1_out[10004] & ~layer1_out[10005];
     layer2_out[11956] <= ~(layer1_out[1805] | layer1_out[1806]);
     layer2_out[11957] <= layer1_out[6484] & ~layer1_out[6485];
     layer2_out[11958] <= ~layer1_out[8547];
     layer2_out[11959] <= layer1_out[7281] ^ layer1_out[7282];
     layer2_out[11960] <= 1'b0;
     layer2_out[11961] <= ~(layer1_out[4412] & layer1_out[4413]);
     layer2_out[11962] <= layer1_out[814] | layer1_out[815];
     layer2_out[11963] <= ~layer1_out[7796] | layer1_out[7797];
     layer2_out[11964] <= ~layer1_out[727] | layer1_out[726];
     layer2_out[11965] <= ~layer1_out[11794];
     layer2_out[11966] <= ~layer1_out[800];
     layer2_out[11967] <= ~(layer1_out[2863] | layer1_out[2864]);
     layer2_out[11968] <= layer1_out[1065] & layer1_out[1066];
     layer2_out[11969] <= layer1_out[9230];
     layer2_out[11970] <= ~layer1_out[6688];
     layer2_out[11971] <= layer1_out[2613] & ~layer1_out[2614];
     layer2_out[11972] <= layer1_out[7852] & ~layer1_out[7853];
     layer2_out[11973] <= ~layer1_out[3319] | layer1_out[3320];
     layer2_out[11974] <= ~layer1_out[8301];
     layer2_out[11975] <= layer1_out[4944];
     layer2_out[11976] <= ~layer1_out[9418] | layer1_out[9419];
     layer2_out[11977] <= ~layer1_out[5096];
     layer2_out[11978] <= ~layer1_out[1595];
     layer2_out[11979] <= layer1_out[9822] & ~layer1_out[9821];
     layer2_out[11980] <= ~layer1_out[11324] | layer1_out[11325];
     layer2_out[11981] <= layer1_out[7002] ^ layer1_out[7003];
     layer2_out[11982] <= layer1_out[5728] & ~layer1_out[5729];
     layer2_out[11983] <= 1'b0;
     layer2_out[11984] <= layer1_out[10312] ^ layer1_out[10313];
     layer2_out[11985] <= ~(layer1_out[7291] ^ layer1_out[7292]);
     layer2_out[11986] <= ~layer1_out[8093];
     layer2_out[11987] <= layer1_out[330] & ~layer1_out[331];
     layer2_out[11988] <= ~layer1_out[2074] | layer1_out[2075];
     layer2_out[11989] <= ~layer1_out[7105] | layer1_out[7106];
     layer2_out[11990] <= layer1_out[10309] ^ layer1_out[10310];
     layer2_out[11991] <= ~(layer1_out[238] & layer1_out[239]);
     layer2_out[11992] <= layer1_out[10933];
     layer2_out[11993] <= ~layer1_out[5770] | layer1_out[5769];
     layer2_out[11994] <= ~(layer1_out[11256] & layer1_out[11257]);
     layer2_out[11995] <= ~layer1_out[4126] | layer1_out[4127];
     layer2_out[11996] <= layer1_out[4307] | layer1_out[4308];
     layer2_out[11997] <= layer1_out[5165] ^ layer1_out[5166];
     layer2_out[11998] <= layer1_out[10562];
     layer2_out[11999] <= ~layer1_out[269] | layer1_out[268];
     layer3_out[0] <= ~layer2_out[831];
     layer3_out[1] <= layer2_out[11173];
     layer3_out[2] <= ~layer2_out[6858] | layer2_out[6857];
     layer3_out[3] <= ~layer2_out[2781];
     layer3_out[4] <= ~layer2_out[8181];
     layer3_out[5] <= layer2_out[2468];
     layer3_out[6] <= ~(layer2_out[1148] ^ layer2_out[1149]);
     layer3_out[7] <= ~layer2_out[10142] | layer2_out[10143];
     layer3_out[8] <= ~(layer2_out[4840] | layer2_out[4841]);
     layer3_out[9] <= ~layer2_out[1109];
     layer3_out[10] <= layer2_out[10928];
     layer3_out[11] <= layer2_out[9622];
     layer3_out[12] <= layer2_out[3392] & ~layer2_out[3393];
     layer3_out[13] <= ~layer2_out[5343];
     layer3_out[14] <= ~layer2_out[11811] | layer2_out[11810];
     layer3_out[15] <= ~layer2_out[6690] | layer2_out[6691];
     layer3_out[16] <= layer2_out[5697] & ~layer2_out[5698];
     layer3_out[17] <= layer2_out[374] ^ layer2_out[375];
     layer3_out[18] <= layer2_out[1388] & ~layer2_out[1387];
     layer3_out[19] <= layer2_out[5874] & ~layer2_out[5875];
     layer3_out[20] <= layer2_out[1102] & ~layer2_out[1101];
     layer3_out[21] <= ~(layer2_out[5884] & layer2_out[5885]);
     layer3_out[22] <= layer2_out[5112] & layer2_out[5113];
     layer3_out[23] <= ~(layer2_out[8521] ^ layer2_out[8522]);
     layer3_out[24] <= ~layer2_out[11353];
     layer3_out[25] <= ~layer2_out[2043];
     layer3_out[26] <= layer2_out[11612];
     layer3_out[27] <= ~(layer2_out[8072] | layer2_out[8073]);
     layer3_out[28] <= ~layer2_out[7720] | layer2_out[7719];
     layer3_out[29] <= ~(layer2_out[1118] | layer2_out[1119]);
     layer3_out[30] <= ~layer2_out[11040];
     layer3_out[31] <= layer2_out[6162] & ~layer2_out[6161];
     layer3_out[32] <= layer2_out[5283];
     layer3_out[33] <= ~layer2_out[9011];
     layer3_out[34] <= ~layer2_out[3286];
     layer3_out[35] <= layer2_out[2419];
     layer3_out[36] <= layer2_out[9948] & ~layer2_out[9947];
     layer3_out[37] <= layer2_out[475];
     layer3_out[38] <= ~(layer2_out[3180] & layer2_out[3181]);
     layer3_out[39] <= ~layer2_out[567] | layer2_out[566];
     layer3_out[40] <= layer2_out[8525] ^ layer2_out[8526];
     layer3_out[41] <= ~layer2_out[182];
     layer3_out[42] <= layer2_out[6300] ^ layer2_out[6301];
     layer3_out[43] <= ~(layer2_out[7298] ^ layer2_out[7299]);
     layer3_out[44] <= ~(layer2_out[2616] ^ layer2_out[2617]);
     layer3_out[45] <= layer2_out[4163];
     layer3_out[46] <= layer2_out[2897] & ~layer2_out[2896];
     layer3_out[47] <= ~layer2_out[4864];
     layer3_out[48] <= ~layer2_out[2128] | layer2_out[2129];
     layer3_out[49] <= ~(layer2_out[11274] | layer2_out[11275]);
     layer3_out[50] <= layer2_out[5755] & ~layer2_out[5756];
     layer3_out[51] <= layer2_out[7126] | layer2_out[7127];
     layer3_out[52] <= ~(layer2_out[355] & layer2_out[356]);
     layer3_out[53] <= ~layer2_out[9323] | layer2_out[9324];
     layer3_out[54] <= ~layer2_out[10875];
     layer3_out[55] <= ~layer2_out[8870] | layer2_out[8871];
     layer3_out[56] <= ~layer2_out[8589];
     layer3_out[57] <= layer2_out[4384] ^ layer2_out[4385];
     layer3_out[58] <= ~(layer2_out[1706] ^ layer2_out[1707]);
     layer3_out[59] <= ~(layer2_out[9866] ^ layer2_out[9867]);
     layer3_out[60] <= ~layer2_out[10631];
     layer3_out[61] <= ~(layer2_out[2094] ^ layer2_out[2095]);
     layer3_out[62] <= ~(layer2_out[10455] | layer2_out[10456]);
     layer3_out[63] <= layer2_out[9561] & ~layer2_out[9560];
     layer3_out[64] <= ~layer2_out[1395];
     layer3_out[65] <= ~layer2_out[10375];
     layer3_out[66] <= ~layer2_out[3091];
     layer3_out[67] <= layer2_out[6082] & ~layer2_out[6083];
     layer3_out[68] <= ~layer2_out[7749] | layer2_out[7748];
     layer3_out[69] <= layer2_out[11175];
     layer3_out[70] <= layer2_out[5135] ^ layer2_out[5136];
     layer3_out[71] <= layer2_out[9068] & ~layer2_out[9067];
     layer3_out[72] <= layer2_out[5017];
     layer3_out[73] <= layer2_out[10294] & layer2_out[10295];
     layer3_out[74] <= ~layer2_out[924];
     layer3_out[75] <= layer2_out[3641];
     layer3_out[76] <= ~(layer2_out[4170] | layer2_out[4171]);
     layer3_out[77] <= layer2_out[6193] & ~layer2_out[6194];
     layer3_out[78] <= ~(layer2_out[2588] | layer2_out[2589]);
     layer3_out[79] <= ~layer2_out[9267] | layer2_out[9268];
     layer3_out[80] <= ~(layer2_out[724] | layer2_out[725]);
     layer3_out[81] <= layer2_out[3249] | layer2_out[3250];
     layer3_out[82] <= layer2_out[11775] & ~layer2_out[11776];
     layer3_out[83] <= layer2_out[8022] & layer2_out[8023];
     layer3_out[84] <= layer2_out[5267];
     layer3_out[85] <= layer2_out[9321] & ~layer2_out[9320];
     layer3_out[86] <= ~layer2_out[1819];
     layer3_out[87] <= layer2_out[4711];
     layer3_out[88] <= ~(layer2_out[8338] | layer2_out[8339]);
     layer3_out[89] <= layer2_out[2769] ^ layer2_out[2770];
     layer3_out[90] <= ~(layer2_out[3429] | layer2_out[3430]);
     layer3_out[91] <= layer2_out[8342] ^ layer2_out[8343];
     layer3_out[92] <= layer2_out[3024] & ~layer2_out[3023];
     layer3_out[93] <= ~layer2_out[9715];
     layer3_out[94] <= layer2_out[4212] & layer2_out[4213];
     layer3_out[95] <= layer2_out[6469] & layer2_out[6470];
     layer3_out[96] <= ~(layer2_out[8255] ^ layer2_out[8256]);
     layer3_out[97] <= layer2_out[7616];
     layer3_out[98] <= ~layer2_out[4110];
     layer3_out[99] <= ~layer2_out[1925];
     layer3_out[100] <= layer2_out[11748];
     layer3_out[101] <= ~(layer2_out[11700] ^ layer2_out[11701]);
     layer3_out[102] <= layer2_out[5503] & ~layer2_out[5502];
     layer3_out[103] <= layer2_out[11912];
     layer3_out[104] <= ~layer2_out[5445];
     layer3_out[105] <= layer2_out[10438] & ~layer2_out[10439];
     layer3_out[106] <= layer2_out[6544] & layer2_out[6545];
     layer3_out[107] <= layer2_out[3904] & layer2_out[3905];
     layer3_out[108] <= ~layer2_out[10201];
     layer3_out[109] <= ~layer2_out[927];
     layer3_out[110] <= layer2_out[7944] & ~layer2_out[7945];
     layer3_out[111] <= ~(layer2_out[3991] ^ layer2_out[3992]);
     layer3_out[112] <= ~layer2_out[2406];
     layer3_out[113] <= layer2_out[8749] & ~layer2_out[8748];
     layer3_out[114] <= layer2_out[4394] & layer2_out[4395];
     layer3_out[115] <= layer2_out[1612];
     layer3_out[116] <= layer2_out[6885];
     layer3_out[117] <= layer2_out[4000] & layer2_out[4001];
     layer3_out[118] <= ~layer2_out[3944];
     layer3_out[119] <= layer2_out[11148] & ~layer2_out[11149];
     layer3_out[120] <= ~layer2_out[6635] | layer2_out[6634];
     layer3_out[121] <= layer2_out[1935];
     layer3_out[122] <= layer2_out[2343] ^ layer2_out[2344];
     layer3_out[123] <= layer2_out[11639] & ~layer2_out[11640];
     layer3_out[124] <= layer2_out[11859];
     layer3_out[125] <= layer2_out[9188];
     layer3_out[126] <= layer2_out[9710] & ~layer2_out[9709];
     layer3_out[127] <= ~(layer2_out[2657] & layer2_out[2658]);
     layer3_out[128] <= layer2_out[4017] & layer2_out[4018];
     layer3_out[129] <= ~(layer2_out[10114] | layer2_out[10115]);
     layer3_out[130] <= ~layer2_out[5833] | layer2_out[5832];
     layer3_out[131] <= layer2_out[500];
     layer3_out[132] <= layer2_out[2360];
     layer3_out[133] <= ~layer2_out[5042];
     layer3_out[134] <= ~(layer2_out[5834] & layer2_out[5835]);
     layer3_out[135] <= ~(layer2_out[7764] | layer2_out[7765]);
     layer3_out[136] <= ~layer2_out[2841];
     layer3_out[137] <= layer2_out[3372] & ~layer2_out[3373];
     layer3_out[138] <= ~layer2_out[11098] | layer2_out[11097];
     layer3_out[139] <= ~layer2_out[303];
     layer3_out[140] <= layer2_out[9020];
     layer3_out[141] <= ~(layer2_out[1967] & layer2_out[1968]);
     layer3_out[142] <= layer2_out[5176];
     layer3_out[143] <= layer2_out[8957] ^ layer2_out[8958];
     layer3_out[144] <= ~layer2_out[6539];
     layer3_out[145] <= ~layer2_out[6098];
     layer3_out[146] <= layer2_out[5327] & layer2_out[5328];
     layer3_out[147] <= ~layer2_out[11819];
     layer3_out[148] <= ~(layer2_out[10832] & layer2_out[10833]);
     layer3_out[149] <= layer2_out[7613] & ~layer2_out[7614];
     layer3_out[150] <= ~(layer2_out[8582] | layer2_out[8583]);
     layer3_out[151] <= ~layer2_out[2625];
     layer3_out[152] <= ~(layer2_out[9164] ^ layer2_out[9165]);
     layer3_out[153] <= layer2_out[11288] & layer2_out[11289];
     layer3_out[154] <= layer2_out[1913] & layer2_out[1914];
     layer3_out[155] <= layer2_out[4474] & layer2_out[4475];
     layer3_out[156] <= ~layer2_out[11785];
     layer3_out[157] <= layer2_out[29] & ~layer2_out[28];
     layer3_out[158] <= layer2_out[6263] & ~layer2_out[6264];
     layer3_out[159] <= layer2_out[6761];
     layer3_out[160] <= ~(layer2_out[9801] | layer2_out[9802]);
     layer3_out[161] <= layer2_out[1747] | layer2_out[1748];
     layer3_out[162] <= ~(layer2_out[767] ^ layer2_out[768]);
     layer3_out[163] <= ~layer2_out[3844];
     layer3_out[164] <= ~layer2_out[2755];
     layer3_out[165] <= ~(layer2_out[3885] ^ layer2_out[3886]);
     layer3_out[166] <= ~layer2_out[6290];
     layer3_out[167] <= ~(layer2_out[5323] | layer2_out[5324]);
     layer3_out[168] <= layer2_out[4341];
     layer3_out[169] <= layer2_out[2275];
     layer3_out[170] <= layer2_out[6491];
     layer3_out[171] <= ~layer2_out[11919] | layer2_out[11918];
     layer3_out[172] <= ~layer2_out[11703];
     layer3_out[173] <= layer2_out[2740];
     layer3_out[174] <= layer2_out[21] & layer2_out[22];
     layer3_out[175] <= layer2_out[6076] & layer2_out[6077];
     layer3_out[176] <= ~layer2_out[10508] | layer2_out[10509];
     layer3_out[177] <= ~layer2_out[3746];
     layer3_out[178] <= layer2_out[11367] & layer2_out[11368];
     layer3_out[179] <= layer2_out[9511] & ~layer2_out[9512];
     layer3_out[180] <= layer2_out[10465] & ~layer2_out[10466];
     layer3_out[181] <= layer2_out[3123] & layer2_out[3124];
     layer3_out[182] <= layer2_out[10838] ^ layer2_out[10839];
     layer3_out[183] <= ~layer2_out[1074];
     layer3_out[184] <= ~layer2_out[3333];
     layer3_out[185] <= layer2_out[651];
     layer3_out[186] <= ~(layer2_out[6177] ^ layer2_out[6178]);
     layer3_out[187] <= ~layer2_out[9166];
     layer3_out[188] <= layer2_out[1325] & ~layer2_out[1326];
     layer3_out[189] <= layer2_out[2526];
     layer3_out[190] <= layer2_out[11439] ^ layer2_out[11440];
     layer3_out[191] <= ~layer2_out[11996];
     layer3_out[192] <= layer2_out[3411] & ~layer2_out[3410];
     layer3_out[193] <= ~layer2_out[11521] | layer2_out[11522];
     layer3_out[194] <= ~layer2_out[119];
     layer3_out[195] <= ~layer2_out[5675] | layer2_out[5676];
     layer3_out[196] <= ~layer2_out[8040] | layer2_out[8041];
     layer3_out[197] <= layer2_out[9182] & ~layer2_out[9183];
     layer3_out[198] <= layer2_out[665];
     layer3_out[199] <= layer2_out[9040];
     layer3_out[200] <= layer2_out[8690] & ~layer2_out[8691];
     layer3_out[201] <= layer2_out[6599] & ~layer2_out[6600];
     layer3_out[202] <= layer2_out[9386];
     layer3_out[203] <= ~layer2_out[7100];
     layer3_out[204] <= ~(layer2_out[9818] ^ layer2_out[9819]);
     layer3_out[205] <= ~layer2_out[2295];
     layer3_out[206] <= layer2_out[10523] & layer2_out[10524];
     layer3_out[207] <= ~layer2_out[1403];
     layer3_out[208] <= layer2_out[3483] & layer2_out[3484];
     layer3_out[209] <= ~layer2_out[7747] | layer2_out[7748];
     layer3_out[210] <= layer2_out[11892] & ~layer2_out[11891];
     layer3_out[211] <= ~layer2_out[1437];
     layer3_out[212] <= ~layer2_out[7225];
     layer3_out[213] <= layer2_out[10154] & ~layer2_out[10153];
     layer3_out[214] <= layer2_out[8504] ^ layer2_out[8505];
     layer3_out[215] <= ~(layer2_out[10336] ^ layer2_out[10337]);
     layer3_out[216] <= layer2_out[2512];
     layer3_out[217] <= layer2_out[11887] & ~layer2_out[11888];
     layer3_out[218] <= ~(layer2_out[9195] ^ layer2_out[9196]);
     layer3_out[219] <= layer2_out[8998];
     layer3_out[220] <= ~layer2_out[9155];
     layer3_out[221] <= layer2_out[1388];
     layer3_out[222] <= layer2_out[3847] ^ layer2_out[3848];
     layer3_out[223] <= layer2_out[5497] & layer2_out[5498];
     layer3_out[224] <= layer2_out[434] & ~layer2_out[433];
     layer3_out[225] <= ~layer2_out[4632];
     layer3_out[226] <= layer2_out[7445] ^ layer2_out[7446];
     layer3_out[227] <= ~layer2_out[11648] | layer2_out[11649];
     layer3_out[228] <= ~(layer2_out[9743] | layer2_out[9744]);
     layer3_out[229] <= layer2_out[2014] & layer2_out[2015];
     layer3_out[230] <= layer2_out[7086] & layer2_out[7087];
     layer3_out[231] <= ~layer2_out[5203];
     layer3_out[232] <= layer2_out[1296];
     layer3_out[233] <= layer2_out[592];
     layer3_out[234] <= ~layer2_out[7875];
     layer3_out[235] <= ~(layer2_out[7412] ^ layer2_out[7413]);
     layer3_out[236] <= layer2_out[11969] & ~layer2_out[11970];
     layer3_out[237] <= layer2_out[2061] ^ layer2_out[2062];
     layer3_out[238] <= ~layer2_out[377];
     layer3_out[239] <= ~(layer2_out[9959] ^ layer2_out[9960]);
     layer3_out[240] <= ~(layer2_out[6299] ^ layer2_out[6300]);
     layer3_out[241] <= ~(layer2_out[7433] | layer2_out[7434]);
     layer3_out[242] <= layer2_out[282];
     layer3_out[243] <= ~(layer2_out[9085] ^ layer2_out[9086]);
     layer3_out[244] <= layer2_out[8960] ^ layer2_out[8961];
     layer3_out[245] <= ~layer2_out[9636];
     layer3_out[246] <= layer2_out[8507];
     layer3_out[247] <= layer2_out[9982] & ~layer2_out[9981];
     layer3_out[248] <= layer2_out[3827];
     layer3_out[249] <= layer2_out[196] & layer2_out[197];
     layer3_out[250] <= layer2_out[3925];
     layer3_out[251] <= ~layer2_out[8845];
     layer3_out[252] <= ~(layer2_out[7022] | layer2_out[7023]);
     layer3_out[253] <= ~layer2_out[11455];
     layer3_out[254] <= ~layer2_out[10701];
     layer3_out[255] <= ~layer2_out[7366];
     layer3_out[256] <= layer2_out[7918] ^ layer2_out[7919];
     layer3_out[257] <= ~(layer2_out[5184] ^ layer2_out[5185]);
     layer3_out[258] <= ~layer2_out[4849];
     layer3_out[259] <= ~layer2_out[9954];
     layer3_out[260] <= ~layer2_out[1918] | layer2_out[1917];
     layer3_out[261] <= layer2_out[3420] ^ layer2_out[3421];
     layer3_out[262] <= ~layer2_out[717];
     layer3_out[263] <= ~layer2_out[4151];
     layer3_out[264] <= ~layer2_out[6065];
     layer3_out[265] <= ~layer2_out[4262];
     layer3_out[266] <= layer2_out[2216] & layer2_out[2217];
     layer3_out[267] <= layer2_out[153] & ~layer2_out[152];
     layer3_out[268] <= layer2_out[9223];
     layer3_out[269] <= layer2_out[8180] & ~layer2_out[8181];
     layer3_out[270] <= layer2_out[9855];
     layer3_out[271] <= layer2_out[3528] & ~layer2_out[3529];
     layer3_out[272] <= layer2_out[8560];
     layer3_out[273] <= layer2_out[8366];
     layer3_out[274] <= layer2_out[10609];
     layer3_out[275] <= ~layer2_out[8697];
     layer3_out[276] <= ~layer2_out[908];
     layer3_out[277] <= layer2_out[1606] ^ layer2_out[1607];
     layer3_out[278] <= layer2_out[3676];
     layer3_out[279] <= ~(layer2_out[1174] & layer2_out[1175]);
     layer3_out[280] <= ~layer2_out[1247];
     layer3_out[281] <= ~(layer2_out[6197] | layer2_out[6198]);
     layer3_out[282] <= layer2_out[3955] & ~layer2_out[3956];
     layer3_out[283] <= ~layer2_out[11992];
     layer3_out[284] <= layer2_out[8531] & ~layer2_out[8530];
     layer3_out[285] <= layer2_out[4612];
     layer3_out[286] <= ~layer2_out[9251];
     layer3_out[287] <= ~layer2_out[7289];
     layer3_out[288] <= ~layer2_out[3007];
     layer3_out[289] <= layer2_out[6549];
     layer3_out[290] <= layer2_out[2569] & ~layer2_out[2570];
     layer3_out[291] <= ~(layer2_out[9429] | layer2_out[9430]);
     layer3_out[292] <= ~layer2_out[8660];
     layer3_out[293] <= ~layer2_out[1237] | layer2_out[1238];
     layer3_out[294] <= layer2_out[7473] & ~layer2_out[7474];
     layer3_out[295] <= layer2_out[5921];
     layer3_out[296] <= layer2_out[6263] & ~layer2_out[6262];
     layer3_out[297] <= ~(layer2_out[4577] | layer2_out[4578]);
     layer3_out[298] <= ~(layer2_out[7140] | layer2_out[7141]);
     layer3_out[299] <= layer2_out[5635] & layer2_out[5636];
     layer3_out[300] <= layer2_out[7878];
     layer3_out[301] <= layer2_out[8980] & layer2_out[8981];
     layer3_out[302] <= layer2_out[5496] & ~layer2_out[5495];
     layer3_out[303] <= layer2_out[168] & layer2_out[169];
     layer3_out[304] <= ~layer2_out[942];
     layer3_out[305] <= layer2_out[7009];
     layer3_out[306] <= layer2_out[731] & ~layer2_out[730];
     layer3_out[307] <= layer2_out[1670];
     layer3_out[308] <= ~layer2_out[11853];
     layer3_out[309] <= layer2_out[6022] & ~layer2_out[6023];
     layer3_out[310] <= ~(layer2_out[4791] ^ layer2_out[4792]);
     layer3_out[311] <= layer2_out[8790] & ~layer2_out[8789];
     layer3_out[312] <= layer2_out[3103];
     layer3_out[313] <= ~layer2_out[1034];
     layer3_out[314] <= layer2_out[3982];
     layer3_out[315] <= ~(layer2_out[552] & layer2_out[553]);
     layer3_out[316] <= layer2_out[7129] ^ layer2_out[7130];
     layer3_out[317] <= layer2_out[10810];
     layer3_out[318] <= layer2_out[4244] & ~layer2_out[4243];
     layer3_out[319] <= ~(layer2_out[7506] | layer2_out[7507]);
     layer3_out[320] <= layer2_out[9331] & ~layer2_out[9332];
     layer3_out[321] <= layer2_out[496] | layer2_out[497];
     layer3_out[322] <= ~layer2_out[7523] | layer2_out[7522];
     layer3_out[323] <= ~layer2_out[6502] | layer2_out[6501];
     layer3_out[324] <= ~layer2_out[6682];
     layer3_out[325] <= layer2_out[2545] & layer2_out[2546];
     layer3_out[326] <= layer2_out[7675];
     layer3_out[327] <= ~layer2_out[2764];
     layer3_out[328] <= layer2_out[4086] & layer2_out[4087];
     layer3_out[329] <= ~(layer2_out[8537] ^ layer2_out[8538]);
     layer3_out[330] <= ~layer2_out[11403];
     layer3_out[331] <= layer2_out[1177] | layer2_out[1178];
     layer3_out[332] <= layer2_out[11414] & ~layer2_out[11415];
     layer3_out[333] <= ~(layer2_out[4635] ^ layer2_out[4636]);
     layer3_out[334] <= ~(layer2_out[2819] | layer2_out[2820]);
     layer3_out[335] <= ~layer2_out[8498];
     layer3_out[336] <= ~(layer2_out[9994] & layer2_out[9995]);
     layer3_out[337] <= layer2_out[345] & ~layer2_out[346];
     layer3_out[338] <= layer2_out[2940] & layer2_out[2941];
     layer3_out[339] <= ~layer2_out[4872] | layer2_out[4871];
     layer3_out[340] <= layer2_out[10760];
     layer3_out[341] <= ~layer2_out[321];
     layer3_out[342] <= layer2_out[2571] & ~layer2_out[2570];
     layer3_out[343] <= layer2_out[9730] & ~layer2_out[9731];
     layer3_out[344] <= ~layer2_out[2103];
     layer3_out[345] <= ~(layer2_out[10575] ^ layer2_out[10576]);
     layer3_out[346] <= ~layer2_out[7954];
     layer3_out[347] <= ~(layer2_out[5553] ^ layer2_out[5554]);
     layer3_out[348] <= ~layer2_out[6167] | layer2_out[6166];
     layer3_out[349] <= ~(layer2_out[10340] | layer2_out[10341]);
     layer3_out[350] <= ~(layer2_out[3734] ^ layer2_out[3735]);
     layer3_out[351] <= layer2_out[4221] & ~layer2_out[4220];
     layer3_out[352] <= layer2_out[6831] & ~layer2_out[6830];
     layer3_out[353] <= ~layer2_out[8600];
     layer3_out[354] <= layer2_out[10756] & ~layer2_out[10755];
     layer3_out[355] <= ~(layer2_out[1733] | layer2_out[1734]);
     layer3_out[356] <= ~layer2_out[370];
     layer3_out[357] <= layer2_out[2539] & layer2_out[2540];
     layer3_out[358] <= ~(layer2_out[622] ^ layer2_out[623]);
     layer3_out[359] <= layer2_out[1580] ^ layer2_out[1581];
     layer3_out[360] <= ~layer2_out[4712] | layer2_out[4713];
     layer3_out[361] <= layer2_out[10848] & layer2_out[10849];
     layer3_out[362] <= layer2_out[11084] & layer2_out[11085];
     layer3_out[363] <= layer2_out[7462];
     layer3_out[364] <= layer2_out[11328] | layer2_out[11329];
     layer3_out[365] <= layer2_out[6074] & ~layer2_out[6073];
     layer3_out[366] <= ~layer2_out[2142];
     layer3_out[367] <= ~(layer2_out[10850] | layer2_out[10851]);
     layer3_out[368] <= layer2_out[7058];
     layer3_out[369] <= layer2_out[2133] & ~layer2_out[2132];
     layer3_out[370] <= layer2_out[3323] & layer2_out[3324];
     layer3_out[371] <= layer2_out[1110] & ~layer2_out[1111];
     layer3_out[372] <= ~(layer2_out[6560] | layer2_out[6561]);
     layer3_out[373] <= ~layer2_out[3581];
     layer3_out[374] <= layer2_out[8652];
     layer3_out[375] <= ~layer2_out[11508] | layer2_out[11509];
     layer3_out[376] <= layer2_out[2368];
     layer3_out[377] <= ~(layer2_out[853] & layer2_out[854]);
     layer3_out[378] <= layer2_out[11110] ^ layer2_out[11111];
     layer3_out[379] <= layer2_out[1825];
     layer3_out[380] <= ~layer2_out[5148] | layer2_out[5149];
     layer3_out[381] <= layer2_out[6583];
     layer3_out[382] <= layer2_out[10232];
     layer3_out[383] <= ~layer2_out[2825] | layer2_out[2826];
     layer3_out[384] <= ~layer2_out[10428];
     layer3_out[385] <= ~layer2_out[9323];
     layer3_out[386] <= layer2_out[7718];
     layer3_out[387] <= ~layer2_out[2169];
     layer3_out[388] <= layer2_out[9590] & layer2_out[9591];
     layer3_out[389] <= ~layer2_out[6446];
     layer3_out[390] <= layer2_out[10977] & ~layer2_out[10976];
     layer3_out[391] <= ~layer2_out[7121] | layer2_out[7120];
     layer3_out[392] <= layer2_out[2897] & ~layer2_out[2898];
     layer3_out[393] <= layer2_out[11175];
     layer3_out[394] <= layer2_out[2854] & ~layer2_out[2853];
     layer3_out[395] <= ~(layer2_out[10946] | layer2_out[10947]);
     layer3_out[396] <= layer2_out[9502];
     layer3_out[397] <= ~(layer2_out[4066] ^ layer2_out[4067]);
     layer3_out[398] <= ~layer2_out[5065];
     layer3_out[399] <= layer2_out[10646] ^ layer2_out[10647];
     layer3_out[400] <= ~layer2_out[3791] | layer2_out[3792];
     layer3_out[401] <= ~layer2_out[525];
     layer3_out[402] <= layer2_out[2335];
     layer3_out[403] <= layer2_out[6983];
     layer3_out[404] <= ~(layer2_out[1003] ^ layer2_out[1004]);
     layer3_out[405] <= ~layer2_out[2845] | layer2_out[2844];
     layer3_out[406] <= layer2_out[10963] & ~layer2_out[10962];
     layer3_out[407] <= layer2_out[5647];
     layer3_out[408] <= layer2_out[7210];
     layer3_out[409] <= layer2_out[6462];
     layer3_out[410] <= layer2_out[7985];
     layer3_out[411] <= layer2_out[11765];
     layer3_out[412] <= ~layer2_out[11754];
     layer3_out[413] <= layer2_out[4928] | layer2_out[4929];
     layer3_out[414] <= layer2_out[905] & ~layer2_out[904];
     layer3_out[415] <= layer2_out[1305];
     layer3_out[416] <= layer2_out[5026] & layer2_out[5027];
     layer3_out[417] <= ~(layer2_out[3029] ^ layer2_out[3030]);
     layer3_out[418] <= ~layer2_out[11180];
     layer3_out[419] <= layer2_out[5005];
     layer3_out[420] <= layer2_out[8193] & ~layer2_out[8194];
     layer3_out[421] <= ~layer2_out[3885] | layer2_out[3884];
     layer3_out[422] <= ~layer2_out[3731] | layer2_out[3732];
     layer3_out[423] <= layer2_out[3331];
     layer3_out[424] <= layer2_out[1239] & layer2_out[1240];
     layer3_out[425] <= ~layer2_out[4576];
     layer3_out[426] <= layer2_out[807];
     layer3_out[427] <= ~(layer2_out[612] & layer2_out[613]);
     layer3_out[428] <= layer2_out[10174];
     layer3_out[429] <= ~(layer2_out[1868] | layer2_out[1869]);
     layer3_out[430] <= layer2_out[87] & layer2_out[88];
     layer3_out[431] <= ~layer2_out[7854];
     layer3_out[432] <= ~layer2_out[7031];
     layer3_out[433] <= layer2_out[6210];
     layer3_out[434] <= layer2_out[11522];
     layer3_out[435] <= layer2_out[9037];
     layer3_out[436] <= layer2_out[86] & ~layer2_out[85];
     layer3_out[437] <= ~(layer2_out[8508] ^ layer2_out[8509]);
     layer3_out[438] <= ~layer2_out[9179];
     layer3_out[439] <= ~(layer2_out[10905] ^ layer2_out[10906]);
     layer3_out[440] <= layer2_out[2044] & layer2_out[2045];
     layer3_out[441] <= layer2_out[7362];
     layer3_out[442] <= ~(layer2_out[3909] ^ layer2_out[3910]);
     layer3_out[443] <= layer2_out[2837] ^ layer2_out[2838];
     layer3_out[444] <= layer2_out[5526] & ~layer2_out[5527];
     layer3_out[445] <= layer2_out[7178] & ~layer2_out[7179];
     layer3_out[446] <= ~(layer2_out[3358] | layer2_out[3359]);
     layer3_out[447] <= ~(layer2_out[11467] ^ layer2_out[11468]);
     layer3_out[448] <= ~layer2_out[10152];
     layer3_out[449] <= layer2_out[11007] & ~layer2_out[11006];
     layer3_out[450] <= ~(layer2_out[5770] ^ layer2_out[5771]);
     layer3_out[451] <= layer2_out[9028];
     layer3_out[452] <= ~layer2_out[772];
     layer3_out[453] <= layer2_out[7654];
     layer3_out[454] <= ~layer2_out[2080];
     layer3_out[455] <= ~(layer2_out[6977] & layer2_out[6978]);
     layer3_out[456] <= ~layer2_out[11320] | layer2_out[11321];
     layer3_out[457] <= ~(layer2_out[11113] | layer2_out[11114]);
     layer3_out[458] <= ~layer2_out[8731] | layer2_out[8732];
     layer3_out[459] <= ~layer2_out[6643];
     layer3_out[460] <= layer2_out[1286] & ~layer2_out[1285];
     layer3_out[461] <= layer2_out[9303];
     layer3_out[462] <= layer2_out[10619];
     layer3_out[463] <= ~(layer2_out[84] & layer2_out[85]);
     layer3_out[464] <= layer2_out[2893];
     layer3_out[465] <= layer2_out[10961] & ~layer2_out[10960];
     layer3_out[466] <= ~layer2_out[1343];
     layer3_out[467] <= ~layer2_out[8399];
     layer3_out[468] <= ~(layer2_out[11861] | layer2_out[11862]);
     layer3_out[469] <= ~(layer2_out[214] | layer2_out[215]);
     layer3_out[470] <= layer2_out[2698];
     layer3_out[471] <= layer2_out[1816] & ~layer2_out[1817];
     layer3_out[472] <= ~(layer2_out[8321] & layer2_out[8322]);
     layer3_out[473] <= layer2_out[4392] & layer2_out[4393];
     layer3_out[474] <= layer2_out[1009] | layer2_out[1010];
     layer3_out[475] <= layer2_out[2929];
     layer3_out[476] <= layer2_out[8937];
     layer3_out[477] <= layer2_out[9317] & ~layer2_out[9318];
     layer3_out[478] <= ~(layer2_out[7387] | layer2_out[7388]);
     layer3_out[479] <= ~layer2_out[9554];
     layer3_out[480] <= layer2_out[4884] & ~layer2_out[4885];
     layer3_out[481] <= ~layer2_out[4499] | layer2_out[4500];
     layer3_out[482] <= ~(layer2_out[6753] ^ layer2_out[6754]);
     layer3_out[483] <= ~(layer2_out[2578] ^ layer2_out[2579]);
     layer3_out[484] <= layer2_out[556];
     layer3_out[485] <= ~layer2_out[4043];
     layer3_out[486] <= layer2_out[8437] & layer2_out[8438];
     layer3_out[487] <= ~layer2_out[9613];
     layer3_out[488] <= ~layer2_out[3870];
     layer3_out[489] <= ~layer2_out[6344] | layer2_out[6343];
     layer3_out[490] <= layer2_out[2861];
     layer3_out[491] <= ~(layer2_out[7802] & layer2_out[7803]);
     layer3_out[492] <= layer2_out[2484];
     layer3_out[493] <= layer2_out[690];
     layer3_out[494] <= ~layer2_out[3349];
     layer3_out[495] <= layer2_out[9605];
     layer3_out[496] <= layer2_out[2242] & ~layer2_out[2243];
     layer3_out[497] <= layer2_out[10849] & ~layer2_out[10850];
     layer3_out[498] <= ~layer2_out[4318];
     layer3_out[499] <= ~layer2_out[2071];
     layer3_out[500] <= layer2_out[11259] & ~layer2_out[11258];
     layer3_out[501] <= layer2_out[6992] & ~layer2_out[6991];
     layer3_out[502] <= layer2_out[299];
     layer3_out[503] <= ~layer2_out[5015];
     layer3_out[504] <= ~layer2_out[9452] | layer2_out[9451];
     layer3_out[505] <= ~(layer2_out[694] ^ layer2_out[695]);
     layer3_out[506] <= layer2_out[2826];
     layer3_out[507] <= ~layer2_out[225];
     layer3_out[508] <= ~layer2_out[2401];
     layer3_out[509] <= ~(layer2_out[7966] | layer2_out[7967]);
     layer3_out[510] <= layer2_out[4473] & layer2_out[4474];
     layer3_out[511] <= layer2_out[592] & ~layer2_out[591];
     layer3_out[512] <= layer2_out[8994] & layer2_out[8995];
     layer3_out[513] <= ~(layer2_out[6941] ^ layer2_out[6942]);
     layer3_out[514] <= layer2_out[3701] & layer2_out[3702];
     layer3_out[515] <= ~layer2_out[10142];
     layer3_out[516] <= layer2_out[5165] & ~layer2_out[5164];
     layer3_out[517] <= ~(layer2_out[10777] ^ layer2_out[10778]);
     layer3_out[518] <= layer2_out[1271] & ~layer2_out[1270];
     layer3_out[519] <= ~layer2_out[9736];
     layer3_out[520] <= layer2_out[8142] & layer2_out[8143];
     layer3_out[521] <= ~layer2_out[4118];
     layer3_out[522] <= layer2_out[2761] ^ layer2_out[2762];
     layer3_out[523] <= ~layer2_out[3156];
     layer3_out[524] <= ~layer2_out[1609];
     layer3_out[525] <= layer2_out[5876] ^ layer2_out[5877];
     layer3_out[526] <= ~layer2_out[5118] | layer2_out[5117];
     layer3_out[527] <= layer2_out[3600] & ~layer2_out[3599];
     layer3_out[528] <= ~layer2_out[10424];
     layer3_out[529] <= ~layer2_out[1092];
     layer3_out[530] <= ~layer2_out[427];
     layer3_out[531] <= ~layer2_out[2051];
     layer3_out[532] <= layer2_out[4395] & ~layer2_out[4396];
     layer3_out[533] <= layer2_out[6451] ^ layer2_out[6452];
     layer3_out[534] <= layer2_out[8240] ^ layer2_out[8241];
     layer3_out[535] <= layer2_out[10425];
     layer3_out[536] <= ~(layer2_out[10112] ^ layer2_out[10113]);
     layer3_out[537] <= ~layer2_out[11686];
     layer3_out[538] <= ~layer2_out[2391];
     layer3_out[539] <= layer2_out[3016] & layer2_out[3017];
     layer3_out[540] <= layer2_out[5325] & layer2_out[5326];
     layer3_out[541] <= layer2_out[10673] & ~layer2_out[10672];
     layer3_out[542] <= layer2_out[11139] ^ layer2_out[11140];
     layer3_out[543] <= layer2_out[8611] & ~layer2_out[8610];
     layer3_out[544] <= ~layer2_out[11665] | layer2_out[11664];
     layer3_out[545] <= layer2_out[1915];
     layer3_out[546] <= ~layer2_out[4800] | layer2_out[4801];
     layer3_out[547] <= ~(layer2_out[2308] ^ layer2_out[2309]);
     layer3_out[548] <= layer2_out[8129];
     layer3_out[549] <= ~layer2_out[6426] | layer2_out[6427];
     layer3_out[550] <= ~(layer2_out[4774] | layer2_out[4775]);
     layer3_out[551] <= ~layer2_out[4562];
     layer3_out[552] <= layer2_out[3613] & ~layer2_out[3612];
     layer3_out[553] <= ~layer2_out[10160];
     layer3_out[554] <= ~(layer2_out[5106] | layer2_out[5107]);
     layer3_out[555] <= layer2_out[8332];
     layer3_out[556] <= layer2_out[9357];
     layer3_out[557] <= layer2_out[10295];
     layer3_out[558] <= ~(layer2_out[10001] | layer2_out[10002]);
     layer3_out[559] <= layer2_out[7350] & ~layer2_out[7351];
     layer3_out[560] <= layer2_out[5576] ^ layer2_out[5577];
     layer3_out[561] <= ~(layer2_out[1423] | layer2_out[1424]);
     layer3_out[562] <= layer2_out[4390];
     layer3_out[563] <= layer2_out[6823] & ~layer2_out[6824];
     layer3_out[564] <= layer2_out[10459];
     layer3_out[565] <= ~layer2_out[8586] | layer2_out[8587];
     layer3_out[566] <= ~(layer2_out[6975] ^ layer2_out[6976]);
     layer3_out[567] <= layer2_out[2675];
     layer3_out[568] <= ~layer2_out[10783];
     layer3_out[569] <= ~layer2_out[9350];
     layer3_out[570] <= layer2_out[9789] & ~layer2_out[9788];
     layer3_out[571] <= layer2_out[7317] ^ layer2_out[7318];
     layer3_out[572] <= ~layer2_out[5554] | layer2_out[5555];
     layer3_out[573] <= layer2_out[9857];
     layer3_out[574] <= ~(layer2_out[348] ^ layer2_out[349]);
     layer3_out[575] <= layer2_out[234] & ~layer2_out[235];
     layer3_out[576] <= layer2_out[769];
     layer3_out[577] <= layer2_out[4874] | layer2_out[4875];
     layer3_out[578] <= ~(layer2_out[119] | layer2_out[120]);
     layer3_out[579] <= layer2_out[11328] & ~layer2_out[11327];
     layer3_out[580] <= ~(layer2_out[2794] ^ layer2_out[2795]);
     layer3_out[581] <= ~layer2_out[11520] | layer2_out[11519];
     layer3_out[582] <= layer2_out[916] & ~layer2_out[917];
     layer3_out[583] <= layer2_out[3411];
     layer3_out[584] <= layer2_out[5672] & ~layer2_out[5673];
     layer3_out[585] <= layer2_out[2201];
     layer3_out[586] <= ~(layer2_out[5537] & layer2_out[5538]);
     layer3_out[587] <= layer2_out[9236];
     layer3_out[588] <= layer2_out[3808] & ~layer2_out[3809];
     layer3_out[589] <= layer2_out[7836] & layer2_out[7837];
     layer3_out[590] <= ~layer2_out[9174] | layer2_out[9175];
     layer3_out[591] <= layer2_out[10846];
     layer3_out[592] <= ~layer2_out[9638];
     layer3_out[593] <= ~(layer2_out[7326] ^ layer2_out[7327]);
     layer3_out[594] <= ~layer2_out[4142];
     layer3_out[595] <= layer2_out[9104];
     layer3_out[596] <= layer2_out[1950] ^ layer2_out[1951];
     layer3_out[597] <= ~layer2_out[6843];
     layer3_out[598] <= ~(layer2_out[5192] ^ layer2_out[5193]);
     layer3_out[599] <= ~layer2_out[3282];
     layer3_out[600] <= layer2_out[3167];
     layer3_out[601] <= ~(layer2_out[10791] & layer2_out[10792]);
     layer3_out[602] <= ~layer2_out[3583];
     layer3_out[603] <= ~(layer2_out[2945] ^ layer2_out[2946]);
     layer3_out[604] <= ~layer2_out[7091] | layer2_out[7090];
     layer3_out[605] <= ~layer2_out[6468] | layer2_out[6467];
     layer3_out[606] <= layer2_out[8937];
     layer3_out[607] <= ~(layer2_out[3142] & layer2_out[3143]);
     layer3_out[608] <= layer2_out[2724] ^ layer2_out[2725];
     layer3_out[609] <= layer2_out[11498];
     layer3_out[610] <= layer2_out[659] & ~layer2_out[660];
     layer3_out[611] <= layer2_out[7926];
     layer3_out[612] <= ~layer2_out[819];
     layer3_out[613] <= ~layer2_out[1132];
     layer3_out[614] <= layer2_out[11252] ^ layer2_out[11253];
     layer3_out[615] <= layer2_out[4821];
     layer3_out[616] <= layer2_out[995] & layer2_out[996];
     layer3_out[617] <= ~layer2_out[6115] | layer2_out[6114];
     layer3_out[618] <= layer2_out[299];
     layer3_out[619] <= ~layer2_out[9609];
     layer3_out[620] <= layer2_out[3050] ^ layer2_out[3051];
     layer3_out[621] <= ~(layer2_out[4533] & layer2_out[4534]);
     layer3_out[622] <= layer2_out[1180];
     layer3_out[623] <= layer2_out[9049];
     layer3_out[624] <= ~(layer2_out[4542] | layer2_out[4543]);
     layer3_out[625] <= layer2_out[8085] & ~layer2_out[8086];
     layer3_out[626] <= layer2_out[466];
     layer3_out[627] <= ~layer2_out[7896];
     layer3_out[628] <= layer2_out[6252] ^ layer2_out[6253];
     layer3_out[629] <= ~layer2_out[1302] | layer2_out[1301];
     layer3_out[630] <= ~(layer2_out[8696] | layer2_out[8697]);
     layer3_out[631] <= ~(layer2_out[878] | layer2_out[879]);
     layer3_out[632] <= layer2_out[4793] & ~layer2_out[4794];
     layer3_out[633] <= layer2_out[3509] ^ layer2_out[3510];
     layer3_out[634] <= ~(layer2_out[9744] & layer2_out[9745]);
     layer3_out[635] <= layer2_out[3416];
     layer3_out[636] <= layer2_out[5241] & ~layer2_out[5242];
     layer3_out[637] <= ~(layer2_out[6698] ^ layer2_out[6699]);
     layer3_out[638] <= layer2_out[4669];
     layer3_out[639] <= ~(layer2_out[6198] | layer2_out[6199]);
     layer3_out[640] <= layer2_out[9998];
     layer3_out[641] <= layer2_out[4238] & ~layer2_out[4239];
     layer3_out[642] <= layer2_out[10365] & layer2_out[10366];
     layer3_out[643] <= ~layer2_out[6083];
     layer3_out[644] <= layer2_out[7773];
     layer3_out[645] <= ~(layer2_out[7955] | layer2_out[7956]);
     layer3_out[646] <= ~(layer2_out[2106] & layer2_out[2107]);
     layer3_out[647] <= ~(layer2_out[6980] & layer2_out[6981]);
     layer3_out[648] <= ~layer2_out[7233] | layer2_out[7232];
     layer3_out[649] <= layer2_out[6593] & ~layer2_out[6592];
     layer3_out[650] <= layer2_out[7974];
     layer3_out[651] <= layer2_out[9632];
     layer3_out[652] <= layer2_out[5644] & layer2_out[5645];
     layer3_out[653] <= layer2_out[10943] & ~layer2_out[10944];
     layer3_out[654] <= layer2_out[3100] & ~layer2_out[3101];
     layer3_out[655] <= ~layer2_out[4939];
     layer3_out[656] <= ~layer2_out[174];
     layer3_out[657] <= layer2_out[2650];
     layer3_out[658] <= ~layer2_out[4683];
     layer3_out[659] <= layer2_out[1410];
     layer3_out[660] <= ~(layer2_out[9624] | layer2_out[9625]);
     layer3_out[661] <= layer2_out[7390];
     layer3_out[662] <= layer2_out[7701] | layer2_out[7702];
     layer3_out[663] <= layer2_out[1197] ^ layer2_out[1198];
     layer3_out[664] <= layer2_out[3368];
     layer3_out[665] <= layer2_out[4672] & layer2_out[4673];
     layer3_out[666] <= ~layer2_out[4814] | layer2_out[4815];
     layer3_out[667] <= layer2_out[4821];
     layer3_out[668] <= ~layer2_out[3098];
     layer3_out[669] <= layer2_out[4214] ^ layer2_out[4215];
     layer3_out[670] <= layer2_out[8313] ^ layer2_out[8314];
     layer3_out[671] <= layer2_out[11762];
     layer3_out[672] <= layer2_out[9227] & ~layer2_out[9228];
     layer3_out[673] <= ~layer2_out[853] | layer2_out[852];
     layer3_out[674] <= ~(layer2_out[7324] | layer2_out[7325]);
     layer3_out[675] <= layer2_out[7625];
     layer3_out[676] <= layer2_out[2950];
     layer3_out[677] <= ~layer2_out[8571];
     layer3_out[678] <= ~layer2_out[5539];
     layer3_out[679] <= layer2_out[4830] | layer2_out[4831];
     layer3_out[680] <= layer2_out[208];
     layer3_out[681] <= ~(layer2_out[0] & layer2_out[2]);
     layer3_out[682] <= layer2_out[10509] | layer2_out[10510];
     layer3_out[683] <= layer2_out[1140];
     layer3_out[684] <= layer2_out[5674];
     layer3_out[685] <= layer2_out[10915] & layer2_out[10916];
     layer3_out[686] <= layer2_out[1134];
     layer3_out[687] <= layer2_out[5976] | layer2_out[5977];
     layer3_out[688] <= layer2_out[4917];
     layer3_out[689] <= layer2_out[6090] & ~layer2_out[6091];
     layer3_out[690] <= layer2_out[11590] ^ layer2_out[11591];
     layer3_out[691] <= ~layer2_out[9807] | layer2_out[9808];
     layer3_out[692] <= ~(layer2_out[1055] ^ layer2_out[1056]);
     layer3_out[693] <= ~(layer2_out[4860] & layer2_out[4861]);
     layer3_out[694] <= layer2_out[1241];
     layer3_out[695] <= layer2_out[1311] ^ layer2_out[1312];
     layer3_out[696] <= ~(layer2_out[4040] ^ layer2_out[4041]);
     layer3_out[697] <= ~layer2_out[7545];
     layer3_out[698] <= ~(layer2_out[8035] | layer2_out[8036]);
     layer3_out[699] <= ~layer2_out[9842];
     layer3_out[700] <= ~(layer2_out[2093] ^ layer2_out[2094]);
     layer3_out[701] <= layer2_out[4964] | layer2_out[4965];
     layer3_out[702] <= ~(layer2_out[310] ^ layer2_out[311]);
     layer3_out[703] <= layer2_out[5964] | layer2_out[5965];
     layer3_out[704] <= ~layer2_out[11043];
     layer3_out[705] <= ~(layer2_out[10695] | layer2_out[10696]);
     layer3_out[706] <= layer2_out[9774];
     layer3_out[707] <= layer2_out[7961] & layer2_out[7962];
     layer3_out[708] <= ~(layer2_out[2513] | layer2_out[2514]);
     layer3_out[709] <= ~layer2_out[3844];
     layer3_out[710] <= layer2_out[6248] ^ layer2_out[6249];
     layer3_out[711] <= ~layer2_out[472];
     layer3_out[712] <= layer2_out[4657];
     layer3_out[713] <= ~layer2_out[854];
     layer3_out[714] <= layer2_out[2596];
     layer3_out[715] <= layer2_out[10883];
     layer3_out[716] <= ~layer2_out[4028];
     layer3_out[717] <= layer2_out[10489] & layer2_out[10490];
     layer3_out[718] <= ~(layer2_out[1712] ^ layer2_out[1713]);
     layer3_out[719] <= ~layer2_out[6094] | layer2_out[6095];
     layer3_out[720] <= layer2_out[3275];
     layer3_out[721] <= ~(layer2_out[3314] ^ layer2_out[3315]);
     layer3_out[722] <= ~layer2_out[8591];
     layer3_out[723] <= ~layer2_out[7031];
     layer3_out[724] <= layer2_out[8549] ^ layer2_out[8550];
     layer3_out[725] <= layer2_out[5449] ^ layer2_out[5450];
     layer3_out[726] <= ~layer2_out[9139];
     layer3_out[727] <= ~layer2_out[3545];
     layer3_out[728] <= layer2_out[10660] | layer2_out[10661];
     layer3_out[729] <= ~layer2_out[11579];
     layer3_out[730] <= ~layer2_out[764];
     layer3_out[731] <= ~(layer2_out[11081] | layer2_out[11082]);
     layer3_out[732] <= ~(layer2_out[6808] | layer2_out[6809]);
     layer3_out[733] <= ~layer2_out[10858] | layer2_out[10857];
     layer3_out[734] <= ~layer2_out[3774];
     layer3_out[735] <= ~layer2_out[10052];
     layer3_out[736] <= layer2_out[2523] ^ layer2_out[2524];
     layer3_out[737] <= layer2_out[7105];
     layer3_out[738] <= layer2_out[5982];
     layer3_out[739] <= layer2_out[4627] | layer2_out[4628];
     layer3_out[740] <= layer2_out[11859];
     layer3_out[741] <= layer2_out[8218];
     layer3_out[742] <= ~layer2_out[7982];
     layer3_out[743] <= ~(layer2_out[10694] | layer2_out[10695]);
     layer3_out[744] <= layer2_out[151];
     layer3_out[745] <= layer2_out[111];
     layer3_out[746] <= layer2_out[1272];
     layer3_out[747] <= layer2_out[1980] ^ layer2_out[1981];
     layer3_out[748] <= layer2_out[11600];
     layer3_out[749] <= ~(layer2_out[693] & layer2_out[694]);
     layer3_out[750] <= ~layer2_out[4330];
     layer3_out[751] <= layer2_out[7868] & layer2_out[7869];
     layer3_out[752] <= layer2_out[10326] & ~layer2_out[10327];
     layer3_out[753] <= layer2_out[937];
     layer3_out[754] <= layer2_out[4422];
     layer3_out[755] <= layer2_out[295] & ~layer2_out[296];
     layer3_out[756] <= layer2_out[1990] & ~layer2_out[1991];
     layer3_out[757] <= layer2_out[1253] & layer2_out[1254];
     layer3_out[758] <= layer2_out[7077] ^ layer2_out[7078];
     layer3_out[759] <= layer2_out[7769];
     layer3_out[760] <= ~(layer2_out[4260] ^ layer2_out[4261]);
     layer3_out[761] <= layer2_out[2913] & ~layer2_out[2914];
     layer3_out[762] <= layer2_out[1531] & ~layer2_out[1530];
     layer3_out[763] <= layer2_out[9478];
     layer3_out[764] <= layer2_out[9192] & layer2_out[9193];
     layer3_out[765] <= layer2_out[3949];
     layer3_out[766] <= ~layer2_out[3760] | layer2_out[3759];
     layer3_out[767] <= layer2_out[9747];
     layer3_out[768] <= ~layer2_out[2274] | layer2_out[2273];
     layer3_out[769] <= ~(layer2_out[7033] & layer2_out[7034]);
     layer3_out[770] <= layer2_out[2484];
     layer3_out[771] <= ~layer2_out[7485];
     layer3_out[772] <= layer2_out[4418];
     layer3_out[773] <= ~layer2_out[9389];
     layer3_out[774] <= ~layer2_out[3247];
     layer3_out[775] <= ~layer2_out[10359] | layer2_out[10358];
     layer3_out[776] <= ~layer2_out[10079];
     layer3_out[777] <= layer2_out[6562] & ~layer2_out[6563];
     layer3_out[778] <= layer2_out[7480] & layer2_out[7481];
     layer3_out[779] <= ~(layer2_out[9332] | layer2_out[9333]);
     layer3_out[780] <= layer2_out[9653] ^ layer2_out[9654];
     layer3_out[781] <= layer2_out[6645];
     layer3_out[782] <= ~layer2_out[10799];
     layer3_out[783] <= ~(layer2_out[11923] | layer2_out[11924]);
     layer3_out[784] <= layer2_out[7654];
     layer3_out[785] <= layer2_out[244] & layer2_out[245];
     layer3_out[786] <= ~(layer2_out[8911] | layer2_out[8912]);
     layer3_out[787] <= ~layer2_out[4189];
     layer3_out[788] <= ~(layer2_out[3543] | layer2_out[3544]);
     layer3_out[789] <= ~layer2_out[6312];
     layer3_out[790] <= ~layer2_out[5719];
     layer3_out[791] <= layer2_out[4235];
     layer3_out[792] <= layer2_out[2242];
     layer3_out[793] <= layer2_out[8863] & ~layer2_out[8862];
     layer3_out[794] <= ~layer2_out[3173];
     layer3_out[795] <= layer2_out[6415] ^ layer2_out[6416];
     layer3_out[796] <= ~(layer2_out[700] | layer2_out[701]);
     layer3_out[797] <= layer2_out[11096];
     layer3_out[798] <= ~layer2_out[1096] | layer2_out[1097];
     layer3_out[799] <= layer2_out[797] & ~layer2_out[796];
     layer3_out[800] <= ~layer2_out[3351];
     layer3_out[801] <= ~(layer2_out[1059] & layer2_out[1060]);
     layer3_out[802] <= ~layer2_out[10841] | layer2_out[10842];
     layer3_out[803] <= ~layer2_out[4683];
     layer3_out[804] <= layer2_out[5286];
     layer3_out[805] <= ~layer2_out[7149] | layer2_out[7150];
     layer3_out[806] <= layer2_out[9728] ^ layer2_out[9729];
     layer3_out[807] <= ~(layer2_out[11935] | layer2_out[11936]);
     layer3_out[808] <= layer2_out[11866];
     layer3_out[809] <= ~layer2_out[10533];
     layer3_out[810] <= layer2_out[9590] & ~layer2_out[9589];
     layer3_out[811] <= layer2_out[1120];
     layer3_out[812] <= layer2_out[5104] ^ layer2_out[5105];
     layer3_out[813] <= layer2_out[10250] ^ layer2_out[10251];
     layer3_out[814] <= layer2_out[7984] | layer2_out[7985];
     layer3_out[815] <= layer2_out[2901];
     layer3_out[816] <= ~(layer2_out[11245] ^ layer2_out[11246]);
     layer3_out[817] <= layer2_out[2958];
     layer3_out[818] <= layer2_out[4152] & ~layer2_out[4151];
     layer3_out[819] <= layer2_out[6061];
     layer3_out[820] <= ~layer2_out[8556];
     layer3_out[821] <= ~(layer2_out[7852] | layer2_out[7853]);
     layer3_out[822] <= ~(layer2_out[2363] | layer2_out[2364]);
     layer3_out[823] <= layer2_out[4886] & ~layer2_out[4885];
     layer3_out[824] <= layer2_out[3659];
     layer3_out[825] <= layer2_out[905];
     layer3_out[826] <= ~(layer2_out[10788] | layer2_out[10789]);
     layer3_out[827] <= ~(layer2_out[6744] | layer2_out[6745]);
     layer3_out[828] <= layer2_out[8326];
     layer3_out[829] <= ~layer2_out[8174];
     layer3_out[830] <= ~layer2_out[6776];
     layer3_out[831] <= layer2_out[4809] & ~layer2_out[4810];
     layer3_out[832] <= ~(layer2_out[11569] & layer2_out[11570]);
     layer3_out[833] <= layer2_out[3908];
     layer3_out[834] <= layer2_out[10926];
     layer3_out[835] <= layer2_out[7054];
     layer3_out[836] <= layer2_out[3371] | layer2_out[3372];
     layer3_out[837] <= layer2_out[4664] | layer2_out[4665];
     layer3_out[838] <= layer2_out[7910] & layer2_out[7911];
     layer3_out[839] <= ~(layer2_out[5289] | layer2_out[5290]);
     layer3_out[840] <= layer2_out[3745] & ~layer2_out[3746];
     layer3_out[841] <= ~(layer2_out[6708] | layer2_out[6709]);
     layer3_out[842] <= ~layer2_out[2604] | layer2_out[2605];
     layer3_out[843] <= layer2_out[5025] & ~layer2_out[5024];
     layer3_out[844] <= layer2_out[3020] & ~layer2_out[3019];
     layer3_out[845] <= layer2_out[9622];
     layer3_out[846] <= ~(layer2_out[6476] | layer2_out[6477]);
     layer3_out[847] <= ~(layer2_out[11011] ^ layer2_out[11012]);
     layer3_out[848] <= layer2_out[5404] ^ layer2_out[5405];
     layer3_out[849] <= ~layer2_out[5518];
     layer3_out[850] <= ~(layer2_out[3129] ^ layer2_out[3130]);
     layer3_out[851] <= ~layer2_out[3019];
     layer3_out[852] <= layer2_out[9098] | layer2_out[9099];
     layer3_out[853] <= ~(layer2_out[5118] & layer2_out[5119]);
     layer3_out[854] <= ~(layer2_out[4201] | layer2_out[4202]);
     layer3_out[855] <= layer2_out[1821] ^ layer2_out[1822];
     layer3_out[856] <= layer2_out[6013];
     layer3_out[857] <= ~(layer2_out[3424] ^ layer2_out[3425]);
     layer3_out[858] <= layer2_out[4801];
     layer3_out[859] <= ~(layer2_out[3628] | layer2_out[3629]);
     layer3_out[860] <= ~layer2_out[4068];
     layer3_out[861] <= layer2_out[1841] & layer2_out[1842];
     layer3_out[862] <= ~layer2_out[1044];
     layer3_out[863] <= layer2_out[4406];
     layer3_out[864] <= ~(layer2_out[9484] ^ layer2_out[9485]);
     layer3_out[865] <= layer2_out[3250] | layer2_out[3251];
     layer3_out[866] <= layer2_out[473] ^ layer2_out[474];
     layer3_out[867] <= layer2_out[5904] | layer2_out[5905];
     layer3_out[868] <= layer2_out[9563] & layer2_out[9564];
     layer3_out[869] <= ~(layer2_out[2085] ^ layer2_out[2086]);
     layer3_out[870] <= ~(layer2_out[5338] & layer2_out[5339]);
     layer3_out[871] <= layer2_out[11454] & ~layer2_out[11455];
     layer3_out[872] <= layer2_out[7236];
     layer3_out[873] <= ~layer2_out[9636];
     layer3_out[874] <= layer2_out[8009];
     layer3_out[875] <= layer2_out[9681] & ~layer2_out[9680];
     layer3_out[876] <= layer2_out[10693];
     layer3_out[877] <= layer2_out[2893] | layer2_out[2894];
     layer3_out[878] <= layer2_out[6685] & layer2_out[6686];
     layer3_out[879] <= layer2_out[950];
     layer3_out[880] <= ~layer2_out[7156];
     layer3_out[881] <= layer2_out[7068] & layer2_out[7069];
     layer3_out[882] <= ~layer2_out[74];
     layer3_out[883] <= ~layer2_out[8068] | layer2_out[8069];
     layer3_out[884] <= ~layer2_out[7775] | layer2_out[7774];
     layer3_out[885] <= layer2_out[4327];
     layer3_out[886] <= layer2_out[5291];
     layer3_out[887] <= ~(layer2_out[6392] & layer2_out[6393]);
     layer3_out[888] <= ~layer2_out[9441];
     layer3_out[889] <= ~(layer2_out[9069] | layer2_out[9070]);
     layer3_out[890] <= layer2_out[9705] & layer2_out[9706];
     layer3_out[891] <= ~(layer2_out[795] ^ layer2_out[796]);
     layer3_out[892] <= ~layer2_out[2655] | layer2_out[2654];
     layer3_out[893] <= ~layer2_out[10163];
     layer3_out[894] <= ~(layer2_out[8098] ^ layer2_out[8099]);
     layer3_out[895] <= ~(layer2_out[11792] | layer2_out[11793]);
     layer3_out[896] <= ~(layer2_out[8054] ^ layer2_out[8055]);
     layer3_out[897] <= ~(layer2_out[8841] ^ layer2_out[8842]);
     layer3_out[898] <= ~layer2_out[8294] | layer2_out[8293];
     layer3_out[899] <= layer2_out[395];
     layer3_out[900] <= ~layer2_out[6031];
     layer3_out[901] <= layer2_out[5749];
     layer3_out[902] <= ~(layer2_out[182] | layer2_out[183]);
     layer3_out[903] <= layer2_out[9822] & ~layer2_out[9823];
     layer3_out[904] <= layer2_out[3526];
     layer3_out[905] <= layer2_out[10809] & ~layer2_out[10808];
     layer3_out[906] <= ~layer2_out[3365];
     layer3_out[907] <= layer2_out[8606] & ~layer2_out[8607];
     layer3_out[908] <= layer2_out[9721];
     layer3_out[909] <= ~(layer2_out[5063] ^ layer2_out[5064]);
     layer3_out[910] <= layer2_out[1163];
     layer3_out[911] <= layer2_out[2053] ^ layer2_out[2054];
     layer3_out[912] <= layer2_out[3856];
     layer3_out[913] <= layer2_out[6400];
     layer3_out[914] <= layer2_out[9000] ^ layer2_out[9001];
     layer3_out[915] <= ~layer2_out[10008] | layer2_out[10009];
     layer3_out[916] <= ~layer2_out[11554];
     layer3_out[917] <= ~layer2_out[1327] | layer2_out[1328];
     layer3_out[918] <= layer2_out[5951];
     layer3_out[919] <= layer2_out[5959] & layer2_out[5960];
     layer3_out[920] <= layer2_out[2233] & ~layer2_out[2234];
     layer3_out[921] <= layer2_out[8703] ^ layer2_out[8704];
     layer3_out[922] <= ~(layer2_out[1158] ^ layer2_out[1159]);
     layer3_out[923] <= layer2_out[4965] | layer2_out[4966];
     layer3_out[924] <= layer2_out[9582] & layer2_out[9583];
     layer3_out[925] <= layer2_out[9498];
     layer3_out[926] <= ~(layer2_out[2669] & layer2_out[2670]);
     layer3_out[927] <= layer2_out[7999];
     layer3_out[928] <= layer2_out[3899] ^ layer2_out[3900];
     layer3_out[929] <= ~(layer2_out[383] | layer2_out[384]);
     layer3_out[930] <= layer2_out[1961] & layer2_out[1962];
     layer3_out[931] <= ~(layer2_out[11795] | layer2_out[11796]);
     layer3_out[932] <= ~layer2_out[7693] | layer2_out[7694];
     layer3_out[933] <= layer2_out[8663] & ~layer2_out[8662];
     layer3_out[934] <= ~(layer2_out[10610] ^ layer2_out[10611]);
     layer3_out[935] <= layer2_out[9800] & ~layer2_out[9801];
     layer3_out[936] <= layer2_out[2226];
     layer3_out[937] <= layer2_out[8809];
     layer3_out[938] <= layer2_out[547];
     layer3_out[939] <= layer2_out[10492] ^ layer2_out[10493];
     layer3_out[940] <= layer2_out[4580] & ~layer2_out[4579];
     layer3_out[941] <= layer2_out[5953] & ~layer2_out[5952];
     layer3_out[942] <= layer2_out[1773];
     layer3_out[943] <= ~(layer2_out[8197] | layer2_out[8198]);
     layer3_out[944] <= ~layer2_out[3832];
     layer3_out[945] <= layer2_out[1418];
     layer3_out[946] <= ~(layer2_out[3860] | layer2_out[3861]);
     layer3_out[947] <= layer2_out[884] & ~layer2_out[885];
     layer3_out[948] <= ~layer2_out[8108];
     layer3_out[949] <= layer2_out[6609];
     layer3_out[950] <= layer2_out[7704];
     layer3_out[951] <= ~layer2_out[11959];
     layer3_out[952] <= ~layer2_out[8061];
     layer3_out[953] <= layer2_out[4360] & ~layer2_out[4359];
     layer3_out[954] <= ~layer2_out[10515];
     layer3_out[955] <= ~(layer2_out[2105] | layer2_out[2106]);
     layer3_out[956] <= ~layer2_out[8568] | layer2_out[8569];
     layer3_out[957] <= layer2_out[3205] & ~layer2_out[3204];
     layer3_out[958] <= ~(layer2_out[6371] | layer2_out[6372]);
     layer3_out[959] <= ~layer2_out[5600];
     layer3_out[960] <= layer2_out[1405];
     layer3_out[961] <= layer2_out[7847];
     layer3_out[962] <= ~(layer2_out[1661] ^ layer2_out[1662]);
     layer3_out[963] <= layer2_out[10891] & ~layer2_out[10890];
     layer3_out[964] <= layer2_out[2560] & ~layer2_out[2561];
     layer3_out[965] <= ~(layer2_out[5726] ^ layer2_out[5727]);
     layer3_out[966] <= layer2_out[9794] & ~layer2_out[9793];
     layer3_out[967] <= ~(layer2_out[3357] | layer2_out[3358]);
     layer3_out[968] <= ~layer2_out[11965];
     layer3_out[969] <= layer2_out[10606] ^ layer2_out[10607];
     layer3_out[970] <= ~layer2_out[10498] | layer2_out[10497];
     layer3_out[971] <= ~layer2_out[5489];
     layer3_out[972] <= layer2_out[3967];
     layer3_out[973] <= ~(layer2_out[8592] & layer2_out[8593]);
     layer3_out[974] <= layer2_out[1742] & layer2_out[1743];
     layer3_out[975] <= ~layer2_out[2634];
     layer3_out[976] <= layer2_out[7000];
     layer3_out[977] <= ~(layer2_out[1094] | layer2_out[1095]);
     layer3_out[978] <= layer2_out[5244];
     layer3_out[979] <= layer2_out[6047] & ~layer2_out[6046];
     layer3_out[980] <= layer2_out[9475] ^ layer2_out[9476];
     layer3_out[981] <= layer2_out[177] & ~layer2_out[178];
     layer3_out[982] <= layer2_out[4152] & layer2_out[4153];
     layer3_out[983] <= layer2_out[6609] & ~layer2_out[6610];
     layer3_out[984] <= ~layer2_out[11517];
     layer3_out[985] <= ~(layer2_out[7309] ^ layer2_out[7310]);
     layer3_out[986] <= layer2_out[10235] ^ layer2_out[10236];
     layer3_out[987] <= layer2_out[7192] ^ layer2_out[7193];
     layer3_out[988] <= layer2_out[3380] & ~layer2_out[3379];
     layer3_out[989] <= ~layer2_out[3240] | layer2_out[3239];
     layer3_out[990] <= ~(layer2_out[8166] ^ layer2_out[8167]);
     layer3_out[991] <= ~layer2_out[11323] | layer2_out[11324];
     layer3_out[992] <= layer2_out[8254] & ~layer2_out[8253];
     layer3_out[993] <= layer2_out[3526];
     layer3_out[994] <= layer2_out[9426];
     layer3_out[995] <= ~layer2_out[11970];
     layer3_out[996] <= layer2_out[2652] ^ layer2_out[2653];
     layer3_out[997] <= ~layer2_out[11274];
     layer3_out[998] <= ~(layer2_out[4759] ^ layer2_out[4760]);
     layer3_out[999] <= ~layer2_out[9474];
     layer3_out[1000] <= ~(layer2_out[9373] & layer2_out[9374]);
     layer3_out[1001] <= layer2_out[6834] & ~layer2_out[6835];
     layer3_out[1002] <= layer2_out[873];
     layer3_out[1003] <= ~layer2_out[7431];
     layer3_out[1004] <= layer2_out[2135] & ~layer2_out[2136];
     layer3_out[1005] <= ~(layer2_out[2159] ^ layer2_out[2160]);
     layer3_out[1006] <= ~(layer2_out[6167] & layer2_out[6168]);
     layer3_out[1007] <= layer2_out[11979];
     layer3_out[1008] <= layer2_out[2616];
     layer3_out[1009] <= ~layer2_out[7750] | layer2_out[7751];
     layer3_out[1010] <= layer2_out[9943] & ~layer2_out[9942];
     layer3_out[1011] <= ~layer2_out[6033];
     layer3_out[1012] <= ~layer2_out[4856];
     layer3_out[1013] <= layer2_out[9020] & ~layer2_out[9021];
     layer3_out[1014] <= ~(layer2_out[6693] | layer2_out[6694]);
     layer3_out[1015] <= ~(layer2_out[10145] ^ layer2_out[10146]);
     layer3_out[1016] <= ~layer2_out[11594];
     layer3_out[1017] <= layer2_out[1840] & layer2_out[1841];
     layer3_out[1018] <= layer2_out[5276] ^ layer2_out[5277];
     layer3_out[1019] <= ~layer2_out[2243];
     layer3_out[1020] <= ~(layer2_out[11812] ^ layer2_out[11813]);
     layer3_out[1021] <= ~layer2_out[7997];
     layer3_out[1022] <= ~layer2_out[9361];
     layer3_out[1023] <= layer2_out[8451];
     layer3_out[1024] <= layer2_out[7933];
     layer3_out[1025] <= ~(layer2_out[8677] & layer2_out[8678]);
     layer3_out[1026] <= ~layer2_out[11295];
     layer3_out[1027] <= layer2_out[2723] ^ layer2_out[2724];
     layer3_out[1028] <= layer2_out[6911] & ~layer2_out[6910];
     layer3_out[1029] <= layer2_out[361];
     layer3_out[1030] <= layer2_out[4929] | layer2_out[4930];
     layer3_out[1031] <= ~layer2_out[9142];
     layer3_out[1032] <= ~(layer2_out[3733] ^ layer2_out[3734]);
     layer3_out[1033] <= ~layer2_out[1098] | layer2_out[1097];
     layer3_out[1034] <= layer2_out[284];
     layer3_out[1035] <= ~layer2_out[11162];
     layer3_out[1036] <= ~layer2_out[8731];
     layer3_out[1037] <= layer2_out[4103] | layer2_out[4104];
     layer3_out[1038] <= ~(layer2_out[398] | layer2_out[399]);
     layer3_out[1039] <= layer2_out[10379];
     layer3_out[1040] <= ~layer2_out[11095];
     layer3_out[1041] <= ~layer2_out[8182];
     layer3_out[1042] <= ~layer2_out[4385] | layer2_out[4386];
     layer3_out[1043] <= layer2_out[1740];
     layer3_out[1044] <= layer2_out[9576] & ~layer2_out[9577];
     layer3_out[1045] <= layer2_out[6510];
     layer3_out[1046] <= layer2_out[1572] ^ layer2_out[1573];
     layer3_out[1047] <= layer2_out[8184] & ~layer2_out[8183];
     layer3_out[1048] <= layer2_out[8889] | layer2_out[8890];
     layer3_out[1049] <= layer2_out[5300] & layer2_out[5301];
     layer3_out[1050] <= layer2_out[2104];
     layer3_out[1051] <= layer2_out[11899] | layer2_out[11900];
     layer3_out[1052] <= layer2_out[3328] | layer2_out[3329];
     layer3_out[1053] <= layer2_out[10497];
     layer3_out[1054] <= layer2_out[3821] & ~layer2_out[3820];
     layer3_out[1055] <= ~layer2_out[6366];
     layer3_out[1056] <= layer2_out[6189] ^ layer2_out[6190];
     layer3_out[1057] <= layer2_out[6672];
     layer3_out[1058] <= ~(layer2_out[6146] | layer2_out[6147]);
     layer3_out[1059] <= ~layer2_out[4799];
     layer3_out[1060] <= layer2_out[9107];
     layer3_out[1061] <= ~(layer2_out[7857] | layer2_out[7858]);
     layer3_out[1062] <= layer2_out[11881];
     layer3_out[1063] <= layer2_out[6052];
     layer3_out[1064] <= ~layer2_out[9741];
     layer3_out[1065] <= layer2_out[4536] | layer2_out[4537];
     layer3_out[1066] <= ~(layer2_out[11338] & layer2_out[11339]);
     layer3_out[1067] <= layer2_out[7519] & layer2_out[7520];
     layer3_out[1068] <= ~layer2_out[8281];
     layer3_out[1069] <= ~layer2_out[2979];
     layer3_out[1070] <= ~layer2_out[10249];
     layer3_out[1071] <= layer2_out[7520] & ~layer2_out[7521];
     layer3_out[1072] <= layer2_out[3641] & layer2_out[3642];
     layer3_out[1073] <= ~layer2_out[8454] | layer2_out[8455];
     layer3_out[1074] <= layer2_out[7905];
     layer3_out[1075] <= ~(layer2_out[9579] | layer2_out[9580]);
     layer3_out[1076] <= ~layer2_out[10730] | layer2_out[10731];
     layer3_out[1077] <= ~(layer2_out[1552] ^ layer2_out[1553]);
     layer3_out[1078] <= layer2_out[10186];
     layer3_out[1079] <= layer2_out[5451];
     layer3_out[1080] <= layer2_out[185] & layer2_out[186];
     layer3_out[1081] <= layer2_out[4252] & ~layer2_out[4253];
     layer3_out[1082] <= layer2_out[11210];
     layer3_out[1083] <= layer2_out[9051];
     layer3_out[1084] <= ~layer2_out[2388] | layer2_out[2387];
     layer3_out[1085] <= layer2_out[10206];
     layer3_out[1086] <= layer2_out[3613];
     layer3_out[1087] <= ~layer2_out[1387];
     layer3_out[1088] <= layer2_out[11070];
     layer3_out[1089] <= layer2_out[6470] & layer2_out[6471];
     layer3_out[1090] <= ~layer2_out[2964];
     layer3_out[1091] <= layer2_out[2026] ^ layer2_out[2027];
     layer3_out[1092] <= ~(layer2_out[8664] ^ layer2_out[8665]);
     layer3_out[1093] <= layer2_out[11835] ^ layer2_out[11836];
     layer3_out[1094] <= layer2_out[9244] & layer2_out[9245];
     layer3_out[1095] <= ~layer2_out[5737];
     layer3_out[1096] <= ~layer2_out[9715];
     layer3_out[1097] <= ~(layer2_out[6260] ^ layer2_out[6261]);
     layer3_out[1098] <= layer2_out[5509];
     layer3_out[1099] <= ~(layer2_out[9408] | layer2_out[9409]);
     layer3_out[1100] <= layer2_out[280] & ~layer2_out[281];
     layer3_out[1101] <= layer2_out[7847];
     layer3_out[1102] <= layer2_out[6134];
     layer3_out[1103] <= layer2_out[1223] ^ layer2_out[1224];
     layer3_out[1104] <= ~layer2_out[9354];
     layer3_out[1105] <= layer2_out[8903];
     layer3_out[1106] <= layer2_out[1622] ^ layer2_out[1623];
     layer3_out[1107] <= layer2_out[2726] & layer2_out[2727];
     layer3_out[1108] <= ~(layer2_out[401] | layer2_out[402]);
     layer3_out[1109] <= ~(layer2_out[7291] | layer2_out[7292]);
     layer3_out[1110] <= layer2_out[10688];
     layer3_out[1111] <= layer2_out[708];
     layer3_out[1112] <= ~(layer2_out[8585] & layer2_out[8586]);
     layer3_out[1113] <= ~(layer2_out[5105] | layer2_out[5106]);
     layer3_out[1114] <= layer2_out[3897] ^ layer2_out[3898];
     layer3_out[1115] <= ~(layer2_out[2712] & layer2_out[2713]);
     layer3_out[1116] <= layer2_out[10693] & ~layer2_out[10694];
     layer3_out[1117] <= layer2_out[8718] ^ layer2_out[8719];
     layer3_out[1118] <= ~layer2_out[9828];
     layer3_out[1119] <= ~(layer2_out[7880] ^ layer2_out[7881]);
     layer3_out[1120] <= layer2_out[9517];
     layer3_out[1121] <= layer2_out[7447];
     layer3_out[1122] <= ~layer2_out[3025];
     layer3_out[1123] <= layer2_out[6656];
     layer3_out[1124] <= ~layer2_out[5447] | layer2_out[5448];
     layer3_out[1125] <= layer2_out[3967] & ~layer2_out[3966];
     layer3_out[1126] <= layer2_out[10619] & ~layer2_out[10620];
     layer3_out[1127] <= layer2_out[4161] & ~layer2_out[4162];
     layer3_out[1128] <= layer2_out[4947];
     layer3_out[1129] <= ~(layer2_out[7199] | layer2_out[7200]);
     layer3_out[1130] <= layer2_out[2342] & layer2_out[2343];
     layer3_out[1131] <= layer2_out[6358] & ~layer2_out[6359];
     layer3_out[1132] <= layer2_out[10638] ^ layer2_out[10639];
     layer3_out[1133] <= layer2_out[3661];
     layer3_out[1134] <= ~layer2_out[9988];
     layer3_out[1135] <= layer2_out[9418];
     layer3_out[1136] <= ~(layer2_out[8683] | layer2_out[8684]);
     layer3_out[1137] <= layer2_out[4302];
     layer3_out[1138] <= layer2_out[7069] & ~layer2_out[7070];
     layer3_out[1139] <= ~(layer2_out[4902] | layer2_out[4903]);
     layer3_out[1140] <= layer2_out[11616];
     layer3_out[1141] <= ~layer2_out[2261];
     layer3_out[1142] <= layer2_out[10573] & ~layer2_out[10574];
     layer3_out[1143] <= layer2_out[9490] ^ layer2_out[9491];
     layer3_out[1144] <= layer2_out[11399];
     layer3_out[1145] <= layer2_out[2661];
     layer3_out[1146] <= layer2_out[475];
     layer3_out[1147] <= ~layer2_out[3612];
     layer3_out[1148] <= layer2_out[2736];
     layer3_out[1149] <= layer2_out[8746];
     layer3_out[1150] <= ~layer2_out[11203];
     layer3_out[1151] <= layer2_out[8650];
     layer3_out[1152] <= layer2_out[2339] & ~layer2_out[2340];
     layer3_out[1153] <= layer2_out[4887] & ~layer2_out[4888];
     layer3_out[1154] <= layer2_out[1357] & layer2_out[1358];
     layer3_out[1155] <= ~layer2_out[7493];
     layer3_out[1156] <= ~(layer2_out[4850] ^ layer2_out[4851]);
     layer3_out[1157] <= ~(layer2_out[11465] | layer2_out[11466]);
     layer3_out[1158] <= layer2_out[8809] & ~layer2_out[8808];
     layer3_out[1159] <= layer2_out[4096] & layer2_out[4097];
     layer3_out[1160] <= layer2_out[11345];
     layer3_out[1161] <= layer2_out[5693];
     layer3_out[1162] <= layer2_out[1453] & layer2_out[1454];
     layer3_out[1163] <= layer2_out[8910] & ~layer2_out[8909];
     layer3_out[1164] <= layer2_out[3910] & layer2_out[3911];
     layer3_out[1165] <= ~(layer2_out[11805] | layer2_out[11806]);
     layer3_out[1166] <= layer2_out[803] & ~layer2_out[804];
     layer3_out[1167] <= ~layer2_out[2902];
     layer3_out[1168] <= ~(layer2_out[4799] & layer2_out[4800]);
     layer3_out[1169] <= ~(layer2_out[5536] & layer2_out[5537]);
     layer3_out[1170] <= layer2_out[5621] ^ layer2_out[5622];
     layer3_out[1171] <= layer2_out[209] ^ layer2_out[210];
     layer3_out[1172] <= layer2_out[6662] & layer2_out[6663];
     layer3_out[1173] <= layer2_out[9094] | layer2_out[9095];
     layer3_out[1174] <= ~(layer2_out[5507] ^ layer2_out[5508]);
     layer3_out[1175] <= layer2_out[11042];
     layer3_out[1176] <= ~(layer2_out[2655] & layer2_out[2656]);
     layer3_out[1177] <= ~layer2_out[2427];
     layer3_out[1178] <= ~(layer2_out[2364] | layer2_out[2365]);
     layer3_out[1179] <= layer2_out[545];
     layer3_out[1180] <= ~(layer2_out[9161] ^ layer2_out[9162]);
     layer3_out[1181] <= layer2_out[5493] & layer2_out[5494];
     layer3_out[1182] <= ~(layer2_out[8527] | layer2_out[8528]);
     layer3_out[1183] <= layer2_out[6398];
     layer3_out[1184] <= layer2_out[2144] & layer2_out[2145];
     layer3_out[1185] <= ~layer2_out[8319];
     layer3_out[1186] <= layer2_out[9255] ^ layer2_out[9256];
     layer3_out[1187] <= layer2_out[6070] & ~layer2_out[6071];
     layer3_out[1188] <= layer2_out[2585];
     layer3_out[1189] <= ~(layer2_out[3539] ^ layer2_out[3540]);
     layer3_out[1190] <= ~layer2_out[3423] | layer2_out[3422];
     layer3_out[1191] <= layer2_out[8225] & layer2_out[8226];
     layer3_out[1192] <= ~layer2_out[6632] | layer2_out[6633];
     layer3_out[1193] <= layer2_out[11452] & layer2_out[11453];
     layer3_out[1194] <= layer2_out[10802] | layer2_out[10803];
     layer3_out[1195] <= ~layer2_out[9927];
     layer3_out[1196] <= ~(layer2_out[10620] & layer2_out[10621]);
     layer3_out[1197] <= ~layer2_out[1866];
     layer3_out[1198] <= layer2_out[9816];
     layer3_out[1199] <= layer2_out[11774] & layer2_out[11775];
     layer3_out[1200] <= ~layer2_out[5200];
     layer3_out[1201] <= ~(layer2_out[1883] ^ layer2_out[1884]);
     layer3_out[1202] <= ~layer2_out[195];
     layer3_out[1203] <= ~layer2_out[9983] | layer2_out[9984];
     layer3_out[1204] <= layer2_out[3309];
     layer3_out[1205] <= ~layer2_out[10937];
     layer3_out[1206] <= layer2_out[4544];
     layer3_out[1207] <= ~layer2_out[6070] | layer2_out[6069];
     layer3_out[1208] <= layer2_out[3354] ^ layer2_out[3355];
     layer3_out[1209] <= layer2_out[5814] ^ layer2_out[5815];
     layer3_out[1210] <= layer2_out[104];
     layer3_out[1211] <= layer2_out[9667] | layer2_out[9668];
     layer3_out[1212] <= layer2_out[6590] & layer2_out[6591];
     layer3_out[1213] <= ~(layer2_out[7182] ^ layer2_out[7183]);
     layer3_out[1214] <= ~layer2_out[5224] | layer2_out[5223];
     layer3_out[1215] <= ~layer2_out[10356];
     layer3_out[1216] <= ~layer2_out[9734];
     layer3_out[1217] <= layer2_out[5935] & layer2_out[5936];
     layer3_out[1218] <= ~(layer2_out[2505] ^ layer2_out[2506]);
     layer3_out[1219] <= ~layer2_out[10339];
     layer3_out[1220] <= layer2_out[944] | layer2_out[945];
     layer3_out[1221] <= ~(layer2_out[3840] | layer2_out[3841]);
     layer3_out[1222] <= ~(layer2_out[9438] & layer2_out[9439]);
     layer3_out[1223] <= layer2_out[3995] & layer2_out[3996];
     layer3_out[1224] <= ~layer2_out[3459];
     layer3_out[1225] <= ~layer2_out[11154];
     layer3_out[1226] <= layer2_out[6432];
     layer3_out[1227] <= layer2_out[5149] | layer2_out[5150];
     layer3_out[1228] <= layer2_out[4655] & layer2_out[4656];
     layer3_out[1229] <= ~layer2_out[2662];
     layer3_out[1230] <= ~layer2_out[4383];
     layer3_out[1231] <= ~layer2_out[4904] | layer2_out[4903];
     layer3_out[1232] <= layer2_out[7083] & ~layer2_out[7084];
     layer3_out[1233] <= ~layer2_out[387] | layer2_out[386];
     layer3_out[1234] <= ~layer2_out[11269] | layer2_out[11268];
     layer3_out[1235] <= layer2_out[1072];
     layer3_out[1236] <= layer2_out[8002] | layer2_out[8003];
     layer3_out[1237] <= layer2_out[4147] & layer2_out[4148];
     layer3_out[1238] <= ~(layer2_out[5375] & layer2_out[5376]);
     layer3_out[1239] <= ~layer2_out[952];
     layer3_out[1240] <= ~(layer2_out[7128] | layer2_out[7129]);
     layer3_out[1241] <= ~layer2_out[11598] | layer2_out[11599];
     layer3_out[1242] <= layer2_out[11646] & ~layer2_out[11647];
     layer3_out[1243] <= ~layer2_out[10016];
     layer3_out[1244] <= layer2_out[6377] ^ layer2_out[6378];
     layer3_out[1245] <= ~layer2_out[6027];
     layer3_out[1246] <= layer2_out[10103];
     layer3_out[1247] <= ~layer2_out[10339];
     layer3_out[1248] <= ~layer2_out[8415];
     layer3_out[1249] <= layer2_out[10156];
     layer3_out[1250] <= layer2_out[2493] ^ layer2_out[2494];
     layer3_out[1251] <= layer2_out[8189] | layer2_out[8190];
     layer3_out[1252] <= ~layer2_out[5383];
     layer3_out[1253] <= layer2_out[8931] | layer2_out[8932];
     layer3_out[1254] <= ~layer2_out[1797];
     layer3_out[1255] <= ~(layer2_out[6521] ^ layer2_out[6522]);
     layer3_out[1256] <= layer2_out[6528];
     layer3_out[1257] <= layer2_out[663] | layer2_out[664];
     layer3_out[1258] <= layer2_out[10496];
     layer3_out[1259] <= ~layer2_out[11157] | layer2_out[11158];
     layer3_out[1260] <= ~layer2_out[2385];
     layer3_out[1261] <= ~layer2_out[7342] | layer2_out[7341];
     layer3_out[1262] <= layer2_out[8188] & layer2_out[8189];
     layer3_out[1263] <= ~(layer2_out[10681] | layer2_out[10682]);
     layer3_out[1264] <= ~layer2_out[4274];
     layer3_out[1265] <= layer2_out[1997] | layer2_out[1998];
     layer3_out[1266] <= ~layer2_out[1277];
     layer3_out[1267] <= layer2_out[5763];
     layer3_out[1268] <= ~layer2_out[7125];
     layer3_out[1269] <= layer2_out[11426];
     layer3_out[1270] <= layer2_out[2037];
     layer3_out[1271] <= layer2_out[3232];
     layer3_out[1272] <= layer2_out[8751];
     layer3_out[1273] <= ~layer2_out[8484];
     layer3_out[1274] <= ~layer2_out[2397];
     layer3_out[1275] <= ~(layer2_out[9383] | layer2_out[9384]);
     layer3_out[1276] <= layer2_out[5694] & ~layer2_out[5693];
     layer3_out[1277] <= layer2_out[2468] | layer2_out[2469];
     layer3_out[1278] <= layer2_out[3224] & ~layer2_out[3223];
     layer3_out[1279] <= ~layer2_out[3883] | layer2_out[3882];
     layer3_out[1280] <= layer2_out[2598];
     layer3_out[1281] <= ~(layer2_out[4292] & layer2_out[4293]);
     layer3_out[1282] <= ~(layer2_out[3921] & layer2_out[3922]);
     layer3_out[1283] <= ~(layer2_out[7546] & layer2_out[7547]);
     layer3_out[1284] <= ~layer2_out[10621] | layer2_out[10622];
     layer3_out[1285] <= ~(layer2_out[2859] ^ layer2_out[2860]);
     layer3_out[1286] <= ~(layer2_out[1044] | layer2_out[1045]);
     layer3_out[1287] <= ~layer2_out[11947];
     layer3_out[1288] <= layer2_out[8824] ^ layer2_out[8825];
     layer3_out[1289] <= ~layer2_out[9028];
     layer3_out[1290] <= layer2_out[5425];
     layer3_out[1291] <= ~(layer2_out[10234] | layer2_out[10235]);
     layer3_out[1292] <= ~(layer2_out[6882] & layer2_out[6883]);
     layer3_out[1293] <= layer2_out[3957] & ~layer2_out[3956];
     layer3_out[1294] <= ~layer2_out[1169];
     layer3_out[1295] <= layer2_out[10955] & layer2_out[10956];
     layer3_out[1296] <= ~layer2_out[9122] | layer2_out[9123];
     layer3_out[1297] <= layer2_out[8379];
     layer3_out[1298] <= layer2_out[2224];
     layer3_out[1299] <= ~layer2_out[5810];
     layer3_out[1300] <= layer2_out[125] & layer2_out[126];
     layer3_out[1301] <= ~layer2_out[11221];
     layer3_out[1302] <= layer2_out[3790] & layer2_out[3791];
     layer3_out[1303] <= ~layer2_out[6186] | layer2_out[6185];
     layer3_out[1304] <= ~(layer2_out[651] | layer2_out[652]);
     layer3_out[1305] <= layer2_out[9945] ^ layer2_out[9946];
     layer3_out[1306] <= ~layer2_out[3679];
     layer3_out[1307] <= ~layer2_out[2880];
     layer3_out[1308] <= ~layer2_out[9944] | layer2_out[9943];
     layer3_out[1309] <= layer2_out[686] & layer2_out[687];
     layer3_out[1310] <= ~layer2_out[4312] | layer2_out[4311];
     layer3_out[1311] <= ~layer2_out[5623];
     layer3_out[1312] <= layer2_out[7589] | layer2_out[7590];
     layer3_out[1313] <= layer2_out[11026] & layer2_out[11027];
     layer3_out[1314] <= layer2_out[764] & ~layer2_out[763];
     layer3_out[1315] <= ~(layer2_out[5221] & layer2_out[5222]);
     layer3_out[1316] <= layer2_out[9200] & ~layer2_out[9199];
     layer3_out[1317] <= layer2_out[11185] & layer2_out[11186];
     layer3_out[1318] <= layer2_out[4297];
     layer3_out[1319] <= ~layer2_out[2697];
     layer3_out[1320] <= ~layer2_out[2020];
     layer3_out[1321] <= layer2_out[8895] & ~layer2_out[8894];
     layer3_out[1322] <= layer2_out[4693];
     layer3_out[1323] <= ~layer2_out[5912] | layer2_out[5911];
     layer3_out[1324] <= ~(layer2_out[5491] ^ layer2_out[5492]);
     layer3_out[1325] <= layer2_out[2975];
     layer3_out[1326] <= layer2_out[2571];
     layer3_out[1327] <= ~layer2_out[5859];
     layer3_out[1328] <= layer2_out[6755];
     layer3_out[1329] <= layer2_out[629];
     layer3_out[1330] <= ~layer2_out[11739];
     layer3_out[1331] <= layer2_out[3287] | layer2_out[3288];
     layer3_out[1332] <= ~layer2_out[11794];
     layer3_out[1333] <= layer2_out[883];
     layer3_out[1334] <= ~layer2_out[889];
     layer3_out[1335] <= ~layer2_out[5505];
     layer3_out[1336] <= ~layer2_out[4870];
     layer3_out[1337] <= layer2_out[10804];
     layer3_out[1338] <= ~layer2_out[1458];
     layer3_out[1339] <= ~layer2_out[5790];
     layer3_out[1340] <= layer2_out[6304] & layer2_out[6305];
     layer3_out[1341] <= layer2_out[285];
     layer3_out[1342] <= layer2_out[7870];
     layer3_out[1343] <= ~layer2_out[4333];
     layer3_out[1344] <= ~layer2_out[4774] | layer2_out[4773];
     layer3_out[1345] <= ~layer2_out[10774];
     layer3_out[1346] <= layer2_out[3111] | layer2_out[3112];
     layer3_out[1347] <= layer2_out[4068] | layer2_out[4069];
     layer3_out[1348] <= layer2_out[2501];
     layer3_out[1349] <= ~layer2_out[1458];
     layer3_out[1350] <= ~layer2_out[2155];
     layer3_out[1351] <= ~(layer2_out[11714] | layer2_out[11715]);
     layer3_out[1352] <= layer2_out[11575];
     layer3_out[1353] <= layer2_out[9390] & ~layer2_out[9391];
     layer3_out[1354] <= ~layer2_out[4251];
     layer3_out[1355] <= ~(layer2_out[10421] | layer2_out[10422]);
     layer3_out[1356] <= ~(layer2_out[6788] & layer2_out[6789]);
     layer3_out[1357] <= ~(layer2_out[7241] & layer2_out[7242]);
     layer3_out[1358] <= layer2_out[11265];
     layer3_out[1359] <= layer2_out[6155];
     layer3_out[1360] <= ~layer2_out[10854];
     layer3_out[1361] <= ~layer2_out[3504] | layer2_out[3505];
     layer3_out[1362] <= layer2_out[3523] ^ layer2_out[3524];
     layer3_out[1363] <= ~layer2_out[8891] | layer2_out[8892];
     layer3_out[1364] <= ~layer2_out[922];
     layer3_out[1365] <= ~layer2_out[2835] | layer2_out[2834];
     layer3_out[1366] <= layer2_out[6997];
     layer3_out[1367] <= ~layer2_out[8512] | layer2_out[8513];
     layer3_out[1368] <= layer2_out[7544] | layer2_out[7545];
     layer3_out[1369] <= layer2_out[7144];
     layer3_out[1370] <= layer2_out[550];
     layer3_out[1371] <= ~layer2_out[3744];
     layer3_out[1372] <= ~layer2_out[9547] | layer2_out[9548];
     layer3_out[1373] <= ~(layer2_out[6918] & layer2_out[6919]);
     layer3_out[1374] <= ~layer2_out[5991];
     layer3_out[1375] <= ~(layer2_out[7562] & layer2_out[7563]);
     layer3_out[1376] <= ~layer2_out[5381] | layer2_out[5380];
     layer3_out[1377] <= ~(layer2_out[3218] ^ layer2_out[3219]);
     layer3_out[1378] <= ~(layer2_out[3481] ^ layer2_out[3482]);
     layer3_out[1379] <= layer2_out[3313] & ~layer2_out[3312];
     layer3_out[1380] <= layer2_out[5406];
     layer3_out[1381] <= ~layer2_out[8687];
     layer3_out[1382] <= layer2_out[9449];
     layer3_out[1383] <= ~(layer2_out[7304] ^ layer2_out[7305]);
     layer3_out[1384] <= ~layer2_out[8496] | layer2_out[8495];
     layer3_out[1385] <= layer2_out[10187];
     layer3_out[1386] <= layer2_out[1625];
     layer3_out[1387] <= ~layer2_out[7408];
     layer3_out[1388] <= ~(layer2_out[2956] ^ layer2_out[2957]);
     layer3_out[1389] <= layer2_out[6478];
     layer3_out[1390] <= layer2_out[5160] & ~layer2_out[5161];
     layer3_out[1391] <= layer2_out[5357];
     layer3_out[1392] <= layer2_out[4185] & ~layer2_out[4186];
     layer3_out[1393] <= ~layer2_out[5460] | layer2_out[5459];
     layer3_out[1394] <= ~layer2_out[1313] | layer2_out[1314];
     layer3_out[1395] <= layer2_out[8412];
     layer3_out[1396] <= layer2_out[4992];
     layer3_out[1397] <= ~layer2_out[11005];
     layer3_out[1398] <= ~layer2_out[8802] | layer2_out[8803];
     layer3_out[1399] <= layer2_out[2375];
     layer3_out[1400] <= ~layer2_out[3002] | layer2_out[3003];
     layer3_out[1401] <= ~layer2_out[5570] | layer2_out[5571];
     layer3_out[1402] <= layer2_out[8913];
     layer3_out[1403] <= layer2_out[8949];
     layer3_out[1404] <= ~(layer2_out[8779] ^ layer2_out[8780]);
     layer3_out[1405] <= layer2_out[6079];
     layer3_out[1406] <= layer2_out[8390] & layer2_out[8391];
     layer3_out[1407] <= ~(layer2_out[9913] | layer2_out[9914]);
     layer3_out[1408] <= layer2_out[3063] & ~layer2_out[3062];
     layer3_out[1409] <= ~layer2_out[3265];
     layer3_out[1410] <= layer2_out[1836] | layer2_out[1837];
     layer3_out[1411] <= ~(layer2_out[4307] & layer2_out[4308]);
     layer3_out[1412] <= ~layer2_out[5500] | layer2_out[5501];
     layer3_out[1413] <= layer2_out[8465];
     layer3_out[1414] <= layer2_out[6891];
     layer3_out[1415] <= ~layer2_out[4419];
     layer3_out[1416] <= ~layer2_out[7410];
     layer3_out[1417] <= ~layer2_out[9698];
     layer3_out[1418] <= ~(layer2_out[4990] ^ layer2_out[4991]);
     layer3_out[1419] <= layer2_out[9343] ^ layer2_out[9344];
     layer3_out[1420] <= ~(layer2_out[1918] ^ layer2_out[1919]);
     layer3_out[1421] <= ~layer2_out[10381] | layer2_out[10380];
     layer3_out[1422] <= layer2_out[7498] ^ layer2_out[7499];
     layer3_out[1423] <= layer2_out[1684];
     layer3_out[1424] <= ~(layer2_out[8648] | layer2_out[8649]);
     layer3_out[1425] <= layer2_out[8374];
     layer3_out[1426] <= ~layer2_out[5048];
     layer3_out[1427] <= layer2_out[10813] | layer2_out[10814];
     layer3_out[1428] <= layer2_out[6128] & ~layer2_out[6127];
     layer3_out[1429] <= ~layer2_out[11451];
     layer3_out[1430] <= layer2_out[4881];
     layer3_out[1431] <= layer2_out[7732];
     layer3_out[1432] <= layer2_out[9002];
     layer3_out[1433] <= ~layer2_out[6703];
     layer3_out[1434] <= ~(layer2_out[10079] | layer2_out[10080]);
     layer3_out[1435] <= ~layer2_out[6967] | layer2_out[6966];
     layer3_out[1436] <= ~layer2_out[7025];
     layer3_out[1437] <= layer2_out[9537] & layer2_out[9538];
     layer3_out[1438] <= layer2_out[10119];
     layer3_out[1439] <= ~layer2_out[10743];
     layer3_out[1440] <= layer2_out[7346];
     layer3_out[1441] <= ~layer2_out[3002] | layer2_out[3001];
     layer3_out[1442] <= layer2_out[5706] | layer2_out[5707];
     layer3_out[1443] <= ~(layer2_out[9660] & layer2_out[9661]);
     layer3_out[1444] <= layer2_out[3624] | layer2_out[3625];
     layer3_out[1445] <= ~(layer2_out[11538] ^ layer2_out[11539]);
     layer3_out[1446] <= ~layer2_out[4089];
     layer3_out[1447] <= ~layer2_out[1524] | layer2_out[1523];
     layer3_out[1448] <= layer2_out[9462] | layer2_out[9463];
     layer3_out[1449] <= ~layer2_out[10582] | layer2_out[10583];
     layer3_out[1450] <= ~layer2_out[884] | layer2_out[883];
     layer3_out[1451] <= ~layer2_out[5605] | layer2_out[5606];
     layer3_out[1452] <= ~layer2_out[1242];
     layer3_out[1453] <= layer2_out[11277];
     layer3_out[1454] <= layer2_out[6892] | layer2_out[6893];
     layer3_out[1455] <= layer2_out[5110] ^ layer2_out[5111];
     layer3_out[1456] <= layer2_out[945] & layer2_out[946];
     layer3_out[1457] <= ~(layer2_out[573] & layer2_out[574]);
     layer3_out[1458] <= layer2_out[10863] & ~layer2_out[10864];
     layer3_out[1459] <= ~(layer2_out[7692] & layer2_out[7693]);
     layer3_out[1460] <= ~layer2_out[1412] | layer2_out[1411];
     layer3_out[1461] <= ~(layer2_out[3489] | layer2_out[3490]);
     layer3_out[1462] <= ~layer2_out[5144];
     layer3_out[1463] <= layer2_out[8500] & ~layer2_out[8501];
     layer3_out[1464] <= layer2_out[2791] | layer2_out[2792];
     layer3_out[1465] <= layer2_out[4238];
     layer3_out[1466] <= ~layer2_out[2520];
     layer3_out[1467] <= ~(layer2_out[7935] & layer2_out[7936]);
     layer3_out[1468] <= layer2_out[10197];
     layer3_out[1469] <= layer2_out[543];
     layer3_out[1470] <= ~layer2_out[3305];
     layer3_out[1471] <= ~layer2_out[6760];
     layer3_out[1472] <= ~layer2_out[3319];
     layer3_out[1473] <= ~layer2_out[9447];
     layer3_out[1474] <= layer2_out[6448] & ~layer2_out[6447];
     layer3_out[1475] <= ~layer2_out[6519];
     layer3_out[1476] <= layer2_out[5721] & ~layer2_out[5722];
     layer3_out[1477] <= ~layer2_out[1184];
     layer3_out[1478] <= ~layer2_out[3371] | layer2_out[3370];
     layer3_out[1479] <= layer2_out[2305];
     layer3_out[1480] <= layer2_out[2107] | layer2_out[2108];
     layer3_out[1481] <= ~(layer2_out[10034] ^ layer2_out[10035]);
     layer3_out[1482] <= layer2_out[11368] ^ layer2_out[11369];
     layer3_out[1483] <= ~layer2_out[4007];
     layer3_out[1484] <= ~layer2_out[10746] | layer2_out[10747];
     layer3_out[1485] <= ~layer2_out[108] | layer2_out[107];
     layer3_out[1486] <= layer2_out[7347] & ~layer2_out[7348];
     layer3_out[1487] <= ~layer2_out[10013];
     layer3_out[1488] <= layer2_out[1205];
     layer3_out[1489] <= ~(layer2_out[3196] | layer2_out[3197]);
     layer3_out[1490] <= ~layer2_out[7917];
     layer3_out[1491] <= ~layer2_out[692];
     layer3_out[1492] <= ~(layer2_out[10625] ^ layer2_out[10626]);
     layer3_out[1493] <= ~layer2_out[1246];
     layer3_out[1494] <= ~(layer2_out[8995] & layer2_out[8996]);
     layer3_out[1495] <= ~layer2_out[10488] | layer2_out[10487];
     layer3_out[1496] <= ~(layer2_out[11692] & layer2_out[11693]);
     layer3_out[1497] <= layer2_out[2048];
     layer3_out[1498] <= layer2_out[8967];
     layer3_out[1499] <= layer2_out[6655];
     layer3_out[1500] <= ~layer2_out[4643];
     layer3_out[1501] <= layer2_out[10450];
     layer3_out[1502] <= layer2_out[2686] & layer2_out[2687];
     layer3_out[1503] <= layer2_out[4397];
     layer3_out[1504] <= layer2_out[1644] ^ layer2_out[1645];
     layer3_out[1505] <= ~layer2_out[11807] | layer2_out[11806];
     layer3_out[1506] <= layer2_out[8146] | layer2_out[8147];
     layer3_out[1507] <= ~layer2_out[1117];
     layer3_out[1508] <= layer2_out[3450];
     layer3_out[1509] <= ~(layer2_out[9634] | layer2_out[9635]);
     layer3_out[1510] <= ~(layer2_out[6009] & layer2_out[6010]);
     layer3_out[1511] <= ~layer2_out[3724] | layer2_out[3723];
     layer3_out[1512] <= layer2_out[10484];
     layer3_out[1513] <= layer2_out[9467] | layer2_out[9468];
     layer3_out[1514] <= layer2_out[9851];
     layer3_out[1515] <= ~(layer2_out[6204] & layer2_out[6205]);
     layer3_out[1516] <= ~layer2_out[6735];
     layer3_out[1517] <= ~(layer2_out[7190] ^ layer2_out[7191]);
     layer3_out[1518] <= layer2_out[1407];
     layer3_out[1519] <= layer2_out[11811];
     layer3_out[1520] <= ~layer2_out[670];
     layer3_out[1521] <= layer2_out[6561];
     layer3_out[1522] <= ~(layer2_out[1006] & layer2_out[1007]);
     layer3_out[1523] <= ~layer2_out[4901] | layer2_out[4902];
     layer3_out[1524] <= layer2_out[3256] ^ layer2_out[3257];
     layer3_out[1525] <= layer2_out[4239] | layer2_out[4240];
     layer3_out[1526] <= ~layer2_out[5386] | layer2_out[5387];
     layer3_out[1527] <= ~layer2_out[7581];
     layer3_out[1528] <= ~layer2_out[7706];
     layer3_out[1529] <= layer2_out[9610];
     layer3_out[1530] <= ~layer2_out[7071];
     layer3_out[1531] <= ~layer2_out[8891] | layer2_out[8890];
     layer3_out[1532] <= ~layer2_out[8064] | layer2_out[8065];
     layer3_out[1533] <= ~layer2_out[6458] | layer2_out[6457];
     layer3_out[1534] <= layer2_out[6624];
     layer3_out[1535] <= layer2_out[11331] & ~layer2_out[11332];
     layer3_out[1536] <= ~layer2_out[7411] | layer2_out[7412];
     layer3_out[1537] <= layer2_out[1766];
     layer3_out[1538] <= layer2_out[11743] & ~layer2_out[11742];
     layer3_out[1539] <= layer2_out[4855] & ~layer2_out[4854];
     layer3_out[1540] <= layer2_out[9776] ^ layer2_out[9777];
     layer3_out[1541] <= ~layer2_out[1702] | layer2_out[1701];
     layer3_out[1542] <= ~layer2_out[6999] | layer2_out[7000];
     layer3_out[1543] <= layer2_out[3232];
     layer3_out[1544] <= ~(layer2_out[9529] ^ layer2_out[9530]);
     layer3_out[1545] <= ~layer2_out[1802];
     layer3_out[1546] <= ~layer2_out[5081];
     layer3_out[1547] <= layer2_out[5241];
     layer3_out[1548] <= ~(layer2_out[3044] | layer2_out[3045]);
     layer3_out[1549] <= layer2_out[365];
     layer3_out[1550] <= ~(layer2_out[9301] ^ layer2_out[9302]);
     layer3_out[1551] <= layer2_out[9005] ^ layer2_out[9006];
     layer3_out[1552] <= layer2_out[4666];
     layer3_out[1553] <= ~layer2_out[5006] | layer2_out[5005];
     layer3_out[1554] <= ~layer2_out[1311];
     layer3_out[1555] <= ~(layer2_out[4390] & layer2_out[4391]);
     layer3_out[1556] <= layer2_out[10615];
     layer3_out[1557] <= layer2_out[1843];
     layer3_out[1558] <= ~(layer2_out[9186] | layer2_out[9187]);
     layer3_out[1559] <= ~(layer2_out[10917] ^ layer2_out[10918]);
     layer3_out[1560] <= ~layer2_out[9296];
     layer3_out[1561] <= layer2_out[3020] ^ layer2_out[3021];
     layer3_out[1562] <= ~layer2_out[11778];
     layer3_out[1563] <= layer2_out[858] | layer2_out[859];
     layer3_out[1564] <= layer2_out[8549];
     layer3_out[1565] <= layer2_out[7062] & ~layer2_out[7061];
     layer3_out[1566] <= layer2_out[3229] ^ layer2_out[3230];
     layer3_out[1567] <= ~layer2_out[5930];
     layer3_out[1568] <= layer2_out[127] ^ layer2_out[128];
     layer3_out[1569] <= layer2_out[11683] & layer2_out[11684];
     layer3_out[1570] <= ~(layer2_out[4407] & layer2_out[4408]);
     layer3_out[1571] <= layer2_out[9294] ^ layer2_out[9295];
     layer3_out[1572] <= ~(layer2_out[10346] ^ layer2_out[10347]);
     layer3_out[1573] <= ~layer2_out[6494];
     layer3_out[1574] <= ~layer2_out[2704];
     layer3_out[1575] <= ~(layer2_out[1944] & layer2_out[1945]);
     layer3_out[1576] <= layer2_out[2857] ^ layer2_out[2858];
     layer3_out[1577] <= ~layer2_out[4535];
     layer3_out[1578] <= layer2_out[2701];
     layer3_out[1579] <= ~(layer2_out[4709] & layer2_out[4710]);
     layer3_out[1580] <= layer2_out[179];
     layer3_out[1581] <= ~layer2_out[3399] | layer2_out[3398];
     layer3_out[1582] <= layer2_out[6503] & ~layer2_out[6504];
     layer3_out[1583] <= ~layer2_out[10360];
     layer3_out[1584] <= layer2_out[2457] | layer2_out[2458];
     layer3_out[1585] <= ~layer2_out[10071];
     layer3_out[1586] <= ~layer2_out[6192];
     layer3_out[1587] <= ~layer2_out[541];
     layer3_out[1588] <= ~layer2_out[11808];
     layer3_out[1589] <= ~layer2_out[7752];
     layer3_out[1590] <= ~(layer2_out[506] ^ layer2_out[507]);
     layer3_out[1591] <= ~layer2_out[10677];
     layer3_out[1592] <= ~(layer2_out[9527] & layer2_out[9528]);
     layer3_out[1593] <= layer2_out[8604];
     layer3_out[1594] <= ~layer2_out[9599];
     layer3_out[1595] <= ~layer2_out[9364] | layer2_out[9365];
     layer3_out[1596] <= layer2_out[202];
     layer3_out[1597] <= layer2_out[927] | layer2_out[928];
     layer3_out[1598] <= ~layer2_out[6414];
     layer3_out[1599] <= layer2_out[8791] | layer2_out[8792];
     layer3_out[1600] <= layer2_out[3799] & ~layer2_out[3800];
     layer3_out[1601] <= ~layer2_out[11863];
     layer3_out[1602] <= layer2_out[6254] & layer2_out[6255];
     layer3_out[1603] <= layer2_out[5168] | layer2_out[5169];
     layer3_out[1604] <= layer2_out[10873];
     layer3_out[1605] <= ~layer2_out[1216];
     layer3_out[1606] <= layer2_out[868];
     layer3_out[1607] <= ~(layer2_out[2062] | layer2_out[2063]);
     layer3_out[1608] <= ~layer2_out[10834] | layer2_out[10835];
     layer3_out[1609] <= ~(layer2_out[8792] ^ layer2_out[8793]);
     layer3_out[1610] <= ~layer2_out[2216];
     layer3_out[1611] <= layer2_out[9614];
     layer3_out[1612] <= layer2_out[9206] & layer2_out[9207];
     layer3_out[1613] <= ~layer2_out[9396];
     layer3_out[1614] <= ~(layer2_out[6895] & layer2_out[6896]);
     layer3_out[1615] <= ~layer2_out[2481];
     layer3_out[1616] <= ~layer2_out[10559] | layer2_out[10560];
     layer3_out[1617] <= layer2_out[11372] | layer2_out[11373];
     layer3_out[1618] <= ~layer2_out[5063];
     layer3_out[1619] <= ~(layer2_out[10074] ^ layer2_out[10075]);
     layer3_out[1620] <= layer2_out[4960] | layer2_out[4961];
     layer3_out[1621] <= layer2_out[10641] ^ layer2_out[10642];
     layer3_out[1622] <= layer2_out[10958] & layer2_out[10959];
     layer3_out[1623] <= ~layer2_out[11253] | layer2_out[11254];
     layer3_out[1624] <= ~layer2_out[7378];
     layer3_out[1625] <= ~layer2_out[9980] | layer2_out[9981];
     layer3_out[1626] <= layer2_out[6332] | layer2_out[6333];
     layer3_out[1627] <= ~layer2_out[1447];
     layer3_out[1628] <= layer2_out[3977] ^ layer2_out[3978];
     layer3_out[1629] <= ~layer2_out[1909] | layer2_out[1910];
     layer3_out[1630] <= layer2_out[3303] | layer2_out[3304];
     layer3_out[1631] <= layer2_out[1228];
     layer3_out[1632] <= layer2_out[966] & ~layer2_out[965];
     layer3_out[1633] <= layer2_out[3722] ^ layer2_out[3723];
     layer3_out[1634] <= layer2_out[8459];
     layer3_out[1635] <= layer2_out[9378];
     layer3_out[1636] <= layer2_out[8796] | layer2_out[8797];
     layer3_out[1637] <= layer2_out[4286] ^ layer2_out[4287];
     layer3_out[1638] <= layer2_out[8449] | layer2_out[8450];
     layer3_out[1639] <= layer2_out[2250] & ~layer2_out[2249];
     layer3_out[1640] <= layer2_out[6104] ^ layer2_out[6105];
     layer3_out[1641] <= ~layer2_out[1929];
     layer3_out[1642] <= layer2_out[4533];
     layer3_out[1643] <= ~layer2_out[3474];
     layer3_out[1644] <= layer2_out[9030];
     layer3_out[1645] <= ~(layer2_out[9773] ^ layer2_out[9774]);
     layer3_out[1646] <= ~layer2_out[9381] | layer2_out[9380];
     layer3_out[1647] <= layer2_out[7909] ^ layer2_out[7910];
     layer3_out[1648] <= layer2_out[8838];
     layer3_out[1649] <= ~layer2_out[192];
     layer3_out[1650] <= layer2_out[11750];
     layer3_out[1651] <= layer2_out[2280] & ~layer2_out[2281];
     layer3_out[1652] <= layer2_out[8513];
     layer3_out[1653] <= ~layer2_out[2089];
     layer3_out[1654] <= ~layer2_out[225];
     layer3_out[1655] <= ~layer2_out[1012] | layer2_out[1013];
     layer3_out[1656] <= layer2_out[11895] & ~layer2_out[11896];
     layer3_out[1657] <= layer2_out[1957];
     layer3_out[1658] <= ~layer2_out[2069];
     layer3_out[1659] <= layer2_out[4734];
     layer3_out[1660] <= layer2_out[11905] | layer2_out[11906];
     layer3_out[1661] <= ~layer2_out[1555] | layer2_out[1554];
     layer3_out[1662] <= layer2_out[7269];
     layer3_out[1663] <= layer2_out[3106];
     layer3_out[1664] <= ~(layer2_out[1846] ^ layer2_out[1847]);
     layer3_out[1665] <= ~(layer2_out[6043] ^ layer2_out[6044]);
     layer3_out[1666] <= layer2_out[7981];
     layer3_out[1667] <= layer2_out[5194];
     layer3_out[1668] <= ~layer2_out[9976] | layer2_out[9977];
     layer3_out[1669] <= layer2_out[7193] & layer2_out[7194];
     layer3_out[1670] <= layer2_out[8086];
     layer3_out[1671] <= layer2_out[4206];
     layer3_out[1672] <= ~layer2_out[6009] | layer2_out[6008];
     layer3_out[1673] <= layer2_out[11059];
     layer3_out[1674] <= ~layer2_out[11346];
     layer3_out[1675] <= ~layer2_out[2398] | layer2_out[2399];
     layer3_out[1676] <= ~(layer2_out[7154] ^ layer2_out[7155]);
     layer3_out[1677] <= ~layer2_out[3133] | layer2_out[3132];
     layer3_out[1678] <= ~(layer2_out[11152] ^ layer2_out[11153]);
     layer3_out[1679] <= ~layer2_out[8516];
     layer3_out[1680] <= layer2_out[2370] | layer2_out[2371];
     layer3_out[1681] <= ~layer2_out[11739];
     layer3_out[1682] <= layer2_out[5824];
     layer3_out[1683] <= ~layer2_out[1152];
     layer3_out[1684] <= ~layer2_out[6072];
     layer3_out[1685] <= layer2_out[1188];
     layer3_out[1686] <= ~layer2_out[2087];
     layer3_out[1687] <= layer2_out[7250] & ~layer2_out[7251];
     layer3_out[1688] <= ~layer2_out[11650] | layer2_out[11649];
     layer3_out[1689] <= layer2_out[10643];
     layer3_out[1690] <= ~layer2_out[11169];
     layer3_out[1691] <= layer2_out[9949];
     layer3_out[1692] <= layer2_out[6766] | layer2_out[6767];
     layer3_out[1693] <= ~layer2_out[2608];
     layer3_out[1694] <= ~layer2_out[3060];
     layer3_out[1695] <= layer2_out[3254] & ~layer2_out[3253];
     layer3_out[1696] <= layer2_out[8024];
     layer3_out[1697] <= ~(layer2_out[7414] | layer2_out[7415]);
     layer3_out[1698] <= ~layer2_out[11007];
     layer3_out[1699] <= ~layer2_out[1848];
     layer3_out[1700] <= layer2_out[5426];
     layer3_out[1701] <= layer2_out[4469] & ~layer2_out[4468];
     layer3_out[1702] <= layer2_out[4086];
     layer3_out[1703] <= layer2_out[5278];
     layer3_out[1704] <= ~(layer2_out[3515] ^ layer2_out[3516]);
     layer3_out[1705] <= ~(layer2_out[1060] & layer2_out[1061]);
     layer3_out[1706] <= layer2_out[11520] & layer2_out[11521];
     layer3_out[1707] <= layer2_out[6829];
     layer3_out[1708] <= layer2_out[9663] | layer2_out[9664];
     layer3_out[1709] <= ~(layer2_out[9778] & layer2_out[9779]);
     layer3_out[1710] <= ~(layer2_out[1105] & layer2_out[1106]);
     layer3_out[1711] <= layer2_out[9970];
     layer3_out[1712] <= ~(layer2_out[1858] | layer2_out[1859]);
     layer3_out[1713] <= ~layer2_out[850];
     layer3_out[1714] <= layer2_out[7886] | layer2_out[7887];
     layer3_out[1715] <= ~(layer2_out[7321] & layer2_out[7322]);
     layer3_out[1716] <= ~(layer2_out[8701] | layer2_out[8702]);
     layer3_out[1717] <= layer2_out[10600];
     layer3_out[1718] <= layer2_out[7338];
     layer3_out[1719] <= layer2_out[3566] | layer2_out[3567];
     layer3_out[1720] <= ~layer2_out[632];
     layer3_out[1721] <= layer2_out[352] & ~layer2_out[351];
     layer3_out[1722] <= layer2_out[5671] ^ layer2_out[5672];
     layer3_out[1723] <= layer2_out[8896] | layer2_out[8897];
     layer3_out[1724] <= layer2_out[4862];
     layer3_out[1725] <= layer2_out[5086] & ~layer2_out[5085];
     layer3_out[1726] <= layer2_out[7957];
     layer3_out[1727] <= layer2_out[5853] | layer2_out[5854];
     layer3_out[1728] <= ~layer2_out[6188];
     layer3_out[1729] <= layer2_out[11222] | layer2_out[11223];
     layer3_out[1730] <= layer2_out[209];
     layer3_out[1731] <= layer2_out[11678] & ~layer2_out[11677];
     layer3_out[1732] <= layer2_out[7038] & layer2_out[7039];
     layer3_out[1733] <= layer2_out[2789] & ~layer2_out[2790];
     layer3_out[1734] <= ~layer2_out[8250];
     layer3_out[1735] <= ~layer2_out[7157];
     layer3_out[1736] <= ~(layer2_out[4723] & layer2_out[4724]);
     layer3_out[1737] <= ~layer2_out[6907] | layer2_out[6908];
     layer3_out[1738] <= ~(layer2_out[577] ^ layer2_out[578]);
     layer3_out[1739] <= ~(layer2_out[7467] ^ layer2_out[7468]);
     layer3_out[1740] <= layer2_out[11971] & ~layer2_out[11972];
     layer3_out[1741] <= ~layer2_out[2227];
     layer3_out[1742] <= layer2_out[423] ^ layer2_out[424];
     layer3_out[1743] <= layer2_out[230] | layer2_out[231];
     layer3_out[1744] <= layer2_out[8163] ^ layer2_out[8164];
     layer3_out[1745] <= layer2_out[3692] ^ layer2_out[3693];
     layer3_out[1746] <= layer2_out[5526];
     layer3_out[1747] <= ~layer2_out[5252];
     layer3_out[1748] <= ~layer2_out[4061] | layer2_out[4062];
     layer3_out[1749] <= ~layer2_out[10539];
     layer3_out[1750] <= ~layer2_out[1549];
     layer3_out[1751] <= ~layer2_out[2823] | layer2_out[2822];
     layer3_out[1752] <= layer2_out[2169] | layer2_out[2170];
     layer3_out[1753] <= ~(layer2_out[7219] & layer2_out[7220]);
     layer3_out[1754] <= layer2_out[7550] | layer2_out[7551];
     layer3_out[1755] <= layer2_out[1658] & layer2_out[1659];
     layer3_out[1756] <= layer2_out[7217];
     layer3_out[1757] <= ~layer2_out[1182];
     layer3_out[1758] <= ~(layer2_out[7609] ^ layer2_out[7610]);
     layer3_out[1759] <= ~layer2_out[10797];
     layer3_out[1760] <= layer2_out[9748] | layer2_out[9749];
     layer3_out[1761] <= layer2_out[7537] | layer2_out[7538];
     layer3_out[1762] <= ~layer2_out[3606] | layer2_out[3605];
     layer3_out[1763] <= ~(layer2_out[10026] ^ layer2_out[10027]);
     layer3_out[1764] <= layer2_out[11834];
     layer3_out[1765] <= layer2_out[4592];
     layer3_out[1766] <= layer2_out[9788];
     layer3_out[1767] <= layer2_out[11246];
     layer3_out[1768] <= layer2_out[1129] | layer2_out[1130];
     layer3_out[1769] <= layer2_out[1526];
     layer3_out[1770] <= ~(layer2_out[10094] ^ layer2_out[10095]);
     layer3_out[1771] <= ~(layer2_out[5468] | layer2_out[5469]);
     layer3_out[1772] <= ~layer2_out[7474] | layer2_out[7475];
     layer3_out[1773] <= ~(layer2_out[7919] ^ layer2_out[7920]);
     layer3_out[1774] <= ~layer2_out[5114];
     layer3_out[1775] <= ~layer2_out[568];
     layer3_out[1776] <= layer2_out[8196] | layer2_out[8197];
     layer3_out[1777] <= layer2_out[9327];
     layer3_out[1778] <= ~layer2_out[9986];
     layer3_out[1779] <= layer2_out[8112] & ~layer2_out[8111];
     layer3_out[1780] <= layer2_out[3326];
     layer3_out[1781] <= layer2_out[5471];
     layer3_out[1782] <= layer2_out[1058];
     layer3_out[1783] <= ~layer2_out[5902];
     layer3_out[1784] <= ~layer2_out[90] | layer2_out[89];
     layer3_out[1785] <= ~(layer2_out[7404] | layer2_out[7405]);
     layer3_out[1786] <= ~layer2_out[10334];
     layer3_out[1787] <= layer2_out[2282] | layer2_out[2283];
     layer3_out[1788] <= layer2_out[8119];
     layer3_out[1789] <= layer2_out[2921] & ~layer2_out[2922];
     layer3_out[1790] <= ~layer2_out[4620];
     layer3_out[1791] <= ~(layer2_out[4905] ^ layer2_out[4906]);
     layer3_out[1792] <= layer2_out[9544] ^ layer2_out[9545];
     layer3_out[1793] <= ~layer2_out[8109] | layer2_out[8108];
     layer3_out[1794] <= layer2_out[54] ^ layer2_out[55];
     layer3_out[1795] <= layer2_out[10862];
     layer3_out[1796] <= ~(layer2_out[5201] ^ layer2_out[5202]);
     layer3_out[1797] <= ~layer2_out[6426];
     layer3_out[1798] <= ~layer2_out[7712];
     layer3_out[1799] <= ~layer2_out[9379] | layer2_out[9380];
     layer3_out[1800] <= ~layer2_out[8278];
     layer3_out[1801] <= layer2_out[6297];
     layer3_out[1802] <= layer2_out[414];
     layer3_out[1803] <= ~(layer2_out[1354] & layer2_out[1355]);
     layer3_out[1804] <= layer2_out[1674];
     layer3_out[1805] <= layer2_out[93];
     layer3_out[1806] <= layer2_out[8295];
     layer3_out[1807] <= layer2_out[10240] ^ layer2_out[10241];
     layer3_out[1808] <= layer2_out[8168];
     layer3_out[1809] <= ~layer2_out[5713];
     layer3_out[1810] <= ~layer2_out[8512] | layer2_out[8511];
     layer3_out[1811] <= layer2_out[7740] & layer2_out[7741];
     layer3_out[1812] <= layer2_out[8878];
     layer3_out[1813] <= layer2_out[11736] & ~layer2_out[11735];
     layer3_out[1814] <= ~layer2_out[736];
     layer3_out[1815] <= layer2_out[5606];
     layer3_out[1816] <= ~(layer2_out[5801] & layer2_out[5802]);
     layer3_out[1817] <= layer2_out[532];
     layer3_out[1818] <= layer2_out[2394] & ~layer2_out[2395];
     layer3_out[1819] <= layer2_out[3251];
     layer3_out[1820] <= layer2_out[4310];
     layer3_out[1821] <= ~layer2_out[5257];
     layer3_out[1822] <= ~(layer2_out[8516] | layer2_out[8517]);
     layer3_out[1823] <= layer2_out[4762];
     layer3_out[1824] <= ~(layer2_out[2101] ^ layer2_out[2102]);
     layer3_out[1825] <= ~layer2_out[6148] | layer2_out[6147];
     layer3_out[1826] <= ~(layer2_out[9177] & layer2_out[9178]);
     layer3_out[1827] <= ~layer2_out[3980] | layer2_out[3981];
     layer3_out[1828] <= ~(layer2_out[3193] | layer2_out[3194]);
     layer3_out[1829] <= ~layer2_out[1935];
     layer3_out[1830] <= layer2_out[5528] | layer2_out[5529];
     layer3_out[1831] <= layer2_out[10978];
     layer3_out[1832] <= ~layer2_out[2256] | layer2_out[2255];
     layer3_out[1833] <= layer2_out[7695] ^ layer2_out[7696];
     layer3_out[1834] <= layer2_out[11909] & layer2_out[11910];
     layer3_out[1835] <= ~layer2_out[3433] | layer2_out[3434];
     layer3_out[1836] <= ~layer2_out[5314];
     layer3_out[1837] <= ~layer2_out[4784];
     layer3_out[1838] <= layer2_out[791];
     layer3_out[1839] <= layer2_out[3994] & layer2_out[3995];
     layer3_out[1840] <= ~(layer2_out[4747] ^ layer2_out[4748]);
     layer3_out[1841] <= ~layer2_out[10227];
     layer3_out[1842] <= layer2_out[9515] & layer2_out[9516];
     layer3_out[1843] <= layer2_out[1016] | layer2_out[1017];
     layer3_out[1844] <= ~layer2_out[4219] | layer2_out[4220];
     layer3_out[1845] <= ~layer2_out[9176] | layer2_out[9175];
     layer3_out[1846] <= ~layer2_out[1947];
     layer3_out[1847] <= layer2_out[937] ^ layer2_out[938];
     layer3_out[1848] <= ~layer2_out[8902];
     layer3_out[1849] <= layer2_out[10407];
     layer3_out[1850] <= ~(layer2_out[4985] | layer2_out[4986]);
     layer3_out[1851] <= layer2_out[2572] & layer2_out[2573];
     layer3_out[1852] <= ~(layer2_out[10572] & layer2_out[10573]);
     layer3_out[1853] <= layer2_out[11798] | layer2_out[11799];
     layer3_out[1854] <= layer2_out[11914];
     layer3_out[1855] <= ~layer2_out[981];
     layer3_out[1856] <= layer2_out[9351] ^ layer2_out[9352];
     layer3_out[1857] <= layer2_out[3005];
     layer3_out[1858] <= layer2_out[374];
     layer3_out[1859] <= layer2_out[2773] | layer2_out[2774];
     layer3_out[1860] <= layer2_out[1454] ^ layer2_out[1455];
     layer3_out[1861] <= ~(layer2_out[9724] | layer2_out[9725]);
     layer3_out[1862] <= layer2_out[6497] | layer2_out[6498];
     layer3_out[1863] <= ~layer2_out[8671];
     layer3_out[1864] <= ~(layer2_out[8251] | layer2_out[8252]);
     layer3_out[1865] <= layer2_out[521];
     layer3_out[1866] <= ~layer2_out[2432];
     layer3_out[1867] <= layer2_out[269] ^ layer2_out[270];
     layer3_out[1868] <= ~layer2_out[10945] | layer2_out[10944];
     layer3_out[1869] <= ~(layer2_out[10724] | layer2_out[10725]);
     layer3_out[1870] <= ~layer2_out[10033];
     layer3_out[1871] <= layer2_out[10503];
     layer3_out[1872] <= ~(layer2_out[91] ^ layer2_out[92]);
     layer3_out[1873] <= ~(layer2_out[1307] ^ layer2_out[1308]);
     layer3_out[1874] <= ~layer2_out[9800] | layer2_out[9799];
     layer3_out[1875] <= layer2_out[9488] ^ layer2_out[9489];
     layer3_out[1876] <= ~(layer2_out[8644] ^ layer2_out[8645]);
     layer3_out[1877] <= layer2_out[8796];
     layer3_out[1878] <= ~(layer2_out[7737] ^ layer2_out[7738]);
     layer3_out[1879] <= layer2_out[8757] & ~layer2_out[8758];
     layer3_out[1880] <= ~(layer2_out[10876] ^ layer2_out[10877]);
     layer3_out[1881] <= ~layer2_out[9670] | layer2_out[9669];
     layer3_out[1882] <= layer2_out[9371];
     layer3_out[1883] <= layer2_out[3352];
     layer3_out[1884] <= ~layer2_out[3196] | layer2_out[3195];
     layer3_out[1885] <= ~layer2_out[2736] | layer2_out[2735];
     layer3_out[1886] <= layer2_out[2767] ^ layer2_out[2768];
     layer3_out[1887] <= layer2_out[4442];
     layer3_out[1888] <= ~layer2_out[3502];
     layer3_out[1889] <= layer2_out[7708];
     layer3_out[1890] <= layer2_out[3705];
     layer3_out[1891] <= layer2_out[10096];
     layer3_out[1892] <= layer2_out[10305];
     layer3_out[1893] <= ~layer2_out[5059];
     layer3_out[1894] <= layer2_out[5415];
     layer3_out[1895] <= ~layer2_out[8260];
     layer3_out[1896] <= layer2_out[9850];
     layer3_out[1897] <= layer2_out[9603];
     layer3_out[1898] <= ~layer2_out[1868];
     layer3_out[1899] <= ~layer2_out[581] | layer2_out[582];
     layer3_out[1900] <= ~layer2_out[8869];
     layer3_out[1901] <= layer2_out[10158];
     layer3_out[1902] <= layer2_out[11608];
     layer3_out[1903] <= ~(layer2_out[11679] | layer2_out[11680]);
     layer3_out[1904] <= ~layer2_out[7794] | layer2_out[7795];
     layer3_out[1905] <= ~layer2_out[5126];
     layer3_out[1906] <= layer2_out[8391] & layer2_out[8392];
     layer3_out[1907] <= layer2_out[11874] ^ layer2_out[11875];
     layer3_out[1908] <= ~layer2_out[11233] | layer2_out[11234];
     layer3_out[1909] <= layer2_out[1072];
     layer3_out[1910] <= ~(layer2_out[11280] ^ layer2_out[11281]);
     layer3_out[1911] <= layer2_out[3041] & layer2_out[3042];
     layer3_out[1912] <= ~layer2_out[11943] | layer2_out[11944];
     layer3_out[1913] <= ~layer2_out[10222] | layer2_out[10221];
     layer3_out[1914] <= ~(layer2_out[4046] & layer2_out[4047]);
     layer3_out[1915] <= ~layer2_out[4042];
     layer3_out[1916] <= ~(layer2_out[1216] & layer2_out[1217]);
     layer3_out[1917] <= layer2_out[9077];
     layer3_out[1918] <= layer2_out[349] | layer2_out[350];
     layer3_out[1919] <= ~(layer2_out[2188] & layer2_out[2189]);
     layer3_out[1920] <= ~layer2_out[6120];
     layer3_out[1921] <= layer2_out[9160];
     layer3_out[1922] <= ~(layer2_out[4839] ^ layer2_out[4840]);
     layer3_out[1923] <= ~layer2_out[9078];
     layer3_out[1924] <= ~layer2_out[1723] | layer2_out[1722];
     layer3_out[1925] <= layer2_out[6126] & ~layer2_out[6127];
     layer3_out[1926] <= layer2_out[3025] & ~layer2_out[3026];
     layer3_out[1927] <= layer2_out[7067];
     layer3_out[1928] <= ~(layer2_out[3796] ^ layer2_out[3797]);
     layer3_out[1929] <= ~(layer2_out[7242] & layer2_out[7243]);
     layer3_out[1930] <= ~layer2_out[10681];
     layer3_out[1931] <= ~layer2_out[5585];
     layer3_out[1932] <= layer2_out[3519] | layer2_out[3520];
     layer3_out[1933] <= layer2_out[9946] ^ layer2_out[9947];
     layer3_out[1934] <= layer2_out[2313];
     layer3_out[1935] <= layer2_out[5663];
     layer3_out[1936] <= layer2_out[6429];
     layer3_out[1937] <= layer2_out[1384] | layer2_out[1385];
     layer3_out[1938] <= ~layer2_out[3830];
     layer3_out[1939] <= layer2_out[11320] & ~layer2_out[11319];
     layer3_out[1940] <= ~(layer2_out[4285] ^ layer2_out[4286]);
     layer3_out[1941] <= layer2_out[1530];
     layer3_out[1942] <= layer2_out[756];
     layer3_out[1943] <= layer2_out[8214] & layer2_out[8215];
     layer3_out[1944] <= layer2_out[1188] | layer2_out[1189];
     layer3_out[1945] <= layer2_out[7809];
     layer3_out[1946] <= layer2_out[7250];
     layer3_out[1947] <= ~layer2_out[7322] | layer2_out[7323];
     layer3_out[1948] <= layer2_out[4692] & layer2_out[4693];
     layer3_out[1949] <= ~layer2_out[9456];
     layer3_out[1950] <= ~layer2_out[574] | layer2_out[575];
     layer3_out[1951] <= ~(layer2_out[7906] & layer2_out[7907]);
     layer3_out[1952] <= layer2_out[11490];
     layer3_out[1953] <= layer2_out[6736];
     layer3_out[1954] <= layer2_out[1645] ^ layer2_out[1646];
     layer3_out[1955] <= layer2_out[8053];
     layer3_out[1956] <= layer2_out[10195] ^ layer2_out[10196];
     layer3_out[1957] <= layer2_out[3092] ^ layer2_out[3093];
     layer3_out[1958] <= layer2_out[11543];
     layer3_out[1959] <= ~layer2_out[3400];
     layer3_out[1960] <= ~layer2_out[7592] | layer2_out[7591];
     layer3_out[1961] <= layer2_out[11433] ^ layer2_out[11434];
     layer3_out[1962] <= layer2_out[3041] & ~layer2_out[3040];
     layer3_out[1963] <= layer2_out[9650] | layer2_out[9651];
     layer3_out[1964] <= ~layer2_out[7935];
     layer3_out[1965] <= layer2_out[6557] ^ layer2_out[6558];
     layer3_out[1966] <= ~layer2_out[6810] | layer2_out[6811];
     layer3_out[1967] <= ~layer2_out[5897];
     layer3_out[1968] <= ~layer2_out[2448];
     layer3_out[1969] <= layer2_out[10546] | layer2_out[10547];
     layer3_out[1970] <= layer2_out[4875];
     layer3_out[1971] <= layer2_out[6916] & ~layer2_out[6915];
     layer3_out[1972] <= ~(layer2_out[956] | layer2_out[957]);
     layer3_out[1973] <= ~layer2_out[9753];
     layer3_out[1974] <= ~layer2_out[2714];
     layer3_out[1975] <= ~layer2_out[10823];
     layer3_out[1976] <= ~(layer2_out[1828] ^ layer2_out[1829]);
     layer3_out[1977] <= ~layer2_out[2922] | layer2_out[2923];
     layer3_out[1978] <= layer2_out[10164];
     layer3_out[1979] <= ~layer2_out[9700] | layer2_out[9699];
     layer3_out[1980] <= layer2_out[8628] & layer2_out[8629];
     layer3_out[1981] <= ~layer2_out[6169];
     layer3_out[1982] <= ~layer2_out[6241];
     layer3_out[1983] <= ~layer2_out[1984] | layer2_out[1985];
     layer3_out[1984] <= layer2_out[8258];
     layer3_out[1985] <= layer2_out[8880] | layer2_out[8881];
     layer3_out[1986] <= layer2_out[7124];
     layer3_out[1987] <= ~(layer2_out[11952] & layer2_out[11953]);
     layer3_out[1988] <= layer2_out[10341];
     layer3_out[1989] <= layer2_out[380];
     layer3_out[1990] <= ~layer2_out[8103];
     layer3_out[1991] <= ~(layer2_out[8560] ^ layer2_out[8561]);
     layer3_out[1992] <= ~layer2_out[166];
     layer3_out[1993] <= layer2_out[9585] | layer2_out[9586];
     layer3_out[1994] <= ~layer2_out[4786] | layer2_out[4785];
     layer3_out[1995] <= layer2_out[9272];
     layer3_out[1996] <= ~layer2_out[5328];
     layer3_out[1997] <= layer2_out[11137];
     layer3_out[1998] <= ~layer2_out[11079];
     layer3_out[1999] <= layer2_out[4108] | layer2_out[4109];
     layer3_out[2000] <= layer2_out[7883];
     layer3_out[2001] <= ~layer2_out[4419] | layer2_out[4420];
     layer3_out[2002] <= layer2_out[5887];
     layer3_out[2003] <= ~layer2_out[1167];
     layer3_out[2004] <= layer2_out[11501] & layer2_out[11502];
     layer3_out[2005] <= ~(layer2_out[10244] ^ layer2_out[10245]);
     layer3_out[2006] <= layer2_out[8476];
     layer3_out[2007] <= ~layer2_out[10726];
     layer3_out[2008] <= layer2_out[5339];
     layer3_out[2009] <= layer2_out[6974];
     layer3_out[2010] <= ~layer2_out[1586];
     layer3_out[2011] <= ~(layer2_out[6705] & layer2_out[6706]);
     layer3_out[2012] <= layer2_out[10278];
     layer3_out[2013] <= layer2_out[9942];
     layer3_out[2014] <= ~layer2_out[5611];
     layer3_out[2015] <= layer2_out[559];
     layer3_out[2016] <= layer2_out[10286] ^ layer2_out[10287];
     layer3_out[2017] <= ~layer2_out[6212];
     layer3_out[2018] <= layer2_out[11457] | layer2_out[11458];
     layer3_out[2019] <= layer2_out[9021] | layer2_out[9022];
     layer3_out[2020] <= ~layer2_out[654] | layer2_out[655];
     layer3_out[2021] <= layer2_out[11689] & layer2_out[11690];
     layer3_out[2022] <= layer2_out[8708];
     layer3_out[2023] <= ~layer2_out[11313];
     layer3_out[2024] <= layer2_out[892];
     layer3_out[2025] <= ~layer2_out[6045] | layer2_out[6046];
     layer3_out[2026] <= layer2_out[8486];
     layer3_out[2027] <= layer2_out[2656] & layer2_out[2657];
     layer3_out[2028] <= ~(layer2_out[5299] & layer2_out[5300]);
     layer3_out[2029] <= layer2_out[5613] & ~layer2_out[5614];
     layer3_out[2030] <= ~layer2_out[9431];
     layer3_out[2031] <= layer2_out[3573] ^ layer2_out[3574];
     layer3_out[2032] <= layer2_out[5056];
     layer3_out[2033] <= ~layer2_out[597];
     layer3_out[2034] <= ~layer2_out[6842];
     layer3_out[2035] <= layer2_out[8262] | layer2_out[8263];
     layer3_out[2036] <= ~layer2_out[6131];
     layer3_out[2037] <= layer2_out[720] | layer2_out[721];
     layer3_out[2038] <= layer2_out[715];
     layer3_out[2039] <= ~layer2_out[2905] | layer2_out[2904];
     layer3_out[2040] <= ~layer2_out[11];
     layer3_out[2041] <= ~layer2_out[6499] | layer2_out[6498];
     layer3_out[2042] <= ~layer2_out[10056] | layer2_out[10057];
     layer3_out[2043] <= layer2_out[8403] & ~layer2_out[8402];
     layer3_out[2044] <= layer2_out[2211] & layer2_out[2212];
     layer3_out[2045] <= ~layer2_out[10787];
     layer3_out[2046] <= ~layer2_out[3049];
     layer3_out[2047] <= ~layer2_out[7815] | layer2_out[7816];
     layer3_out[2048] <= layer2_out[6451];
     layer3_out[2049] <= layer2_out[824] | layer2_out[825];
     layer3_out[2050] <= ~layer2_out[9203];
     layer3_out[2051] <= layer2_out[10314] & layer2_out[10315];
     layer3_out[2052] <= layer2_out[6662];
     layer3_out[2053] <= ~layer2_out[4663];
     layer3_out[2054] <= ~layer2_out[7073];
     layer3_out[2055] <= ~(layer2_out[10538] | layer2_out[10539]);
     layer3_out[2056] <= layer2_out[1668];
     layer3_out[2057] <= layer2_out[8929];
     layer3_out[2058] <= layer2_out[2568];
     layer3_out[2059] <= layer2_out[10285];
     layer3_out[2060] <= layer2_out[8574];
     layer3_out[2061] <= ~(layer2_out[10654] & layer2_out[10655]);
     layer3_out[2062] <= ~(layer2_out[8874] ^ layer2_out[8875]);
     layer3_out[2063] <= ~(layer2_out[525] & layer2_out[526]);
     layer3_out[2064] <= ~layer2_out[2432];
     layer3_out[2065] <= layer2_out[4588] & ~layer2_out[4589];
     layer3_out[2066] <= layer2_out[11856] & layer2_out[11857];
     layer3_out[2067] <= layer2_out[11308];
     layer3_out[2068] <= layer2_out[10730];
     layer3_out[2069] <= ~layer2_out[7555];
     layer3_out[2070] <= layer2_out[4106] ^ layer2_out[4107];
     layer3_out[2071] <= ~layer2_out[10086];
     layer3_out[2072] <= ~layer2_out[10033];
     layer3_out[2073] <= layer2_out[5441] & layer2_out[5442];
     layer3_out[2074] <= layer2_out[6989];
     layer3_out[2075] <= layer2_out[6924] & ~layer2_out[6925];
     layer3_out[2076] <= ~layer2_out[6773];
     layer3_out[2077] <= ~layer2_out[5100];
     layer3_out[2078] <= layer2_out[2982] | layer2_out[2983];
     layer3_out[2079] <= layer2_out[6203];
     layer3_out[2080] <= ~layer2_out[2377] | layer2_out[2378];
     layer3_out[2081] <= layer2_out[4647] ^ layer2_out[4648];
     layer3_out[2082] <= ~layer2_out[4110] | layer2_out[4111];
     layer3_out[2083] <= ~layer2_out[6783] | layer2_out[6782];
     layer3_out[2084] <= ~layer2_out[369] | layer2_out[368];
     layer3_out[2085] <= layer2_out[6042];
     layer3_out[2086] <= ~(layer2_out[6653] ^ layer2_out[6654]);
     layer3_out[2087] <= ~(layer2_out[8298] & layer2_out[8299]);
     layer3_out[2088] <= layer2_out[6002] & ~layer2_out[6003];
     layer3_out[2089] <= ~layer2_out[5842] | layer2_out[5843];
     layer3_out[2090] <= layer2_out[10128] & ~layer2_out[10127];
     layer3_out[2091] <= layer2_out[10656];
     layer3_out[2092] <= ~layer2_out[11469];
     layer3_out[2093] <= ~layer2_out[9675];
     layer3_out[2094] <= layer2_out[6933] | layer2_out[6934];
     layer3_out[2095] <= layer2_out[11776];
     layer3_out[2096] <= layer2_out[1335];
     layer3_out[2097] <= layer2_out[11561] & ~layer2_out[11562];
     layer3_out[2098] <= layer2_out[5065];
     layer3_out[2099] <= ~layer2_out[6363];
     layer3_out[2100] <= ~(layer2_out[1469] ^ layer2_out[1470]);
     layer3_out[2101] <= layer2_out[4553];
     layer3_out[2102] <= ~layer2_out[4795];
     layer3_out[2103] <= ~layer2_out[4653];
     layer3_out[2104] <= ~(layer2_out[5460] & layer2_out[5461]);
     layer3_out[2105] <= layer2_out[9417];
     layer3_out[2106] <= ~(layer2_out[1556] & layer2_out[1557]);
     layer3_out[2107] <= layer2_out[6512] & ~layer2_out[6511];
     layer3_out[2108] <= ~(layer2_out[5087] | layer2_out[5088]);
     layer3_out[2109] <= layer2_out[7434] | layer2_out[7435];
     layer3_out[2110] <= ~layer2_out[2473] | layer2_out[2472];
     layer3_out[2111] <= ~layer2_out[3772];
     layer3_out[2112] <= ~layer2_out[1131] | layer2_out[1130];
     layer3_out[2113] <= layer2_out[5744];
     layer3_out[2114] <= ~layer2_out[7755] | layer2_out[7756];
     layer3_out[2115] <= ~(layer2_out[979] & layer2_out[980]);
     layer3_out[2116] <= layer2_out[3881] | layer2_out[3882];
     layer3_out[2117] <= layer2_out[9664] | layer2_out[9665];
     layer3_out[2118] <= ~(layer2_out[977] & layer2_out[978]);
     layer3_out[2119] <= ~layer2_out[3027];
     layer3_out[2120] <= ~(layer2_out[5190] & layer2_out[5191]);
     layer3_out[2121] <= layer2_out[2038];
     layer3_out[2122] <= layer2_out[10919];
     layer3_out[2123] <= layer2_out[4617];
     layer3_out[2124] <= layer2_out[11393];
     layer3_out[2125] <= ~layer2_out[10754];
     layer3_out[2126] <= ~layer2_out[8032];
     layer3_out[2127] <= layer2_out[4987] | layer2_out[4988];
     layer3_out[2128] <= ~layer2_out[2948] | layer2_out[2949];
     layer3_out[2129] <= layer2_out[4230] & ~layer2_out[4231];
     layer3_out[2130] <= ~(layer2_out[779] ^ layer2_out[780]);
     layer3_out[2131] <= ~(layer2_out[2876] | layer2_out[2877]);
     layer3_out[2132] <= ~(layer2_out[3026] | layer2_out[3027]);
     layer3_out[2133] <= layer2_out[2835] ^ layer2_out[2836];
     layer3_out[2134] <= ~layer2_out[9464] | layer2_out[9463];
     layer3_out[2135] <= layer2_out[3118];
     layer3_out[2136] <= ~layer2_out[9239];
     layer3_out[2137] <= layer2_out[431] ^ layer2_out[432];
     layer3_out[2138] <= layer2_out[5789] & ~layer2_out[5788];
     layer3_out[2139] <= layer2_out[10078] & ~layer2_out[10077];
     layer3_out[2140] <= ~layer2_out[3585];
     layer3_out[2141] <= ~layer2_out[7];
     layer3_out[2142] <= layer2_out[6986];
     layer3_out[2143] <= ~layer2_out[2842];
     layer3_out[2144] <= ~(layer2_out[10017] ^ layer2_out[10018]);
     layer3_out[2145] <= ~(layer2_out[546] ^ layer2_out[547]);
     layer3_out[2146] <= layer2_out[6335];
     layer3_out[2147] <= layer2_out[4858] & layer2_out[4859];
     layer3_out[2148] <= layer2_out[11963];
     layer3_out[2149] <= layer2_out[6432] & ~layer2_out[6431];
     layer3_out[2150] <= layer2_out[5514];
     layer3_out[2151] <= layer2_out[2210];
     layer3_out[2152] <= layer2_out[4851] ^ layer2_out[4852];
     layer3_out[2153] <= ~(layer2_out[9725] ^ layer2_out[9726]);
     layer3_out[2154] <= layer2_out[9272];
     layer3_out[2155] <= layer2_out[5485] | layer2_out[5486];
     layer3_out[2156] <= ~layer2_out[298];
     layer3_out[2157] <= ~layer2_out[11212] | layer2_out[11213];
     layer3_out[2158] <= ~layer2_out[1515];
     layer3_out[2159] <= ~(layer2_out[6611] ^ layer2_out[6612]);
     layer3_out[2160] <= layer2_out[5109] | layer2_out[5110];
     layer3_out[2161] <= ~(layer2_out[1417] & layer2_out[1418]);
     layer3_out[2162] <= layer2_out[8041];
     layer3_out[2163] <= layer2_out[6135] & layer2_out[6136];
     layer3_out[2164] <= ~layer2_out[4753] | layer2_out[4752];
     layer3_out[2165] <= ~(layer2_out[10166] & layer2_out[10167]);
     layer3_out[2166] <= layer2_out[2701] & layer2_out[2702];
     layer3_out[2167] <= layer2_out[7845] | layer2_out[7846];
     layer3_out[2168] <= ~(layer2_out[8355] & layer2_out[8356]);
     layer3_out[2169] <= ~layer2_out[509];
     layer3_out[2170] <= layer2_out[7553];
     layer3_out[2171] <= layer2_out[4931];
     layer3_out[2172] <= ~layer2_out[698];
     layer3_out[2173] <= ~layer2_out[1288];
     layer3_out[2174] <= ~layer2_out[7306];
     layer3_out[2175] <= ~(layer2_out[4613] | layer2_out[4614]);
     layer3_out[2176] <= ~layer2_out[6714] | layer2_out[6715];
     layer3_out[2177] <= layer2_out[7136];
     layer3_out[2178] <= layer2_out[3970] & ~layer2_out[3971];
     layer3_out[2179] <= layer2_out[463] ^ layer2_out[464];
     layer3_out[2180] <= ~layer2_out[9345];
     layer3_out[2181] <= layer2_out[7016] & ~layer2_out[7017];
     layer3_out[2182] <= ~layer2_out[2254] | layer2_out[2255];
     layer3_out[2183] <= layer2_out[8510];
     layer3_out[2184] <= layer2_out[743] | layer2_out[744];
     layer3_out[2185] <= layer2_out[672];
     layer3_out[2186] <= ~(layer2_out[1226] ^ layer2_out[1227]);
     layer3_out[2187] <= layer2_out[5044];
     layer3_out[2188] <= ~layer2_out[4329];
     layer3_out[2189] <= layer2_out[11789];
     layer3_out[2190] <= layer2_out[10055];
     layer3_out[2191] <= layer2_out[3705] & layer2_out[3706];
     layer3_out[2192] <= ~layer2_out[4380];
     layer3_out[2193] <= layer2_out[4832];
     layer3_out[2194] <= layer2_out[4290];
     layer3_out[2195] <= layer2_out[3438] | layer2_out[3439];
     layer3_out[2196] <= ~layer2_out[11364];
     layer3_out[2197] <= layer2_out[10851] & ~layer2_out[10852];
     layer3_out[2198] <= ~layer2_out[9915];
     layer3_out[2199] <= layer2_out[9169] ^ layer2_out[9170];
     layer3_out[2200] <= ~layer2_out[3974] | layer2_out[3975];
     layer3_out[2201] <= ~layer2_out[8044];
     layer3_out[2202] <= layer2_out[3160];
     layer3_out[2203] <= ~(layer2_out[3347] & layer2_out[3348]);
     layer3_out[2204] <= layer2_out[3198] & layer2_out[3199];
     layer3_out[2205] <= ~layer2_out[28];
     layer3_out[2206] <= layer2_out[3865];
     layer3_out[2207] <= layer2_out[11167] | layer2_out[11168];
     layer3_out[2208] <= layer2_out[11102];
     layer3_out[2209] <= ~layer2_out[4639] | layer2_out[4638];
     layer3_out[2210] <= layer2_out[10281];
     layer3_out[2211] <= ~(layer2_out[6938] ^ layer2_out[6939]);
     layer3_out[2212] <= ~(layer2_out[2236] & layer2_out[2237]);
     layer3_out[2213] <= ~layer2_out[4333];
     layer3_out[2214] <= ~layer2_out[4843];
     layer3_out[2215] <= layer2_out[1207] | layer2_out[1208];
     layer3_out[2216] <= ~layer2_out[4998];
     layer3_out[2217] <= ~(layer2_out[1962] ^ layer2_out[1963]);
     layer3_out[2218] <= layer2_out[10790];
     layer3_out[2219] <= ~(layer2_out[11183] ^ layer2_out[11184]);
     layer3_out[2220] <= ~layer2_out[11295];
     layer3_out[2221] <= ~(layer2_out[5311] ^ layer2_out[5312]);
     layer3_out[2222] <= layer2_out[9859];
     layer3_out[2223] <= layer2_out[3652];
     layer3_out[2224] <= layer2_out[8005];
     layer3_out[2225] <= ~(layer2_out[7621] ^ layer2_out[7622]);
     layer3_out[2226] <= ~layer2_out[7906];
     layer3_out[2227] <= ~layer2_out[11589];
     layer3_out[2228] <= layer2_out[11603];
     layer3_out[2229] <= layer2_out[8941];
     layer3_out[2230] <= ~layer2_out[9211] | layer2_out[9212];
     layer3_out[2231] <= ~(layer2_out[6368] & layer2_out[6369]);
     layer3_out[2232] <= layer2_out[1598];
     layer3_out[2233] <= ~(layer2_out[5591] & layer2_out[5592]);
     layer3_out[2234] <= layer2_out[761] & ~layer2_out[760];
     layer3_out[2235] <= layer2_out[380] & ~layer2_out[379];
     layer3_out[2236] <= layer2_out[7114];
     layer3_out[2237] <= ~layer2_out[8928] | layer2_out[8929];
     layer3_out[2238] <= layer2_out[9062];
     layer3_out[2239] <= ~(layer2_out[4558] & layer2_out[4559]);
     layer3_out[2240] <= layer2_out[9490];
     layer3_out[2241] <= layer2_out[6587] | layer2_out[6588];
     layer3_out[2242] <= layer2_out[4435];
     layer3_out[2243] <= ~layer2_out[2839];
     layer3_out[2244] <= ~(layer2_out[2300] | layer2_out[2301]);
     layer3_out[2245] <= ~layer2_out[8074] | layer2_out[8073];
     layer3_out[2246] <= layer2_out[11118] | layer2_out[11119];
     layer3_out[2247] <= ~layer2_out[9930];
     layer3_out[2248] <= layer2_out[10093];
     layer3_out[2249] <= layer2_out[11672];
     layer3_out[2250] <= ~(layer2_out[2437] & layer2_out[2438]);
     layer3_out[2251] <= ~(layer2_out[11360] & layer2_out[11361]);
     layer3_out[2252] <= layer2_out[6863];
     layer3_out[2253] <= layer2_out[6545];
     layer3_out[2254] <= layer2_out[2291];
     layer3_out[2255] <= ~(layer2_out[3436] & layer2_out[3437]);
     layer3_out[2256] <= layer2_out[2113];
     layer3_out[2257] <= ~layer2_out[7179];
     layer3_out[2258] <= layer2_out[9773];
     layer3_out[2259] <= layer2_out[10990] & ~layer2_out[10989];
     layer3_out[2260] <= layer2_out[2558];
     layer3_out[2261] <= ~layer2_out[8232];
     layer3_out[2262] <= layer2_out[3665];
     layer3_out[2263] <= layer2_out[4430];
     layer3_out[2264] <= layer2_out[8222] | layer2_out[8223];
     layer3_out[2265] <= ~layer2_out[4485];
     layer3_out[2266] <= ~layer2_out[4686];
     layer3_out[2267] <= ~(layer2_out[2556] & layer2_out[2557]);
     layer3_out[2268] <= ~layer2_out[11285] | layer2_out[11284];
     layer3_out[2269] <= layer2_out[3594] | layer2_out[3595];
     layer3_out[2270] <= layer2_out[11498];
     layer3_out[2271] <= ~layer2_out[2619] | layer2_out[2618];
     layer3_out[2272] <= ~(layer2_out[369] & layer2_out[370]);
     layer3_out[2273] <= ~layer2_out[10774];
     layer3_out[2274] <= layer2_out[8675] ^ layer2_out[8676];
     layer3_out[2275] <= layer2_out[399];
     layer3_out[2276] <= layer2_out[7260] & ~layer2_out[7259];
     layer3_out[2277] <= layer2_out[5035] | layer2_out[5036];
     layer3_out[2278] <= ~layer2_out[563] | layer2_out[564];
     layer3_out[2279] <= ~layer2_out[11064] | layer2_out[11065];
     layer3_out[2280] <= layer2_out[8670];
     layer3_out[2281] <= ~layer2_out[11493] | layer2_out[11492];
     layer3_out[2282] <= layer2_out[2935];
     layer3_out[2283] <= layer2_out[742] | layer2_out[743];
     layer3_out[2284] <= ~layer2_out[315] | layer2_out[316];
     layer3_out[2285] <= ~layer2_out[3685];
     layer3_out[2286] <= ~(layer2_out[6967] & layer2_out[6968]);
     layer3_out[2287] <= layer2_out[1778] ^ layer2_out[1779];
     layer3_out[2288] <= layer2_out[2379] ^ layer2_out[2380];
     layer3_out[2289] <= layer2_out[7344] & ~layer2_out[7345];
     layer3_out[2290] <= layer2_out[9441] & layer2_out[9442];
     layer3_out[2291] <= ~layer2_out[3958] | layer2_out[3957];
     layer3_out[2292] <= ~layer2_out[2884] | layer2_out[2883];
     layer3_out[2293] <= ~layer2_out[1248];
     layer3_out[2294] <= ~layer2_out[7916];
     layer3_out[2295] <= layer2_out[8646];
     layer3_out[2296] <= ~(layer2_out[8487] ^ layer2_out[8488]);
     layer3_out[2297] <= layer2_out[8494] & layer2_out[8495];
     layer3_out[2298] <= ~layer2_out[7496];
     layer3_out[2299] <= layer2_out[7577] | layer2_out[7578];
     layer3_out[2300] <= layer2_out[9891];
     layer3_out[2301] <= layer2_out[5551];
     layer3_out[2302] <= layer2_out[3758] | layer2_out[3759];
     layer3_out[2303] <= layer2_out[1484] | layer2_out[1485];
     layer3_out[2304] <= layer2_out[7602];
     layer3_out[2305] <= layer2_out[1473];
     layer3_out[2306] <= ~layer2_out[5029] | layer2_out[5028];
     layer3_out[2307] <= layer2_out[10448] | layer2_out[10449];
     layer3_out[2308] <= ~layer2_out[337];
     layer3_out[2309] <= ~(layer2_out[3072] | layer2_out[3073]);
     layer3_out[2310] <= ~layer2_out[7278] | layer2_out[7279];
     layer3_out[2311] <= layer2_out[11576] | layer2_out[11577];
     layer3_out[2312] <= layer2_out[4747] & ~layer2_out[4746];
     layer3_out[2313] <= ~(layer2_out[4567] ^ layer2_out[4568]);
     layer3_out[2314] <= ~layer2_out[4565];
     layer3_out[2315] <= ~layer2_out[6840];
     layer3_out[2316] <= layer2_out[10604] & ~layer2_out[10605];
     layer3_out[2317] <= ~(layer2_out[8100] ^ layer2_out[8101]);
     layer3_out[2318] <= ~layer2_out[4795];
     layer3_out[2319] <= ~(layer2_out[9269] | layer2_out[9270]);
     layer3_out[2320] <= ~layer2_out[11313];
     layer3_out[2321] <= layer2_out[9071];
     layer3_out[2322] <= ~layer2_out[2931];
     layer3_out[2323] <= ~layer2_out[5956];
     layer3_out[2324] <= ~(layer2_out[9234] ^ layer2_out[9235]);
     layer3_out[2325] <= ~layer2_out[3357] | layer2_out[3356];
     layer3_out[2326] <= layer2_out[11052];
     layer3_out[2327] <= layer2_out[10557];
     layer3_out[2328] <= ~(layer2_out[5940] & layer2_out[5941]);
     layer3_out[2329] <= ~layer2_out[1695];
     layer3_out[2330] <= layer2_out[2294] | layer2_out[2295];
     layer3_out[2331] <= ~(layer2_out[3] ^ layer2_out[4]);
     layer3_out[2332] <= ~layer2_out[6133];
     layer3_out[2333] <= ~(layer2_out[9304] & layer2_out[9305]);
     layer3_out[2334] <= ~(layer2_out[6378] & layer2_out[6379]);
     layer3_out[2335] <= layer2_out[5492] ^ layer2_out[5493];
     layer3_out[2336] <= ~layer2_out[4490] | layer2_out[4491];
     layer3_out[2337] <= layer2_out[7499] ^ layer2_out[7500];
     layer3_out[2338] <= layer2_out[4777] ^ layer2_out[4778];
     layer3_out[2339] <= ~(layer2_out[7244] & layer2_out[7245]);
     layer3_out[2340] <= layer2_out[1089] & layer2_out[1090];
     layer3_out[2341] <= ~(layer2_out[1264] & layer2_out[1265]);
     layer3_out[2342] <= ~(layer2_out[2245] ^ layer2_out[2246]);
     layer3_out[2343] <= layer2_out[5776];
     layer3_out[2344] <= ~layer2_out[2878];
     layer3_out[2345] <= layer2_out[8865] & ~layer2_out[8864];
     layer3_out[2346] <= layer2_out[8210] | layer2_out[8211];
     layer3_out[2347] <= ~layer2_out[8992];
     layer3_out[2348] <= layer2_out[2956] & ~layer2_out[2955];
     layer3_out[2349] <= ~layer2_out[8687];
     layer3_out[2350] <= layer2_out[1595] | layer2_out[1596];
     layer3_out[2351] <= layer2_out[1849];
     layer3_out[2352] <= ~(layer2_out[3327] | layer2_out[3328]);
     layer3_out[2353] <= ~layer2_out[3115];
     layer3_out[2354] <= ~layer2_out[476];
     layer3_out[2355] <= layer2_out[571];
     layer3_out[2356] <= ~(layer2_out[10399] & layer2_out[10400]);
     layer3_out[2357] <= layer2_out[8364];
     layer3_out[2358] <= layer2_out[8405];
     layer3_out[2359] <= ~(layer2_out[593] & layer2_out[594]);
     layer3_out[2360] <= ~(layer2_out[8793] & layer2_out[8794]);
     layer3_out[2361] <= ~(layer2_out[10702] ^ layer2_out[10703]);
     layer3_out[2362] <= ~(layer2_out[6663] ^ layer2_out[6664]);
     layer3_out[2363] <= ~(layer2_out[6301] ^ layer2_out[6302]);
     layer3_out[2364] <= ~layer2_out[11844] | layer2_out[11845];
     layer3_out[2365] <= layer2_out[304];
     layer3_out[2366] <= layer2_out[6381] | layer2_out[6382];
     layer3_out[2367] <= layer2_out[6283];
     layer3_out[2368] <= layer2_out[3550];
     layer3_out[2369] <= ~layer2_out[6058];
     layer3_out[2370] <= layer2_out[7888] | layer2_out[7889];
     layer3_out[2371] <= ~(layer2_out[5534] ^ layer2_out[5535]);
     layer3_out[2372] <= layer2_out[4399];
     layer3_out[2373] <= ~(layer2_out[3341] | layer2_out[3342]);
     layer3_out[2374] <= ~layer2_out[6101] | layer2_out[6102];
     layer3_out[2375] <= ~(layer2_out[8553] | layer2_out[8554]);
     layer3_out[2376] <= layer2_out[9601] ^ layer2_out[9602];
     layer3_out[2377] <= ~layer2_out[3841] | layer2_out[3842];
     layer3_out[2378] <= ~layer2_out[11666];
     layer3_out[2379] <= ~layer2_out[8690];
     layer3_out[2380] <= layer2_out[7596] | layer2_out[7597];
     layer3_out[2381] <= ~layer2_out[10744];
     layer3_out[2382] <= ~layer2_out[9258];
     layer3_out[2383] <= layer2_out[3166];
     layer3_out[2384] <= ~layer2_out[4465];
     layer3_out[2385] <= ~layer2_out[10922] | layer2_out[10921];
     layer3_out[2386] <= layer2_out[7374];
     layer3_out[2387] <= layer2_out[2909] | layer2_out[2910];
     layer3_out[2388] <= ~layer2_out[3635] | layer2_out[3636];
     layer3_out[2389] <= ~(layer2_out[3184] | layer2_out[3185]);
     layer3_out[2390] <= ~layer2_out[11679] | layer2_out[11678];
     layer3_out[2391] <= ~layer2_out[11783];
     layer3_out[2392] <= ~layer2_out[588];
     layer3_out[2393] <= layer2_out[9349] | layer2_out[9350];
     layer3_out[2394] <= layer2_out[4500] | layer2_out[4501];
     layer3_out[2395] <= ~layer2_out[9211];
     layer3_out[2396] <= layer2_out[11771] ^ layer2_out[11772];
     layer3_out[2397] <= ~(layer2_out[561] & layer2_out[562]);
     layer3_out[2398] <= ~layer2_out[5908];
     layer3_out[2399] <= ~(layer2_out[3294] ^ layer2_out[3295]);
     layer3_out[2400] <= layer2_out[10949] ^ layer2_out[10950];
     layer3_out[2401] <= ~(layer2_out[10699] ^ layer2_out[10700]);
     layer3_out[2402] <= layer2_out[5973] | layer2_out[5974];
     layer3_out[2403] <= layer2_out[2919];
     layer3_out[2404] <= ~(layer2_out[6190] ^ layer2_out[6191]);
     layer3_out[2405] <= layer2_out[10143];
     layer3_out[2406] <= layer2_out[2763] ^ layer2_out[2764];
     layer3_out[2407] <= ~layer2_out[9125];
     layer3_out[2408] <= layer2_out[2421] & ~layer2_out[2420];
     layer3_out[2409] <= layer2_out[3794] & ~layer2_out[3793];
     layer3_out[2410] <= ~layer2_out[9156];
     layer3_out[2411] <= ~(layer2_out[6891] | layer2_out[6892]);
     layer3_out[2412] <= ~(layer2_out[8756] & layer2_out[8757]);
     layer3_out[2413] <= layer2_out[5416] & ~layer2_out[5417];
     layer3_out[2414] <= ~(layer2_out[2719] ^ layer2_out[2720]);
     layer3_out[2415] <= ~layer2_out[10275];
     layer3_out[2416] <= ~(layer2_out[8702] | layer2_out[8703]);
     layer3_out[2417] <= layer2_out[4485] & ~layer2_out[4484];
     layer3_out[2418] <= layer2_out[1895] & ~layer2_out[1896];
     layer3_out[2419] <= ~layer2_out[7429];
     layer3_out[2420] <= ~layer2_out[10065];
     layer3_out[2421] <= layer2_out[10712];
     layer3_out[2422] <= ~layer2_out[11685];
     layer3_out[2423] <= layer2_out[11013];
     layer3_out[2424] <= layer2_out[1467] & ~layer2_out[1468];
     layer3_out[2425] <= layer2_out[11669] & ~layer2_out[11670];
     layer3_out[2426] <= ~layer2_out[2497] | layer2_out[2498];
     layer3_out[2427] <= layer2_out[9326] & ~layer2_out[9325];
     layer3_out[2428] <= layer2_out[5354] ^ layer2_out[5355];
     layer3_out[2429] <= layer2_out[8271] & ~layer2_out[8270];
     layer3_out[2430] <= layer2_out[3760] ^ layer2_out[3761];
     layer3_out[2431] <= ~layer2_out[10368];
     layer3_out[2432] <= layer2_out[2360] ^ layer2_out[2361];
     layer3_out[2433] <= layer2_out[1257];
     layer3_out[2434] <= ~(layer2_out[5125] ^ layer2_out[5126]);
     layer3_out[2435] <= layer2_out[10889] & ~layer2_out[10890];
     layer3_out[2436] <= ~layer2_out[7380];
     layer3_out[2437] <= layer2_out[534];
     layer3_out[2438] <= ~layer2_out[8591];
     layer3_out[2439] <= ~(layer2_out[11794] ^ layer2_out[11795]);
     layer3_out[2440] <= ~layer2_out[2198];
     layer3_out[2441] <= ~layer2_out[8756];
     layer3_out[2442] <= layer2_out[2126] & layer2_out[2127];
     layer3_out[2443] <= ~(layer2_out[8561] | layer2_out[8562]);
     layer3_out[2444] <= ~(layer2_out[11149] | layer2_out[11150]);
     layer3_out[2445] <= layer2_out[3766] ^ layer2_out[3767];
     layer3_out[2446] <= ~layer2_out[4166];
     layer3_out[2447] <= layer2_out[2912] & ~layer2_out[2913];
     layer3_out[2448] <= ~layer2_out[1992];
     layer3_out[2449] <= layer2_out[5261] ^ layer2_out[5262];
     layer3_out[2450] <= layer2_out[10413];
     layer3_out[2451] <= layer2_out[10586] ^ layer2_out[10587];
     layer3_out[2452] <= layer2_out[2175] ^ layer2_out[2176];
     layer3_out[2453] <= ~layer2_out[9016];
     layer3_out[2454] <= layer2_out[11129] ^ layer2_out[11130];
     layer3_out[2455] <= ~(layer2_out[1804] ^ layer2_out[1805]);
     layer3_out[2456] <= ~(layer2_out[2593] | layer2_out[2594]);
     layer3_out[2457] <= layer2_out[7312] & layer2_out[7313];
     layer3_out[2458] <= layer2_out[11893];
     layer3_out[2459] <= layer2_out[5577] & layer2_out[5578];
     layer3_out[2460] <= ~(layer2_out[4650] ^ layer2_out[4651]);
     layer3_out[2461] <= layer2_out[10706] & layer2_out[10707];
     layer3_out[2462] <= layer2_out[807];
     layer3_out[2463] <= ~layer2_out[9910];
     layer3_out[2464] <= layer2_out[1250] & ~layer2_out[1251];
     layer3_out[2465] <= ~(layer2_out[3963] ^ layer2_out[3964]);
     layer3_out[2466] <= layer2_out[4143];
     layer3_out[2467] <= ~(layer2_out[7745] ^ layer2_out[7746]);
     layer3_out[2468] <= layer2_out[2348];
     layer3_out[2469] <= ~layer2_out[1642] | layer2_out[1643];
     layer3_out[2470] <= ~layer2_out[1565] | layer2_out[1566];
     layer3_out[2471] <= layer2_out[4790] & ~layer2_out[4791];
     layer3_out[2472] <= layer2_out[5046] | layer2_out[5047];
     layer3_out[2473] <= layer2_out[10293] & layer2_out[10294];
     layer3_out[2474] <= layer2_out[3335] | layer2_out[3336];
     layer3_out[2475] <= ~layer2_out[9553];
     layer3_out[2476] <= layer2_out[10986] ^ layer2_out[10987];
     layer3_out[2477] <= layer2_out[4303] | layer2_out[4304];
     layer3_out[2478] <= layer2_out[8765] & ~layer2_out[8764];
     layer3_out[2479] <= layer2_out[4303] & ~layer2_out[4302];
     layer3_out[2480] <= layer2_out[5668] & layer2_out[5669];
     layer3_out[2481] <= ~(layer2_out[5129] | layer2_out[5130]);
     layer3_out[2482] <= ~(layer2_out[8879] | layer2_out[8880]);
     layer3_out[2483] <= ~layer2_out[1190];
     layer3_out[2484] <= layer2_out[974];
     layer3_out[2485] <= ~(layer2_out[3049] ^ layer2_out[3050]);
     layer3_out[2486] <= ~(layer2_out[3625] | layer2_out[3626]);
     layer3_out[2487] <= ~layer2_out[9629];
     layer3_out[2488] <= layer2_out[5721] & ~layer2_out[5720];
     layer3_out[2489] <= layer2_out[10812] & ~layer2_out[10813];
     layer3_out[2490] <= ~(layer2_out[8747] | layer2_out[8748]);
     layer3_out[2491] <= ~layer2_out[3144];
     layer3_out[2492] <= layer2_out[11562] & layer2_out[11563];
     layer3_out[2493] <= layer2_out[4877] & ~layer2_out[4876];
     layer3_out[2494] <= layer2_out[501];
     layer3_out[2495] <= layer2_out[11115] ^ layer2_out[11116];
     layer3_out[2496] <= layer2_out[3275] & ~layer2_out[3274];
     layer3_out[2497] <= ~(layer2_out[4127] ^ layer2_out[4128]);
     layer3_out[2498] <= layer2_out[4661] & ~layer2_out[4660];
     layer3_out[2499] <= layer2_out[6302] & layer2_out[6303];
     layer3_out[2500] <= layer2_out[11483];
     layer3_out[2501] <= layer2_out[581];
     layer3_out[2502] <= layer2_out[7004];
     layer3_out[2503] <= ~(layer2_out[1219] | layer2_out[1220]);
     layer3_out[2504] <= ~layer2_out[6540];
     layer3_out[2505] <= ~layer2_out[10505] | layer2_out[10504];
     layer3_out[2506] <= layer2_out[4337];
     layer3_out[2507] <= ~layer2_out[2972] | layer2_out[2971];
     layer3_out[2508] <= layer2_out[1182] & ~layer2_out[1183];
     layer3_out[2509] <= layer2_out[844];
     layer3_out[2510] <= layer2_out[8526] ^ layer2_out[8527];
     layer3_out[2511] <= ~(layer2_out[10420] ^ layer2_out[10421]);
     layer3_out[2512] <= ~(layer2_out[3460] ^ layer2_out[3461]);
     layer3_out[2513] <= ~layer2_out[2643];
     layer3_out[2514] <= layer2_out[7461];
     layer3_out[2515] <= ~(layer2_out[6020] & layer2_out[6021]);
     layer3_out[2516] <= layer2_out[2848] & layer2_out[2849];
     layer3_out[2517] <= layer2_out[11985];
     layer3_out[2518] <= ~(layer2_out[7330] ^ layer2_out[7331]);
     layer3_out[2519] <= layer2_out[5310];
     layer3_out[2520] <= layer2_out[7527];
     layer3_out[2521] <= ~(layer2_out[5237] ^ layer2_out[5238]);
     layer3_out[2522] <= ~(layer2_out[8099] ^ layer2_out[8100]);
     layer3_out[2523] <= layer2_out[1760] & layer2_out[1761];
     layer3_out[2524] <= ~(layer2_out[7094] ^ layer2_out[7095]);
     layer3_out[2525] <= layer2_out[9817];
     layer3_out[2526] <= layer2_out[334] & ~layer2_out[333];
     layer3_out[2527] <= layer2_out[2434] & ~layer2_out[2435];
     layer3_out[2528] <= ~layer2_out[3801];
     layer3_out[2529] <= ~(layer2_out[994] ^ layer2_out[995]);
     layer3_out[2530] <= layer2_out[38] & layer2_out[39];
     layer3_out[2531] <= ~layer2_out[4858];
     layer3_out[2532] <= layer2_out[7466] & ~layer2_out[7467];
     layer3_out[2533] <= ~layer2_out[5108];
     layer3_out[2534] <= layer2_out[4648] & ~layer2_out[4649];
     layer3_out[2535] <= layer2_out[2783] & ~layer2_out[2782];
     layer3_out[2536] <= ~(layer2_out[9514] ^ layer2_out[9515]);
     layer3_out[2537] <= layer2_out[4657] ^ layer2_out[4658];
     layer3_out[2538] <= layer2_out[1442];
     layer3_out[2539] <= ~layer2_out[11317] | layer2_out[11316];
     layer3_out[2540] <= layer2_out[6971];
     layer3_out[2541] <= ~(layer2_out[1662] ^ layer2_out[1663]);
     layer3_out[2542] <= ~layer2_out[3176];
     layer3_out[2543] <= layer2_out[7071] & ~layer2_out[7070];
     layer3_out[2544] <= layer2_out[5050];
     layer3_out[2545] <= ~layer2_out[10444];
     layer3_out[2546] <= layer2_out[4191] & ~layer2_out[4190];
     layer3_out[2547] <= layer2_out[8718] & ~layer2_out[8717];
     layer3_out[2548] <= layer2_out[5988];
     layer3_out[2549] <= ~(layer2_out[4361] | layer2_out[4362]);
     layer3_out[2550] <= layer2_out[1275] & layer2_out[1276];
     layer3_out[2551] <= ~(layer2_out[610] | layer2_out[611]);
     layer3_out[2552] <= layer2_out[2074] ^ layer2_out[2075];
     layer3_out[2553] <= layer2_out[5729];
     layer3_out[2554] <= layer2_out[8419] ^ layer2_out[8420];
     layer3_out[2555] <= layer2_out[11145] & layer2_out[11146];
     layer3_out[2556] <= ~(layer2_out[4969] | layer2_out[4970]);
     layer3_out[2557] <= ~layer2_out[1114] | layer2_out[1115];
     layer3_out[2558] <= layer2_out[5249] & ~layer2_out[5250];
     layer3_out[2559] <= layer2_out[10030] & ~layer2_out[10029];
     layer3_out[2560] <= layer2_out[2003] ^ layer2_out[2004];
     layer3_out[2561] <= ~layer2_out[271];
     layer3_out[2562] <= ~(layer2_out[6745] ^ layer2_out[6746]);
     layer3_out[2563] <= ~layer2_out[2614];
     layer3_out[2564] <= layer2_out[7145] | layer2_out[7146];
     layer3_out[2565] <= layer2_out[8776] & ~layer2_out[8775];
     layer3_out[2566] <= ~layer2_out[6141];
     layer3_out[2567] <= layer2_out[7405] | layer2_out[7406];
     layer3_out[2568] <= layer2_out[11636] & ~layer2_out[11635];
     layer3_out[2569] <= layer2_out[8712] & ~layer2_out[8713];
     layer3_out[2570] <= ~(layer2_out[10248] | layer2_out[10249]);
     layer3_out[2571] <= ~layer2_out[1992];
     layer3_out[2572] <= layer2_out[11958] & ~layer2_out[11959];
     layer3_out[2573] <= layer2_out[6816] & ~layer2_out[6815];
     layer3_out[2574] <= layer2_out[4837];
     layer3_out[2575] <= layer2_out[4661] & ~layer2_out[4662];
     layer3_out[2576] <= ~(layer2_out[7787] ^ layer2_out[7788]);
     layer3_out[2577] <= layer2_out[3920] ^ layer2_out[3921];
     layer3_out[2578] <= layer2_out[2160];
     layer3_out[2579] <= ~layer2_out[7173];
     layer3_out[2580] <= layer2_out[10869] | layer2_out[10870];
     layer3_out[2581] <= ~layer2_out[5996] | layer2_out[5995];
     layer3_out[2582] <= ~(layer2_out[7187] | layer2_out[7188]);
     layer3_out[2583] <= layer2_out[11409];
     layer3_out[2584] <= ~layer2_out[5521];
     layer3_out[2585] <= layer2_out[1077] ^ layer2_out[1078];
     layer3_out[2586] <= ~(layer2_out[491] | layer2_out[492]);
     layer3_out[2587] <= ~layer2_out[863];
     layer3_out[2588] <= layer2_out[1248];
     layer3_out[2589] <= layer2_out[3362] ^ layer2_out[3363];
     layer3_out[2590] <= layer2_out[5121] & ~layer2_out[5122];
     layer3_out[2591] <= ~(layer2_out[6344] ^ layer2_out[6345]);
     layer3_out[2592] <= ~layer2_out[7978];
     layer3_out[2593] <= layer2_out[8749];
     layer3_out[2594] <= layer2_out[7023] ^ layer2_out[7024];
     layer3_out[2595] <= ~(layer2_out[11504] | layer2_out[11505]);
     layer3_out[2596] <= layer2_out[2100];
     layer3_out[2597] <= ~(layer2_out[9760] | layer2_out[9761]);
     layer3_out[2598] <= ~layer2_out[5466];
     layer3_out[2599] <= ~(layer2_out[11624] ^ layer2_out[11625]);
     layer3_out[2600] <= ~(layer2_out[702] | layer2_out[703]);
     layer3_out[2601] <= layer2_out[7410] & layer2_out[7411];
     layer3_out[2602] <= layer2_out[837] ^ layer2_out[838];
     layer3_out[2603] <= ~layer2_out[11788];
     layer3_out[2604] <= ~(layer2_out[344] ^ layer2_out[345]);
     layer3_out[2605] <= ~layer2_out[1820];
     layer3_out[2606] <= layer2_out[6703] & ~layer2_out[6704];
     layer3_out[2607] <= layer2_out[1846] & ~layer2_out[1845];
     layer3_out[2608] <= layer2_out[11541] & ~layer2_out[11540];
     layer3_out[2609] <= layer2_out[6917];
     layer3_out[2610] <= layer2_out[5696] & ~layer2_out[5697];
     layer3_out[2611] <= layer2_out[6669];
     layer3_out[2612] <= layer2_out[3229] & ~layer2_out[3228];
     layer3_out[2613] <= layer2_out[10846] & layer2_out[10847];
     layer3_out[2614] <= layer2_out[11821];
     layer3_out[2615] <= ~layer2_out[5129];
     layer3_out[2616] <= layer2_out[5167] & layer2_out[5168];
     layer3_out[2617] <= layer2_out[649];
     layer3_out[2618] <= ~layer2_out[11111] | layer2_out[11112];
     layer3_out[2619] <= ~(layer2_out[6325] ^ layer2_out[6326]);
     layer3_out[2620] <= ~(layer2_out[766] ^ layer2_out[767]);
     layer3_out[2621] <= ~(layer2_out[1741] ^ layer2_out[1742]);
     layer3_out[2622] <= layer2_out[4154] ^ layer2_out[4155];
     layer3_out[2623] <= ~(layer2_out[10419] | layer2_out[10420]);
     layer3_out[2624] <= ~layer2_out[6893];
     layer3_out[2625] <= layer2_out[7162] & layer2_out[7163];
     layer3_out[2626] <= layer2_out[9135] & layer2_out[9136];
     layer3_out[2627] <= ~layer2_out[8119];
     layer3_out[2628] <= ~layer2_out[728] | layer2_out[729];
     layer3_out[2629] <= layer2_out[7579] & ~layer2_out[7580];
     layer3_out[2630] <= layer2_out[2258] ^ layer2_out[2259];
     layer3_out[2631] <= layer2_out[5785];
     layer3_out[2632] <= layer2_out[9034];
     layer3_out[2633] <= ~(layer2_out[5084] ^ layer2_out[5085]);
     layer3_out[2634] <= layer2_out[7780];
     layer3_out[2635] <= ~(layer2_out[8215] | layer2_out[8216]);
     layer3_out[2636] <= layer2_out[8085];
     layer3_out[2637] <= layer2_out[8063];
     layer3_out[2638] <= layer2_out[277] & ~layer2_out[276];
     layer3_out[2639] <= layer2_out[8548];
     layer3_out[2640] <= ~layer2_out[4228] | layer2_out[4227];
     layer3_out[2641] <= ~(layer2_out[3755] ^ layer2_out[3756]);
     layer3_out[2642] <= layer2_out[5984] | layer2_out[5985];
     layer3_out[2643] <= ~(layer2_out[1542] | layer2_out[1543]);
     layer3_out[2644] <= layer2_out[11554];
     layer3_out[2645] <= layer2_out[5929];
     layer3_out[2646] <= layer2_out[5023];
     layer3_out[2647] <= layer2_out[1069] ^ layer2_out[1070];
     layer3_out[2648] <= ~layer2_out[7055];
     layer3_out[2649] <= ~layer2_out[10535];
     layer3_out[2650] <= layer2_out[6472] ^ layer2_out[6473];
     layer3_out[2651] <= layer2_out[10556] & ~layer2_out[10557];
     layer3_out[2652] <= layer2_out[7784] ^ layer2_out[7785];
     layer3_out[2653] <= layer2_out[9948];
     layer3_out[2654] <= layer2_out[8473];
     layer3_out[2655] <= ~(layer2_out[9710] ^ layer2_out[9711]);
     layer3_out[2656] <= layer2_out[1185];
     layer3_out[2657] <= ~layer2_out[3508];
     layer3_out[2658] <= ~(layer2_out[7652] ^ layer2_out[7653]);
     layer3_out[2659] <= ~(layer2_out[2854] | layer2_out[2855]);
     layer3_out[2660] <= layer2_out[7227] | layer2_out[7228];
     layer3_out[2661] <= layer2_out[7471] ^ layer2_out[7472];
     layer3_out[2662] <= layer2_out[10478] & ~layer2_out[10477];
     layer3_out[2663] <= layer2_out[11200] & layer2_out[11201];
     layer3_out[2664] <= layer2_out[7165] & ~layer2_out[7164];
     layer3_out[2665] <= ~layer2_out[11626];
     layer3_out[2666] <= layer2_out[6716] ^ layer2_out[6717];
     layer3_out[2667] <= ~layer2_out[4257] | layer2_out[4258];
     layer3_out[2668] <= ~(layer2_out[9824] ^ layer2_out[9825]);
     layer3_out[2669] <= layer2_out[10894];
     layer3_out[2670] <= layer2_out[11918] & ~layer2_out[11917];
     layer3_out[2671] <= ~layer2_out[3592] | layer2_out[3593];
     layer3_out[2672] <= layer2_out[4118] & layer2_out[4119];
     layer3_out[2673] <= layer2_out[10894];
     layer3_out[2674] <= ~layer2_out[4079];
     layer3_out[2675] <= layer2_out[1986] ^ layer2_out[1987];
     layer3_out[2676] <= layer2_out[6886];
     layer3_out[2677] <= ~layer2_out[886] | layer2_out[887];
     layer3_out[2678] <= layer2_out[1632];
     layer3_out[2679] <= ~layer2_out[2206] | layer2_out[2207];
     layer3_out[2680] <= layer2_out[3834];
     layer3_out[2681] <= ~(layer2_out[3127] | layer2_out[3128]);
     layer3_out[2682] <= layer2_out[4457] ^ layer2_out[4458];
     layer3_out[2683] <= layer2_out[5173] & layer2_out[5174];
     layer3_out[2684] <= ~(layer2_out[5036] | layer2_out[5037]);
     layer3_out[2685] <= ~(layer2_out[11736] & layer2_out[11737]);
     layer3_out[2686] <= layer2_out[8681] & ~layer2_out[8680];
     layer3_out[2687] <= layer2_out[9705];
     layer3_out[2688] <= layer2_out[309] ^ layer2_out[310];
     layer3_out[2689] <= layer2_out[8199] & layer2_out[8200];
     layer3_out[2690] <= layer2_out[7773];
     layer3_out[2691] <= layer2_out[5335] & ~layer2_out[5334];
     layer3_out[2692] <= layer2_out[2977] & ~layer2_out[2976];
     layer3_out[2693] <= layer2_out[26] & layer2_out[27];
     layer3_out[2694] <= ~(layer2_out[4942] ^ layer2_out[4943]);
     layer3_out[2695] <= layer2_out[4838];
     layer3_out[2696] <= ~layer2_out[5925] | layer2_out[5926];
     layer3_out[2697] <= layer2_out[2059] ^ layer2_out[2060];
     layer3_out[2698] <= ~layer2_out[7296];
     layer3_out[2699] <= ~(layer2_out[3803] | layer2_out[3804]);
     layer3_out[2700] <= ~(layer2_out[3208] | layer2_out[3209]);
     layer3_out[2701] <= layer2_out[382] & ~layer2_out[381];
     layer3_out[2702] <= ~layer2_out[1348];
     layer3_out[2703] <= layer2_out[57];
     layer3_out[2704] <= layer2_out[4571] | layer2_out[4572];
     layer3_out[2705] <= ~layer2_out[730] | layer2_out[729];
     layer3_out[2706] <= layer2_out[9414] & ~layer2_out[9415];
     layer3_out[2707] <= layer2_out[9922] & ~layer2_out[9921];
     layer3_out[2708] <= ~(layer2_out[8849] ^ layer2_out[8850]);
     layer3_out[2709] <= layer2_out[7509] ^ layer2_out[7510];
     layer3_out[2710] <= layer2_out[4071];
     layer3_out[2711] <= ~layer2_out[3244];
     layer3_out[2712] <= layer2_out[6036];
     layer3_out[2713] <= layer2_out[826] & ~layer2_out[825];
     layer3_out[2714] <= layer2_out[7449];
     layer3_out[2715] <= layer2_out[134] & layer2_out[135];
     layer3_out[2716] <= ~(layer2_out[6764] & layer2_out[6765]);
     layer3_out[2717] <= ~(layer2_out[789] ^ layer2_out[790]);
     layer3_out[2718] <= ~layer2_out[4967] | layer2_out[4968];
     layer3_out[2719] <= ~layer2_out[1881] | layer2_out[1880];
     layer3_out[2720] <= layer2_out[3238];
     layer3_out[2721] <= ~layer2_out[7114];
     layer3_out[2722] <= layer2_out[8587] ^ layer2_out[8588];
     layer3_out[2723] <= ~layer2_out[10215];
     layer3_out[2724] <= ~(layer2_out[8782] & layer2_out[8783]);
     layer3_out[2725] <= ~layer2_out[8431];
     layer3_out[2726] <= layer2_out[5646] & ~layer2_out[5645];
     layer3_out[2727] <= ~(layer2_out[815] | layer2_out[816]);
     layer3_out[2728] <= ~layer2_out[2496] | layer2_out[2495];
     layer3_out[2729] <= layer2_out[2645];
     layer3_out[2730] <= layer2_out[2714] | layer2_out[2715];
     layer3_out[2731] <= layer2_out[4979] & ~layer2_out[4978];
     layer3_out[2732] <= layer2_out[11389] & ~layer2_out[11388];
     layer3_out[2733] <= layer2_out[9221] & layer2_out[9222];
     layer3_out[2734] <= ~layer2_out[8608];
     layer3_out[2735] <= layer2_out[10251];
     layer3_out[2736] <= ~(layer2_out[7354] ^ layer2_out[7355]);
     layer3_out[2737] <= layer2_out[1365];
     layer3_out[2738] <= layer2_out[8934];
     layer3_out[2739] <= layer2_out[4569] ^ layer2_out[4570];
     layer3_out[2740] <= ~(layer2_out[9363] | layer2_out[9364]);
     layer3_out[2741] <= ~(layer2_out[3477] | layer2_out[3478]);
     layer3_out[2742] <= ~(layer2_out[9055] | layer2_out[9056]);
     layer3_out[2743] <= layer2_out[4815] ^ layer2_out[4816];
     layer3_out[2744] <= ~(layer2_out[11403] ^ layer2_out[11404]);
     layer3_out[2745] <= ~(layer2_out[847] | layer2_out[848]);
     layer3_out[2746] <= layer2_out[3834] & ~layer2_out[3835];
     layer3_out[2747] <= ~layer2_out[1053] | layer2_out[1052];
     layer3_out[2748] <= ~(layer2_out[7806] | layer2_out[7807]);
     layer3_out[2749] <= layer2_out[932] & ~layer2_out[931];
     layer3_out[2750] <= ~layer2_out[4369];
     layer3_out[2751] <= layer2_out[978] & layer2_out[979];
     layer3_out[2752] <= ~(layer2_out[8967] ^ layer2_out[8968]);
     layer3_out[2753] <= ~(layer2_out[3729] & layer2_out[3730]);
     layer3_out[2754] <= ~(layer2_out[5366] ^ layer2_out[5367]);
     layer3_out[2755] <= layer2_out[6873] & layer2_out[6874];
     layer3_out[2756] <= layer2_out[7990] & ~layer2_out[7989];
     layer3_out[2757] <= layer2_out[2481];
     layer3_out[2758] <= layer2_out[3177] & ~layer2_out[3178];
     layer3_out[2759] <= layer2_out[9808];
     layer3_out[2760] <= ~(layer2_out[6067] ^ layer2_out[6068]);
     layer3_out[2761] <= layer2_out[10782];
     layer3_out[2762] <= layer2_out[2007] & layer2_out[2008];
     layer3_out[2763] <= ~(layer2_out[1169] ^ layer2_out[1170]);
     layer3_out[2764] <= ~(layer2_out[11879] | layer2_out[11880]);
     layer3_out[2765] <= layer2_out[4316] & ~layer2_out[4315];
     layer3_out[2766] <= ~layer2_out[10470];
     layer3_out[2767] <= ~layer2_out[10534];
     layer3_out[2768] <= layer2_out[2208];
     layer3_out[2769] <= layer2_out[8049] & ~layer2_out[8048];
     layer3_out[2770] <= layer2_out[9707];
     layer3_out[2771] <= layer2_out[5540] & ~layer2_out[5539];
     layer3_out[2772] <= layer2_out[10527];
     layer3_out[2773] <= layer2_out[8360];
     layer3_out[2774] <= layer2_out[1990] & ~layer2_out[1989];
     layer3_out[2775] <= layer2_out[8543];
     layer3_out[2776] <= layer2_out[8772] & ~layer2_out[8771];
     layer3_out[2777] <= layer2_out[11332] & layer2_out[11333];
     layer3_out[2778] <= ~(layer2_out[5331] ^ layer2_out[5332]);
     layer3_out[2779] <= ~(layer2_out[9200] & layer2_out[9201]);
     layer3_out[2780] <= ~(layer2_out[9645] ^ layer2_out[9646]);
     layer3_out[2781] <= layer2_out[11192];
     layer3_out[2782] <= ~(layer2_out[7512] | layer2_out[7513]);
     layer3_out[2783] <= ~(layer2_out[10038] ^ layer2_out[10039]);
     layer3_out[2784] <= layer2_out[3479] & ~layer2_out[3478];
     layer3_out[2785] <= ~layer2_out[10714];
     layer3_out[2786] <= ~(layer2_out[1800] ^ layer2_out[1801]);
     layer3_out[2787] <= ~layer2_out[7556];
     layer3_out[2788] <= layer2_out[1101];
     layer3_out[2789] <= ~layer2_out[3077];
     layer3_out[2790] <= ~layer2_out[3530];
     layer3_out[2791] <= layer2_out[2757];
     layer3_out[2792] <= layer2_out[8632] ^ layer2_out[8633];
     layer3_out[2793] <= ~(layer2_out[3484] ^ layer2_out[3485]);
     layer3_out[2794] <= ~(layer2_out[6724] & layer2_out[6725]);
     layer3_out[2795] <= ~(layer2_out[8327] ^ layer2_out[8328]);
     layer3_out[2796] <= ~layer2_out[4605];
     layer3_out[2797] <= layer2_out[5120];
     layer3_out[2798] <= layer2_out[5025] & layer2_out[5026];
     layer3_out[2799] <= layer2_out[4321] | layer2_out[4322];
     layer3_out[2800] <= layer2_out[11164];
     layer3_out[2801] <= ~(layer2_out[100] ^ layer2_out[101]);
     layer3_out[2802] <= layer2_out[5293] & ~layer2_out[5292];
     layer3_out[2803] <= layer2_out[11002];
     layer3_out[2804] <= layer2_out[5083] & ~layer2_out[5084];
     layer3_out[2805] <= layer2_out[5546] ^ layer2_out[5547];
     layer3_out[2806] <= layer2_out[8050] ^ layer2_out[8051];
     layer3_out[2807] <= ~layer2_out[1558];
     layer3_out[2808] <= layer2_out[77] | layer2_out[78];
     layer3_out[2809] <= ~(layer2_out[5666] ^ layer2_out[5667]);
     layer3_out[2810] <= ~(layer2_out[7610] ^ layer2_out[7611]);
     layer3_out[2811] <= ~layer2_out[8072] | layer2_out[8071];
     layer3_out[2812] <= ~layer2_out[6474];
     layer3_out[2813] <= ~(layer2_out[6487] | layer2_out[6488]);
     layer3_out[2814] <= ~layer2_out[439];
     layer3_out[2815] <= layer2_out[2077] & ~layer2_out[2078];
     layer3_out[2816] <= layer2_out[4432] ^ layer2_out[4433];
     layer3_out[2817] <= layer2_out[5387] & ~layer2_out[5388];
     layer3_out[2818] <= layer2_out[10722] ^ layer2_out[10723];
     layer3_out[2819] <= ~(layer2_out[6316] | layer2_out[6317]);
     layer3_out[2820] <= ~(layer2_out[489] | layer2_out[490]);
     layer3_out[2821] <= layer2_out[11256] & ~layer2_out[11255];
     layer3_out[2822] <= layer2_out[5746];
     layer3_out[2823] <= ~(layer2_out[2754] | layer2_out[2755]);
     layer3_out[2824] <= layer2_out[10716] & ~layer2_out[10717];
     layer3_out[2825] <= ~(layer2_out[2104] ^ layer2_out[2105]);
     layer3_out[2826] <= layer2_out[10021] & layer2_out[10022];
     layer3_out[2827] <= ~layer2_out[5583];
     layer3_out[2828] <= layer2_out[11875] & ~layer2_out[11876];
     layer3_out[2829] <= ~(layer2_out[11418] | layer2_out[11419]);
     layer3_out[2830] <= layer2_out[3278] ^ layer2_out[3279];
     layer3_out[2831] <= layer2_out[3911] ^ layer2_out[3912];
     layer3_out[2832] <= ~layer2_out[6175];
     layer3_out[2833] <= ~layer2_out[2509];
     layer3_out[2834] <= layer2_out[242] ^ layer2_out[243];
     layer3_out[2835] <= ~layer2_out[467] | layer2_out[468];
     layer3_out[2836] <= layer2_out[2649] & layer2_out[2650];
     layer3_out[2837] <= ~(layer2_out[4233] ^ layer2_out[4234]);
     layer3_out[2838] <= ~layer2_out[2408] | layer2_out[2407];
     layer3_out[2839] <= layer2_out[4733];
     layer3_out[2840] <= layer2_out[5511];
     layer3_out[2841] <= layer2_out[3217];
     layer3_out[2842] <= layer2_out[8208] ^ layer2_out[8209];
     layer3_out[2843] <= ~(layer2_out[11566] ^ layer2_out[11567]);
     layer3_out[2844] <= layer2_out[5715] & ~layer2_out[5714];
     layer3_out[2845] <= ~(layer2_out[7358] & layer2_out[7359]);
     layer3_out[2846] <= layer2_out[9387] & layer2_out[9388];
     layer3_out[2847] <= ~layer2_out[9820];
     layer3_out[2848] <= ~(layer2_out[723] | layer2_out[724]);
     layer3_out[2849] <= ~layer2_out[3554] | layer2_out[3553];
     layer3_out[2850] <= ~layer2_out[1513];
     layer3_out[2851] <= layer2_out[4561] ^ layer2_out[4562];
     layer3_out[2852] <= ~(layer2_out[2961] ^ layer2_out[2962]);
     layer3_out[2853] <= ~layer2_out[1329] | layer2_out[1328];
     layer3_out[2854] <= layer2_out[9566] & ~layer2_out[9567];
     layer3_out[2855] <= ~layer2_out[7626];
     layer3_out[2856] <= layer2_out[7921];
     layer3_out[2857] <= layer2_out[6324] & ~layer2_out[6325];
     layer3_out[2858] <= ~(layer2_out[9505] & layer2_out[9506]);
     layer3_out[2859] <= layer2_out[9539] ^ layer2_out[9540];
     layer3_out[2860] <= layer2_out[5869] & ~layer2_out[5868];
     layer3_out[2861] <= ~layer2_out[1263];
     layer3_out[2862] <= ~layer2_out[5188];
     layer3_out[2863] <= layer2_out[2417] & ~layer2_out[2416];
     layer3_out[2864] <= layer2_out[5434];
     layer3_out[2865] <= ~layer2_out[2091];
     layer3_out[2866] <= ~(layer2_out[5179] ^ layer2_out[5180]);
     layer3_out[2867] <= layer2_out[8241] & ~layer2_out[8242];
     layer3_out[2868] <= ~(layer2_out[4927] ^ layer2_out[4928]);
     layer3_out[2869] <= ~layer2_out[1552] | layer2_out[1551];
     layer3_out[2870] <= ~layer2_out[2965] | layer2_out[2966];
     layer3_out[2871] <= ~layer2_out[11491];
     layer3_out[2872] <= ~(layer2_out[3664] ^ layer2_out[3665]);
     layer3_out[2873] <= layer2_out[5871] & ~layer2_out[5872];
     layer3_out[2874] <= layer2_out[3453] | layer2_out[3454];
     layer3_out[2875] <= ~(layer2_out[2829] ^ layer2_out[2830]);
     layer3_out[2876] <= layer2_out[4782] ^ layer2_out[4783];
     layer3_out[2877] <= ~layer2_out[2386] | layer2_out[2387];
     layer3_out[2878] <= layer2_out[5866] ^ layer2_out[5867];
     layer3_out[2879] <= ~(layer2_out[7549] | layer2_out[7550]);
     layer3_out[2880] <= ~(layer2_out[9026] ^ layer2_out[9027]);
     layer3_out[2881] <= layer2_out[102];
     layer3_out[2882] <= layer2_out[9804] & ~layer2_out[9803];
     layer3_out[2883] <= ~(layer2_out[10673] | layer2_out[10674]);
     layer3_out[2884] <= layer2_out[8449];
     layer3_out[2885] <= layer2_out[4515];
     layer3_out[2886] <= layer2_out[9262];
     layer3_out[2887] <= layer2_out[6241];
     layer3_out[2888] <= layer2_out[124] & ~layer2_out[125];
     layer3_out[2889] <= layer2_out[2122];
     layer3_out[2890] <= layer2_out[2053];
     layer3_out[2891] <= layer2_out[10888] & ~layer2_out[10887];
     layer3_out[2892] <= layer2_out[7837];
     layer3_out[2893] <= layer2_out[6954];
     layer3_out[2894] <= layer2_out[1765];
     layer3_out[2895] <= ~(layer2_out[11688] & layer2_out[11689]);
     layer3_out[2896] <= layer2_out[2717] ^ layer2_out[2718];
     layer3_out[2897] <= layer2_out[4673];
     layer3_out[2898] <= layer2_out[6123];
     layer3_out[2899] <= layer2_out[4529];
     layer3_out[2900] <= ~layer2_out[7230] | layer2_out[7229];
     layer3_out[2901] <= layer2_out[2739];
     layer3_out[2902] <= layer2_out[10833] & layer2_out[10834];
     layer3_out[2903] <= layer2_out[6517];
     layer3_out[2904] <= layer2_out[4354];
     layer3_out[2905] <= ~(layer2_out[8350] | layer2_out[8351]);
     layer3_out[2906] <= ~(layer2_out[11961] & layer2_out[11962]);
     layer3_out[2907] <= layer2_out[2741] & ~layer2_out[2742];
     layer3_out[2908] <= ~layer2_out[7110];
     layer3_out[2909] <= layer2_out[6027];
     layer3_out[2910] <= ~(layer2_out[2442] ^ layer2_out[2443]);
     layer3_out[2911] <= ~(layer2_out[5597] | layer2_out[5598]);
     layer3_out[2912] <= ~layer2_out[4899];
     layer3_out[2913] <= ~layer2_out[11908];
     layer3_out[2914] <= ~layer2_out[385] | layer2_out[384];
     layer3_out[2915] <= layer2_out[243] ^ layer2_out[244];
     layer3_out[2916] <= layer2_out[7376] & ~layer2_out[7377];
     layer3_out[2917] <= ~layer2_out[4164];
     layer3_out[2918] <= ~layer2_out[9429] | layer2_out[9428];
     layer3_out[2919] <= layer2_out[5054] & ~layer2_out[5055];
     layer3_out[2920] <= ~layer2_out[3071];
     layer3_out[2921] <= ~(layer2_out[7726] ^ layer2_out[7727]);
     layer3_out[2922] <= layer2_out[5766] & ~layer2_out[5765];
     layer3_out[2923] <= layer2_out[11565] & ~layer2_out[11564];
     layer3_out[2924] <= layer2_out[4228] ^ layer2_out[4229];
     layer3_out[2925] <= layer2_out[11483];
     layer3_out[2926] <= ~layer2_out[1597];
     layer3_out[2927] <= ~layer2_out[4636] | layer2_out[4637];
     layer3_out[2928] <= layer2_out[1235] ^ layer2_out[1236];
     layer3_out[2929] <= layer2_out[1860] & ~layer2_out[1861];
     layer3_out[2930] <= layer2_out[10381] & ~layer2_out[10382];
     layer3_out[2931] <= ~layer2_out[2435];
     layer3_out[2932] <= ~(layer2_out[3450] ^ layer2_out[3451]);
     layer3_out[2933] <= layer2_out[4999] ^ layer2_out[5000];
     layer3_out[2934] <= ~layer2_out[253] | layer2_out[254];
     layer3_out[2935] <= layer2_out[8380] | layer2_out[8381];
     layer3_out[2936] <= ~layer2_out[2195];
     layer3_out[2937] <= layer2_out[8030] & ~layer2_out[8029];
     layer3_out[2938] <= layer2_out[10395] & layer2_out[10396];
     layer3_out[2939] <= layer2_out[4548];
     layer3_out[2940] <= ~layer2_out[2910];
     layer3_out[2941] <= ~layer2_out[3473];
     layer3_out[2942] <= ~(layer2_out[10601] | layer2_out[10602]);
     layer3_out[2943] <= layer2_out[10592] ^ layer2_out[10593];
     layer3_out[2944] <= ~layer2_out[5523];
     layer3_out[2945] <= layer2_out[2041] & ~layer2_out[2040];
     layer3_out[2946] <= layer2_out[9130] & ~layer2_out[9129];
     layer3_out[2947] <= layer2_out[4608] | layer2_out[4609];
     layer3_out[2948] <= ~(layer2_out[7718] ^ layer2_out[7719]);
     layer3_out[2949] <= ~(layer2_out[7608] ^ layer2_out[7609]);
     layer3_out[2950] <= layer2_out[4475];
     layer3_out[2951] <= layer2_out[5994];
     layer3_out[2952] <= layer2_out[5094];
     layer3_out[2953] <= layer2_out[5405] & ~layer2_out[5406];
     layer3_out[2954] <= ~(layer2_out[8176] | layer2_out[8177]);
     layer3_out[2955] <= ~layer2_out[6652];
     layer3_out[2956] <= layer2_out[953];
     layer3_out[2957] <= ~layer2_out[10029];
     layer3_out[2958] <= layer2_out[6016] & layer2_out[6017];
     layer3_out[2959] <= layer2_out[6405];
     layer3_out[2960] <= ~layer2_out[4950];
     layer3_out[2961] <= ~layer2_out[4424];
     layer3_out[2962] <= layer2_out[10751];
     layer3_out[2963] <= layer2_out[11413] & layer2_out[11414];
     layer3_out[2964] <= ~layer2_out[7134];
     layer3_out[2965] <= ~layer2_out[4566] | layer2_out[4565];
     layer3_out[2966] <= ~layer2_out[9592];
     layer3_out[2967] <= layer2_out[9767] | layer2_out[9768];
     layer3_out[2968] <= ~(layer2_out[4525] ^ layer2_out[4526]);
     layer3_out[2969] <= layer2_out[3367];
     layer3_out[2970] <= ~(layer2_out[2674] | layer2_out[2675]);
     layer3_out[2971] <= layer2_out[9328] ^ layer2_out[9329];
     layer3_out[2972] <= ~layer2_out[3716];
     layer3_out[2973] <= ~(layer2_out[8698] ^ layer2_out[8699]);
     layer3_out[2974] <= ~layer2_out[10426] | layer2_out[10427];
     layer3_out[2975] <= layer2_out[10218] ^ layer2_out[10219];
     layer3_out[2976] <= layer2_out[11698] & ~layer2_out[11697];
     layer3_out[2977] <= layer2_out[260];
     layer3_out[2978] <= ~layer2_out[1253];
     layer3_out[2979] <= ~layer2_out[4833];
     layer3_out[2980] <= layer2_out[1179];
     layer3_out[2981] <= layer2_out[1277] ^ layer2_out[1278];
     layer3_out[2982] <= layer2_out[4507];
     layer3_out[2983] <= layer2_out[1469] & ~layer2_out[1468];
     layer3_out[2984] <= ~layer2_out[746] | layer2_out[745];
     layer3_out[2985] <= layer2_out[2930];
     layer3_out[2986] <= layer2_out[5971] & ~layer2_out[5970];
     layer3_out[2987] <= ~(layer2_out[6961] & layer2_out[6962]);
     layer3_out[2988] <= layer2_out[3056];
     layer3_out[2989] <= layer2_out[11512];
     layer3_out[2990] <= ~(layer2_out[7247] & layer2_out[7248]);
     layer3_out[2991] <= ~(layer2_out[2733] ^ layer2_out[2734]);
     layer3_out[2992] <= layer2_out[7830] & layer2_out[7831];
     layer3_out[2993] <= layer2_out[4541] & ~layer2_out[4542];
     layer3_out[2994] <= layer2_out[10532];
     layer3_out[2995] <= layer2_out[1740];
     layer3_out[2996] <= layer2_out[7275];
     layer3_out[2997] <= layer2_out[1025] & ~layer2_out[1026];
     layer3_out[2998] <= layer2_out[1164] ^ layer2_out[1165];
     layer3_out[2999] <= layer2_out[8969] & ~layer2_out[8970];
     layer3_out[3000] <= ~layer2_out[19];
     layer3_out[3001] <= layer2_out[7928];
     layer3_out[3002] <= ~layer2_out[1642];
     layer3_out[3003] <= layer2_out[677] & layer2_out[678];
     layer3_out[3004] <= ~(layer2_out[11662] | layer2_out[11663]);
     layer3_out[3005] <= layer2_out[9040] ^ layer2_out[9041];
     layer3_out[3006] <= layer2_out[3639] ^ layer2_out[3640];
     layer3_out[3007] <= layer2_out[8203] & layer2_out[8204];
     layer3_out[3008] <= layer2_out[4071];
     layer3_out[3009] <= ~layer2_out[10331];
     layer3_out[3010] <= layer2_out[4784] & ~layer2_out[4785];
     layer3_out[3011] <= layer2_out[8958] & layer2_out[8959];
     layer3_out[3012] <= ~layer2_out[7783];
     layer3_out[3013] <= layer2_out[11798] & ~layer2_out[11797];
     layer3_out[3014] <= layer2_out[4622] & ~layer2_out[4621];
     layer3_out[3015] <= layer2_out[10727];
     layer3_out[3016] <= layer2_out[5034] & ~layer2_out[5035];
     layer3_out[3017] <= layer2_out[4744] ^ layer2_out[4745];
     layer3_out[3018] <= layer2_out[6508];
     layer3_out[3019] <= ~(layer2_out[10411] ^ layer2_out[10412]);
     layer3_out[3020] <= ~layer2_out[10314];
     layer3_out[3021] <= layer2_out[8584] ^ layer2_out[8585];
     layer3_out[3022] <= ~layer2_out[2634];
     layer3_out[3023] <= layer2_out[154];
     layer3_out[3024] <= layer2_out[783];
     layer3_out[3025] <= ~(layer2_out[7381] ^ layer2_out[7382]);
     layer3_out[3026] <= layer2_out[6802] ^ layer2_out[6803];
     layer3_out[3027] <= ~layer2_out[5122];
     layer3_out[3028] <= ~(layer2_out[4961] ^ layer2_out[4962]);
     layer3_out[3029] <= layer2_out[5971] & layer2_out[5972];
     layer3_out[3030] <= layer2_out[1414];
     layer3_out[3031] <= layer2_out[11448] | layer2_out[11449];
     layer3_out[3032] <= ~layer2_out[9257] | layer2_out[9258];
     layer3_out[3033] <= layer2_out[1871] | layer2_out[1872];
     layer3_out[3034] <= ~(layer2_out[5077] | layer2_out[5078]);
     layer3_out[3035] <= ~layer2_out[2862];
     layer3_out[3036] <= layer2_out[160];
     layer3_out[3037] <= layer2_out[11085] & layer2_out[11086];
     layer3_out[3038] <= ~layer2_out[8338];
     layer3_out[3039] <= layer2_out[7761];
     layer3_out[3040] <= layer2_out[9340] | layer2_out[9341];
     layer3_out[3041] <= layer2_out[3893] ^ layer2_out[3894];
     layer3_out[3042] <= ~layer2_out[7153];
     layer3_out[3043] <= ~layer2_out[3163];
     layer3_out[3044] <= ~(layer2_out[7286] & layer2_out[7287]);
     layer3_out[3045] <= ~layer2_out[4911];
     layer3_out[3046] <= layer2_out[1894] & layer2_out[1895];
     layer3_out[3047] <= ~layer2_out[519];
     layer3_out[3048] <= layer2_out[11752] & ~layer2_out[11753];
     layer3_out[3049] <= ~layer2_out[7301];
     layer3_out[3050] <= layer2_out[8760];
     layer3_out[3051] <= ~(layer2_out[3373] & layer2_out[3374]);
     layer3_out[3052] <= ~layer2_out[7375] | layer2_out[7376];
     layer3_out[3053] <= layer2_out[8772];
     layer3_out[3054] <= layer2_out[4887] & ~layer2_out[4886];
     layer3_out[3055] <= layer2_out[2919] & ~layer2_out[2918];
     layer3_out[3056] <= ~(layer2_out[9498] | layer2_out[9499]);
     layer3_out[3057] <= layer2_out[7118] ^ layer2_out[7119];
     layer3_out[3058] <= layer2_out[9058];
     layer3_out[3059] <= layer2_out[7911] | layer2_out[7912];
     layer3_out[3060] <= ~layer2_out[6585];
     layer3_out[3061] <= layer2_out[5529] ^ layer2_out[5530];
     layer3_out[3062] <= layer2_out[8829];
     layer3_out[3063] <= ~(layer2_out[5181] | layer2_out[5182]);
     layer3_out[3064] <= ~layer2_out[6805];
     layer3_out[3065] <= ~layer2_out[8165];
     layer3_out[3066] <= ~(layer2_out[3560] | layer2_out[3561]);
     layer3_out[3067] <= ~layer2_out[3434];
     layer3_out[3068] <= ~(layer2_out[3387] | layer2_out[3388]);
     layer3_out[3069] <= layer2_out[5399];
     layer3_out[3070] <= ~(layer2_out[1925] | layer2_out[1926]);
     layer3_out[3071] <= layer2_out[9912] ^ layer2_out[9913];
     layer3_out[3072] <= ~layer2_out[8372];
     layer3_out[3073] <= layer2_out[2944] | layer2_out[2945];
     layer3_out[3074] <= ~(layer2_out[5958] ^ layer2_out[5959]);
     layer3_out[3075] <= ~(layer2_out[7531] ^ layer2_out[7532]);
     layer3_out[3076] <= layer2_out[2745] ^ layer2_out[2746];
     layer3_out[3077] <= layer2_out[6552] & layer2_out[6553];
     layer3_out[3078] <= ~(layer2_out[9691] ^ layer2_out[9692]);
     layer3_out[3079] <= layer2_out[4438] ^ layer2_out[4439];
     layer3_out[3080] <= layer2_out[2353];
     layer3_out[3081] <= ~(layer2_out[1922] ^ layer2_out[1923]);
     layer3_out[3082] <= layer2_out[4365] | layer2_out[4366];
     layer3_out[3083] <= ~(layer2_out[1506] | layer2_out[1507]);
     layer3_out[3084] <= ~layer2_out[11691];
     layer3_out[3085] <= layer2_out[3405];
     layer3_out[3086] <= layer2_out[1415];
     layer3_out[3087] <= ~(layer2_out[11694] | layer2_out[11695]);
     layer3_out[3088] <= ~layer2_out[4149];
     layer3_out[3089] <= layer2_out[9139] & ~layer2_out[9138];
     layer3_out[3090] <= layer2_out[3593] & ~layer2_out[3594];
     layer3_out[3091] <= layer2_out[10596] ^ layer2_out[10597];
     layer3_out[3092] <= ~(layer2_out[9062] ^ layer2_out[9063]);
     layer3_out[3093] <= layer2_out[7707] & ~layer2_out[7708];
     layer3_out[3094] <= ~(layer2_out[11680] ^ layer2_out[11681]);
     layer3_out[3095] <= layer2_out[4808];
     layer3_out[3096] <= ~layer2_out[11569] | layer2_out[11568];
     layer3_out[3097] <= ~layer2_out[2851] | layer2_out[2852];
     layer3_out[3098] <= layer2_out[1143];
     layer3_out[3099] <= ~(layer2_out[6758] ^ layer2_out[6759]);
     layer3_out[3100] <= ~layer2_out[7924];
     layer3_out[3101] <= ~layer2_out[6141];
     layer3_out[3102] <= ~layer2_out[3421];
     layer3_out[3103] <= ~(layer2_out[11389] ^ layer2_out[11390]);
     layer3_out[3104] <= layer2_out[2002] ^ layer2_out[2003];
     layer3_out[3105] <= ~(layer2_out[5558] ^ layer2_out[5559]);
     layer3_out[3106] <= layer2_out[11421];
     layer3_out[3107] <= layer2_out[6874] & layer2_out[6875];
     layer3_out[3108] <= layer2_out[11383] & ~layer2_out[11382];
     layer3_out[3109] <= ~layer2_out[8825];
     layer3_out[3110] <= layer2_out[9153] ^ layer2_out[9154];
     layer3_out[3111] <= ~layer2_out[3108];
     layer3_out[3112] <= layer2_out[11064] & ~layer2_out[11063];
     layer3_out[3113] <= ~(layer2_out[9652] | layer2_out[9653]);
     layer3_out[3114] <= ~layer2_out[667];
     layer3_out[3115] <= layer2_out[2441];
     layer3_out[3116] <= layer2_out[5207];
     layer3_out[3117] <= ~layer2_out[11230];
     layer3_out[3118] <= ~(layer2_out[725] | layer2_out[726]);
     layer3_out[3119] <= ~(layer2_out[1090] ^ layer2_out[1091]);
     layer3_out[3120] <= ~(layer2_out[3872] ^ layer2_out[3873]);
     layer3_out[3121] <= layer2_out[7907] & layer2_out[7908];
     layer3_out[3122] <= layer2_out[4571];
     layer3_out[3123] <= layer2_out[7185];
     layer3_out[3124] <= layer2_out[5611];
     layer3_out[3125] <= ~layer2_out[6676];
     layer3_out[3126] <= layer2_out[425];
     layer3_out[3127] <= layer2_out[7252] ^ layer2_out[7253];
     layer3_out[3128] <= layer2_out[2411];
     layer3_out[3129] <= ~layer2_out[116];
     layer3_out[3130] <= ~layer2_out[7331];
     layer3_out[3131] <= layer2_out[1058] ^ layer2_out[1059];
     layer3_out[3132] <= layer2_out[8481];
     layer3_out[3133] <= layer2_out[4616] & ~layer2_out[4615];
     layer3_out[3134] <= ~(layer2_out[8479] & layer2_out[8480]);
     layer3_out[3135] <= layer2_out[2828] & ~layer2_out[2829];
     layer3_out[3136] <= ~layer2_out[10956];
     layer3_out[3137] <= layer2_out[6781] & ~layer2_out[6780];
     layer3_out[3138] <= layer2_out[889];
     layer3_out[3139] <= layer2_out[9219] ^ layer2_out[9220];
     layer3_out[3140] <= layer2_out[6350] & ~layer2_out[6351];
     layer3_out[3141] <= ~layer2_out[7979];
     layer3_out[3142] <= ~(layer2_out[3600] ^ layer2_out[3601]);
     layer3_out[3143] <= ~layer2_out[6074];
     layer3_out[3144] <= ~(layer2_out[1677] | layer2_out[1678]);
     layer3_out[3145] <= layer2_out[10148];
     layer3_out[3146] <= ~(layer2_out[6062] ^ layer2_out[6063]);
     layer3_out[3147] <= layer2_out[5813];
     layer3_out[3148] <= layer2_out[1] & ~layer2_out[2];
     layer3_out[3149] <= layer2_out[8076] & ~layer2_out[8075];
     layer3_out[3150] <= ~layer2_out[10062] | layer2_out[10061];
     layer3_out[3151] <= ~(layer2_out[2270] | layer2_out[2271]);
     layer3_out[3152] <= ~(layer2_out[3201] | layer2_out[3202]);
     layer3_out[3153] <= layer2_out[9798] & ~layer2_out[9797];
     layer3_out[3154] <= ~layer2_out[7137];
     layer3_out[3155] <= layer2_out[8204] & layer2_out[8205];
     layer3_out[3156] <= layer2_out[9348] & ~layer2_out[9349];
     layer3_out[3157] <= layer2_out[3720];
     layer3_out[3158] <= ~(layer2_out[2750] | layer2_out[2751]);
     layer3_out[3159] <= layer2_out[7172] & ~layer2_out[7171];
     layer3_out[3160] <= layer2_out[8227];
     layer3_out[3161] <= layer2_out[2606];
     layer3_out[3162] <= 1'b0;
     layer3_out[3163] <= ~(layer2_out[8456] | layer2_out[8457]);
     layer3_out[3164] <= layer2_out[1414] | layer2_out[1415];
     layer3_out[3165] <= ~(layer2_out[2124] ^ layer2_out[2125]);
     layer3_out[3166] <= ~layer2_out[11108];
     layer3_out[3167] <= layer2_out[5819] & ~layer2_out[5818];
     layer3_out[3168] <= ~(layer2_out[1260] ^ layer2_out[1261]);
     layer3_out[3169] <= layer2_out[11952];
     layer3_out[3170] <= layer2_out[3822] & ~layer2_out[3823];
     layer3_out[3171] <= layer2_out[1012] & ~layer2_out[1011];
     layer3_out[3172] <= ~(layer2_out[9064] | layer2_out[9065]);
     layer3_out[3173] <= ~(layer2_out[9936] & layer2_out[9937]);
     layer3_out[3174] <= ~(layer2_out[10969] ^ layer2_out[10970]);
     layer3_out[3175] <= layer2_out[1257];
     layer3_out[3176] <= ~layer2_out[8787];
     layer3_out[3177] <= ~layer2_out[3865];
     layer3_out[3178] <= ~layer2_out[7754];
     layer3_out[3179] <= layer2_out[9214] & ~layer2_out[9213];
     layer3_out[3180] <= ~(layer2_out[2784] & layer2_out[2785]);
     layer3_out[3181] <= ~(layer2_out[4018] | layer2_out[4019]);
     layer3_out[3182] <= layer2_out[4724] & layer2_out[4725];
     layer3_out[3183] <= ~layer2_out[8116];
     layer3_out[3184] <= layer2_out[10060] & layer2_out[10061];
     layer3_out[3185] <= ~(layer2_out[7040] | layer2_out[7041]);
     layer3_out[3186] <= layer2_out[2990] & ~layer2_out[2989];
     layer3_out[3187] <= layer2_out[7430] & ~layer2_out[7429];
     layer3_out[3188] <= ~layer2_out[6265];
     layer3_out[3189] <= ~(layer2_out[630] ^ layer2_out[631]);
     layer3_out[3190] <= ~layer2_out[5516];
     layer3_out[3191] <= ~(layer2_out[3043] ^ layer2_out[3044]);
     layer3_out[3192] <= layer2_out[2366] & ~layer2_out[2367];
     layer3_out[3193] <= layer2_out[8566] & ~layer2_out[8567];
     layer3_out[3194] <= ~layer2_out[9586];
     layer3_out[3195] <= layer2_out[11374] & ~layer2_out[11373];
     layer3_out[3196] <= ~(layer2_out[470] ^ layer2_out[471]);
     layer3_out[3197] <= ~layer2_out[10450];
     layer3_out[3198] <= layer2_out[11430] & ~layer2_out[11429];
     layer3_out[3199] <= ~(layer2_out[9567] | layer2_out[9568]);
     layer3_out[3200] <= layer2_out[9565] ^ layer2_out[9566];
     layer3_out[3201] <= layer2_out[7133] & ~layer2_out[7132];
     layer3_out[3202] <= ~layer2_out[6533];
     layer3_out[3203] <= ~(layer2_out[2933] | layer2_out[2934]);
     layer3_out[3204] <= layer2_out[2056] ^ layer2_out[2057];
     layer3_out[3205] <= ~(layer2_out[8161] | layer2_out[8162]);
     layer3_out[3206] <= layer2_out[7641] ^ layer2_out[7642];
     layer3_out[3207] <= ~layer2_out[3814];
     layer3_out[3208] <= layer2_out[11506];
     layer3_out[3209] <= layer2_out[1212] & ~layer2_out[1211];
     layer3_out[3210] <= layer2_out[42] ^ layer2_out[43];
     layer3_out[3211] <= ~(layer2_out[10282] ^ layer2_out[10283]);
     layer3_out[3212] <= ~layer2_out[5386];
     layer3_out[3213] <= layer2_out[4501] & ~layer2_out[4502];
     layer3_out[3214] <= ~layer2_out[7867] | layer2_out[7868];
     layer3_out[3215] <= layer2_out[10985] & ~layer2_out[10984];
     layer3_out[3216] <= ~(layer2_out[5303] & layer2_out[5304]);
     layer3_out[3217] <= layer2_out[11410] ^ layer2_out[11411];
     layer3_out[3218] <= layer2_out[3336];
     layer3_out[3219] <= ~layer2_out[1712];
     layer3_out[3220] <= layer2_out[2307] ^ layer2_out[2308];
     layer3_out[3221] <= ~(layer2_out[5259] ^ layer2_out[5260]);
     layer3_out[3222] <= layer2_out[1930] & ~layer2_out[1931];
     layer3_out[3223] <= layer2_out[5306];
     layer3_out[3224] <= layer2_out[11616] | layer2_out[11617];
     layer3_out[3225] <= ~layer2_out[2989];
     layer3_out[3226] <= ~layer2_out[9997] | layer2_out[9996];
     layer3_out[3227] <= layer2_out[6479];
     layer3_out[3228] <= layer2_out[251] & ~layer2_out[252];
     layer3_out[3229] <= layer2_out[9546] & ~layer2_out[9545];
     layer3_out[3230] <= layer2_out[4222];
     layer3_out[3231] <= layer2_out[3787] & layer2_out[3788];
     layer3_out[3232] <= ~(layer2_out[184] ^ layer2_out[185]);
     layer3_out[3233] <= layer2_out[5360];
     layer3_out[3234] <= ~layer2_out[5658];
     layer3_out[3235] <= ~(layer2_out[5643] ^ layer2_out[5644]);
     layer3_out[3236] <= ~layer2_out[3577];
     layer3_out[3237] <= layer2_out[9662] | layer2_out[9663];
     layer3_out[3238] <= ~layer2_out[5142];
     layer3_out[3239] <= ~layer2_out[76] | layer2_out[77];
     layer3_out[3240] <= layer2_out[2533] ^ layer2_out[2534];
     layer3_out[3241] <= layer2_out[8264] & ~layer2_out[8265];
     layer3_out[3242] <= layer2_out[10085] & ~layer2_out[10084];
     layer3_out[3243] <= layer2_out[3116];
     layer3_out[3244] <= layer2_out[10551] ^ layer2_out[10552];
     layer3_out[3245] <= layer2_out[302] ^ layer2_out[303];
     layer3_out[3246] <= ~layer2_out[8908];
     layer3_out[3247] <= ~layer2_out[7026];
     layer3_out[3248] <= ~layer2_out[11075];
     layer3_out[3249] <= ~layer2_out[9022];
     layer3_out[3250] <= layer2_out[2942];
     layer3_out[3251] <= ~layer2_out[1479];
     layer3_out[3252] <= ~layer2_out[9536];
     layer3_out[3253] <= ~(layer2_out[6787] | layer2_out[6788]);
     layer3_out[3254] <= ~layer2_out[6624] | layer2_out[6625];
     layer3_out[3255] <= layer2_out[11435];
     layer3_out[3256] <= layer2_out[6697];
     layer3_out[3257] <= layer2_out[10236];
     layer3_out[3258] <= ~layer2_out[5101];
     layer3_out[3259] <= layer2_out[3453] & ~layer2_out[3452];
     layer3_out[3260] <= layer2_out[8284];
     layer3_out[3261] <= layer2_out[10120];
     layer3_out[3262] <= layer2_out[11421] & ~layer2_out[11420];
     layer3_out[3263] <= ~(layer2_out[9764] & layer2_out[9765]);
     layer3_out[3264] <= ~layer2_out[10392] | layer2_out[10393];
     layer3_out[3265] <= ~layer2_out[4584] | layer2_out[4583];
     layer3_out[3266] <= ~layer2_out[6764];
     layer3_out[3267] <= layer2_out[4089] & layer2_out[4090];
     layer3_out[3268] <= layer2_out[1316] & ~layer2_out[1315];
     layer3_out[3269] <= layer2_out[1307];
     layer3_out[3270] <= layer2_out[3685];
     layer3_out[3271] <= layer2_out[3471];
     layer3_out[3272] <= ~(layer2_out[3131] | layer2_out[3132]);
     layer3_out[3273] <= ~layer2_out[10817];
     layer3_out[3274] <= layer2_out[7018] ^ layer2_out[7019];
     layer3_out[3275] <= layer2_out[5477];
     layer3_out[3276] <= ~layer2_out[3221];
     layer3_out[3277] <= layer2_out[6653] & ~layer2_out[6652];
     layer3_out[3278] <= layer2_out[9968] ^ layer2_out[9969];
     layer3_out[3279] <= layer2_out[733];
     layer3_out[3280] <= layer2_out[9376];
     layer3_out[3281] <= ~layer2_out[2867];
     layer3_out[3282] <= ~layer2_out[542] | layer2_out[541];
     layer3_out[3283] <= ~(layer2_out[4100] ^ layer2_out[4101]);
     layer3_out[3284] <= layer2_out[8979] & layer2_out[8980];
     layer3_out[3285] <= layer2_out[1647] ^ layer2_out[1648];
     layer3_out[3286] <= ~layer2_out[7095] | layer2_out[7096];
     layer3_out[3287] <= layer2_out[8171] & layer2_out[8172];
     layer3_out[3288] <= layer2_out[8673] | layer2_out[8674];
     layer3_out[3289] <= layer2_out[8315] & layer2_out[8316];
     layer3_out[3290] <= layer2_out[9712] & ~layer2_out[9713];
     layer3_out[3291] <= layer2_out[4167] & layer2_out[4168];
     layer3_out[3292] <= layer2_out[8493];
     layer3_out[3293] <= layer2_out[11594] & layer2_out[11595];
     layer3_out[3294] <= layer2_out[10925] & ~layer2_out[10924];
     layer3_out[3295] <= ~(layer2_out[6372] | layer2_out[6373]);
     layer3_out[3296] <= ~layer2_out[203];
     layer3_out[3297] <= layer2_out[6680] & ~layer2_out[6681];
     layer3_out[3298] <= layer2_out[11667];
     layer3_out[3299] <= layer2_out[11821];
     layer3_out[3300] <= layer2_out[11390] & ~layer2_out[11391];
     layer3_out[3301] <= layer2_out[11235] ^ layer2_out[11236];
     layer3_out[3302] <= layer2_out[9966] ^ layer2_out[9967];
     layer3_out[3303] <= layer2_out[7017] | layer2_out[7018];
     layer3_out[3304] <= layer2_out[6670] & layer2_out[6671];
     layer3_out[3305] <= layer2_out[7634] & ~layer2_out[7633];
     layer3_out[3306] <= layer2_out[814] & ~layer2_out[815];
     layer3_out[3307] <= layer2_out[8273] & ~layer2_out[8272];
     layer3_out[3308] <= ~(layer2_out[3823] | layer2_out[3824]);
     layer3_out[3309] <= layer2_out[9091];
     layer3_out[3310] <= layer2_out[10247] & ~layer2_out[10248];
     layer3_out[3311] <= ~(layer2_out[3697] & layer2_out[3698]);
     layer3_out[3312] <= layer2_out[3315] & layer2_out[3316];
     layer3_out[3313] <= layer2_out[9105] & ~layer2_out[9106];
     layer3_out[3314] <= layer2_out[653] & layer2_out[654];
     layer3_out[3315] <= layer2_out[7651] ^ layer2_out[7652];
     layer3_out[3316] <= layer2_out[11532] & layer2_out[11533];
     layer3_out[3317] <= ~(layer2_out[9046] ^ layer2_out[9047]);
     layer3_out[3318] <= ~layer2_out[7314];
     layer3_out[3319] <= ~layer2_out[6234] | layer2_out[6235];
     layer3_out[3320] <= ~(layer2_out[1728] ^ layer2_out[1729]);
     layer3_out[3321] <= layer2_out[8784] | layer2_out[8785];
     layer3_out[3322] <= ~(layer2_out[5503] ^ layer2_out[5504]);
     layer3_out[3323] <= ~layer2_out[1946];
     layer3_out[3324] <= ~(layer2_out[8556] | layer2_out[8557]);
     layer3_out[3325] <= ~(layer2_out[2683] | layer2_out[2684]);
     layer3_out[3326] <= layer2_out[1529] & ~layer2_out[1528];
     layer3_out[3327] <= ~layer2_out[3817];
     layer3_out[3328] <= layer2_out[2809] & ~layer2_out[2808];
     layer3_out[3329] <= layer2_out[5822] & ~layer2_out[5821];
     layer3_out[3330] <= ~layer2_out[9092] | layer2_out[9091];
     layer3_out[3331] <= layer2_out[9281];
     layer3_out[3332] <= layer2_out[9134] & ~layer2_out[9133];
     layer3_out[3333] <= ~layer2_out[963];
     layer3_out[3334] <= ~(layer2_out[7508] ^ layer2_out[7509]);
     layer3_out[3335] <= layer2_out[3757] & ~layer2_out[3758];
     layer3_out[3336] <= ~(layer2_out[3642] | layer2_out[3643]);
     layer3_out[3337] <= layer2_out[8340];
     layer3_out[3338] <= ~layer2_out[6362];
     layer3_out[3339] <= ~(layer2_out[10611] | layer2_out[10612]);
     layer3_out[3340] <= layer2_out[6032];
     layer3_out[3341] <= ~(layer2_out[2742] & layer2_out[2743]);
     layer3_out[3342] <= layer2_out[8867] ^ layer2_out[8868];
     layer3_out[3343] <= layer2_out[8124] & ~layer2_out[8125];
     layer3_out[3344] <= layer2_out[11710];
     layer3_out[3345] <= layer2_out[7700];
     layer3_out[3346] <= ~(layer2_out[10580] | layer2_out[10581]);
     layer3_out[3347] <= layer2_out[8292] & ~layer2_out[8293];
     layer3_out[3348] <= layer2_out[2404] & layer2_out[2405];
     layer3_out[3349] <= layer2_out[11385] & ~layer2_out[11384];
     layer3_out[3350] <= ~layer2_out[9820];
     layer3_out[3351] <= ~layer2_out[9853] | layer2_out[9854];
     layer3_out[3352] <= ~layer2_out[8162];
     layer3_out[3353] <= layer2_out[4227];
     layer3_out[3354] <= layer2_out[3492] ^ layer2_out[3493];
     layer3_out[3355] <= ~layer2_out[9394];
     layer3_out[3356] <= ~(layer2_out[11528] ^ layer2_out[11529]);
     layer3_out[3357] <= ~layer2_out[10090];
     layer3_out[3358] <= ~layer2_out[2909];
     layer3_out[3359] <= layer2_out[9865];
     layer3_out[3360] <= ~layer2_out[10548];
     layer3_out[3361] <= layer2_out[1775] & ~layer2_out[1774];
     layer3_out[3362] <= layer2_out[2809] | layer2_out[2810];
     layer3_out[3363] <= layer2_out[7630];
     layer3_out[3364] <= layer2_out[6364] ^ layer2_out[6365];
     layer3_out[3365] <= ~layer2_out[10975] | layer2_out[10974];
     layer3_out[3366] <= layer2_out[8037];
     layer3_out[3367] <= layer2_out[893];
     layer3_out[3368] <= ~(layer2_out[1428] | layer2_out[1429]);
     layer3_out[3369] <= layer2_out[11888] | layer2_out[11889];
     layer3_out[3370] <= ~layer2_out[1435];
     layer3_out[3371] <= layer2_out[254] ^ layer2_out[255];
     layer3_out[3372] <= layer2_out[9342] & ~layer2_out[9343];
     layer3_out[3373] <= ~layer2_out[11932];
     layer3_out[3374] <= ~(layer2_out[9447] ^ layer2_out[9448]);
     layer3_out[3375] <= ~(layer2_out[6068] | layer2_out[6069]);
     layer3_out[3376] <= layer2_out[6714];
     layer3_out[3377] <= ~layer2_out[5166];
     layer3_out[3378] <= layer2_out[10793] & layer2_out[10794];
     layer3_out[3379] <= layer2_out[5220] & layer2_out[5221];
     layer3_out[3380] <= ~layer2_out[8751] | layer2_out[8750];
     layer3_out[3381] <= layer2_out[4953];
     layer3_out[3382] <= layer2_out[4841] & layer2_out[4842];
     layer3_out[3383] <= layer2_out[8613];
     layer3_out[3384] <= ~(layer2_out[3404] ^ layer2_out[3405]);
     layer3_out[3385] <= ~layer2_out[10039];
     layer3_out[3386] <= layer2_out[3226] & ~layer2_out[3227];
     layer3_out[3387] <= layer2_out[2153];
     layer3_out[3388] <= layer2_out[4641] & layer2_out[4642];
     layer3_out[3389] <= ~layer2_out[4284];
     layer3_out[3390] <= layer2_out[7169];
     layer3_out[3391] <= ~(layer2_out[4094] ^ layer2_out[4095]);
     layer3_out[3392] <= ~layer2_out[3035];
     layer3_out[3393] <= ~layer2_out[3533];
     layer3_out[3394] <= layer2_out[11843];
     layer3_out[3395] <= ~layer2_out[2400];
     layer3_out[3396] <= ~layer2_out[7965];
     layer3_out[3397] <= ~(layer2_out[10184] ^ layer2_out[10185]);
     layer3_out[3398] <= ~layer2_out[11121];
     layer3_out[3399] <= layer2_out[5820] & ~layer2_out[5821];
     layer3_out[3400] <= ~layer2_out[5225];
     layer3_out[3401] <= ~layer2_out[7215];
     layer3_out[3402] <= ~layer2_out[11099];
     layer3_out[3403] <= ~(layer2_out[1135] ^ layer2_out[1136]);
     layer3_out[3404] <= layer2_out[5545] ^ layer2_out[5546];
     layer3_out[3405] <= layer2_out[6510] ^ layer2_out[6511];
     layer3_out[3406] <= ~(layer2_out[3402] | layer2_out[3403]);
     layer3_out[3407] <= layer2_out[6699] & ~layer2_out[6700];
     layer3_out[3408] <= ~(layer2_out[10408] | layer2_out[10409]);
     layer3_out[3409] <= layer2_out[11379];
     layer3_out[3410] <= layer2_out[7665];
     layer3_out[3411] <= ~layer2_out[9355];
     layer3_out[3412] <= ~layer2_out[9016];
     layer3_out[3413] <= ~(layer2_out[1305] ^ layer2_out[1306]);
     layer3_out[3414] <= ~(layer2_out[10923] | layer2_out[10924]);
     layer3_out[3415] <= layer2_out[5984] & ~layer2_out[5983];
     layer3_out[3416] <= layer2_out[2820] & layer2_out[2821];
     layer3_out[3417] <= layer2_out[8273] & layer2_out[8274];
     layer3_out[3418] <= layer2_out[3634] & ~layer2_out[3633];
     layer3_out[3419] <= ~(layer2_out[10632] ^ layer2_out[10633]);
     layer3_out[3420] <= layer2_out[1492] & ~layer2_out[1493];
     layer3_out[3421] <= layer2_out[5634] & layer2_out[5635];
     layer3_out[3422] <= layer2_out[7494] & layer2_out[7495];
     layer3_out[3423] <= layer2_out[8554];
     layer3_out[3424] <= ~layer2_out[1239] | layer2_out[1238];
     layer3_out[3425] <= layer2_out[10010];
     layer3_out[3426] <= ~(layer2_out[11592] ^ layer2_out[11593]);
     layer3_out[3427] <= layer2_out[8916] ^ layer2_out[8917];
     layer3_out[3428] <= ~(layer2_out[8475] & layer2_out[8476]);
     layer3_out[3429] <= layer2_out[5196] ^ layer2_out[5197];
     layer3_out[3430] <= ~layer2_out[6727];
     layer3_out[3431] <= layer2_out[3324] & layer2_out[3325];
     layer3_out[3432] <= layer2_out[10793];
     layer3_out[3433] <= ~layer2_out[7649];
     layer3_out[3434] <= layer2_out[6783] ^ layer2_out[6784];
     layer3_out[3435] <= layer2_out[4463] ^ layer2_out[4464];
     layer3_out[3436] <= layer2_out[1232] & ~layer2_out[1231];
     layer3_out[3437] <= ~layer2_out[714];
     layer3_out[3438] <= ~layer2_out[7789];
     layer3_out[3439] <= layer2_out[5019] & ~layer2_out[5018];
     layer3_out[3440] <= ~(layer2_out[2331] ^ layer2_out[2332]);
     layer3_out[3441] <= layer2_out[6687];
     layer3_out[3442] <= layer2_out[4391];
     layer3_out[3443] <= layer2_out[9574] & ~layer2_out[9575];
     layer3_out[3444] <= layer2_out[11003] ^ layer2_out[11004];
     layer3_out[3445] <= ~layer2_out[2013];
     layer3_out[3446] <= layer2_out[11947] & ~layer2_out[11946];
     layer3_out[3447] <= layer2_out[10344];
     layer3_out[3448] <= ~(layer2_out[10683] ^ layer2_out[10684]);
     layer3_out[3449] <= layer2_out[3815] & ~layer2_out[3816];
     layer3_out[3450] <= ~layer2_out[8082];
     layer3_out[3451] <= ~layer2_out[4411] | layer2_out[4412];
     layer3_out[3452] <= ~(layer2_out[1603] ^ layer2_out[1604]);
     layer3_out[3453] <= layer2_out[3119] ^ layer2_out[3120];
     layer3_out[3454] <= ~(layer2_out[7496] ^ layer2_out[7497]);
     layer3_out[3455] <= layer2_out[10478] & ~layer2_out[10479];
     layer3_out[3456] <= layer2_out[102] & ~layer2_out[103];
     layer3_out[3457] <= layer2_out[4619] | layer2_out[4620];
     layer3_out[3458] <= ~(layer2_out[5286] ^ layer2_out[5287]);
     layer3_out[3459] <= layer2_out[2971] & ~layer2_out[2970];
     layer3_out[3460] <= layer2_out[5511] & ~layer2_out[5510];
     layer3_out[3461] <= ~layer2_out[5658];
     layer3_out[3462] <= layer2_out[9224] ^ layer2_out[9225];
     layer3_out[3463] <= layer2_out[210] & layer2_out[211];
     layer3_out[3464] <= layer2_out[3442] & layer2_out[3443];
     layer3_out[3465] <= ~(layer2_out[7875] & layer2_out[7876]);
     layer3_out[3466] <= ~(layer2_out[3397] | layer2_out[3398]);
     layer3_out[3467] <= ~layer2_out[9654];
     layer3_out[3468] <= layer2_out[2055] ^ layer2_out[2056];
     layer3_out[3469] <= layer2_out[9708] ^ layer2_out[9709];
     layer3_out[3470] <= layer2_out[11630];
     layer3_out[3471] <= layer2_out[7842] & ~layer2_out[7841];
     layer3_out[3472] <= layer2_out[2987] & ~layer2_out[2988];
     layer3_out[3473] <= layer2_out[8743] & layer2_out[8744];
     layer3_out[3474] <= layer2_out[10899];
     layer3_out[3475] <= ~layer2_out[11501];
     layer3_out[3476] <= layer2_out[10393] & layer2_out[10394];
     layer3_out[3477] <= layer2_out[8722] & ~layer2_out[8723];
     layer3_out[3478] <= ~layer2_out[9733];
     layer3_out[3479] <= layer2_out[11060] & layer2_out[11061];
     layer3_out[3480] <= layer2_out[7311];
     layer3_out[3481] <= layer2_out[1015];
     layer3_out[3482] <= ~layer2_out[9141] | layer2_out[9140];
     layer3_out[3483] <= ~layer2_out[1698] | layer2_out[1697];
     layer3_out[3484] <= layer2_out[691] & layer2_out[692];
     layer3_out[3485] <= layer2_out[10545] & ~layer2_out[10546];
     layer3_out[3486] <= layer2_out[10125];
     layer3_out[3487] <= ~(layer2_out[3444] | layer2_out[3445]);
     layer3_out[3488] <= ~(layer2_out[11490] | layer2_out[11491]);
     layer3_out[3489] <= layer2_out[6428];
     layer3_out[3490] <= layer2_out[7157];
     layer3_out[3491] <= layer2_out[8127] & layer2_out[8128];
     layer3_out[3492] <= layer2_out[6416];
     layer3_out[3493] <= ~layer2_out[7010];
     layer3_out[3494] <= layer2_out[3425] & ~layer2_out[3426];
     layer3_out[3495] <= layer2_out[8016];
     layer3_out[3496] <= layer2_out[7366] & layer2_out[7367];
     layer3_out[3497] <= layer2_out[5822] | layer2_out[5823];
     layer3_out[3498] <= layer2_out[9403] ^ layer2_out[9404];
     layer3_out[3499] <= ~(layer2_out[8630] ^ layer2_out[8631]);
     layer3_out[3500] <= layer2_out[3493] ^ layer2_out[3494];
     layer3_out[3501] <= layer2_out[1038];
     layer3_out[3502] <= layer2_out[7014];
     layer3_out[3503] <= ~layer2_out[5653];
     layer3_out[3504] <= layer2_out[3679] ^ layer2_out[3680];
     layer3_out[3505] <= ~layer2_out[6353];
     layer3_out[3506] <= layer2_out[2832] ^ layer2_out[2833];
     layer3_out[3507] <= layer2_out[1835] & ~layer2_out[1836];
     layer3_out[3508] <= ~(layer2_out[2489] ^ layer2_out[2490]);
     layer3_out[3509] <= ~layer2_out[7626];
     layer3_out[3510] <= layer2_out[8206] ^ layer2_out[8207];
     layer3_out[3511] <= ~layer2_out[9631];
     layer3_out[3512] <= layer2_out[2125] ^ layer2_out[2126];
     layer3_out[3513] <= layer2_out[3918] & ~layer2_out[3917];
     layer3_out[3514] <= ~layer2_out[8911];
     layer3_out[3515] <= layer2_out[7057] & layer2_out[7058];
     layer3_out[3516] <= ~layer2_out[5214];
     layer3_out[3517] <= ~(layer2_out[10484] | layer2_out[10485]);
     layer3_out[3518] <= ~(layer2_out[7672] ^ layer2_out[7673]);
     layer3_out[3519] <= layer2_out[8159];
     layer3_out[3520] <= layer2_out[6563] & layer2_out[6564];
     layer3_out[3521] <= ~layer2_out[7010];
     layer3_out[3522] <= ~(layer2_out[10993] ^ layer2_out[10994]);
     layer3_out[3523] <= layer2_out[4405] & ~layer2_out[4404];
     layer3_out[3524] <= layer2_out[7285] & ~layer2_out[7284];
     layer3_out[3525] <= ~(layer2_out[8471] ^ layer2_out[8472]);
     layer3_out[3526] <= ~layer2_out[11232];
     layer3_out[3527] <= layer2_out[2410];
     layer3_out[3528] <= layer2_out[6475] & ~layer2_out[6476];
     layer3_out[3529] <= layer2_out[939];
     layer3_out[3530] <= layer2_out[2002];
     layer3_out[3531] <= layer2_out[11067] ^ layer2_out[11068];
     layer3_out[3532] <= layer2_out[10043] & layer2_out[10044];
     layer3_out[3533] <= ~layer2_out[10210];
     layer3_out[3534] <= layer2_out[10243] & ~layer2_out[10242];
     layer3_out[3535] <= ~layer2_out[1981];
     layer3_out[3536] <= layer2_out[11636] & layer2_out[11637];
     layer3_out[3537] <= ~(layer2_out[4423] | layer2_out[4424]);
     layer3_out[3538] <= layer2_out[11825] | layer2_out[11826];
     layer3_out[3539] <= layer2_out[4671] ^ layer2_out[4672];
     layer3_out[3540] <= layer2_out[9569] & ~layer2_out[9568];
     layer3_out[3541] <= layer2_out[661] & ~layer2_out[660];
     layer3_out[3542] <= layer2_out[4757] & layer2_out[4758];
     layer3_out[3543] <= layer2_out[4819];
     layer3_out[3544] <= layer2_out[8218];
     layer3_out[3545] <= layer2_out[1159] ^ layer2_out[1160];
     layer3_out[3546] <= layer2_out[15] & layer2_out[16];
     layer3_out[3547] <= ~layer2_out[173];
     layer3_out[3548] <= layer2_out[2635] ^ layer2_out[2636];
     layer3_out[3549] <= layer2_out[798] ^ layer2_out[799];
     layer3_out[3550] <= ~(layer2_out[6328] & layer2_out[6329]);
     layer3_out[3551] <= layer2_out[1167] & layer2_out[1168];
     layer3_out[3552] <= layer2_out[2836] | layer2_out[2837];
     layer3_out[3553] <= ~(layer2_out[8536] ^ layer2_out[8537]);
     layer3_out[3554] <= layer2_out[452];
     layer3_out[3555] <= ~layer2_out[8497];
     layer3_out[3556] <= layer2_out[7384];
     layer3_out[3557] <= layer2_out[3292] ^ layer2_out[3293];
     layer3_out[3558] <= ~(layer2_out[11924] ^ layer2_out[11925]);
     layer3_out[3559] <= ~layer2_out[5684];
     layer3_out[3560] <= layer2_out[4209] ^ layer2_out[4210];
     layer3_out[3561] <= ~layer2_out[3487];
     layer3_out[3562] <= layer2_out[1983];
     layer3_out[3563] <= layer2_out[1409];
     layer3_out[3564] <= layer2_out[1489] | layer2_out[1490];
     layer3_out[3565] <= layer2_out[3476] & ~layer2_out[3477];
     layer3_out[3566] <= layer2_out[3498] & ~layer2_out[3497];
     layer3_out[3567] <= layer2_out[11631];
     layer3_out[3568] <= layer2_out[11050] ^ layer2_out[11051];
     layer3_out[3569] <= ~(layer2_out[11046] | layer2_out[11047]);
     layer3_out[3570] <= ~(layer2_out[2469] ^ layer2_out[2470]);
     layer3_out[3571] <= layer2_out[5344];
     layer3_out[3572] <= layer2_out[343];
     layer3_out[3573] <= ~layer2_out[5724];
     layer3_out[3574] <= layer2_out[4977] & ~layer2_out[4978];
     layer3_out[3575] <= ~layer2_out[1002];
     layer3_out[3576] <= layer2_out[170] & ~layer2_out[171];
     layer3_out[3577] <= ~layer2_out[4160];
     layer3_out[3578] <= ~layer2_out[5637];
     layer3_out[3579] <= layer2_out[8246] & ~layer2_out[8247];
     layer3_out[3580] <= layer2_out[9314] & ~layer2_out[9313];
     layer3_out[3581] <= ~layer2_out[3986] | layer2_out[3985];
     layer3_out[3582] <= layer2_out[1564] & ~layer2_out[1565];
     layer3_out[3583] <= ~layer2_out[2116] | layer2_out[2117];
     layer3_out[3584] <= layer2_out[10823] & ~layer2_out[10822];
     layer3_out[3585] <= layer2_out[1724] ^ layer2_out[1725];
     layer3_out[3586] <= ~layer2_out[6747];
     layer3_out[3587] <= layer2_out[3770] & layer2_out[3771];
     layer3_out[3588] <= layer2_out[11238];
     layer3_out[3589] <= layer2_out[3574];
     layer3_out[3590] <= ~layer2_out[2426];
     layer3_out[3591] <= layer2_out[918] ^ layer2_out[919];
     layer3_out[3592] <= ~(layer2_out[6461] & layer2_out[6462]);
     layer3_out[3593] <= layer2_out[5847] ^ layer2_out[5848];
     layer3_out[3594] <= ~(layer2_out[2186] ^ layer2_out[2187]);
     layer3_out[3595] <= layer2_out[1620] & ~layer2_out[1621];
     layer3_out[3596] <= layer2_out[10501] & ~layer2_out[10500];
     layer3_out[3597] <= ~layer2_out[5239];
     layer3_out[3598] <= layer2_out[6421] & ~layer2_out[6422];
     layer3_out[3599] <= ~(layer2_out[4491] | layer2_out[4492]);
     layer3_out[3600] <= layer2_out[8625] & ~layer2_out[8624];
     layer3_out[3601] <= ~layer2_out[9087];
     layer3_out[3602] <= ~(layer2_out[3346] ^ layer2_out[3347]);
     layer3_out[3603] <= ~(layer2_out[10705] & layer2_out[10706]);
     layer3_out[3604] <= ~layer2_out[8921];
     layer3_out[3605] <= layer2_out[3623] & layer2_out[3624];
     layer3_out[3606] <= layer2_out[3253];
     layer3_out[3607] <= layer2_out[9411] | layer2_out[9412];
     layer3_out[3608] <= layer2_out[6626] & layer2_out[6627];
     layer3_out[3609] <= layer2_out[10281] ^ layer2_out[10282];
     layer3_out[3610] <= layer2_out[2522] | layer2_out[2523];
     layer3_out[3611] <= layer2_out[10351] & ~layer2_out[10352];
     layer3_out[3612] <= layer2_out[8774];
     layer3_out[3613] <= layer2_out[2672] | layer2_out[2673];
     layer3_out[3614] <= ~(layer2_out[8861] | layer2_out[8862]);
     layer3_out[3615] <= layer2_out[2323];
     layer3_out[3616] <= layer2_out[4999] & ~layer2_out[4998];
     layer3_out[3617] <= ~layer2_out[3664];
     layer3_out[3618] <= layer2_out[2412];
     layer3_out[3619] <= ~(layer2_out[1519] | layer2_out[1520]);
     layer3_out[3620] <= layer2_out[4034];
     layer3_out[3621] <= layer2_out[6357] ^ layer2_out[6358];
     layer3_out[3622] <= layer2_out[11163] ^ layer2_out[11164];
     layer3_out[3623] <= layer2_out[2120] & ~layer2_out[2121];
     layer3_out[3624] <= ~layer2_out[662] | layer2_out[663];
     layer3_out[3625] <= layer2_out[1358] ^ layer2_out[1359];
     layer3_out[3626] <= ~(layer2_out[4399] & layer2_out[4400]);
     layer3_out[3627] <= ~(layer2_out[8413] & layer2_out[8414]);
     layer3_out[3628] <= layer2_out[3431];
     layer3_out[3629] <= layer2_out[5320] & ~layer2_out[5319];
     layer3_out[3630] <= layer2_out[6336] & ~layer2_out[6337];
     layer3_out[3631] <= layer2_out[6456];
     layer3_out[3632] <= layer2_out[11365];
     layer3_out[3633] <= layer2_out[9115];
     layer3_out[3634] <= ~layer2_out[2457];
     layer3_out[3635] <= ~(layer2_out[1838] ^ layer2_out[1839]);
     layer3_out[3636] <= ~layer2_out[838] | layer2_out[839];
     layer3_out[3637] <= ~(layer2_out[3465] | layer2_out[3466]);
     layer3_out[3638] <= layer2_out[10637] ^ layer2_out[10638];
     layer3_out[3639] <= layer2_out[7801] ^ layer2_out[7802];
     layer3_out[3640] <= ~(layer2_out[10967] & layer2_out[10968]);
     layer3_out[3641] <= layer2_out[1343] & layer2_out[1344];
     layer3_out[3642] <= layer2_out[11938];
     layer3_out[3643] <= ~layer2_out[11076] | layer2_out[11075];
     layer3_out[3644] <= ~(layer2_out[11634] & layer2_out[11635]);
     layer3_out[3645] <= ~layer2_out[4455];
     layer3_out[3646] <= layer2_out[4014] & layer2_out[4015];
     layer3_out[3647] <= layer2_out[1726] & layer2_out[1727];
     layer3_out[3648] <= layer2_out[2670] & ~layer2_out[2671];
     layer3_out[3649] <= ~(layer2_out[11837] ^ layer2_out[11838]);
     layer3_out[3650] <= ~layer2_out[247];
     layer3_out[3651] <= layer2_out[7398] & layer2_out[7399];
     layer3_out[3652] <= ~layer2_out[6946];
     layer3_out[3653] <= ~layer2_out[3121] | layer2_out[3122];
     layer3_out[3654] <= ~layer2_out[628] | layer2_out[627];
     layer3_out[3655] <= layer2_out[6275] & ~layer2_out[6274];
     layer3_out[3656] <= layer2_out[7011] ^ layer2_out[7012];
     layer3_out[3657] <= ~layer2_out[4188];
     layer3_out[3658] <= ~layer2_out[2074];
     layer3_out[3659] <= ~(layer2_out[2303] & layer2_out[2304]);
     layer3_out[3660] <= ~layer2_out[2799];
     layer3_out[3661] <= layer2_out[6182];
     layer3_out[3662] <= layer2_out[6106] ^ layer2_out[6107];
     layer3_out[3663] <= layer2_out[3879];
     layer3_out[3664] <= ~layer2_out[9706];
     layer3_out[3665] <= ~layer2_out[11060];
     layer3_out[3666] <= layer2_out[4507];
     layer3_out[3667] <= layer2_out[1988] & ~layer2_out[1989];
     layer3_out[3668] <= layer2_out[3638] & ~layer2_out[3639];
     layer3_out[3669] <= layer2_out[9922] & layer2_out[9923];
     layer3_out[3670] <= layer2_out[1220];
     layer3_out[3671] <= layer2_out[3439];
     layer3_out[3672] <= ~(layer2_out[7216] ^ layer2_out[7217]);
     layer3_out[3673] <= ~(layer2_out[8069] | layer2_out[8070]);
     layer3_out[3674] <= layer2_out[3413];
     layer3_out[3675] <= ~layer2_out[8370] | layer2_out[8371];
     layer3_out[3676] <= layer2_out[6489] & ~layer2_out[6490];
     layer3_out[3677] <= ~layer2_out[2771];
     layer3_out[3678] <= ~(layer2_out[1770] ^ layer2_out[1771]);
     layer3_out[3679] <= ~layer2_out[638] | layer2_out[639];
     layer3_out[3680] <= layer2_out[5502] & ~layer2_out[5501];
     layer3_out[3681] <= layer2_out[456];
     layer3_out[3682] <= ~(layer2_out[4477] & layer2_out[4478]);
     layer3_out[3683] <= layer2_out[1032] & ~layer2_out[1033];
     layer3_out[3684] <= ~(layer2_out[6400] | layer2_out[6401]);
     layer3_out[3685] <= layer2_out[3545] & ~layer2_out[3546];
     layer3_out[3686] <= ~(layer2_out[7795] ^ layer2_out[7796]);
     layer3_out[3687] <= ~layer2_out[9371] | layer2_out[9370];
     layer3_out[3688] <= ~(layer2_out[11535] ^ layer2_out[11536]);
     layer3_out[3689] <= ~(layer2_out[4278] | layer2_out[4279]);
     layer3_out[3690] <= ~layer2_out[4597];
     layer3_out[3691] <= layer2_out[4336] | layer2_out[4337];
     layer3_out[3692] <= layer2_out[7760] | layer2_out[7761];
     layer3_out[3693] <= ~layer2_out[3329];
     layer3_out[3694] <= layer2_out[8216];
     layer3_out[3695] <= ~(layer2_out[4515] | layer2_out[4516]);
     layer3_out[3696] <= layer2_out[3012] ^ layer2_out[3013];
     layer3_out[3697] <= ~(layer2_out[9248] & layer2_out[9249]);
     layer3_out[3698] <= layer2_out[1043];
     layer3_out[3699] <= layer2_out[11997];
     layer3_out[3700] <= ~(layer2_out[1939] ^ layer2_out[1940]);
     layer3_out[3701] <= ~layer2_out[4521];
     layer3_out[3702] <= ~(layer2_out[5043] | layer2_out[5044]);
     layer3_out[3703] <= ~layer2_out[3171];
     layer3_out[3704] <= ~(layer2_out[1455] ^ layer2_out[1456]);
     layer3_out[3705] <= layer2_out[1121] ^ layer2_out[1122];
     layer3_out[3706] <= ~(layer2_out[3825] ^ layer2_out[3826]);
     layer3_out[3707] <= layer2_out[11727] & ~layer2_out[11726];
     layer3_out[3708] <= ~layer2_out[10350] | layer2_out[10349];
     layer3_out[3709] <= layer2_out[490] ^ layer2_out[491];
     layer3_out[3710] <= ~layer2_out[3511] | layer2_out[3512];
     layer3_out[3711] <= layer2_out[3228] & ~layer2_out[3227];
     layer3_out[3712] <= layer2_out[8655] ^ layer2_out[8656];
     layer3_out[3713] <= layer2_out[821];
     layer3_out[3714] <= layer2_out[8990] & ~layer2_out[8989];
     layer3_out[3715] <= layer2_out[2748];
     layer3_out[3716] <= layer2_out[63] ^ layer2_out[64];
     layer3_out[3717] <= layer2_out[813];
     layer3_out[3718] <= layer2_out[6507];
     layer3_out[3719] <= layer2_out[9392];
     layer3_out[3720] <= layer2_out[4696];
     layer3_out[3721] <= ~layer2_out[689] | layer2_out[688];
     layer3_out[3722] <= layer2_out[9971];
     layer3_out[3723] <= ~layer2_out[4713];
     layer3_out[3724] <= layer2_out[7952] ^ layer2_out[7953];
     layer3_out[3725] <= ~layer2_out[2923];
     layer3_out[3726] <= layer2_out[10273] ^ layer2_out[10274];
     layer3_out[3727] <= layer2_out[320];
     layer3_out[3728] <= ~layer2_out[10669];
     layer3_out[3729] <= layer2_out[11560];
     layer3_out[3730] <= layer2_out[7048];
     layer3_out[3731] <= ~layer2_out[4121] | layer2_out[4120];
     layer3_out[3732] <= ~(layer2_out[8130] ^ layer2_out[8131]);
     layer3_out[3733] <= ~layer2_out[5302];
     layer3_out[3734] <= ~(layer2_out[10468] | layer2_out[10469]);
     layer3_out[3735] <= layer2_out[7254] | layer2_out[7255];
     layer3_out[3736] <= layer2_out[5232];
     layer3_out[3737] <= layer2_out[8110];
     layer3_out[3738] <= ~layer2_out[10642] | layer2_out[10643];
     layer3_out[3739] <= layer2_out[2129] ^ layer2_out[2130];
     layer3_out[3740] <= layer2_out[6993];
     layer3_out[3741] <= layer2_out[7986] & ~layer2_out[7987];
     layer3_out[3742] <= layer2_out[4586];
     layer3_out[3743] <= ~(layer2_out[1791] ^ layer2_out[1792]);
     layer3_out[3744] <= ~(layer2_out[1736] & layer2_out[1737]);
     layer3_out[3745] <= ~layer2_out[5079];
     layer3_out[3746] <= layer2_out[4050] ^ layer2_out[4051];
     layer3_out[3747] <= ~layer2_out[10874];
     layer3_out[3748] <= ~(layer2_out[11487] | layer2_out[11488]);
     layer3_out[3749] <= layer2_out[8384] ^ layer2_out[8385];
     layer3_out[3750] <= ~(layer2_out[7698] ^ layer2_out[7699]);
     layer3_out[3751] <= layer2_out[9153];
     layer3_out[3752] <= layer2_out[5136] | layer2_out[5137];
     layer3_out[3753] <= layer2_out[5864];
     layer3_out[3754] <= layer2_out[5298] & layer2_out[5299];
     layer3_out[3755] <= layer2_out[4250] & ~layer2_out[4251];
     layer3_out[3756] <= layer2_out[329];
     layer3_out[3757] <= layer2_out[11035];
     layer3_out[3758] <= ~layer2_out[3666];
     layer3_out[3759] <= ~layer2_out[7124] | layer2_out[7125];
     layer3_out[3760] <= ~layer2_out[95];
     layer3_out[3761] <= layer2_out[4294];
     layer3_out[3762] <= ~(layer2_out[2299] ^ layer2_out[2300]);
     layer3_out[3763] <= layer2_out[7980] ^ layer2_out[7981];
     layer3_out[3764] <= layer2_out[5059];
     layer3_out[3765] <= ~layer2_out[6791];
     layer3_out[3766] <= ~layer2_out[11106];
     layer3_out[3767] <= layer2_out[7968];
     layer3_out[3768] <= layer2_out[2575] ^ layer2_out[2576];
     layer3_out[3769] <= ~layer2_out[2600] | layer2_out[2601];
     layer3_out[3770] <= ~layer2_out[684];
     layer3_out[3771] <= ~layer2_out[8157];
     layer3_out[3772] <= layer2_out[7657];
     layer3_out[3773] <= ~(layer2_out[2895] | layer2_out[2896]);
     layer3_out[3774] <= ~layer2_out[450];
     layer3_out[3775] <= ~layer2_out[2667] | layer2_out[2668];
     layer3_out[3776] <= ~layer2_out[1686];
     layer3_out[3777] <= layer2_out[7353] & layer2_out[7354];
     layer3_out[3778] <= layer2_out[11348];
     layer3_out[3779] <= layer2_out[11984] & layer2_out[11985];
     layer3_out[3780] <= ~layer2_out[4178];
     layer3_out[3781] <= layer2_out[9009] & ~layer2_out[9010];
     layer3_out[3782] <= layer2_out[5815] & ~layer2_out[5816];
     layer3_out[3783] <= ~(layer2_out[10311] ^ layer2_out[10312]);
     layer3_out[3784] <= ~layer2_out[2463];
     layer3_out[3785] <= ~(layer2_out[6878] & layer2_out[6879]);
     layer3_out[3786] <= ~layer2_out[4847] | layer2_out[4846];
     layer3_out[3787] <= ~layer2_out[441] | layer2_out[440];
     layer3_out[3788] <= ~layer2_out[947] | layer2_out[948];
     layer3_out[3789] <= layer2_out[123];
     layer3_out[3790] <= layer2_out[11296] & ~layer2_out[11297];
     layer3_out[3791] <= layer2_out[11394];
     layer3_out[3792] <= ~(layer2_out[4704] & layer2_out[4705]);
     layer3_out[3793] <= ~layer2_out[4327];
     layer3_out[3794] <= layer2_out[8778];
     layer3_out[3795] <= ~(layer2_out[430] ^ layer2_out[431]);
     layer3_out[3796] <= layer2_out[1491] & ~layer2_out[1492];
     layer3_out[3797] <= ~layer2_out[3961];
     layer3_out[3798] <= ~layer2_out[9135] | layer2_out[9134];
     layer3_out[3799] <= ~layer2_out[4866];
     layer3_out[3800] <= ~(layer2_out[1748] | layer2_out[1749]);
     layer3_out[3801] <= layer2_out[9181] & ~layer2_out[9180];
     layer3_out[3802] <= ~(layer2_out[3386] ^ layer2_out[3387]);
     layer3_out[3803] <= layer2_out[2446] ^ layer2_out[2447];
     layer3_out[3804] <= ~layer2_out[8392] | layer2_out[8393];
     layer3_out[3805] <= ~(layer2_out[4360] | layer2_out[4361]);
     layer3_out[3806] <= ~layer2_out[2219];
     layer3_out[3807] <= ~(layer2_out[8429] | layer2_out[8430]);
     layer3_out[3808] <= layer2_out[9118] & layer2_out[9119];
     layer3_out[3809] <= layer2_out[11333] & ~layer2_out[11334];
     layer3_out[3810] <= ~(layer2_out[5550] & layer2_out[5551]);
     layer3_out[3811] <= layer2_out[5283] ^ layer2_out[5284];
     layer3_out[3812] <= ~layer2_out[10880];
     layer3_out[3813] <= layer2_out[4123] | layer2_out[4124];
     layer3_out[3814] <= ~layer2_out[5777];
     layer3_out[3815] <= ~(layer2_out[3058] | layer2_out[3059]);
     layer3_out[3816] <= ~(layer2_out[5631] & layer2_out[5632]);
     layer3_out[3817] <= layer2_out[9719];
     layer3_out[3818] <= ~(layer2_out[4751] | layer2_out[4752]);
     layer3_out[3819] <= layer2_out[5041] ^ layer2_out[5042];
     layer3_out[3820] <= ~(layer2_out[9185] ^ layer2_out[9186]);
     layer3_out[3821] <= layer2_out[6038];
     layer3_out[3822] <= layer2_out[5465];
     layer3_out[3823] <= ~(layer2_out[10513] & layer2_out[10514]);
     layer3_out[3824] <= layer2_out[3115] & ~layer2_out[3114];
     layer3_out[3825] <= layer2_out[11413] & ~layer2_out[11412];
     layer3_out[3826] <= layer2_out[958] & layer2_out[959];
     layer3_out[3827] <= ~layer2_out[10665];
     layer3_out[3828] <= layer2_out[10219];
     layer3_out[3829] <= ~layer2_out[2778] | layer2_out[2777];
     layer3_out[3830] <= ~layer2_out[4113] | layer2_out[4112];
     layer3_out[3831] <= ~layer2_out[3191];
     layer3_out[3832] <= layer2_out[11579];
     layer3_out[3833] <= ~layer2_out[4698] | layer2_out[4699];
     layer3_out[3834] <= ~layer2_out[2640];
     layer3_out[3835] <= ~layer2_out[2771];
     layer3_out[3836] <= ~layer2_out[845] | layer2_out[846];
     layer3_out[3837] <= ~(layer2_out[10424] & layer2_out[10425]);
     layer3_out[3838] <= layer2_out[1696] ^ layer2_out[1697];
     layer3_out[3839] <= layer2_out[2120] & ~layer2_out[2119];
     layer3_out[3840] <= ~layer2_out[766];
     layer3_out[3841] <= ~(layer2_out[1794] | layer2_out[1795]);
     layer3_out[3842] <= ~layer2_out[11836];
     layer3_out[3843] <= layer2_out[8066];
     layer3_out[3844] <= ~layer2_out[3931] | layer2_out[3930];
     layer3_out[3845] <= layer2_out[10742];
     layer3_out[3846] <= ~layer2_out[1205];
     layer3_out[3847] <= ~(layer2_out[11047] ^ layer2_out[11048]);
     layer3_out[3848] <= ~layer2_out[1514] | layer2_out[1515];
     layer3_out[3849] <= layer2_out[5541] ^ layer2_out[5542];
     layer3_out[3850] <= ~layer2_out[10608];
     layer3_out[3851] <= ~(layer2_out[7303] ^ layer2_out[7304]);
     layer3_out[3852] <= layer2_out[7792] ^ layer2_out[7793];
     layer3_out[3853] <= ~(layer2_out[5823] | layer2_out[5824]);
     layer3_out[3854] <= layer2_out[11371] & ~layer2_out[11372];
     layer3_out[3855] <= ~(layer2_out[5838] ^ layer2_out[5839]);
     layer3_out[3856] <= ~layer2_out[4726];
     layer3_out[3857] <= layer2_out[7272] & ~layer2_out[7273];
     layer3_out[3858] <= ~layer2_out[5991];
     layer3_out[3859] <= ~layer2_out[7827];
     layer3_out[3860] <= layer2_out[7518];
     layer3_out[3861] <= ~layer2_out[10050];
     layer3_out[3862] <= layer2_out[7146] | layer2_out[7147];
     layer3_out[3863] <= ~layer2_out[6155];
     layer3_out[3864] <= layer2_out[2619];
     layer3_out[3865] <= ~(layer2_out[9512] ^ layer2_out[9513]);
     layer3_out[3866] <= layer2_out[1425] & ~layer2_out[1426];
     layer3_out[3867] <= ~(layer2_out[9643] ^ layer2_out[9644]);
     layer3_out[3868] <= layer2_out[3081];
     layer3_out[3869] <= ~(layer2_out[10886] ^ layer2_out[10887]);
     layer3_out[3870] <= layer2_out[9042];
     layer3_out[3871] <= layer2_out[8462];
     layer3_out[3872] <= layer2_out[9672] & ~layer2_out[9673];
     layer3_out[3873] <= layer2_out[5910] ^ layer2_out[5911];
     layer3_out[3874] <= ~(layer2_out[861] ^ layer2_out[862]);
     layer3_out[3875] <= layer2_out[1544];
     layer3_out[3876] <= layer2_out[8280] & ~layer2_out[8279];
     layer3_out[3877] <= ~(layer2_out[11210] | layer2_out[11211]);
     layer3_out[3878] <= ~layer2_out[7965];
     layer3_out[3879] <= layer2_out[6686] ^ layer2_out[6687];
     layer3_out[3880] <= layer2_out[10046] & layer2_out[10047];
     layer3_out[3881] <= ~(layer2_out[3987] | layer2_out[3988]);
     layer3_out[3882] <= ~(layer2_out[3269] ^ layer2_out[3270]);
     layer3_out[3883] <= ~layer2_out[6536];
     layer3_out[3884] <= layer2_out[2879] & layer2_out[2880];
     layer3_out[3885] <= layer2_out[10710] & ~layer2_out[10711];
     layer3_out[3886] <= ~(layer2_out[9692] | layer2_out[9693]);
     layer3_out[3887] <= ~layer2_out[7184];
     layer3_out[3888] <= ~layer2_out[9084];
     layer3_out[3889] <= layer2_out[4057];
     layer3_out[3890] <= layer2_out[1490];
     layer3_out[3891] <= ~(layer2_out[10378] | layer2_out[10379]);
     layer3_out[3892] <= ~layer2_out[8088];
     layer3_out[3893] <= layer2_out[4690];
     layer3_out[3894] <= layer2_out[2780];
     layer3_out[3895] <= ~layer2_out[2733] | layer2_out[2732];
     layer3_out[3896] <= layer2_out[1590] & ~layer2_out[1591];
     layer3_out[3897] <= layer2_out[11570] & layer2_out[11571];
     layer3_out[3898] <= ~layer2_out[4604];
     layer3_out[3899] <= layer2_out[10208] & ~layer2_out[10209];
     layer3_out[3900] <= ~(layer2_out[10953] ^ layer2_out[10954]);
     layer3_out[3901] <= ~(layer2_out[2145] ^ layer2_out[2146]);
     layer3_out[3902] <= ~layer2_out[603];
     layer3_out[3903] <= ~layer2_out[7276];
     layer3_out[3904] <= layer2_out[6712];
     layer3_out[3905] <= layer2_out[3141] & layer2_out[3142];
     layer3_out[3906] <= layer2_out[4082];
     layer3_out[3907] <= layer2_out[9243];
     layer3_out[3908] <= ~layer2_out[7222] | layer2_out[7223];
     layer3_out[3909] <= ~layer2_out[5998];
     layer3_out[3910] <= ~layer2_out[10631];
     layer3_out[3911] <= layer2_out[7262];
     layer3_out[3912] <= layer2_out[3989];
     layer3_out[3913] <= ~layer2_out[5504];
     layer3_out[3914] <= layer2_out[10762] & ~layer2_out[10761];
     layer3_out[3915] <= ~layer2_out[268];
     layer3_out[3916] <= ~layer2_out[8193] | layer2_out[8192];
     layer3_out[3917] <= layer2_out[5152] ^ layer2_out[5153];
     layer3_out[3918] <= layer2_out[6096] & ~layer2_out[6095];
     layer3_out[3919] <= layer2_out[6153];
     layer3_out[3920] <= ~(layer2_out[4378] | layer2_out[4379]);
     layer3_out[3921] <= ~layer2_out[6876];
     layer3_out[3922] <= layer2_out[751];
     layer3_out[3923] <= ~layer2_out[4381];
     layer3_out[3924] <= layer2_out[9471] & ~layer2_out[9472];
     layer3_out[3925] <= ~(layer2_out[8336] | layer2_out[8337]);
     layer3_out[3926] <= ~layer2_out[10161];
     layer3_out[3927] <= ~(layer2_out[6213] | layer2_out[6214]);
     layer3_out[3928] <= layer2_out[5937] ^ layer2_out[5938];
     layer3_out[3929] <= ~layer2_out[4895] | layer2_out[4896];
     layer3_out[3930] <= layer2_out[8873];
     layer3_out[3931] <= ~layer2_out[11282];
     layer3_out[3932] <= layer2_out[5845] & ~layer2_out[5844];
     layer3_out[3933] <= layer2_out[3913] & ~layer2_out[3912];
     layer3_out[3934] <= ~(layer2_out[5494] | layer2_out[5495]);
     layer3_out[3935] <= ~layer2_out[4059];
     layer3_out[3936] <= layer2_out[5464];
     layer3_out[3937] <= layer2_out[519] & ~layer2_out[520];
     layer3_out[3938] <= ~(layer2_out[2591] & layer2_out[2592]);
     layer3_out[3939] <= layer2_out[11005] ^ layer2_out[11006];
     layer3_out[3940] <= ~(layer2_out[6814] ^ layer2_out[6815]);
     layer3_out[3941] <= ~layer2_out[8704];
     layer3_out[3942] <= layer2_out[6223] ^ layer2_out[6224];
     layer3_out[3943] <= ~layer2_out[9964] | layer2_out[9965];
     layer3_out[3944] <= ~layer2_out[1500];
     layer3_out[3945] <= layer2_out[778] & ~layer2_out[779];
     layer3_out[3946] <= ~(layer2_out[10664] & layer2_out[10665]);
     layer3_out[3947] <= ~(layer2_out[3182] | layer2_out[3183]);
     layer3_out[3948] <= layer2_out[2334] & layer2_out[2335];
     layer3_out[3949] <= ~(layer2_out[2935] ^ layer2_out[2936]);
     layer3_out[3950] <= ~layer2_out[6629];
     layer3_out[3951] <= layer2_out[1769];
     layer3_out[3952] <= ~layer2_out[2594];
     layer3_out[3953] <= ~layer2_out[2032];
     layer3_out[3954] <= ~(layer2_out[11023] | layer2_out[11024]);
     layer3_out[3955] <= ~layer2_out[3904] | layer2_out[3903];
     layer3_out[3956] <= layer2_out[7541] ^ layer2_out[7542];
     layer3_out[3957] <= layer2_out[318];
     layer3_out[3958] <= layer2_out[11550] ^ layer2_out[11551];
     layer3_out[3959] <= layer2_out[590] | layer2_out[591];
     layer3_out[3960] <= ~layer2_out[3892] | layer2_out[3891];
     layer3_out[3961] <= layer2_out[5617];
     layer3_out[3962] <= ~layer2_out[2984];
     layer3_out[3963] <= ~(layer2_out[6162] | layer2_out[6163]);
     layer3_out[3964] <= ~layer2_out[2475];
     layer3_out[3965] <= ~layer2_out[5141];
     layer3_out[3966] <= ~(layer2_out[2166] & layer2_out[2167]);
     layer3_out[3967] <= ~layer2_out[3739];
     layer3_out[3968] <= layer2_out[11380];
     layer3_out[3969] <= layer2_out[3836];
     layer3_out[3970] <= ~(layer2_out[9193] | layer2_out[9194]);
     layer3_out[3971] <= ~layer2_out[1330];
     layer3_out[3972] <= ~layer2_out[7786];
     layer3_out[3973] <= layer2_out[5761];
     layer3_out[3974] <= ~layer2_out[5041] | layer2_out[5040];
     layer3_out[3975] <= layer2_out[6281];
     layer3_out[3976] <= layer2_out[383];
     layer3_out[3977] <= layer2_out[7941];
     layer3_out[3978] <= layer2_out[5443];
     layer3_out[3979] <= ~layer2_out[9961] | layer2_out[9962];
     layer3_out[3980] <= ~layer2_out[4099] | layer2_out[4100];
     layer3_out[3981] <= layer2_out[9063] & layer2_out[9064];
     layer3_out[3982] <= layer2_out[3749] | layer2_out[3750];
     layer3_out[3983] <= ~layer2_out[6439];
     layer3_out[3984] <= ~layer2_out[2421];
     layer3_out[3985] <= ~layer2_out[5156];
     layer3_out[3986] <= layer2_out[6144] ^ layer2_out[6145];
     layer3_out[3987] <= layer2_out[7401];
     layer3_out[3988] <= ~(layer2_out[5518] ^ layer2_out[5519]);
     layer3_out[3989] <= ~layer2_out[7931];
     layer3_out[3990] <= ~(layer2_out[4342] ^ layer2_out[4343]);
     layer3_out[3991] <= layer2_out[5317] ^ layer2_out[5318];
     layer3_out[3992] <= layer2_out[11431] | layer2_out[11432];
     layer3_out[3993] <= layer2_out[9381] & ~layer2_out[9382];
     layer3_out[3994] <= layer2_out[7082] & layer2_out[7083];
     layer3_out[3995] <= layer2_out[10434] ^ layer2_out[10435];
     layer3_out[3996] <= layer2_out[5263];
     layer3_out[3997] <= layer2_out[2205];
     layer3_out[3998] <= layer2_out[6453] & ~layer2_out[6452];
     layer3_out[3999] <= ~layer2_out[2552];
     layer3_out[4000] <= ~(layer2_out[7558] ^ layer2_out[7559]);
     layer3_out[4001] <= ~layer2_out[4722];
     layer3_out[4002] <= layer2_out[1851];
     layer3_out[4003] <= ~(layer2_out[8357] & layer2_out[8358]);
     layer3_out[4004] <= layer2_out[11151] ^ layer2_out[11152];
     layer3_out[4005] <= ~layer2_out[2015];
     layer3_out[4006] <= ~layer2_out[10705];
     layer3_out[4007] <= layer2_out[1657];
     layer3_out[4008] <= ~(layer2_out[4945] ^ layer2_out[4946]);
     layer3_out[4009] <= ~(layer2_out[2267] ^ layer2_out[2268]);
     layer3_out[4010] <= ~layer2_out[1736] | layer2_out[1735];
     layer3_out[4011] <= layer2_out[5158];
     layer3_out[4012] <= layer2_out[11380];
     layer3_out[4013] <= layer2_out[5915] & ~layer2_out[5916];
     layer3_out[4014] <= ~layer2_out[10254];
     layer3_out[4015] <= layer2_out[139] ^ layer2_out[140];
     layer3_out[4016] <= ~layer2_out[3496];
     layer3_out[4017] <= ~layer2_out[4812] | layer2_out[4811];
     layer3_out[4018] <= layer2_out[5797];
     layer3_out[4019] <= layer2_out[8122] ^ layer2_out[8123];
     layer3_out[4020] <= ~layer2_out[2163];
     layer3_out[4021] <= ~layer2_out[350];
     layer3_out[4022] <= layer2_out[6824] & layer2_out[6825];
     layer3_out[4023] <= ~(layer2_out[10027] ^ layer2_out[10028]);
     layer3_out[4024] <= ~layer2_out[9084];
     layer3_out[4025] <= ~layer2_out[5038];
     layer3_out[4026] <= ~layer2_out[8051];
     layer3_out[4027] <= layer2_out[6538];
     layer3_out[4028] <= ~layer2_out[3495];
     layer3_out[4029] <= ~(layer2_out[992] ^ layer2_out[993]);
     layer3_out[4030] <= layer2_out[11596] & layer2_out[11597];
     layer3_out[4031] <= ~layer2_out[354];
     layer3_out[4032] <= layer2_out[6902];
     layer3_out[4033] <= layer2_out[5947];
     layer3_out[4034] <= ~(layer2_out[8406] & layer2_out[8407]);
     layer3_out[4035] <= ~layer2_out[538];
     layer3_out[4036] <= ~(layer2_out[9333] ^ layer2_out[9334]);
     layer3_out[4037] <= ~(layer2_out[9973] ^ layer2_out[9974]);
     layer3_out[4038] <= ~(layer2_out[1694] ^ layer2_out[1695]);
     layer3_out[4039] <= ~layer2_out[217];
     layer3_out[4040] <= ~(layer2_out[2037] | layer2_out[2038]);
     layer3_out[4041] <= layer2_out[10863];
     layer3_out[4042] <= layer2_out[11046];
     layer3_out[4043] <= ~(layer2_out[10747] | layer2_out[10748]);
     layer3_out[4044] <= ~(layer2_out[2512] ^ layer2_out[2513]);
     layer3_out[4045] <= ~(layer2_out[4255] | layer2_out[4256]);
     layer3_out[4046] <= ~(layer2_out[3618] ^ layer2_out[3619]);
     layer3_out[4047] <= layer2_out[7147] | layer2_out[7148];
     layer3_out[4048] <= layer2_out[6113] ^ layer2_out[6114];
     layer3_out[4049] <= layer2_out[1261];
     layer3_out[4050] <= ~layer2_out[9522] | layer2_out[9523];
     layer3_out[4051] <= ~layer2_out[63];
     layer3_out[4052] <= ~(layer2_out[6833] & layer2_out[6834]);
     layer3_out[4053] <= layer2_out[8300] ^ layer2_out[8301];
     layer3_out[4054] <= ~layer2_out[2921];
     layer3_out[4055] <= ~layer2_out[4284];
     layer3_out[4056] <= layer2_out[5687];
     layer3_out[4057] <= layer2_out[1656] ^ layer2_out[1657];
     layer3_out[4058] <= ~layer2_out[8532] | layer2_out[8531];
     layer3_out[4059] <= ~layer2_out[11671];
     layer3_out[4060] <= layer2_out[759];
     layer3_out[4061] <= ~(layer2_out[8220] ^ layer2_out[8221]);
     layer3_out[4062] <= ~layer2_out[2763] | layer2_out[2762];
     layer3_out[4063] <= layer2_out[11926];
     layer3_out[4064] <= ~layer2_out[11505];
     layer3_out[4065] <= ~(layer2_out[10824] ^ layer2_out[10825]);
     layer3_out[4066] <= layer2_out[10320] & layer2_out[10321];
     layer3_out[4067] <= layer2_out[9962] ^ layer2_out[9963];
     layer3_out[4068] <= ~layer2_out[11043];
     layer3_out[4069] <= ~layer2_out[2592];
     layer3_out[4070] <= ~(layer2_out[8817] & layer2_out[8818]);
     layer3_out[4071] <= layer2_out[3369] ^ layer2_out[3370];
     layer3_out[4072] <= ~layer2_out[674];
     layer3_out[4073] <= layer2_out[6807];
     layer3_out[4074] <= ~layer2_out[4996];
     layer3_out[4075] <= ~layer2_out[10715];
     layer3_out[4076] <= layer2_out[9883] ^ layer2_out[9884];
     layer3_out[4077] <= ~(layer2_out[6593] & layer2_out[6594]);
     layer3_out[4078] <= layer2_out[5863] | layer2_out[5864];
     layer3_out[4079] <= layer2_out[4053];
     layer3_out[4080] <= ~layer2_out[11014];
     layer3_out[4081] <= ~(layer2_out[11138] ^ layer2_out[11139]);
     layer3_out[4082] <= ~(layer2_out[10521] & layer2_out[10522]);
     layer3_out[4083] <= layer2_out[7060] ^ layer2_out[7061];
     layer3_out[4084] <= ~layer2_out[1676];
     layer3_out[4085] <= layer2_out[11658] & ~layer2_out[11657];
     layer3_out[4086] <= ~layer2_out[5213];
     layer3_out[4087] <= layer2_out[1177];
     layer3_out[4088] <= ~layer2_out[7959];
     layer3_out[4089] <= ~layer2_out[1142];
     layer3_out[4090] <= ~(layer2_out[11303] | layer2_out[11304]);
     layer3_out[4091] <= layer2_out[7511] ^ layer2_out[7512];
     layer3_out[4092] <= layer2_out[9604] & ~layer2_out[9605];
     layer3_out[4093] <= ~layer2_out[1361];
     layer3_out[4094] <= layer2_out[9717] & ~layer2_out[9716];
     layer3_out[4095] <= ~layer2_out[3972] | layer2_out[3971];
     layer3_out[4096] <= ~layer2_out[11293];
     layer3_out[4097] <= layer2_out[10473];
     layer3_out[4098] <= layer2_out[3531] & ~layer2_out[3532];
     layer3_out[4099] <= layer2_out[9168] ^ layer2_out[9169];
     layer3_out[4100] <= layer2_out[9934] ^ layer2_out[9935];
     layer3_out[4101] <= layer2_out[2256];
     layer3_out[4102] <= ~layer2_out[8761] | layer2_out[8760];
     layer3_out[4103] <= ~layer2_out[4682];
     layer3_out[4104] <= ~layer2_out[2639];
     layer3_out[4105] <= ~(layer2_out[4308] & layer2_out[4309]);
     layer3_out[4106] <= ~(layer2_out[9685] & layer2_out[9686]);
     layer3_out[4107] <= ~layer2_out[589] | layer2_out[590];
     layer3_out[4108] <= layer2_out[11348];
     layer3_out[4109] <= layer2_out[2503] ^ layer2_out[2504];
     layer3_out[4110] <= layer2_out[7824];
     layer3_out[4111] <= layer2_out[4025] | layer2_out[4026];
     layer3_out[4112] <= ~layer2_out[6367];
     layer3_out[4113] <= layer2_out[4203];
     layer3_out[4114] <= layer2_out[804] | layer2_out[805];
     layer3_out[4115] <= layer2_out[3469] & ~layer2_out[3470];
     layer3_out[4116] <= layer2_out[11886] | layer2_out[11887];
     layer3_out[4117] <= ~layer2_out[8266];
     layer3_out[4118] <= layer2_out[10431];
     layer3_out[4119] <= layer2_out[9478];
     layer3_out[4120] <= ~(layer2_out[1901] | layer2_out[1902]);
     layer3_out[4121] <= ~layer2_out[10526];
     layer3_out[4122] <= ~(layer2_out[9309] ^ layer2_out[9310]);
     layer3_out[4123] <= ~layer2_out[6810] | layer2_out[6809];
     layer3_out[4124] <= layer2_out[11474];
     layer3_out[4125] <= ~(layer2_out[4044] & layer2_out[4045]);
     layer3_out[4126] <= ~(layer2_out[4771] & layer2_out[4772]);
     layer3_out[4127] <= layer2_out[10082] ^ layer2_out[10083];
     layer3_out[4128] <= ~layer2_out[4910] | layer2_out[4911];
     layer3_out[4129] <= ~layer2_out[2100];
     layer3_out[4130] <= ~layer2_out[4448];
     layer3_out[4131] <= ~(layer2_out[3301] | layer2_out[3302]);
     layer3_out[4132] <= ~layer2_out[10848];
     layer3_out[4133] <= layer2_out[9339] & ~layer2_out[9338];
     layer3_out[4134] <= ~(layer2_out[8940] | layer2_out[8941]);
     layer3_out[4135] <= ~layer2_out[3031];
     layer3_out[4136] <= layer2_out[10835] & ~layer2_out[10836];
     layer3_out[4137] <= layer2_out[4340];
     layer3_out[4138] <= layer2_out[6081];
     layer3_out[4139] <= layer2_out[10208];
     layer3_out[4140] <= layer2_out[1230] | layer2_out[1231];
     layer3_out[4141] <= layer2_out[10561] ^ layer2_out[10562];
     layer3_out[4142] <= layer2_out[5862];
     layer3_out[4143] <= ~layer2_out[1008];
     layer3_out[4144] <= ~layer2_out[1889] | layer2_out[1890];
     layer3_out[4145] <= ~layer2_out[1672];
     layer3_out[4146] <= ~layer2_out[7840];
     layer3_out[4147] <= layer2_out[10829] & ~layer2_out[10828];
     layer3_out[4148] <= layer2_out[11306] ^ layer2_out[11307];
     layer3_out[4149] <= layer2_out[10135];
     layer3_out[4150] <= ~layer2_out[11656] | layer2_out[11655];
     layer3_out[4151] <= ~layer2_out[5112] | layer2_out[5111];
     layer3_out[4152] <= ~layer2_out[11916];
     layer3_out[4153] <= ~layer2_out[2127];
     layer3_out[4154] <= layer2_out[11319];
     layer3_out[4155] <= layer2_out[10090] ^ layer2_out[10091];
     layer3_out[4156] <= ~layer2_out[9722];
     layer3_out[4157] <= layer2_out[6560];
     layer3_out[4158] <= layer2_out[57];
     layer3_out[4159] <= ~layer2_out[6316];
     layer3_out[4160] <= ~(layer2_out[5293] ^ layer2_out[5294]);
     layer3_out[4161] <= ~layer2_out[6094] | layer2_out[6093];
     layer3_out[4162] <= layer2_out[3368] ^ layer2_out[3369];
     layer3_out[4163] <= ~layer2_out[192];
     layer3_out[4164] <= ~layer2_out[9824] | layer2_out[9823];
     layer3_out[4165] <= layer2_out[10276] & ~layer2_out[10277];
     layer3_out[4166] <= layer2_out[2454];
     layer3_out[4167] <= ~layer2_out[4736];
     layer3_out[4168] <= layer2_out[4685];
     layer3_out[4169] <= layer2_out[9783];
     layer3_out[4170] <= layer2_out[6530] ^ layer2_out[6531];
     layer3_out[4171] <= ~layer2_out[10784] | layer2_out[10783];
     layer3_out[4172] <= ~(layer2_out[11217] ^ layer2_out[11218]);
     layer3_out[4173] <= layer2_out[9374];
     layer3_out[4174] <= layer2_out[7335] & ~layer2_out[7336];
     layer3_out[4175] <= ~layer2_out[10312] | layer2_out[10313];
     layer3_out[4176] <= ~layer2_out[8382];
     layer3_out[4177] <= ~layer2_out[2793] | layer2_out[2794];
     layer3_out[4178] <= ~(layer2_out[11511] | layer2_out[11512]);
     layer3_out[4179] <= ~layer2_out[1813];
     layer3_out[4180] <= layer2_out[10203];
     layer3_out[4181] <= layer2_out[7196];
     layer3_out[4182] <= layer2_out[421];
     layer3_out[4183] <= ~layer2_out[3261];
     layer3_out[4184] <= ~layer2_out[201];
     layer3_out[4185] <= layer2_out[7355] & layer2_out[7356];
     layer3_out[4186] <= layer2_out[9201];
     layer3_out[4187] <= layer2_out[7453];
     layer3_out[4188] <= ~(layer2_out[6294] | layer2_out[6295]);
     layer3_out[4189] <= ~layer2_out[1498];
     layer3_out[4190] <= layer2_out[6216] & layer2_out[6217];
     layer3_out[4191] <= ~layer2_out[6617];
     layer3_out[4192] <= ~(layer2_out[6286] | layer2_out[6287]);
     layer3_out[4193] <= ~layer2_out[8492];
     layer3_out[4194] <= ~layer2_out[5570] | layer2_out[5569];
     layer3_out[4195] <= ~layer2_out[11951];
     layer3_out[4196] <= layer2_out[8055] & layer2_out[8056];
     layer3_out[4197] <= ~(layer2_out[2115] ^ layer2_out[2116]);
     layer3_out[4198] <= layer2_out[9897] ^ layer2_out[9898];
     layer3_out[4199] <= layer2_out[10952];
     layer3_out[4200] <= ~layer2_out[5651];
     layer3_out[4201] <= ~layer2_out[10784] | layer2_out[10785];
     layer3_out[4202] <= ~layer2_out[6879] | layer2_out[6880];
     layer3_out[4203] <= ~layer2_out[10857] | layer2_out[10856];
     layer3_out[4204] <= layer2_out[2330] & ~layer2_out[2329];
     layer3_out[4205] <= ~layer2_out[1210];
     layer3_out[4206] <= ~layer2_out[10768] | layer2_out[10769];
     layer3_out[4207] <= ~layer2_out[7592] | layer2_out[7593];
     layer3_out[4208] <= ~layer2_out[2832];
     layer3_out[4209] <= ~layer2_out[1102];
     layer3_out[4210] <= ~(layer2_out[11377] ^ layer2_out[11378]);
     layer3_out[4211] <= layer2_out[6719];
     layer3_out[4212] <= ~layer2_out[11800] | layer2_out[11801];
     layer3_out[4213] <= layer2_out[4176] | layer2_out[4177];
     layer3_out[4214] <= layer2_out[4314];
     layer3_out[4215] <= ~layer2_out[5574] | layer2_out[5575];
     layer3_out[4216] <= ~layer2_out[9571];
     layer3_out[4217] <= ~layer2_out[403];
     layer3_out[4218] <= layer2_out[6763];
     layer3_out[4219] <= layer2_out[2230] ^ layer2_out[2231];
     layer3_out[4220] <= layer2_out[2453] | layer2_out[2454];
     layer3_out[4221] <= ~layer2_out[11014];
     layer3_out[4222] <= ~layer2_out[24];
     layer3_out[4223] <= layer2_out[9179] & ~layer2_out[9180];
     layer3_out[4224] <= ~(layer2_out[644] | layer2_out[645]);
     layer3_out[4225] <= layer2_out[606] & ~layer2_out[607];
     layer3_out[4226] <= layer2_out[3555] & ~layer2_out[3554];
     layer3_out[4227] <= ~(layer2_out[6012] | layer2_out[6013]);
     layer3_out[4228] <= ~(layer2_out[1758] | layer2_out[1759]);
     layer3_out[4229] <= layer2_out[585] & layer2_out[586];
     layer3_out[4230] <= layer2_out[9166] ^ layer2_out[9167];
     layer3_out[4231] <= ~layer2_out[462];
     layer3_out[4232] <= layer2_out[6993] & ~layer2_out[6992];
     layer3_out[4233] <= ~layer2_out[5950];
     layer3_out[4234] <= ~(layer2_out[11786] ^ layer2_out[11787]);
     layer3_out[4235] <= ~(layer2_out[2515] | layer2_out[2516]);
     layer3_out[4236] <= layer2_out[4258];
     layer3_out[4237] <= ~(layer2_out[3634] & layer2_out[3635]);
     layer3_out[4238] <= layer2_out[9577] & layer2_out[9578];
     layer3_out[4239] <= layer2_out[2781] ^ layer2_out[2782];
     layer3_out[4240] <= ~layer2_out[6890];
     layer3_out[4241] <= layer2_out[10243];
     layer3_out[4242] <= ~layer2_out[10728];
     layer3_out[4243] <= ~layer2_out[667] | layer2_out[668];
     layer3_out[4244] <= ~(layer2_out[2184] ^ layer2_out[2185]);
     layer3_out[4245] <= ~layer2_out[8907] | layer2_out[8906];
     layer3_out[4246] <= ~(layer2_out[4589] ^ layer2_out[4590]);
     layer3_out[4247] <= ~(layer2_out[2008] & layer2_out[2009]);
     layer3_out[4248] <= ~layer2_out[10502];
     layer3_out[4249] <= layer2_out[9081];
     layer3_out[4250] <= layer2_out[925] | layer2_out[926];
     layer3_out[4251] <= ~(layer2_out[3537] | layer2_out[3538]);
     layer3_out[4252] <= layer2_out[10106] & layer2_out[10107];
     layer3_out[4253] <= ~layer2_out[7978];
     layer3_out[4254] <= layer2_out[5837];
     layer3_out[4255] <= layer2_out[11153] & layer2_out[11154];
     layer3_out[4256] <= ~layer2_out[6743];
     layer3_out[4257] <= layer2_out[6853];
     layer3_out[4258] <= ~layer2_out[6478];
     layer3_out[4259] <= layer2_out[5246];
     layer3_out[4260] <= layer2_out[5699] ^ layer2_out[5700];
     layer3_out[4261] <= layer2_out[9265] & ~layer2_out[9264];
     layer3_out[4262] <= ~layer2_out[3919];
     layer3_out[4263] <= ~(layer2_out[6365] ^ layer2_out[6366]);
     layer3_out[4264] <= ~layer2_out[8989];
     layer3_out[4265] <= ~(layer2_out[5455] & layer2_out[5456]);
     layer3_out[4266] <= ~(layer2_out[5291] & layer2_out[5292]);
     layer3_out[4267] <= layer2_out[3077] | layer2_out[3078];
     layer3_out[4268] <= layer2_out[3459];
     layer3_out[4269] <= ~(layer2_out[5102] ^ layer2_out[5103]);
     layer3_out[4270] <= layer2_out[5022] ^ layer2_out[5023];
     layer3_out[4271] <= ~(layer2_out[8430] | layer2_out[8431]);
     layer3_out[4272] <= ~layer2_out[4347];
     layer3_out[4273] <= layer2_out[9415] & layer2_out[9416];
     layer3_out[4274] <= ~layer2_out[4351] | layer2_out[4352];
     layer3_out[4275] <= ~layer2_out[4601];
     layer3_out[4276] <= layer2_out[862] & ~layer2_out[863];
     layer3_out[4277] <= ~layer2_out[5781];
     layer3_out[4278] <= ~layer2_out[4334];
     layer3_out[4279] <= ~(layer2_out[8518] ^ layer2_out[8519]);
     layer3_out[4280] <= ~(layer2_out[9742] ^ layer2_out[9743]);
     layer3_out[4281] <= ~layer2_out[6411];
     layer3_out[4282] <= ~layer2_out[9612] | layer2_out[9613];
     layer3_out[4283] <= ~layer2_out[2581];
     layer3_out[4284] <= layer2_out[6706] & ~layer2_out[6707];
     layer3_out[4285] <= layer2_out[996] ^ layer2_out[997];
     layer3_out[4286] <= layer2_out[7339] & ~layer2_out[7340];
     layer3_out[4287] <= ~(layer2_out[11241] | layer2_out[11242]);
     layer3_out[4288] <= ~layer2_out[10457] | layer2_out[10458];
     layer3_out[4289] <= ~layer2_out[5335] | layer2_out[5336];
     layer3_out[4290] <= ~(layer2_out[10024] ^ layer2_out[10025]);
     layer3_out[4291] <= ~(layer2_out[872] ^ layer2_out[873]);
     layer3_out[4292] <= layer2_out[11541] ^ layer2_out[11542];
     layer3_out[4293] <= ~(layer2_out[9682] ^ layer2_out[9683]);
     layer3_out[4294] <= ~(layer2_out[569] & layer2_out[570]);
     layer3_out[4295] <= layer2_out[6948] ^ layer2_out[6949];
     layer3_out[4296] <= ~layer2_out[1739];
     layer3_out[4297] <= layer2_out[3637] & layer2_out[3638];
     layer3_out[4298] <= ~layer2_out[3320];
     layer3_out[4299] <= ~(layer2_out[3014] ^ layer2_out[3015]);
     layer3_out[4300] <= layer2_out[7829];
     layer3_out[4301] <= ~layer2_out[7130];
     layer3_out[4302] <= ~layer2_out[3999];
     layer3_out[4303] <= layer2_out[8546];
     layer3_out[4304] <= ~layer2_out[6958];
     layer3_out[4305] <= layer2_out[10758];
     layer3_out[4306] <= layer2_out[7348] ^ layer2_out[7349];
     layer3_out[4307] <= layer2_out[4211];
     layer3_out[4308] <= ~(layer2_out[2332] | layer2_out[2333]);
     layer3_out[4309] <= ~layer2_out[10548];
     layer3_out[4310] <= ~layer2_out[8742];
     layer3_out[4311] <= ~(layer2_out[7855] | layer2_out[7856]);
     layer3_out[4312] <= ~layer2_out[11190];
     layer3_out[4313] <= layer2_out[9649] & ~layer2_out[9650];
     layer3_out[4314] <= layer2_out[5003] | layer2_out[5004];
     layer3_out[4315] <= ~layer2_out[9812];
     layer3_out[4316] <= ~layer2_out[11124];
     layer3_out[4317] <= layer2_out[4922] & ~layer2_out[4923];
     layer3_out[4318] <= layer2_out[7374];
     layer3_out[4319] <= ~layer2_out[5980];
     layer3_out[4320] <= layer2_out[1336] | layer2_out[1337];
     layer3_out[4321] <= layer2_out[11712] ^ layer2_out[11713];
     layer3_out[4322] <= layer2_out[264];
     layer3_out[4323] <= layer2_out[3946];
     layer3_out[4324] <= layer2_out[10130] & ~layer2_out[10131];
     layer3_out[4325] <= ~(layer2_out[9540] ^ layer2_out[9541]);
     layer3_out[4326] <= ~(layer2_out[7490] & layer2_out[7491]);
     layer3_out[4327] <= layer2_out[985] ^ layer2_out[986];
     layer3_out[4328] <= layer2_out[10766];
     layer3_out[4329] <= layer2_out[2192];
     layer3_out[4330] <= ~layer2_out[7143];
     layer3_out[4331] <= layer2_out[8501] | layer2_out[8502];
     layer3_out[4332] <= ~layer2_out[5686] | layer2_out[5685];
     layer3_out[4333] <= layer2_out[2427] ^ layer2_out[2428];
     layer3_out[4334] <= ~(layer2_out[8776] & layer2_out[8777]);
     layer3_out[4335] <= ~(layer2_out[3471] | layer2_out[3472]);
     layer3_out[4336] <= ~layer2_out[9493];
     layer3_out[4337] <= layer2_out[1020] ^ layer2_out[1021];
     layer3_out[4338] <= layer2_out[6729] ^ layer2_out[6730];
     layer3_out[4339] <= layer2_out[11084];
     layer3_out[4340] <= layer2_out[5704] & layer2_out[5705];
     layer3_out[4341] <= layer2_out[1473] & ~layer2_out[1472];
     layer3_out[4342] <= ~(layer2_out[4288] | layer2_out[4289]);
     layer3_out[4343] <= ~layer2_out[7628];
     layer3_out[4344] <= ~(layer2_out[11249] ^ layer2_out[11250]);
     layer3_out[4345] <= ~layer2_out[7668];
     layer3_out[4346] <= ~(layer2_out[9312] | layer2_out[9313]);
     layer3_out[4347] <= ~layer2_out[2082];
     layer3_out[4348] <= layer2_out[8904];
     layer3_out[4349] <= ~(layer2_out[9909] | layer2_out[9910]);
     layer3_out[4350] <= ~layer2_out[10757];
     layer3_out[4351] <= layer2_out[5341];
     layer3_out[4352] <= ~layer2_out[6820];
     layer3_out[4353] <= ~layer2_out[314];
     layer3_out[4354] <= layer2_out[6855] ^ layer2_out[6856];
     layer3_out[4355] <= layer2_out[6721] ^ layer2_out[6722];
     layer3_out[4356] <= ~(layer2_out[3158] ^ layer2_out[3159]);
     layer3_out[4357] <= ~layer2_out[4982];
     layer3_out[4358] <= layer2_out[1024];
     layer3_out[4359] <= ~(layer2_out[9665] ^ layer2_out[9666]);
     layer3_out[4360] <= ~(layer2_out[10383] ^ layer2_out[10384]);
     layer3_out[4361] <= layer2_out[5228];
     layer3_out[4362] <= ~(layer2_out[9302] & layer2_out[9303]);
     layer3_out[4363] <= layer2_out[11256];
     layer3_out[4364] <= layer2_out[8136];
     layer3_out[4365] <= layer2_out[899];
     layer3_out[4366] <= layer2_out[379];
     layer3_out[4367] <= ~layer2_out[1390] | layer2_out[1391];
     layer3_out[4368] <= layer2_out[2540] & ~layer2_out[2541];
     layer3_out[4369] <= layer2_out[1549] ^ layer2_out[1550];
     layer3_out[4370] <= layer2_out[8663] ^ layer2_out[8664];
     layer3_out[4371] <= layer2_out[10759] ^ layer2_out[10760];
     layer3_out[4372] <= ~layer2_out[11022];
     layer3_out[4373] <= layer2_out[1691];
     layer3_out[4374] <= ~(layer2_out[4653] ^ layer2_out[4654]);
     layer3_out[4375] <= layer2_out[10941] & ~layer2_out[10940];
     layer3_out[4376] <= ~layer2_out[7618];
     layer3_out[4377] <= layer2_out[2525] | layer2_out[2526];
     layer3_out[4378] <= layer2_out[1397] ^ layer2_out[1398];
     layer3_out[4379] <= ~layer2_out[4608];
     layer3_out[4380] <= ~layer2_out[6379];
     layer3_out[4381] <= ~(layer2_out[2028] & layer2_out[2029]);
     layer3_out[4382] <= ~layer2_out[4108];
     layer3_out[4383] <= ~layer2_out[10541] | layer2_out[10540];
     layer3_out[4384] <= layer2_out[2248] & ~layer2_out[2247];
     layer3_out[4385] <= ~layer2_out[6781];
     layer3_out[4386] <= ~layer2_out[6218];
     layer3_out[4387] <= ~(layer2_out[6937] | layer2_out[6938]);
     layer3_out[4388] <= layer2_out[8768] | layer2_out[8769];
     layer3_out[4389] <= layer2_out[8324] & ~layer2_out[8325];
     layer3_out[4390] <= layer2_out[898];
     layer3_out[4391] <= layer2_out[5308] ^ layer2_out[5309];
     layer3_out[4392] <= ~layer2_out[4825];
     layer3_out[4393] <= ~layer2_out[6518] | layer2_out[6517];
     layer3_out[4394] <= ~layer2_out[9884];
     layer3_out[4395] <= layer2_out[4663] | layer2_out[4664];
     layer3_out[4396] <= layer2_out[10866] | layer2_out[10867];
     layer3_out[4397] <= ~(layer2_out[8863] ^ layer2_out[8864]);
     layer3_out[4398] <= ~(layer2_out[8001] ^ layer2_out[8002]);
     layer3_out[4399] <= layer2_out[5542] | layer2_out[5543];
     layer3_out[4400] <= ~layer2_out[10378];
     layer3_out[4401] <= ~layer2_out[8078];
     layer3_out[4402] <= ~layer2_out[4705] | layer2_out[4706];
     layer3_out[4403] <= layer2_out[10852];
     layer3_out[4404] <= layer2_out[10126];
     layer3_out[4405] <= ~layer2_out[7133];
     layer3_out[4406] <= ~layer2_out[4881];
     layer3_out[4407] <= ~(layer2_out[5872] ^ layer2_out[5873]);
     layer3_out[4408] <= layer2_out[4431];
     layer3_out[4409] <= ~layer2_out[7067];
     layer3_out[4410] <= ~layer2_out[1790];
     layer3_out[4411] <= layer2_out[6362] | layer2_out[6363];
     layer3_out[4412] <= ~layer2_out[2708];
     layer3_out[4413] <= layer2_out[4429];
     layer3_out[4414] <= ~(layer2_out[1526] ^ layer2_out[1527]);
     layer3_out[4415] <= layer2_out[6720] ^ layer2_out[6721];
     layer3_out[4416] <= layer2_out[7655];
     layer3_out[4417] <= ~layer2_out[6572] | layer2_out[6571];
     layer3_out[4418] <= layer2_out[7403] | layer2_out[7404];
     layer3_out[4419] <= ~(layer2_out[5008] ^ layer2_out[5009]);
     layer3_out[4420] <= ~layer2_out[6846] | layer2_out[6847];
     layer3_out[4421] <= ~(layer2_out[11291] | layer2_out[11292]);
     layer3_out[4422] <= layer2_out[2611] & ~layer2_out[2612];
     layer3_out[4423] <= ~layer2_out[5321];
     layer3_out[4424] <= layer2_out[5637] | layer2_out[5638];
     layer3_out[4425] <= ~(layer2_out[7727] ^ layer2_out[7728]);
     layer3_out[4426] <= ~layer2_out[6351];
     layer3_out[4427] <= ~layer2_out[9065] | layer2_out[9066];
     layer3_out[4428] <= layer2_out[7714] ^ layer2_out[7715];
     layer3_out[4429] <= layer2_out[3631] & ~layer2_out[3630];
     layer3_out[4430] <= layer2_out[5829] & ~layer2_out[5830];
     layer3_out[4431] <= ~(layer2_out[8364] ^ layer2_out[8365]);
     layer3_out[4432] <= ~layer2_out[1402];
     layer3_out[4433] <= layer2_out[9103];
     layer3_out[4434] <= layer2_out[6349];
     layer3_out[4435] <= ~layer2_out[411];
     layer3_out[4436] <= ~(layer2_out[3276] ^ layer2_out[3277]);
     layer3_out[4437] <= ~(layer2_out[6584] ^ layer2_out[6585]);
     layer3_out[4438] <= ~layer2_out[9787];
     layer3_out[4439] <= ~layer2_out[951];
     layer3_out[4440] <= ~layer2_out[10233] | layer2_out[10234];
     layer3_out[4441] <= layer2_out[601] ^ layer2_out[602];
     layer3_out[4442] <= ~layer2_out[1021];
     layer3_out[4443] <= layer2_out[2660] & ~layer2_out[2659];
     layer3_out[4444] <= layer2_out[2486] ^ layer2_out[2487];
     layer3_out[4445] <= ~layer2_out[10579];
     layer3_out[4446] <= ~layer2_out[6294] | layer2_out[6293];
     layer3_out[4447] <= layer2_out[9523];
     layer3_out[4448] <= ~(layer2_out[8114] ^ layer2_out[8115]);
     layer3_out[4449] <= layer2_out[10610];
     layer3_out[4450] <= layer2_out[8845];
     layer3_out[4451] <= layer2_out[7201] ^ layer2_out[7202];
     layer3_out[4452] <= layer2_out[11572] & ~layer2_out[11573];
     layer3_out[4453] <= ~layer2_out[2901];
     layer3_out[4454] <= layer2_out[4] & layer2_out[5];
     layer3_out[4455] <= ~layer2_out[4122] | layer2_out[4123];
     layer3_out[4456] <= layer2_out[4849] ^ layer2_out[4850];
     layer3_out[4457] <= layer2_out[3385] & layer2_out[3386];
     layer3_out[4458] <= layer2_out[9409] & layer2_out[9410];
     layer3_out[4459] <= ~layer2_out[11539];
     layer3_out[4460] <= ~(layer2_out[4946] & layer2_out[4947]);
     layer3_out[4461] <= ~(layer2_out[6410] | layer2_out[6411]);
     layer3_out[4462] <= layer2_out[10223] & ~layer2_out[10222];
     layer3_out[4463] <= ~(layer2_out[1471] ^ layer2_out[1472]);
     layer3_out[4464] <= ~(layer2_out[3673] & layer2_out[3674]);
     layer3_out[4465] <= layer2_out[6115] & ~layer2_out[6116];
     layer3_out[4466] <= ~layer2_out[5412];
     layer3_out[4467] <= ~(layer2_out[178] ^ layer2_out[179]);
     layer3_out[4468] <= ~layer2_out[8596] | layer2_out[8595];
     layer3_out[4469] <= layer2_out[10303] & ~layer2_out[10304];
     layer3_out[4470] <= ~layer2_out[7577];
     layer3_out[4471] <= ~layer2_out[11020];
     layer3_out[4472] <= ~(layer2_out[10628] ^ layer2_out[10629]);
     layer3_out[4473] <= ~(layer2_out[10801] ^ layer2_out[10802]);
     layer3_out[4474] <= layer2_out[6088] & ~layer2_out[6089];
     layer3_out[4475] <= layer2_out[9144] & ~layer2_out[9143];
     layer3_out[4476] <= layer2_out[7741] ^ layer2_out[7742];
     layer3_out[4477] <= layer2_out[11141];
     layer3_out[4478] <= layer2_out[3891];
     layer3_out[4479] <= layer2_out[2996] ^ layer2_out[2997];
     layer3_out[4480] <= layer2_out[6738] & ~layer2_out[6739];
     layer3_out[4481] <= layer2_out[3601] ^ layer2_out[3602];
     layer3_out[4482] <= layer2_out[6006];
     layer3_out[4483] <= layer2_out[10390] ^ layer2_out[10391];
     layer3_out[4484] <= layer2_out[1479];
     layer3_out[4485] <= ~layer2_out[1208];
     layer3_out[4486] <= layer2_out[1709];
     layer3_out[4487] <= layer2_out[6807];
     layer3_out[4488] <= ~layer2_out[1654];
     layer3_out[4489] <= layer2_out[6434] ^ layer2_out[6435];
     layer3_out[4490] <= layer2_out[11462];
     layer3_out[4491] <= ~layer2_out[1075] | layer2_out[1074];
     layer3_out[4492] <= ~layer2_out[7379];
     layer3_out[4493] <= ~layer2_out[5001] | layer2_out[5002];
     layer3_out[4494] <= ~layer2_out[3075];
     layer3_out[4495] <= ~(layer2_out[9376] & layer2_out[9377]);
     layer3_out[4496] <= ~layer2_out[7492];
     layer3_out[4497] <= ~layer2_out[3929] | layer2_out[3930];
     layer3_out[4498] <= layer2_out[8888];
     layer3_out[4499] <= ~layer2_out[5345];
     layer3_out[4500] <= layer2_out[1381];
     layer3_out[4501] <= ~layer2_out[8567];
     layer3_out[4502] <= layer2_out[8852];
     layer3_out[4503] <= ~(layer2_out[4113] & layer2_out[4114]);
     layer3_out[4504] <= layer2_out[5798] | layer2_out[5799];
     layer3_out[4505] <= layer2_out[1979] ^ layer2_out[1980];
     layer3_out[4506] <= ~layer2_out[8857];
     layer3_out[4507] <= ~(layer2_out[6261] ^ layer2_out[6262]);
     layer3_out[4508] <= ~(layer2_out[6150] & layer2_out[6151]);
     layer3_out[4509] <= layer2_out[2620] & ~layer2_out[2621];
     layer3_out[4510] <= layer2_out[8609];
     layer3_out[4511] <= layer2_out[9339] | layer2_out[9340];
     layer3_out[4512] <= ~layer2_out[10254];
     layer3_out[4513] <= layer2_out[2692] ^ layer2_out[2693];
     layer3_out[4514] <= ~layer2_out[9895];
     layer3_out[4515] <= layer2_out[6635] & layer2_out[6636];
     layer3_out[4516] <= layer2_out[454];
     layer3_out[4517] <= ~(layer2_out[6863] | layer2_out[6864]);
     layer3_out[4518] <= ~(layer2_out[9954] ^ layer2_out[9955]);
     layer3_out[4519] <= ~layer2_out[3954];
     layer3_out[4520] <= ~(layer2_out[10144] ^ layer2_out[10145]);
     layer3_out[4521] <= ~layer2_out[7364] | layer2_out[7363];
     layer3_out[4522] <= layer2_out[7469] & layer2_out[7470];
     layer3_out[4523] <= ~layer2_out[7390];
     layer3_out[4524] <= ~layer2_out[2028];
     layer3_out[4525] <= ~layer2_out[2506];
     layer3_out[4526] <= ~layer2_out[9252];
     layer3_out[4527] <= ~layer2_out[1671] | layer2_out[1670];
     layer3_out[4528] <= layer2_out[130] | layer2_out[131];
     layer3_out[4529] <= ~layer2_out[6287];
     layer3_out[4530] <= layer2_out[3494] & ~layer2_out[3495];
     layer3_out[4531] <= ~layer2_out[10988];
     layer3_out[4532] <= layer2_out[1068];
     layer3_out[4533] <= ~layer2_out[11453] | layer2_out[11454];
     layer3_out[4534] <= layer2_out[5029] & layer2_out[5030];
     layer3_out[4535] <= ~layer2_out[1995] | layer2_out[1996];
     layer3_out[4536] <= layer2_out[5473] & ~layer2_out[5472];
     layer3_out[4537] <= layer2_out[1111];
     layer3_out[4538] <= layer2_out[3219] ^ layer2_out[3220];
     layer3_out[4539] <= ~(layer2_out[4345] | layer2_out[4346]);
     layer3_out[4540] <= ~(layer2_out[167] & layer2_out[168]);
     layer3_out[4541] <= ~layer2_out[11769];
     layer3_out[4542] <= layer2_out[7137] & ~layer2_out[7136];
     layer3_out[4543] <= ~(layer2_out[2711] ^ layer2_out[2712]);
     layer3_out[4544] <= ~layer2_out[8078];
     layer3_out[4545] <= ~layer2_out[2485] | layer2_out[2486];
     layer3_out[4546] <= layer2_out[3352] ^ layer2_out[3353];
     layer3_out[4547] <= layer2_out[4020] ^ layer2_out[4021];
     layer3_out[4548] <= ~layer2_out[1015];
     layer3_out[4549] <= ~(layer2_out[7587] | layer2_out[7588]);
     layer3_out[4550] <= ~layer2_out[2872] | layer2_out[2871];
     layer3_out[4551] <= layer2_out[3289] & ~layer2_out[3288];
     layer3_out[4552] <= ~layer2_out[4825];
     layer3_out[4553] <= layer2_out[4490];
     layer3_out[4554] <= layer2_out[8376] ^ layer2_out[8377];
     layer3_out[4555] <= ~layer2_out[9045];
     layer3_out[4556] <= ~(layer2_out[147] ^ layer2_out[148]);
     layer3_out[4557] <= layer2_out[7548] ^ layer2_out[7549];
     layer3_out[4558] <= layer2_out[3105] | layer2_out[3106];
     layer3_out[4559] <= layer2_out[2357];
     layer3_out[4560] <= ~(layer2_out[4781] | layer2_out[4782]);
     layer3_out[4561] <= layer2_out[641] & ~layer2_out[642];
     layer3_out[4562] <= ~(layer2_out[4049] | layer2_out[4050]);
     layer3_out[4563] <= layer2_out[6619] ^ layer2_out[6620];
     layer3_out[4564] <= layer2_out[2297] | layer2_out[2298];
     layer3_out[4565] <= ~layer2_out[1660];
     layer3_out[4566] <= ~layer2_out[5562];
     layer3_out[4567] <= ~layer2_out[1640];
     layer3_out[4568] <= layer2_out[585] & ~layer2_out[584];
     layer3_out[4569] <= ~layer2_out[9502];
     layer3_out[4570] <= layer2_out[10041] & ~layer2_out[10042];
     layer3_out[4571] <= ~layer2_out[7949] | layer2_out[7950];
     layer3_out[4572] <= ~layer2_out[8724] | layer2_out[8725];
     layer3_out[4573] <= layer2_out[5883];
     layer3_out[4574] <= ~layer2_out[679] | layer2_out[678];
     layer3_out[4575] <= ~layer2_out[455] | layer2_out[454];
     layer3_out[4576] <= ~(layer2_out[1793] | layer2_out[1794]);
     layer3_out[4577] <= layer2_out[9054] | layer2_out[9055];
     layer3_out[4578] <= layer2_out[10443];
     layer3_out[4579] <= layer2_out[6948];
     layer3_out[4580] <= layer2_out[9842];
     layer3_out[4581] <= layer2_out[1320] & ~layer2_out[1319];
     layer3_out[4582] <= ~layer2_out[4777];
     layer3_out[4583] <= layer2_out[10410] | layer2_out[10411];
     layer3_out[4584] <= layer2_out[2030] ^ layer2_out[2031];
     layer3_out[4585] <= layer2_out[2548];
     layer3_out[4586] <= layer2_out[3817] & ~layer2_out[3816];
     layer3_out[4587] <= layer2_out[3712];
     layer3_out[4588] <= ~layer2_out[213];
     layer3_out[4589] <= ~(layer2_out[11863] | layer2_out[11864]);
     layer3_out[4590] <= ~layer2_out[5509];
     layer3_out[4591] <= ~layer2_out[11645];
     layer3_out[4592] <= ~layer2_out[11528] | layer2_out[11527];
     layer3_out[4593] <= layer2_out[7574];
     layer3_out[4594] <= ~layer2_out[5001];
     layer3_out[4595] <= ~layer2_out[1753];
     layer3_out[4596] <= ~(layer2_out[6238] ^ layer2_out[6239]);
     layer3_out[4597] <= layer2_out[8705] ^ layer2_out[8706];
     layer3_out[4598] <= ~layer2_out[8624];
     layer3_out[4599] <= ~(layer2_out[809] | layer2_out[810]);
     layer3_out[4600] <= layer2_out[11349];
     layer3_out[4601] <= ~(layer2_out[643] | layer2_out[644]);
     layer3_out[4602] <= ~layer2_out[6206];
     layer3_out[4603] <= ~layer2_out[10998] | layer2_out[10999];
     layer3_out[4604] <= ~(layer2_out[11128] ^ layer2_out[11129]);
     layer3_out[4605] <= layer2_out[5589] ^ layer2_out[5590];
     layer3_out[4606] <= layer2_out[172] ^ layer2_out[173];
     layer3_out[4607] <= ~layer2_out[1688];
     layer3_out[4608] <= ~layer2_out[1799] | layer2_out[1798];
     layer3_out[4609] <= ~(layer2_out[1076] & layer2_out[1077]);
     layer3_out[4610] <= layer2_out[5603] & ~layer2_out[5604];
     layer3_out[4611] <= layer2_out[4325] ^ layer2_out[4326];
     layer3_out[4612] <= layer2_out[10255] & layer2_out[10256];
     layer3_out[4613] <= ~layer2_out[9335];
     layer3_out[4614] <= layer2_out[6524];
     layer3_out[4615] <= ~(layer2_out[794] ^ layer2_out[795]);
     layer3_out[4616] <= ~layer2_out[3042];
     layer3_out[4617] <= layer2_out[10879] & ~layer2_out[10878];
     layer3_out[4618] <= ~layer2_out[7143];
     layer3_out[4619] <= ~(layer2_out[8090] | layer2_out[8091]);
     layer3_out[4620] <= layer2_out[5883];
     layer3_out[4621] <= ~(layer2_out[1844] | layer2_out[1845]);
     layer3_out[4622] <= ~layer2_out[2134];
     layer3_out[4623] <= ~layer2_out[9479];
     layer3_out[4624] <= layer2_out[1434];
     layer3_out[4625] <= ~(layer2_out[7542] & layer2_out[7543]);
     layer3_out[4626] <= ~(layer2_out[2066] | layer2_out[2067]);
     layer3_out[4627] <= ~layer2_out[10980];
     layer3_out[4628] <= ~layer2_out[9214] | layer2_out[9215];
     layer3_out[4629] <= layer2_out[10316] ^ layer2_out[10317];
     layer3_out[4630] <= layer2_out[4133];
     layer3_out[4631] <= layer2_out[9588] ^ layer2_out[9589];
     layer3_out[4632] <= ~(layer2_out[8943] & layer2_out[8944]);
     layer3_out[4633] <= layer2_out[9874] & ~layer2_out[9873];
     layer3_out[4634] <= ~layer2_out[8376] | layer2_out[8375];
     layer3_out[4635] <= layer2_out[3039];
     layer3_out[4636] <= ~layer2_out[10663];
     layer3_out[4637] <= layer2_out[7274] ^ layer2_out[7275];
     layer3_out[4638] <= layer2_out[9835];
     layer3_out[4639] <= ~layer2_out[8325];
     layer3_out[4640] <= ~(layer2_out[11772] ^ layer2_out[11773]);
     layer3_out[4641] <= layer2_out[5905] & layer2_out[5906];
     layer3_out[4642] <= ~layer2_out[4289];
     layer3_out[4643] <= ~(layer2_out[11247] | layer2_out[11248]);
     layer3_out[4644] <= layer2_out[4955] & layer2_out[4956];
     layer3_out[4645] <= layer2_out[4754];
     layer3_out[4646] <= layer2_out[10622] & layer2_out[10623];
     layer3_out[4647] <= layer2_out[9354] & ~layer2_out[9353];
     layer3_out[4648] <= ~layer2_out[912];
     layer3_out[4649] <= ~layer2_out[2661];
     layer3_out[4650] <= ~(layer2_out[6732] | layer2_out[6733]);
     layer3_out[4651] <= ~layer2_out[9248];
     layer3_out[4652] <= ~layer2_out[9087];
     layer3_out[4653] <= layer2_out[9793];
     layer3_out[4654] <= layer2_out[3707] ^ layer2_out[3708];
     layer3_out[4655] <= layer2_out[3849];
     layer3_out[4656] <= layer2_out[11069] | layer2_out[11070];
     layer3_out[4657] <= layer2_out[9237];
     layer3_out[4658] <= ~(layer2_out[9089] ^ layer2_out[9090]);
     layer3_out[4659] <= layer2_out[8774] & ~layer2_out[8775];
     layer3_out[4660] <= ~(layer2_out[8805] ^ layer2_out[8806]);
     layer3_out[4661] <= ~(layer2_out[10398] ^ layer2_out[10399]);
     layer3_out[4662] <= ~(layer2_out[9196] | layer2_out[9197]);
     layer3_out[4663] <= layer2_out[5804] & ~layer2_out[5805];
     layer3_out[4664] <= ~(layer2_out[11400] ^ layer2_out[11401]);
     layer3_out[4665] <= ~layer2_out[5773];
     layer3_out[4666] <= layer2_out[6054];
     layer3_out[4667] <= layer2_out[464] ^ layer2_out[465];
     layer3_out[4668] <= layer2_out[1538] ^ layer2_out[1539];
     layer3_out[4669] <= ~(layer2_out[7265] ^ layer2_out[7266]);
     layer3_out[4670] <= ~(layer2_out[710] ^ layer2_out[711]);
     layer3_out[4671] <= layer2_out[11220];
     layer3_out[4672] <= ~layer2_out[7268] | layer2_out[7267];
     layer3_out[4673] <= ~(layer2_out[10652] ^ layer2_out[10653]);
     layer3_out[4674] <= layer2_out[632];
     layer3_out[4675] <= ~layer2_out[10737];
     layer3_out[4676] <= layer2_out[4810];
     layer3_out[4677] <= ~(layer2_out[9483] | layer2_out[9484]);
     layer3_out[4678] <= layer2_out[2524] & layer2_out[2525];
     layer3_out[4679] <= layer2_out[2158];
     layer3_out[4680] <= ~layer2_out[2612] | layer2_out[2613];
     layer3_out[4681] <= ~layer2_out[1559] | layer2_out[1560];
     layer3_out[4682] <= ~layer2_out[9436];
     layer3_out[4683] <= layer2_out[7271];
     layer3_out[4684] <= layer2_out[10401];
     layer3_out[4685] <= layer2_out[5359] & layer2_out[5360];
     layer3_out[4686] <= ~layer2_out[857] | layer2_out[856];
     layer3_out[4687] <= layer2_out[1575] | layer2_out[1576];
     layer3_out[4688] <= layer2_out[11386] | layer2_out[11387];
     layer3_out[4689] <= ~layer2_out[2784];
     layer3_out[4690] <= ~layer2_out[11370] | layer2_out[11369];
     layer3_out[4691] <= ~(layer2_out[7002] ^ layer2_out[7003]);
     layer3_out[4692] <= layer2_out[166] & ~layer2_out[167];
     layer3_out[4693] <= ~(layer2_out[871] | layer2_out[872]);
     layer3_out[4694] <= layer2_out[653];
     layer3_out[4695] <= ~layer2_out[11244];
     layer3_out[4696] <= layer2_out[2875];
     layer3_out[4697] <= ~layer2_out[1147] | layer2_out[1146];
     layer3_out[4698] <= ~layer2_out[4048];
     layer3_out[4699] <= layer2_out[4409];
     layer3_out[4700] <= layer2_out[5867];
     layer3_out[4701] <= ~(layer2_out[4988] ^ layer2_out[4989]);
     layer3_out[4702] <= layer2_out[1447] ^ layer2_out[1448];
     layer3_out[4703] <= layer2_out[10172] ^ layer2_out[10173];
     layer3_out[4704] <= layer2_out[4805] | layer2_out[4806];
     layer3_out[4705] <= ~layer2_out[2731];
     layer3_out[4706] <= ~layer2_out[5514] | layer2_out[5515];
     layer3_out[4707] <= layer2_out[4863] | layer2_out[4864];
     layer3_out[4708] <= layer2_out[7682] ^ layer2_out[7683];
     layer3_out[4709] <= ~layer2_out[11117];
     layer3_out[4710] <= layer2_out[2801];
     layer3_out[4711] <= layer2_out[8113] & ~layer2_out[8112];
     layer3_out[4712] <= layer2_out[48] & ~layer2_out[47];
     layer3_out[4713] <= layer2_out[4531];
     layer3_out[4714] <= layer2_out[9957];
     layer3_out[4715] <= ~(layer2_out[3703] | layer2_out[3704]);
     layer3_out[4716] <= ~layer2_out[7732];
     layer3_out[4717] <= layer2_out[2917];
     layer3_out[4718] <= ~layer2_out[8313] | layer2_out[8312];
     layer3_out[4719] <= ~(layer2_out[7644] & layer2_out[7645]);
     layer3_out[4720] <= ~(layer2_out[10302] ^ layer2_out[10303]);
     layer3_out[4721] <= layer2_out[4206];
     layer3_out[4722] <= ~layer2_out[3388];
     layer3_out[4723] <= layer2_out[3859] | layer2_out[3860];
     layer3_out[4724] <= ~layer2_out[6850];
     layer3_out[4725] <= layer2_out[6376];
     layer3_out[4726] <= ~layer2_out[4505] | layer2_out[4506];
     layer3_out[4727] <= layer2_out[10007] & layer2_out[10008];
     layer3_out[4728] <= ~(layer2_out[146] ^ layer2_out[147]);
     layer3_out[4729] <= layer2_out[11044] ^ layer2_out[11045];
     layer3_out[4730] <= layer2_out[274] & ~layer2_out[275];
     layer3_out[4731] <= ~(layer2_out[7396] & layer2_out[7397]);
     layer3_out[4732] <= ~layer2_out[4229];
     layer3_out[4733] <= layer2_out[1383] & ~layer2_out[1384];
     layer3_out[4734] <= layer2_out[11627];
     layer3_out[4735] <= layer2_out[9160] & ~layer2_out[9161];
     layer3_out[4736] <= ~layer2_out[11641] | layer2_out[11642];
     layer3_out[4737] <= ~layer2_out[10363] | layer2_out[10362];
     layer3_out[4738] <= layer2_out[1540] & ~layer2_out[1541];
     layer3_out[4739] <= ~layer2_out[3902] | layer2_out[3903];
     layer3_out[4740] <= ~(layer2_out[9002] ^ layer2_out[9003]);
     layer3_out[4741] <= layer2_out[10963] | layer2_out[10964];
     layer3_out[4742] <= layer2_out[8523] & ~layer2_out[8524];
     layer3_out[4743] <= layer2_out[11127];
     layer3_out[4744] <= ~layer2_out[6790];
     layer3_out[4745] <= layer2_out[11359] ^ layer2_out[11360];
     layer3_out[4746] <= layer2_out[586] | layer2_out[587];
     layer3_out[4747] <= ~(layer2_out[2112] & layer2_out[2113]);
     layer3_out[4748] <= layer2_out[3406] | layer2_out[3407];
     layer3_out[4749] <= ~(layer2_out[10598] ^ layer2_out[10599]);
     layer3_out[4750] <= layer2_out[6666];
     layer3_out[4751] <= layer2_out[1888];
     layer3_out[4752] <= layer2_out[2172];
     layer3_out[4753] <= layer2_out[4900];
     layer3_out[4754] <= ~layer2_out[8520] | layer2_out[8519];
     layer3_out[4755] <= layer2_out[6281];
     layer3_out[4756] <= layer2_out[11948] ^ layer2_out[11949];
     layer3_out[4757] <= ~(layer2_out[2916] ^ layer2_out[2917]);
     layer3_out[4758] <= ~layer2_out[9443] | layer2_out[9442];
     layer3_out[4759] <= layer2_out[8674] | layer2_out[8675];
     layer3_out[4760] <= ~(layer2_out[740] | layer2_out[741]);
     layer3_out[4761] <= ~layer2_out[1263];
     layer3_out[4762] <= ~layer2_out[8603];
     layer3_out[4763] <= ~layer2_out[9907] | layer2_out[9906];
     layer3_out[4764] <= ~layer2_out[5499];
     layer3_out[4765] <= ~(layer2_out[6731] ^ layer2_out[6732]);
     layer3_out[4766] <= layer2_out[6396];
     layer3_out[4767] <= ~(layer2_out[1600] ^ layer2_out[1601]);
     layer3_out[4768] <= layer2_out[2870];
     layer3_out[4769] <= layer2_out[9832] & layer2_out[9833];
     layer3_out[4770] <= ~layer2_out[3108];
     layer3_out[4771] <= layer2_out[1403] | layer2_out[1404];
     layer3_out[4772] <= layer2_out[8060];
     layer3_out[4773] <= layer2_out[7638] & ~layer2_out[7639];
     layer3_out[4774] <= ~layer2_out[752] | layer2_out[753];
     layer3_out[4775] <= layer2_out[9007];
     layer3_out[4776] <= ~layer2_out[803];
     layer3_out[4777] <= ~layer2_out[258];
     layer3_out[4778] <= layer2_out[2344] & ~layer2_out[2345];
     layer3_out[4779] <= layer2_out[4744];
     layer3_out[4780] <= ~(layer2_out[5382] ^ layer2_out[5383]);
     layer3_out[4781] <= ~layer2_out[7486];
     layer3_out[4782] <= ~(layer2_out[2130] ^ layer2_out[2131]);
     layer3_out[4783] <= layer2_out[1886] & layer2_out[1887];
     layer3_out[4784] <= ~layer2_out[4634];
     layer3_out[4785] <= ~layer2_out[4245] | layer2_out[4246];
     layer3_out[4786] <= layer2_out[9671] & layer2_out[9672];
     layer3_out[4787] <= ~(layer2_out[6214] ^ layer2_out[6215]);
     layer3_out[4788] <= layer2_out[2301] | layer2_out[2302];
     layer3_out[4789] <= layer2_out[10123] & ~layer2_out[10124];
     layer3_out[4790] <= ~(layer2_out[8984] ^ layer2_out[8985]);
     layer3_out[4791] <= layer2_out[3861];
     layer3_out[4792] <= layer2_out[2959];
     layer3_out[4793] <= layer2_out[3060] & layer2_out[3061];
     layer3_out[4794] <= ~(layer2_out[8417] ^ layer2_out[8418]);
     layer3_out[4795] <= ~layer2_out[2677];
     layer3_out[4796] <= ~layer2_out[7371];
     layer3_out[4797] <= ~(layer2_out[5795] & layer2_out[5796]);
     layer3_out[4798] <= layer2_out[3900] ^ layer2_out[3901];
     layer3_out[4799] <= ~layer2_out[10485];
     layer3_out[4800] <= ~layer2_out[11370] | layer2_out[11371];
     layer3_out[4801] <= layer2_out[4156] ^ layer2_out[4157];
     layer3_out[4802] <= ~layer2_out[7117];
     layer3_out[4803] <= ~(layer2_out[9659] ^ layer2_out[9660]);
     layer3_out[4804] <= ~(layer2_out[6573] & layer2_out[6574]);
     layer3_out[4805] <= layer2_out[6348] ^ layer2_out[6349];
     layer3_out[4806] <= ~(layer2_out[64] ^ layer2_out[65]);
     layer3_out[4807] <= layer2_out[7382];
     layer3_out[4808] <= layer2_out[11089] & layer2_out[11090];
     layer3_out[4809] <= layer2_out[1274] ^ layer2_out[1275];
     layer3_out[4810] <= layer2_out[10519] ^ layer2_out[10520];
     layer3_out[4811] <= layer2_out[9437];
     layer3_out[4812] <= layer2_out[7200] & layer2_out[7201];
     layer3_out[4813] <= layer2_out[9838];
     layer3_out[4814] <= layer2_out[3849] & ~layer2_out[3850];
     layer3_out[4815] <= layer2_out[2962] & layer2_out[2963];
     layer3_out[4816] <= layer2_out[2482] & ~layer2_out[2483];
     layer3_out[4817] <= layer2_out[7014] & ~layer2_out[7015];
     layer3_out[4818] <= ~(layer2_out[6710] ^ layer2_out[6711]);
     layer3_out[4819] <= layer2_out[7563] & layer2_out[7564];
     layer3_out[4820] <= layer2_out[8577];
     layer3_out[4821] <= ~(layer2_out[2050] | layer2_out[2051]);
     layer3_out[4822] <= layer2_out[2352] | layer2_out[2353];
     layer3_out[4823] <= layer2_out[2681];
     layer3_out[4824] <= ~(layer2_out[973] & layer2_out[974]);
     layer3_out[4825] <= layer2_out[11376];
     layer3_out[4826] <= layer2_out[2549] & ~layer2_out[2550];
     layer3_out[4827] <= ~(layer2_out[676] ^ layer2_out[677]);
     layer3_out[4828] <= layer2_out[2143];
     layer3_out[4829] <= ~layer2_out[1638];
     layer3_out[4830] <= ~(layer2_out[6979] ^ layer2_out[6980]);
     layer3_out[4831] <= ~(layer2_out[8761] ^ layer2_out[8762]);
     layer3_out[4832] <= layer2_out[6383] ^ layer2_out[6384];
     layer3_out[4833] <= ~(layer2_out[9327] | layer2_out[9328]);
     layer3_out[4834] <= layer2_out[4470] & layer2_out[4471];
     layer3_out[4835] <= layer2_out[3169] & ~layer2_out[3170];
     layer3_out[4836] <= layer2_out[10567] & ~layer2_out[10568];
     layer3_out[4837] <= ~layer2_out[7344] | layer2_out[7343];
     layer3_out[4838] <= ~layer2_out[8669] | layer2_out[8668];
     layer3_out[4839] <= ~layer2_out[11867];
     layer3_out[4840] <= layer2_out[2004] | layer2_out[2005];
     layer3_out[4841] <= ~(layer2_out[10568] | layer2_out[10569]);
     layer3_out[4842] <= ~layer2_out[975];
     layer3_out[4843] <= layer2_out[6936] & ~layer2_out[6935];
     layer3_out[4844] <= ~(layer2_out[2690] ^ layer2_out[2691]);
     layer3_out[4845] <= layer2_out[2693] ^ layer2_out[2694];
     layer3_out[4846] <= layer2_out[8946];
     layer3_out[4847] <= ~layer2_out[10200];
     layer3_out[4848] <= ~(layer2_out[2089] | layer2_out[2090]);
     layer3_out[4849] <= ~(layer2_out[8422] ^ layer2_out[8423]);
     layer3_out[4850] <= ~(layer2_out[8736] & layer2_out[8737]);
     layer3_out[4851] <= ~(layer2_out[2816] ^ layer2_out[2817]);
     layer3_out[4852] <= ~layer2_out[10050];
     layer3_out[4853] <= ~(layer2_out[9623] | layer2_out[9624]);
     layer3_out[4854] <= layer2_out[5138];
     layer3_out[4855] <= ~(layer2_out[10301] ^ layer2_out[10302]);
     layer3_out[4856] <= ~layer2_out[847];
     layer3_out[4857] <= layer2_out[10900] & ~layer2_out[10901];
     layer3_out[4858] <= layer2_out[3978] & ~layer2_out[3979];
     layer3_out[4859] <= layer2_out[2165] & layer2_out[2166];
     layer3_out[4860] <= ~(layer2_out[5946] | layer2_out[5947]);
     layer3_out[4861] <= layer2_out[10997] & layer2_out[10998];
     layer3_out[4862] <= ~layer2_out[6785];
     layer3_out[4863] <= layer2_out[50] & layer2_out[51];
     layer3_out[4864] <= layer2_out[6207] & ~layer2_out[6208];
     layer3_out[4865] <= ~(layer2_out[6109] | layer2_out[6110]);
     layer3_out[4866] <= ~(layer2_out[10387] ^ layer2_out[10388]);
     layer3_out[4867] <= layer2_out[741] | layer2_out[742];
     layer3_out[4868] <= layer2_out[5600] & layer2_out[5601];
     layer3_out[4869] <= layer2_out[7709] & ~layer2_out[7710];
     layer3_out[4870] <= layer2_out[5033] & layer2_out[5034];
     layer3_out[4871] <= layer2_out[5056];
     layer3_out[4872] <= ~layer2_out[1002];
     layer3_out[4873] <= ~(layer2_out[10859] ^ layer2_out[10860]);
     layer3_out[4874] <= ~(layer2_out[8361] ^ layer2_out[8362]);
     layer3_out[4875] <= layer2_out[3767] & layer2_out[3768];
     layer3_out[4876] <= layer2_out[1599] & ~layer2_out[1600];
     layer3_out[4877] <= ~layer2_out[10231];
     layer3_out[4878] <= ~layer2_out[7607];
     layer3_out[4879] <= ~layer2_out[10543] | layer2_out[10544];
     layer3_out[4880] <= layer2_out[267] & ~layer2_out[266];
     layer3_out[4881] <= layer2_out[10685] & ~layer2_out[10686];
     layer3_out[4882] <= ~layer2_out[529];
     layer3_out[4883] <= ~layer2_out[7508];
     layer3_out[4884] <= layer2_out[7207] & layer2_out[7208];
     layer3_out[4885] <= layer2_out[640];
     layer3_out[4886] <= layer2_out[5792] & ~layer2_out[5793];
     layer3_out[4887] <= layer2_out[1086];
     layer3_out[4888] <= layer2_out[7220] & ~layer2_out[7221];
     layer3_out[4889] <= ~layer2_out[4305];
     layer3_out[4890] <= layer2_out[5585];
     layer3_out[4891] <= ~(layer2_out[11696] ^ layer2_out[11697]);
     layer3_out[4892] <= ~(layer2_out[948] | layer2_out[949]);
     layer3_out[4893] <= layer2_out[11417] & ~layer2_out[11418];
     layer3_out[4894] <= layer2_out[7285];
     layer3_out[4895] <= ~layer2_out[963];
     layer3_out[4896] <= layer2_out[3899];
     layer3_out[4897] <= layer2_out[8979] & ~layer2_out[8978];
     layer3_out[4898] <= ~(layer2_out[10308] | layer2_out[10309]);
     layer3_out[4899] <= ~(layer2_out[5103] ^ layer2_out[5104]);
     layer3_out[4900] <= layer2_out[7678] & layer2_out[7679];
     layer3_out[4901] <= ~(layer2_out[10431] | layer2_out[10432]);
     layer3_out[4902] <= layer2_out[1538] & ~layer2_out[1537];
     layer3_out[4903] <= ~layer2_out[6064];
     layer3_out[4904] <= layer2_out[3747] ^ layer2_out[3748];
     layer3_out[4905] <= layer2_out[9171] & layer2_out[9172];
     layer3_out[4906] <= layer2_out[3691];
     layer3_out[4907] <= layer2_out[620] ^ layer2_out[621];
     layer3_out[4908] <= layer2_out[7851] & ~layer2_out[7850];
     layer3_out[4909] <= layer2_out[3263];
     layer3_out[4910] <= ~(layer2_out[757] | layer2_out[758]);
     layer3_out[4911] <= ~layer2_out[11527];
     layer3_out[4912] <= layer2_out[9073] & ~layer2_out[9072];
     layer3_out[4913] <= layer2_out[6153] | layer2_out[6154];
     layer3_out[4914] <= ~(layer2_out[7186] | layer2_out[7187]);
     layer3_out[4915] <= layer2_out[4293] & ~layer2_out[4294];
     layer3_out[4916] <= layer2_out[618] & ~layer2_out[619];
     layer3_out[4917] <= ~(layer2_out[1668] & layer2_out[1669]);
     layer3_out[4918] <= layer2_out[1449];
     layer3_out[4919] <= layer2_out[1324] & layer2_out[1325];
     layer3_out[4920] <= ~(layer2_out[1863] | layer2_out[1864]);
     layer3_out[4921] <= ~(layer2_out[9572] | layer2_out[9573]);
     layer3_out[4922] <= layer2_out[10109];
     layer3_out[4923] <= ~(layer2_out[7427] | layer2_out[7428]);
     layer3_out[4924] <= layer2_out[2279];
     layer3_out[4925] <= layer2_out[7243] & layer2_out[7244];
     layer3_out[4926] <= ~layer2_out[4104];
     layer3_out[4927] <= ~(layer2_out[8065] | layer2_out[8066]);
     layer3_out[4928] <= ~(layer2_out[6145] ^ layer2_out[6146]);
     layer3_out[4929] <= ~layer2_out[4313];
     layer3_out[4930] <= layer2_out[4854] & ~layer2_out[4853];
     layer3_out[4931] <= layer2_out[5936] ^ layer2_out[5937];
     layer3_out[4932] <= layer2_out[522] & layer2_out[523];
     layer3_out[4933] <= ~(layer2_out[6905] | layer2_out[6906]);
     layer3_out[4934] <= layer2_out[793] & ~layer2_out[794];
     layer3_out[4935] <= layer2_out[10662];
     layer3_out[4936] <= layer2_out[3959] & ~layer2_out[3960];
     layer3_out[4937] <= ~layer2_out[3752] | layer2_out[3753];
     layer3_out[4938] <= ~layer2_out[8186];
     layer3_out[4939] <= layer2_out[5032] & ~layer2_out[5031];
     layer3_out[4940] <= layer2_out[6509] & ~layer2_out[6508];
     layer3_out[4941] <= layer2_out[1290] & ~layer2_out[1289];
     layer3_out[4942] <= layer2_out[4093];
     layer3_out[4943] <= ~(layer2_out[8223] | layer2_out[8224]);
     layer3_out[4944] <= ~layer2_out[6321];
     layer3_out[4945] <= layer2_out[7679] & ~layer2_out[7680];
     layer3_out[4946] <= layer2_out[947] & ~layer2_out[946];
     layer3_out[4947] <= ~layer2_out[7225];
     layer3_out[4948] <= layer2_out[5163];
     layer3_out[4949] <= layer2_out[1815] ^ layer2_out[1816];
     layer3_out[4950] <= layer2_out[7341] & ~layer2_out[7340];
     layer3_out[4951] <= layer2_out[10020] & ~layer2_out[10019];
     layer3_out[4952] <= ~layer2_out[11958];
     layer3_out[4953] <= layer2_out[3032] & ~layer2_out[3033];
     layer3_out[4954] <= ~layer2_out[4806];
     layer3_out[4955] <= layer2_out[6250] & ~layer2_out[6251];
     layer3_out[4956] <= layer2_out[2266] & layer2_out[2267];
     layer3_out[4957] <= layer2_out[2758] & ~layer2_out[2759];
     layer3_out[4958] <= layer2_out[2990];
     layer3_out[4959] <= ~(layer2_out[340] ^ layer2_out[341]);
     layer3_out[4960] <= ~layer2_out[9994];
     layer3_out[4961] <= layer2_out[8615];
     layer3_out[4962] <= ~(layer2_out[9378] ^ layer2_out[9379]);
     layer3_out[4963] <= layer2_out[11608] & layer2_out[11609];
     layer3_out[4964] <= layer2_out[11941] & ~layer2_out[11942];
     layer3_out[4965] <= layer2_out[9273] ^ layer2_out[9274];
     layer3_out[4966] <= ~(layer2_out[7256] ^ layer2_out[7257]);
     layer3_out[4967] <= ~(layer2_out[5740] ^ layer2_out[5741]);
     layer3_out[4968] <= ~layer2_out[4859] | layer2_out[4860];
     layer3_out[4969] <= ~layer2_out[2455];
     layer3_out[4970] <= layer2_out[674];
     layer3_out[4971] <= layer2_out[314];
     layer3_out[4972] <= ~(layer2_out[3644] ^ layer2_out[3645]);
     layer3_out[4973] <= ~(layer2_out[2193] ^ layer2_out[2194]);
     layer3_out[4974] <= layer2_out[829];
     layer3_out[4975] <= layer2_out[4559];
     layer3_out[4976] <= layer2_out[5156] & layer2_out[5157];
     layer3_out[4977] <= layer2_out[1265] ^ layer2_out[1266];
     layer3_out[4978] <= layer2_out[5314];
     layer3_out[4979] <= layer2_out[9274] & ~layer2_out[9275];
     layer3_out[4980] <= ~(layer2_out[6765] | layer2_out[6766]);
     layer3_out[4981] <= layer2_out[11001] | layer2_out[11002];
     layer3_out[4982] <= ~(layer2_out[6230] | layer2_out[6231]);
     layer3_out[4983] <= layer2_out[9093] & ~layer2_out[9092];
     layer3_out[4984] <= ~layer2_out[596];
     layer3_out[4985] <= layer2_out[8225] & ~layer2_out[8224];
     layer3_out[4986] <= layer2_out[6613] ^ layer2_out[6614];
     layer3_out[4987] <= ~layer2_out[222];
     layer3_out[4988] <= ~(layer2_out[3332] ^ layer2_out[3333]);
     layer3_out[4989] <= layer2_out[8528] ^ layer2_out[8529];
     layer3_out[4990] <= ~layer2_out[3810];
     layer3_out[4991] <= layer2_out[1942] & layer2_out[1943];
     layer3_out[4992] <= ~layer2_out[5754];
     layer3_out[4993] <= ~layer2_out[5372] | layer2_out[5373];
     layer3_out[4994] <= ~(layer2_out[4420] & layer2_out[4421]);
     layer3_out[4995] <= layer2_out[11179];
     layer3_out[4996] <= ~layer2_out[257];
     layer3_out[4997] <= ~layer2_out[4101];
     layer3_out[4998] <= ~layer2_out[9690];
     layer3_out[4999] <= ~layer2_out[10287];
     layer3_out[5000] <= ~(layer2_out[7765] ^ layer2_out[7766]);
     layer3_out[5001] <= layer2_out[5073];
     layer3_out[5002] <= layer2_out[9953] & ~layer2_out[9952];
     layer3_out[5003] <= layer2_out[4165] & ~layer2_out[4166];
     layer3_out[5004] <= ~layer2_out[5939];
     layer3_out[5005] <= ~(layer2_out[2311] ^ layer2_out[2312]);
     layer3_out[5006] <= ~layer2_out[5273];
     layer3_out[5007] <= ~(layer2_out[11575] | layer2_out[11576]);
     layer3_out[5008] <= layer2_out[11261] & ~layer2_out[11260];
     layer3_out[5009] <= ~(layer2_out[2490] | layer2_out[2491]);
     layer3_out[5010] <= ~(layer2_out[5011] | layer2_out[5012]);
     layer3_out[5011] <= layer2_out[549] & ~layer2_out[550];
     layer3_out[5012] <= ~(layer2_out[301] | layer2_out[302]);
     layer3_out[5013] <= ~layer2_out[6955];
     layer3_out[5014] <= ~(layer2_out[3147] | layer2_out[3148]);
     layer3_out[5015] <= layer2_out[5593] & layer2_out[5594];
     layer3_out[5016] <= ~(layer2_out[1298] | layer2_out[1299]);
     layer3_out[5017] <= layer2_out[8794] & layer2_out[8795];
     layer3_out[5018] <= layer2_out[5432];
     layer3_out[5019] <= ~layer2_out[3939] | layer2_out[3938];
     layer3_out[5020] <= ~(layer2_out[10870] | layer2_out[10871]);
     layer3_out[5021] <= layer2_out[4075] & ~layer2_out[4074];
     layer3_out[5022] <= ~layer2_out[4740];
     layer3_out[5023] <= layer2_out[4397] & layer2_out[4398];
     layer3_out[5024] <= layer2_out[2049] & ~layer2_out[2050];
     layer3_out[5025] <= layer2_out[10319] | layer2_out[10320];
     layer3_out[5026] <= ~layer2_out[10697] | layer2_out[10696];
     layer3_out[5027] <= ~layer2_out[1601];
     layer3_out[5028] <= layer2_out[4619] & ~layer2_out[4618];
     layer3_out[5029] <= layer2_out[5716] & ~layer2_out[5717];
     layer3_out[5030] <= ~layer2_out[3773] | layer2_out[3772];
     layer3_out[5031] <= ~layer2_out[9335];
     layer3_out[5032] <= ~(layer2_out[11196] | layer2_out[11197]);
     layer3_out[5033] <= ~layer2_out[3700] | layer2_out[3699];
     layer3_out[5034] <= ~(layer2_out[11008] & layer2_out[11009]);
     layer3_out[5035] <= layer2_out[1943] & layer2_out[1944];
     layer3_out[5036] <= layer2_out[3888] ^ layer2_out[3889];
     layer3_out[5037] <= layer2_out[11897] & ~layer2_out[11898];
     layer3_out[5038] <= ~(layer2_out[5159] ^ layer2_out[5160]);
     layer3_out[5039] <= layer2_out[3915] & ~layer2_out[3916];
     layer3_out[5040] <= ~layer2_out[6285];
     layer3_out[5041] <= layer2_out[2799] & ~layer2_out[2800];
     layer3_out[5042] <= layer2_out[6707] & layer2_out[6708];
     layer3_out[5043] <= layer2_out[10416] & ~layer2_out[10417];
     layer3_out[5044] <= ~(layer2_out[11484] | layer2_out[11485]);
     layer3_out[5045] <= ~(layer2_out[2602] | layer2_out[2603]);
     layer3_out[5046] <= ~(layer2_out[11289] | layer2_out[11290]);
     layer3_out[5047] <= layer2_out[616] ^ layer2_out[617];
     layer3_out[5048] <= layer2_out[6157] & ~layer2_out[6156];
     layer3_out[5049] <= ~(layer2_out[1505] & layer2_out[1506]);
     layer3_out[5050] <= layer2_out[6226];
     layer3_out[5051] <= layer2_out[10967];
     layer3_out[5052] <= layer2_out[6412] & layer2_out[6413];
     layer3_out[5053] <= ~layer2_out[9331] | layer2_out[9330];
     layer3_out[5054] <= ~layer2_out[6176];
     layer3_out[5055] <= layer2_out[3384];
     layer3_out[5056] <= layer2_out[6334];
     layer3_out[5057] <= layer2_out[1327] & ~layer2_out[1326];
     layer3_out[5058] <= layer2_out[750];
     layer3_out[5059] <= ~layer2_out[3908];
     layer3_out[5060] <= ~layer2_out[7897];
     layer3_out[5061] <= layer2_out[1786] & ~layer2_out[1787];
     layer3_out[5062] <= ~(layer2_out[8737] | layer2_out[8738]);
     layer3_out[5063] <= layer2_out[6149] ^ layer2_out[6150];
     layer3_out[5064] <= layer2_out[516] & ~layer2_out[515];
     layer3_out[5065] <= layer2_out[7728];
     layer3_out[5066] <= ~layer2_out[1890];
     layer3_out[5067] <= ~layer2_out[8463];
     layer3_out[5068] <= ~(layer2_out[484] | layer2_out[485]);
     layer3_out[5069] <= layer2_out[4512] & layer2_out[4513];
     layer3_out[5070] <= layer2_out[9908] & ~layer2_out[9909];
     layer3_out[5071] <= layer2_out[10710];
     layer3_out[5072] <= layer2_out[4270] & ~layer2_out[4271];
     layer3_out[5073] <= layer2_out[10559];
     layer3_out[5074] <= layer2_out[2938] & ~layer2_out[2939];
     layer3_out[5075] <= layer2_out[10713] & ~layer2_out[10714];
     layer3_out[5076] <= ~(layer2_out[6268] | layer2_out[6269]);
     layer3_out[5077] <= ~(layer2_out[10091] ^ layer2_out[10092]);
     layer3_out[5078] <= layer2_out[5532] & ~layer2_out[5533];
     layer3_out[5079] <= ~(layer2_out[10407] | layer2_out[10408]);
     layer3_out[5080] <= layer2_out[11566];
     layer3_out[5081] <= layer2_out[10415] & layer2_out[10416];
     layer3_out[5082] <= layer2_out[906];
     layer3_out[5083] <= layer2_out[3673] & ~layer2_out[3672];
     layer3_out[5084] <= ~(layer2_out[8676] ^ layer2_out[8677]);
     layer3_out[5085] <= layer2_out[5013] & ~layer2_out[5012];
     layer3_out[5086] <= layer2_out[3596] & ~layer2_out[3597];
     layer3_out[5087] <= layer2_out[3584];
     layer3_out[5088] <= ~layer2_out[6355];
     layer3_out[5089] <= ~layer2_out[7591];
     layer3_out[5090] <= ~(layer2_out[10844] ^ layer2_out[10845]);
     layer3_out[5091] <= layer2_out[11033] & ~layer2_out[11032];
     layer3_out[5092] <= layer2_out[842] & ~layer2_out[841];
     layer3_out[5093] <= layer2_out[1088];
     layer3_out[5094] <= layer2_out[1166];
     layer3_out[5095] <= ~(layer2_out[1369] ^ layer2_out[1370]);
     layer3_out[5096] <= layer2_out[2722] ^ layer2_out[2723];
     layer3_out[5097] <= layer2_out[1872] & ~layer2_out[1873];
     layer3_out[5098] <= layer2_out[7565] | layer2_out[7566];
     layer3_out[5099] <= layer2_out[4469] & layer2_out[4470];
     layer3_out[5100] <= layer2_out[6305] & ~layer2_out[6306];
     layer3_out[5101] <= layer2_out[6864] & ~layer2_out[6865];
     layer3_out[5102] <= ~(layer2_out[7177] | layer2_out[7178]);
     layer3_out[5103] <= layer2_out[7139];
     layer3_out[5104] <= layer2_out[8227] & ~layer2_out[8228];
     layer3_out[5105] <= ~(layer2_out[5890] & layer2_out[5891]);
     layer3_out[5106] <= layer2_out[6697] & layer2_out[6698];
     layer3_out[5107] <= ~layer2_out[2796];
     layer3_out[5108] <= ~(layer2_out[7844] | layer2_out[7845]);
     layer3_out[5109] <= layer2_out[11819];
     layer3_out[5110] <= ~layer2_out[2587] | layer2_out[2586];
     layer3_out[5111] <= layer2_out[4037];
     layer3_out[5112] <= layer2_out[8271] & ~layer2_out[8272];
     layer3_out[5113] <= layer2_out[5655];
     layer3_out[5114] <= layer2_out[1972];
     layer3_out[5115] <= ~layer2_out[4453];
     layer3_out[5116] <= layer2_out[11261] ^ layer2_out[11262];
     layer3_out[5117] <= layer2_out[4524] | layer2_out[4525];
     layer3_out[5118] <= layer2_out[3334] & ~layer2_out[3335];
     layer3_out[5119] <= layer2_out[9899] & ~layer2_out[9900];
     layer3_out[5120] <= ~(layer2_out[215] ^ layer2_out[216]);
     layer3_out[5121] <= ~layer2_out[5134];
     layer3_out[5122] <= layer2_out[461];
     layer3_out[5123] <= ~layer2_out[5357];
     layer3_out[5124] <= layer2_out[10226] & layer2_out[10227];
     layer3_out[5125] <= layer2_out[4355];
     layer3_out[5126] <= layer2_out[10516] & ~layer2_out[10517];
     layer3_out[5127] <= ~layer2_out[10482] | layer2_out[10483];
     layer3_out[5128] <= layer2_out[9786];
     layer3_out[5129] <= layer2_out[5266] & ~layer2_out[5265];
     layer3_out[5130] <= ~layer2_out[11867];
     layer3_out[5131] <= ~layer2_out[7620] | layer2_out[7619];
     layer3_out[5132] <= ~(layer2_out[457] | layer2_out[458]);
     layer3_out[5133] <= layer2_out[2716] & layer2_out[2717];
     layer3_out[5134] <= layer2_out[3629];
     layer3_out[5135] <= layer2_out[2926] & ~layer2_out[2925];
     layer3_out[5136] <= ~layer2_out[914];
     layer3_out[5137] <= layer2_out[1471];
     layer3_out[5138] <= layer2_out[2252];
     layer3_out[5139] <= layer2_out[8637];
     layer3_out[5140] <= ~layer2_out[8210];
     layer3_out[5141] <= layer2_out[8276] & ~layer2_out[8277];
     layer3_out[5142] <= layer2_out[5626] ^ layer2_out[5627];
     layer3_out[5143] <= ~(layer2_out[9215] | layer2_out[9216]);
     layer3_out[5144] <= layer2_out[3878];
     layer3_out[5145] <= layer2_out[623] ^ layer2_out[624];
     layer3_out[5146] <= layer2_out[9024] & layer2_out[9025];
     layer3_out[5147] <= layer2_out[10749] & ~layer2_out[10748];
     layer3_out[5148] <= layer2_out[1542] & ~layer2_out[1541];
     layer3_out[5149] <= layer2_out[4375];
     layer3_out[5150] <= layer2_out[2072] ^ layer2_out[2073];
     layer3_out[5151] <= layer2_out[5302];
     layer3_out[5152] <= layer2_out[4770] & ~layer2_out[4769];
     layer3_out[5153] <= ~layer2_out[762];
     layer3_out[5154] <= layer2_out[8580];
     layer3_out[5155] <= layer2_out[6525] & layer2_out[6526];
     layer3_out[5156] <= ~layer2_out[4241];
     layer3_out[5157] <= layer2_out[8623] & ~layer2_out[8622];
     layer3_out[5158] <= layer2_out[7598] ^ layer2_out[7599];
     layer3_out[5159] <= layer2_out[117] & ~layer2_out[116];
     layer3_out[5160] <= layer2_out[128] & layer2_out[129];
     layer3_out[5161] <= layer2_out[8246];
     layer3_out[5162] <= layer2_out[8353];
     layer3_out[5163] <= layer2_out[1595] & ~layer2_out[1594];
     layer3_out[5164] <= ~(layer2_out[8080] ^ layer2_out[8081]);
     layer3_out[5165] <= ~layer2_out[7117];
     layer3_out[5166] <= ~(layer2_out[5216] | layer2_out[5217]);
     layer3_out[5167] <= layer2_out[10217] & ~layer2_out[10216];
     layer3_out[5168] <= ~layer2_out[7055];
     layer3_out[5169] <= ~layer2_out[11489];
     layer3_out[5170] <= layer2_out[7020];
     layer3_out[5171] <= layer2_out[8156] & ~layer2_out[8155];
     layer3_out[5172] <= ~layer2_out[8009] | layer2_out[8010];
     layer3_out[5173] <= layer2_out[3140] & ~layer2_out[3141];
     layer3_out[5174] <= layer2_out[4402] & ~layer2_out[4401];
     layer3_out[5175] <= layer2_out[1745] & layer2_out[1746];
     layer3_out[5176] <= ~layer2_out[10670];
     layer3_out[5177] <= ~(layer2_out[10428] | layer2_out[10429]);
     layer3_out[5178] <= layer2_out[11653] ^ layer2_out[11654];
     layer3_out[5179] <= ~(layer2_out[1955] | layer2_out[1956]);
     layer3_out[5180] <= ~layer2_out[8214];
     layer3_out[5181] <= layer2_out[445] & layer2_out[446];
     layer3_out[5182] <= layer2_out[3457] ^ layer2_out[3458];
     layer3_out[5183] <= ~layer2_out[11615];
     layer3_out[5184] <= ~layer2_out[5583] | layer2_out[5584];
     layer3_out[5185] <= ~(layer2_out[488] | layer2_out[489]);
     layer3_out[5186] <= ~layer2_out[11186];
     layer3_out[5187] <= ~(layer2_out[560] | layer2_out[561]);
     layer3_out[5188] <= ~layer2_out[8826] | layer2_out[8827];
     layer3_out[5189] <= layer2_out[10649] & ~layer2_out[10650];
     layer3_out[5190] <= ~layer2_out[2001];
     layer3_out[5191] <= layer2_out[911] & layer2_out[912];
     layer3_out[5192] <= layer2_out[9739] & ~layer2_out[9740];
     layer3_out[5193] <= ~layer2_out[3120];
     layer3_out[5194] <= layer2_out[7212] & layer2_out[7213];
     layer3_out[5195] <= layer2_out[8315] & ~layer2_out[8314];
     layer3_out[5196] <= layer2_out[6595] & layer2_out[6596];
     layer3_out[5197] <= layer2_out[8572] & layer2_out[8573];
     layer3_out[5198] <= layer2_out[5718] & ~layer2_out[5717];
     layer3_out[5199] <= ~(layer2_out[1392] ^ layer2_out[1393]);
     layer3_out[5200] <= ~(layer2_out[7862] | layer2_out[7863]);
     layer3_out[5201] <= ~(layer2_out[7392] | layer2_out[7393]);
     layer3_out[5202] <= ~layer2_out[4198];
     layer3_out[5203] <= layer2_out[3337] & layer2_out[3338];
     layer3_out[5204] <= ~(layer2_out[3925] & layer2_out[3926]);
     layer3_out[5205] <= layer2_out[1751];
     layer3_out[5206] <= ~(layer2_out[9868] ^ layer2_out[9869]);
     layer3_out[5207] <= ~layer2_out[11564];
     layer3_out[5208] <= ~(layer2_out[10299] ^ layer2_out[10300]);
     layer3_out[5209] <= ~layer2_out[9688];
     layer3_out[5210] <= layer2_out[8021];
     layer3_out[5211] <= layer2_out[9849];
     layer3_out[5212] <= layer2_out[9067] & ~layer2_out[9066];
     layer3_out[5213] <= ~(layer2_out[7529] | layer2_out[7530]);
     layer3_out[5214] <= ~layer2_out[5710];
     layer3_out[5215] <= layer2_out[11764] & layer2_out[11765];
     layer3_out[5216] <= layer2_out[3997] & ~layer2_out[3998];
     layer3_out[5217] <= ~(layer2_out[1643] ^ layer2_out[1644]);
     layer3_out[5218] <= layer2_out[10571] & layer2_out[10572];
     layer3_out[5219] <= layer2_out[1201] & ~layer2_out[1200];
     layer3_out[5220] <= layer2_out[3917] & ~layer2_out[3916];
     layer3_out[5221] <= layer2_out[6199] & layer2_out[6200];
     layer3_out[5222] <= ~layer2_out[3795];
     layer3_out[5223] <= layer2_out[10529] & ~layer2_out[10530];
     layer3_out[5224] <= layer2_out[11904] & ~layer2_out[11905];
     layer3_out[5225] <= ~(layer2_out[2283] ^ layer2_out[2284]);
     layer3_out[5226] <= layer2_out[7500] & layer2_out[7501];
     layer3_out[5227] <= layer2_out[5469] & layer2_out[5470];
     layer3_out[5228] <= layer2_out[6159];
     layer3_out[5229] <= layer2_out[10262];
     layer3_out[5230] <= ~(layer2_out[10807] ^ layer2_out[10808]);
     layer3_out[5231] <= layer2_out[7842] & layer2_out[7843];
     layer3_out[5232] <= layer2_out[5097];
     layer3_out[5233] <= ~(layer2_out[8088] ^ layer2_out[8089]);
     layer3_out[5234] <= layer2_out[8632];
     layer3_out[5235] <= ~(layer2_out[5340] | layer2_out[5341]);
     layer3_out[5236] <= ~layer2_out[10274];
     layer3_out[5237] <= ~layer2_out[8270];
     layer3_out[5238] <= layer2_out[10137] | layer2_out[10138];
     layer3_out[5239] <= layer2_out[5758] ^ layer2_out[5759];
     layer3_out[5240] <= layer2_out[11486];
     layer3_out[5241] <= layer2_out[10724];
     layer3_out[5242] <= layer2_out[1608] & layer2_out[1609];
     layer3_out[5243] <= layer2_out[5759] & ~layer2_out[5760];
     layer3_out[5244] <= layer2_out[7995] & layer2_out[7996];
     layer3_out[5245] <= ~layer2_out[4287];
     layer3_out[5246] <= layer2_out[7198] & layer2_out[7199];
     layer3_out[5247] <= layer2_out[4556] & ~layer2_out[4557];
     layer3_out[5248] <= layer2_out[6600] & layer2_out[6601];
     layer3_out[5249] <= ~(layer2_out[11239] | layer2_out[11240]);
     layer3_out[5250] <= layer2_out[4497];
     layer3_out[5251] <= ~layer2_out[1953];
     layer3_out[5252] <= ~layer2_out[10200];
     layer3_out[5253] <= layer2_out[8729] & ~layer2_out[8730];
     layer3_out[5254] <= layer2_out[11721];
     layer3_out[5255] <= ~layer2_out[9077];
     layer3_out[5256] <= ~(layer2_out[163] ^ layer2_out[164]);
     layer3_out[5257] <= layer2_out[4907];
     layer3_out[5258] <= layer2_out[10345];
     layer3_out[5259] <= ~(layer2_out[6092] | layer2_out[6093]);
     layer3_out[5260] <= ~layer2_out[250];
     layer3_out[5261] <= ~(layer2_out[11724] | layer2_out[11725]);
     layer3_out[5262] <= layer2_out[152] & ~layer2_out[151];
     layer3_out[5263] <= layer2_out[1067] & ~layer2_out[1068];
     layer3_out[5264] <= ~layer2_out[8682] | layer2_out[8681];
     layer3_out[5265] <= layer2_out[34] & layer2_out[35];
     layer3_out[5266] <= ~layer2_out[1194];
     layer3_out[5267] <= ~(layer2_out[6242] | layer2_out[6243]);
     layer3_out[5268] <= ~(layer2_out[3009] ^ layer2_out[3010]);
     layer3_out[5269] <= ~layer2_out[2018];
     layer3_out[5270] <= ~(layer2_out[4298] & layer2_out[4299]);
     layer3_out[5271] <= layer2_out[10354];
     layer3_out[5272] <= layer2_out[11525] ^ layer2_out[11526];
     layer3_out[5273] <= ~layer2_out[8220] | layer2_out[8219];
     layer3_out[5274] <= ~layer2_out[8518] | layer2_out[8517];
     layer3_out[5275] <= layer2_out[9626] & layer2_out[9627];
     layer3_out[5276] <= layer2_out[10059] & layer2_out[10060];
     layer3_out[5277] <= ~(layer2_out[533] ^ layer2_out[534]);
     layer3_out[5278] <= layer2_out[11199];
     layer3_out[5279] <= layer2_out[9845] & layer2_out[9846];
     layer3_out[5280] <= layer2_out[3038] ^ layer2_out[3039];
     layer3_out[5281] <= layer2_out[504];
     layer3_out[5282] <= layer2_out[211];
     layer3_out[5283] <= layer2_out[1433] | layer2_out[1434];
     layer3_out[5284] <= layer2_out[189] & ~layer2_out[188];
     layer3_out[5285] <= layer2_out[30] & ~layer2_out[31];
     layer3_out[5286] <= layer2_out[2033] ^ layer2_out[2034];
     layer3_out[5287] <= layer2_out[9938];
     layer3_out[5288] <= layer2_out[10892] & ~layer2_out[10893];
     layer3_out[5289] <= ~layer2_out[6259];
     layer3_out[5290] <= layer2_out[11509] & ~layer2_out[11510];
     layer3_out[5291] <= layer2_out[11584];
     layer3_out[5292] <= ~layer2_out[9288];
     layer3_out[5293] <= ~(layer2_out[10964] | layer2_out[10965]);
     layer3_out[5294] <= layer2_out[8993] | layer2_out[8994];
     layer3_out[5295] <= layer2_out[10602] ^ layer2_out[10603];
     layer3_out[5296] <= layer2_out[4979] & layer2_out[4980];
     layer3_out[5297] <= ~layer2_out[6761] | layer2_out[6762];
     layer3_out[5298] <= layer2_out[5942] ^ layer2_out[5943];
     layer3_out[5299] <= layer2_out[3235];
     layer3_out[5300] <= layer2_out[10776] ^ layer2_out[10777];
     layer3_out[5301] <= ~layer2_out[7357];
     layer3_out[5302] <= layer2_out[11802] & ~layer2_out[11801];
     layer3_out[5303] <= layer2_out[3079] & ~layer2_out[3078];
     layer3_out[5304] <= layer2_out[6872];
     layer3_out[5305] <= layer2_out[6143] & ~layer2_out[6144];
     layer3_out[5306] <= layer2_out[7052];
     layer3_out[5307] <= ~(layer2_out[8478] & layer2_out[8479]);
     layer3_out[5308] <= layer2_out[8332] & layer2_out[8333];
     layer3_out[5309] <= ~(layer2_out[3565] ^ layer2_out[3566]);
     layer3_out[5310] <= ~layer2_out[7526];
     layer3_out[5311] <= layer2_out[4677] & ~layer2_out[4678];
     layer3_out[5312] <= ~layer2_out[7093];
     layer3_out[5313] <= layer2_out[7706];
     layer3_out[5314] <= layer2_out[5371] & ~layer2_out[5370];
     layer3_out[5315] <= layer2_out[5820];
     layer3_out[5316] <= layer2_out[6078];
     layer3_out[5317] <= ~layer2_out[7189];
     layer3_out[5318] <= layer2_out[9552] & ~layer2_out[9553];
     layer3_out[5319] <= ~layer2_out[9410];
     layer3_out[5320] <= ~layer2_out[11232];
     layer3_out[5321] <= layer2_out[9897] & ~layer2_out[9896];
     layer3_out[5322] <= ~layer2_out[10627];
     layer3_out[5323] <= layer2_out[1949];
     layer3_out[5324] <= ~(layer2_out[4711] | layer2_out[4712]);
     layer3_out[5325] <= layer2_out[10159] & ~layer2_out[10158];
     layer3_out[5326] <= ~layer2_out[11447];
     layer3_out[5327] <= layer2_out[717] & ~layer2_out[716];
     layer3_out[5328] <= layer2_out[4641] & ~layer2_out[4640];
     layer3_out[5329] <= ~(layer2_out[1783] & layer2_out[1784]);
     layer3_out[5330] <= ~layer2_out[1079];
     layer3_out[5331] <= ~layer2_out[5377];
     layer3_out[5332] <= ~layer2_out[6558] | layer2_out[6559];
     layer3_out[5333] <= layer2_out[6025] ^ layer2_out[6026];
     layer3_out[5334] <= ~layer2_out[10640];
     layer3_out[5335] <= ~layer2_out[6377];
     layer3_out[5336] <= layer2_out[11416] & layer2_out[11417];
     layer3_out[5337] <= layer2_out[6018];
     layer3_out[5338] <= ~(layer2_out[7391] | layer2_out[7392]);
     layer3_out[5339] <= ~(layer2_out[7021] | layer2_out[7022]);
     layer3_out[5340] <= ~layer2_out[61] | layer2_out[62];
     layer3_out[5341] <= ~layer2_out[1466];
     layer3_out[5342] <= ~(layer2_out[7686] | layer2_out[7687]);
     layer3_out[5343] <= layer2_out[6118] & ~layer2_out[6119];
     layer3_out[5344] <= layer2_out[8201] & layer2_out[8202];
     layer3_out[5345] <= ~layer2_out[498];
     layer3_out[5346] <= ~(layer2_out[2861] | layer2_out[2862]);
     layer3_out[5347] <= layer2_out[2704] & ~layer2_out[2705];
     layer3_out[5348] <= layer2_out[799] & ~layer2_out[800];
     layer3_out[5349] <= layer2_out[968] & layer2_out[969];
     layer3_out[5350] <= ~(layer2_out[5981] ^ layer2_out[5982]);
     layer3_out[5351] <= layer2_out[7442];
     layer3_out[5352] <= ~layer2_out[1544];
     layer3_out[5353] <= ~layer2_out[1801] | layer2_out[1802];
     layer3_out[5354] <= ~(layer2_out[4684] | layer2_out[4685]);
     layer3_out[5355] <= layer2_out[5879] & ~layer2_out[5878];
     layer3_out[5356] <= ~(layer2_out[2023] | layer2_out[2024]);
     layer3_out[5357] <= ~(layer2_out[1119] | layer2_out[1120]);
     layer3_out[5358] <= layer2_out[4320] | layer2_out[4321];
     layer3_out[5359] <= layer2_out[3815] & ~layer2_out[3814];
     layer3_out[5360] <= ~layer2_out[7914];
     layer3_out[5361] <= ~(layer2_out[8883] | layer2_out[8884]);
     layer3_out[5362] <= layer2_out[9482] ^ layer2_out[9483];
     layer3_out[5363] <= ~(layer2_out[7088] | layer2_out[7089]);
     layer3_out[5364] <= layer2_out[3021] & layer2_out[3022];
     layer3_out[5365] <= layer2_out[1686] & ~layer2_out[1685];
     layer3_out[5366] <= layer2_out[3952];
     layer3_out[5367] <= layer2_out[4409] ^ layer2_out[4410];
     layer3_out[5368] <= ~layer2_out[5957] | layer2_out[5958];
     layer3_out[5369] <= ~(layer2_out[5315] | layer2_out[5316]);
     layer3_out[5370] <= ~(layer2_out[3568] | layer2_out[3569]);
     layer3_out[5371] <= ~(layer2_out[10479] ^ layer2_out[10480]);
     layer3_out[5372] <= ~(layer2_out[562] | layer2_out[563]);
     layer3_out[5373] <= layer2_out[7669];
     layer3_out[5374] <= layer2_out[6792];
     layer3_out[5375] <= ~layer2_out[3215];
     layer3_out[5376] <= layer2_out[468];
     layer3_out[5377] <= layer2_out[6625];
     layer3_out[5378] <= ~layer2_out[111];
     layer3_out[5379] <= layer2_out[5481] & layer2_out[5482];
     layer3_out[5380] <= ~layer2_out[5480] | layer2_out[5481];
     layer3_out[5381] <= ~layer2_out[1148] | layer2_out[1147];
     layer3_out[5382] <= layer2_out[10974];
     layer3_out[5383] <= layer2_out[6228] ^ layer2_out[6229];
     layer3_out[5384] <= layer2_out[5751] & ~layer2_out[5750];
     layer3_out[5385] <= layer2_out[4437] & ~layer2_out[4438];
     layer3_out[5386] <= ~(layer2_out[1432] ^ layer2_out[1433]);
     layer3_out[5387] <= ~layer2_out[1419] | layer2_out[1420];
     layer3_out[5388] <= ~layer2_out[9879];
     layer3_out[5389] <= ~layer2_out[7076];
     layer3_out[5390] <= layer2_out[10044];
     layer3_out[5391] <= layer2_out[9518] | layer2_out[9519];
     layer3_out[5392] <= ~(layer2_out[10635] ^ layer2_out[10636]);
     layer3_out[5393] <= layer2_out[1449];
     layer3_out[5394] <= layer2_out[2219];
     layer3_out[5395] <= layer2_out[8134];
     layer3_out[5396] <= ~layer2_out[10112];
     layer3_out[5397] <= ~(layer2_out[2046] | layer2_out[2047]);
     layer3_out[5398] <= layer2_out[8095];
     layer3_out[5399] <= layer2_out[11925] & layer2_out[11926];
     layer3_out[5400] <= ~layer2_out[659];
     layer3_out[5401] <= layer2_out[4098] & layer2_out[4099];
     layer3_out[5402] <= layer2_out[7420] & ~layer2_out[7421];
     layer3_out[5403] <= layer2_out[6266];
     layer3_out[5404] <= layer2_out[2877] & ~layer2_out[2878];
     layer3_out[5405] <= ~layer2_out[3164] | layer2_out[3165];
     layer3_out[5406] <= ~layer2_out[8153];
     layer3_out[5407] <= ~layer2_out[8400];
     layer3_out[5408] <= layer2_out[5563] ^ layer2_out[5564];
     layer3_out[5409] <= ~(layer2_out[8265] | layer2_out[8266]);
     layer3_out[5410] <= layer2_out[7426] & ~layer2_out[7427];
     layer3_out[5411] <= layer2_out[8083] ^ layer2_out[8084];
     layer3_out[5412] <= layer2_out[2131] ^ layer2_out[2132];
     layer3_out[5413] <= layer2_out[877] & layer2_out[878];
     layer3_out[5414] <= layer2_out[8854] & layer2_out[8855];
     layer3_out[5415] <= layer2_out[3068] ^ layer2_out[3069];
     layer3_out[5416] <= layer2_out[8385];
     layer3_out[5417] <= ~layer2_out[1904];
     layer3_out[5418] <= ~(layer2_out[1422] | layer2_out[1423]);
     layer3_out[5419] <= layer2_out[4981];
     layer3_out[5420] <= layer2_out[5756] & layer2_out[5757];
     layer3_out[5421] <= layer2_out[976] | layer2_out[977];
     layer3_out[5422] <= layer2_out[2500];
     layer3_out[5423] <= ~layer2_out[1268];
     layer3_out[5424] <= layer2_out[6015] & layer2_out[6016];
     layer3_out[5425] <= ~(layer2_out[9470] | layer2_out[9471]);
     layer3_out[5426] <= ~layer2_out[3808] | layer2_out[3807];
     layer3_out[5427] <= layer2_out[2181] & ~layer2_out[2180];
     layer3_out[5428] <= ~(layer2_out[11684] | layer2_out[11685]);
     layer3_out[5429] <= ~(layer2_out[11480] ^ layer2_out[11481]);
     layer3_out[5430] <= layer2_out[6238] & ~layer2_out[6237];
     layer3_out[5431] <= layer2_out[1180];
     layer3_out[5432] <= layer2_out[2986] & ~layer2_out[2987];
     layer3_out[5433] <= layer2_out[11015] & ~layer2_out[11016];
     layer3_out[5434] <= layer2_out[11031] & ~layer2_out[11032];
     layer3_out[5435] <= layer2_out[7131] & ~layer2_out[7132];
     layer3_out[5436] <= ~layer2_out[9325];
     layer3_out[5437] <= ~layer2_out[11902];
     layer3_out[5438] <= layer2_out[4154];
     layer3_out[5439] <= layer2_out[10978] & ~layer2_out[10979];
     layer3_out[5440] <= ~layer2_out[4436];
     layer3_out[5441] <= ~layer2_out[8812];
     layer3_out[5442] <= layer2_out[5985] ^ layer2_out[5986];
     layer3_out[5443] <= layer2_out[1489];
     layer3_out[5444] <= layer2_out[6165] & ~layer2_out[6166];
     layer3_out[5445] <= ~(layer2_out[4716] | layer2_out[4717]);
     layer3_out[5446] <= ~layer2_out[751];
     layer3_out[5447] <= layer2_out[8423] & ~layer2_out[8424];
     layer3_out[5448] <= ~(layer2_out[11362] | layer2_out[11363]);
     layer3_out[5449] <= ~layer2_out[427];
     layer3_out[5450] <= layer2_out[4530];
     layer3_out[5451] <= layer2_out[4187];
     layer3_out[5452] <= layer2_out[4358];
     layer3_out[5453] <= layer2_out[7367] & layer2_out[7368];
     layer3_out[5454] <= layer2_out[5140] & ~layer2_out[5139];
     layer3_out[5455] <= ~layer2_out[1191] | layer2_out[1192];
     layer3_out[5456] <= ~layer2_out[4602];
     layer3_out[5457] <= ~layer2_out[11898];
     layer3_out[5458] <= layer2_out[2766];
     layer3_out[5459] <= ~(layer2_out[10764] | layer2_out[10765]);
     layer3_out[5460] <= ~(layer2_out[3360] | layer2_out[3361]);
     layer3_out[5461] <= layer2_out[4868] & ~layer2_out[4869];
     layer3_out[5462] <= ~(layer2_out[2194] ^ layer2_out[2195]);
     layer3_out[5463] <= layer2_out[5176] & layer2_out[5177];
     layer3_out[5464] <= ~layer2_out[4368];
     layer3_out[5465] <= layer2_out[9130] & ~layer2_out[9131];
     layer3_out[5466] <= layer2_out[1095] & ~layer2_out[1096];
     layer3_out[5467] <= ~layer2_out[9807];
     layer3_out[5468] <= ~(layer2_out[2111] & layer2_out[2112]);
     layer3_out[5469] <= ~layer2_out[1476];
     layer3_out[5470] <= ~(layer2_out[9991] ^ layer2_out[9992]);
     layer3_out[5471] <= layer2_out[2952];
     layer3_out[5472] <= layer2_out[421] & ~layer2_out[420];
     layer3_out[5473] <= layer2_out[6303] & layer2_out[6304];
     layer3_out[5474] <= layer2_out[10467] | layer2_out[10468];
     layer3_out[5475] <= ~(layer2_out[10898] ^ layer2_out[10899]);
     layer3_out[5476] <= ~(layer2_out[6389] | layer2_out[6390]);
     layer3_out[5477] <= ~layer2_out[8249];
     layer3_out[5478] <= layer2_out[5182];
     layer3_out[5479] <= layer2_out[3208] & ~layer2_out[3207];
     layer3_out[5480] <= ~(layer2_out[3233] ^ layer2_out[3234]);
     layer3_out[5481] <= layer2_out[1675] ^ layer2_out[1676];
     layer3_out[5482] <= layer2_out[11609] & ~layer2_out[11610];
     layer3_out[5483] <= layer2_out[10500] & ~layer2_out[10499];
     layer3_out[5484] <= layer2_out[9239];
     layer3_out[5485] <= layer2_out[2209];
     layer3_out[5486] <= layer2_out[1933] & ~layer2_out[1932];
     layer3_out[5487] <= layer2_out[625] & layer2_out[626];
     layer3_out[5488] <= layer2_out[786] & layer2_out[787];
     layer3_out[5489] <= layer2_out[6550] & layer2_out[6551];
     layer3_out[5490] <= layer2_out[7280] ^ layer2_out[7281];
     layer3_out[5491] <= layer2_out[8091] ^ layer2_out[8092];
     layer3_out[5492] <= ~layer2_out[11737];
     layer3_out[5493] <= layer2_out[4135] & ~layer2_out[4134];
     layer3_out[5494] <= layer2_out[8532] & ~layer2_out[8533];
     layer3_out[5495] <= ~(layer2_out[3302] | layer2_out[3303]);
     layer3_out[5496] <= layer2_out[10576] & layer2_out[10577];
     layer3_out[5497] <= layer2_out[9347] & ~layer2_out[9346];
     layer3_out[5498] <= ~layer2_out[2969];
     layer3_out[5499] <= ~(layer2_out[10957] ^ layer2_out[10958]);
     layer3_out[5500] <= layer2_out[860] & layer2_out[861];
     layer3_out[5501] <= ~layer2_out[6849];
     layer3_out[5502] <= layer2_out[7757] & ~layer2_out[7756];
     layer3_out[5503] <= ~layer2_out[1701];
     layer3_out[5504] <= layer2_out[3068] & ~layer2_out[3067];
     layer3_out[5505] <= layer2_out[1555] & layer2_out[1556];
     layer3_out[5506] <= layer2_out[1134] & layer2_out[1135];
     layer3_out[5507] <= ~layer2_out[11838];
     layer3_out[5508] <= layer2_out[1034];
     layer3_out[5509] <= ~layer2_out[1079];
     layer3_out[5510] <= ~(layer2_out[9990] ^ layer2_out[9991]);
     layer3_out[5511] <= layer2_out[11017] & layer2_out[11018];
     layer3_out[5512] <= layer2_out[1596] ^ layer2_out[1597];
     layer3_out[5513] <= layer2_out[6309] ^ layer2_out[6310];
     layer3_out[5514] <= ~layer2_out[1000];
     layer3_out[5515] <= ~layer2_out[4235];
     layer3_out[5516] <= layer2_out[8309] & layer2_out[8310];
     layer3_out[5517] <= layer2_out[7660] & ~layer2_out[7661];
     layer3_out[5518] <= ~layer2_out[9168];
     layer3_out[5519] <= layer2_out[8710] ^ layer2_out[8711];
     layer3_out[5520] <= layer2_out[8721];
     layer3_out[5521] <= layer2_out[3152] & layer2_out[3153];
     layer3_out[5522] <= ~(layer2_out[5295] | layer2_out[5296]);
     layer3_out[5523] <= ~(layer2_out[2855] | layer2_out[2856]);
     layer3_out[5524] <= ~(layer2_out[8467] & layer2_out[8468]);
     layer3_out[5525] <= ~(layer2_out[2012] | layer2_out[2013]);
     layer3_out[5526] <= ~(layer2_out[126] ^ layer2_out[127]);
     layer3_out[5527] <= layer2_out[8502] & ~layer2_out[8503];
     layer3_out[5528] <= ~(layer2_out[4972] ^ layer2_out[4973]);
     layer3_out[5529] <= layer2_out[11304] | layer2_out[11305];
     layer3_out[5530] <= ~layer2_out[4644];
     layer3_out[5531] <= layer2_out[2275] ^ layer2_out[2276];
     layer3_out[5532] <= ~(layer2_out[6458] ^ layer2_out[6459]);
     layer3_out[5533] <= ~(layer2_out[2641] | layer2_out[2642]);
     layer3_out[5534] <= ~(layer2_out[2815] ^ layer2_out[2816]);
     layer3_out[5535] <= layer2_out[4719];
     layer3_out[5536] <= layer2_out[7540];
     layer3_out[5537] <= ~(layer2_out[10550] | layer2_out[10551]);
     layer3_out[5538] <= layer2_out[11829] & ~layer2_out[11828];
     layer3_out[5539] <= layer2_out[9766];
     layer3_out[5540] <= ~layer2_out[5858];
     layer3_out[5541] <= layer2_out[8026];
     layer3_out[5542] <= layer2_out[6388];
     layer3_out[5543] <= ~(layer2_out[3339] ^ layer2_out[3340]);
     layer3_out[5544] <= layer2_out[4856] & ~layer2_out[4857];
     layer3_out[5545] <= ~layer2_out[4372];
     layer3_out[5546] <= layer2_out[4808] & layer2_out[4809];
     layer3_out[5547] <= layer2_out[2292];
     layer3_out[5548] <= layer2_out[277] & ~layer2_out[278];
     layer3_out[5549] <= layer2_out[8346] & ~layer2_out[8347];
     layer3_out[5550] <= layer2_out[5330] & ~layer2_out[5331];
     layer3_out[5551] <= ~layer2_out[7524] | layer2_out[7523];
     layer3_out[5552] <= ~(layer2_out[7945] | layer2_out[7946]);
     layer3_out[5553] <= layer2_out[8408] ^ layer2_out[8409];
     layer3_out[5554] <= ~(layer2_out[3520] | layer2_out[3521]);
     layer3_out[5555] <= layer2_out[1583] ^ layer2_out[1584];
     layer3_out[5556] <= layer2_out[4139];
     layer3_out[5557] <= layer2_out[9232];
     layer3_out[5558] <= layer2_out[10372] & ~layer2_out[10371];
     layer3_out[5559] <= layer2_out[11929] ^ layer2_out[11930];
     layer3_out[5560] <= layer2_out[3807];
     layer3_out[5561] <= layer2_out[3364] & ~layer2_out[3363];
     layer3_out[5562] <= ~(layer2_out[5665] | layer2_out[5666]);
     layer3_out[5563] <= ~layer2_out[5273];
     layer3_out[5564] <= layer2_out[5338];
     layer3_out[5565] <= layer2_out[3291] & ~layer2_out[3292];
     layer3_out[5566] <= layer2_out[8284] & ~layer2_out[8283];
     layer3_out[5567] <= layer2_out[4972] & ~layer2_out[4971];
     layer3_out[5568] <= layer2_out[10018] & ~layer2_out[10019];
     layer3_out[5569] <= ~layer2_out[4716];
     layer3_out[5570] <= layer2_out[11346] & layer2_out[11347];
     layer3_out[5571] <= layer2_out[11572];
     layer3_out[5572] <= ~(layer2_out[3654] | layer2_out[3655]);
     layer3_out[5573] <= layer2_out[3878];
     layer3_out[5574] <= ~(layer2_out[11945] | layer2_out[11946]);
     layer3_out[5575] <= layer2_out[6598] & layer2_out[6599];
     layer3_out[5576] <= ~(layer2_out[903] ^ layer2_out[904]);
     layer3_out[5577] <= layer2_out[6752] ^ layer2_out[6753];
     layer3_out[5578] <= ~(layer2_out[11860] ^ layer2_out[11861]);
     layer3_out[5579] <= layer2_out[4081];
     layer3_out[5580] <= layer2_out[10088] & ~layer2_out[10087];
     layer3_out[5581] <= layer2_out[11864] ^ layer2_out[11865];
     layer3_out[5582] <= layer2_out[2076] & layer2_out[2077];
     layer3_out[5583] <= layer2_out[9310] ^ layer2_out[9311];
     layer3_out[5584] <= layer2_out[2520] & layer2_out[2521];
     layer3_out[5585] <= layer2_out[11394] & ~layer2_out[11395];
     layer3_out[5586] <= ~(layer2_out[1822] | layer2_out[1823]);
     layer3_out[5587] <= layer2_out[6375];
     layer3_out[5588] <= ~(layer2_out[8798] | layer2_out[8799]);
     layer3_out[5589] <= layer2_out[9580];
     layer3_out[5590] <= layer2_out[6272] & ~layer2_out[6271];
     layer3_out[5591] <= ~layer2_out[7801];
     layer3_out[5592] <= layer2_out[1106];
     layer3_out[5593] <= ~(layer2_out[9308] | layer2_out[9309]);
     layer3_out[5594] <= layer2_out[2776] | layer2_out[2777];
     layer3_out[5595] <= layer2_out[8140] & layer2_out[8141];
     layer3_out[5596] <= layer2_out[6797];
     layer3_out[5597] <= layer2_out[11928] & layer2_out[11929];
     layer3_out[5598] <= ~(layer2_out[9385] ^ layer2_out[9386]);
     layer3_out[5599] <= ~layer2_out[9539];
     layer3_out[5600] <= layer2_out[5235] & layer2_out[5236];
     layer3_out[5601] <= layer2_out[11237];
     layer3_out[5602] <= ~(layer2_out[332] | layer2_out[333]);
     layer3_out[5603] <= layer2_out[7960];
     layer3_out[5604] <= ~(layer2_out[11942] ^ layer2_out[11943]);
     layer3_out[5605] <= ~(layer2_out[7902] & layer2_out[7903]);
     layer3_out[5606] <= layer2_out[10912] & ~layer2_out[10913];
     layer3_out[5607] <= ~(layer2_out[718] ^ layer2_out[719]);
     layer3_out[5608] <= ~(layer2_out[11036] | layer2_out[11037]);
     layer3_out[5609] <= ~(layer2_out[1224] | layer2_out[1225]);
     layer3_out[5610] <= ~layer2_out[1587];
     layer3_out[5611] <= layer2_out[139] & ~layer2_out[138];
     layer3_out[5612] <= layer2_out[9990] & ~layer2_out[9989];
     layer3_out[5613] <= ~layer2_out[7122];
     layer3_out[5614] <= layer2_out[1972];
     layer3_out[5615] <= ~layer2_out[439];
     layer3_out[5616] <= layer2_out[11698] & layer2_out[11699];
     layer3_out[5617] <= ~(layer2_out[3764] | layer2_out[3765]);
     layer3_out[5618] <= layer2_out[9790] ^ layer2_out[9791];
     layer3_out[5619] <= layer2_out[3565] & ~layer2_out[3564];
     layer3_out[5620] <= ~layer2_out[9532];
     layer3_out[5621] <= layer2_out[10179] & ~layer2_out[10178];
     layer3_out[5622] <= layer2_out[10241] & layer2_out[10242];
     layer3_out[5623] <= ~layer2_out[7553];
     layer3_out[5624] <= ~(layer2_out[11855] | layer2_out[11856]);
     layer3_out[5625] <= layer2_out[9205] & ~layer2_out[9204];
     layer3_out[5626] <= ~layer2_out[2025];
     layer3_out[5627] <= layer2_out[8992] ^ layer2_out[8993];
     layer3_out[5628] <= layer2_out[5690] & layer2_out[5691];
     layer3_out[5629] <= layer2_out[3313] ^ layer2_out[3314];
     layer3_out[5630] <= ~(layer2_out[1189] ^ layer2_out[1190]);
     layer3_out[5631] <= layer2_out[308];
     layer3_out[5632] <= layer2_out[6324] & ~layer2_out[6323];
     layer3_out[5633] <= ~layer2_out[3750];
     layer3_out[5634] <= layer2_out[10389];
     layer3_out[5635] <= layer2_out[4191];
     layer3_out[5636] <= ~(layer2_out[3510] & layer2_out[3511]);
     layer3_out[5637] <= layer2_out[7313];
     layer3_out[5638] <= ~(layer2_out[4511] ^ layer2_out[4512]);
     layer3_out[5639] <= layer2_out[9735] & layer2_out[9736];
     layer3_out[5640] <= ~layer2_out[11809];
     layer3_out[5641] <= ~layer2_out[9668] | layer2_out[9669];
     layer3_out[5642] <= layer2_out[11088] ^ layer2_out[11089];
     layer3_out[5643] <= ~layer2_out[4267] | layer2_out[4268];
     layer3_out[5644] <= layer2_out[11493] & ~layer2_out[11494];
     layer3_out[5645] <= ~(layer2_out[5986] ^ layer2_out[5987]);
     layer3_out[5646] <= layer2_out[1571] ^ layer2_out[1572];
     layer3_out[5647] <= layer2_out[9320];
     layer3_out[5648] <= ~(layer2_out[5943] ^ layer2_out[5944]);
     layer3_out[5649] <= layer2_out[11087];
     layer3_out[5650] <= layer2_out[8470];
     layer3_out[5651] <= ~layer2_out[11799];
     layer3_out[5652] <= layer2_out[4222];
     layer3_out[5653] <= layer2_out[1788] & ~layer2_out[1787];
     layer3_out[5654] <= layer2_out[82] ^ layer2_out[83];
     layer3_out[5655] <= layer2_out[10188] & ~layer2_out[10187];
     layer3_out[5656] <= layer2_out[4659];
     layer3_out[5657] <= ~layer2_out[8173];
     layer3_out[5658] <= layer2_out[1893] & layer2_out[1894];
     layer3_out[5659] <= layer2_out[9941] & ~layer2_out[9940];
     layer3_out[5660] <= ~layer2_out[10604];
     layer3_out[5661] <= layer2_out[7505];
     layer3_out[5662] <= layer2_out[6277] ^ layer2_out[6278];
     layer3_out[5663] <= layer2_out[3942] ^ layer2_out[3943];
     layer3_out[5664] <= ~(layer2_out[6181] | layer2_out[6182]);
     layer3_out[5665] <= layer2_out[600] & layer2_out[601];
     layer3_out[5666] <= ~(layer2_out[1648] ^ layer2_out[1649]);
     layer3_out[5667] <= ~layer2_out[6176];
     layer3_out[5668] <= ~(layer2_out[11330] ^ layer2_out[11331]);
     layer3_out[5669] <= ~layer2_out[7589] | layer2_out[7588];
     layer3_out[5670] <= layer2_out[8925] & ~layer2_out[8926];
     layer3_out[5671] <= ~(layer2_out[3423] | layer2_out[3424]);
     layer3_out[5672] <= layer2_out[6768] & ~layer2_out[6767];
     layer3_out[5673] <= layer2_out[2385];
     layer3_out[5674] <= ~layer2_out[9779];
     layer3_out[5675] <= layer2_out[8553];
     layer3_out[5676] <= layer2_out[10375] & ~layer2_out[10374];
     layer3_out[5677] <= layer2_out[11515];
     layer3_out[5678] <= ~(layer2_out[8190] | layer2_out[8191]);
     layer3_out[5679] <= ~layer2_out[9128];
     layer3_out[5680] <= layer2_out[1334] ^ layer2_out[1335];
     layer3_out[5681] <= ~(layer2_out[11141] ^ layer2_out[11142]);
     layer3_out[5682] <= layer2_out[10968] ^ layer2_out[10969];
     layer3_out[5683] <= ~(layer2_out[11841] ^ layer2_out[11842]);
     layer3_out[5684] <= layer2_out[9888] & layer2_out[9889];
     layer3_out[5685] <= ~layer2_out[8812];
     layer3_out[5686] <= layer2_out[8522] & ~layer2_out[8523];
     layer3_out[5687] <= ~(layer2_out[141] | layer2_out[142]);
     layer3_out[5688] <= ~(layer2_out[11827] | layer2_out[11828]);
     layer3_out[5689] <= layer2_out[7044] ^ layer2_out[7045];
     layer3_out[5690] <= ~layer2_out[8604];
     layer3_out[5691] <= ~layer2_out[7572] | layer2_out[7573];
     layer3_out[5692] <= layer2_out[1041] & ~layer2_out[1042];
     layer3_out[5693] <= ~(layer2_out[613] | layer2_out[614]);
     layer3_out[5694] <= layer2_out[10239];
     layer3_out[5695] <= layer2_out[1838];
     layer3_out[5696] <= ~layer2_out[1827];
     layer3_out[5697] <= ~(layer2_out[7920] | layer2_out[7921]);
     layer3_out[5698] <= layer2_out[11928];
     layer3_out[5699] <= ~(layer2_out[9869] ^ layer2_out[9870]);
     layer3_out[5700] <= layer2_out[1871];
     layer3_out[5701] <= layer2_out[6917] & ~layer2_out[6916];
     layer3_out[5702] <= layer2_out[887] ^ layer2_out[888];
     layer3_out[5703] <= layer2_out[10553] & ~layer2_out[10554];
     layer3_out[5704] <= layer2_out[1321] & ~layer2_out[1322];
     layer3_out[5705] <= ~layer2_out[5901];
     layer3_out[5706] <= ~layer2_out[10283];
     layer3_out[5707] <= layer2_out[2507] & layer2_out[2508];
     layer3_out[5708] <= ~layer2_out[4094] | layer2_out[4093];
     layer3_out[5709] <= layer2_out[5942];
     layer3_out[5710] <= ~layer2_out[4852];
     layer3_out[5711] <= layer2_out[9781];
     layer3_out[5712] <= layer2_out[3442] & ~layer2_out[3441];
     layer3_out[5713] <= layer2_out[1982] & layer2_out[1983];
     layer3_out[5714] <= layer2_out[4779];
     layer3_out[5715] <= ~(layer2_out[4456] & layer2_out[4457]);
     layer3_out[5716] <= ~layer2_out[1271];
     layer3_out[5717] <= layer2_out[636] & ~layer2_out[637];
     layer3_out[5718] <= layer2_out[6990] & layer2_out[6991];
     layer3_out[5719] <= layer2_out[8740];
     layer3_out[5720] <= ~(layer2_out[10401] ^ layer2_out[10402]);
     layer3_out[5721] <= layer2_out[10567] & ~layer2_out[10566];
     layer3_out[5722] <= layer2_out[51] & layer2_out[52];
     layer3_out[5723] <= layer2_out[10842] ^ layer2_out[10843];
     layer3_out[5724] <= ~(layer2_out[6014] ^ layer2_out[6015]);
     layer3_out[5725] <= ~(layer2_out[159] ^ layer2_out[160]);
     layer3_out[5726] <= ~layer2_out[7762];
     layer3_out[5727] <= layer2_out[317];
     layer3_out[5728] <= layer2_out[11268];
     layer3_out[5729] <= layer2_out[9593] ^ layer2_out[9594];
     layer3_out[5730] <= ~layer2_out[2064];
     layer3_out[5731] <= layer2_out[10691] | layer2_out[10692];
     layer3_out[5732] <= layer2_out[6530] & ~layer2_out[6529];
     layer3_out[5733] <= layer2_out[11936];
     layer3_out[5734] <= layer2_out[5779] & layer2_out[5780];
     layer3_out[5735] <= layer2_out[6549];
     layer3_out[5736] <= ~(layer2_out[7195] | layer2_out[7196]);
     layer3_out[5737] <= ~layer2_out[9401];
     layer3_out[5738] <= ~layer2_out[2802];
     layer3_out[5739] <= ~(layer2_out[7793] ^ layer2_out[7794]);
     layer3_out[5740] <= ~layer2_out[5579];
     layer3_out[5741] <= layer2_out[4674];
     layer3_out[5742] <= layer2_out[11442] & layer2_out[11443];
     layer3_out[5743] <= layer2_out[2395] & ~layer2_out[2396];
     layer3_out[5744] <= layer2_out[1933];
     layer3_out[5745] <= ~(layer2_out[6075] ^ layer2_out[6076]);
     layer3_out[5746] <= ~layer2_out[5670] | layer2_out[5671];
     layer3_out[5747] <= ~(layer2_out[1737] | layer2_out[1738]);
     layer3_out[5748] <= ~(layer2_out[8450] | layer2_out[8451]);
     layer3_out[5749] <= layer2_out[7994] & ~layer2_out[7993];
     layer3_out[5750] <= layer2_out[4789] ^ layer2_out[4790];
     layer3_out[5751] <= layer2_out[6816] & ~layer2_out[6817];
     layer3_out[5752] <= layer2_out[10195] & ~layer2_out[10194];
     layer3_out[5753] <= ~(layer2_out[8328] ^ layer2_out[8329]);
     layer3_out[5754] <= layer2_out[1578] & ~layer2_out[1577];
     layer3_out[5755] <= layer2_out[17] & ~layer2_out[16];
     layer3_out[5756] <= layer2_out[1048] & ~layer2_out[1049];
     layer3_out[5757] <= ~(layer2_out[1531] ^ layer2_out[1532]);
     layer3_out[5758] <= layer2_out[3375] & layer2_out[3376];
     layer3_out[5759] <= ~(layer2_out[7046] | layer2_out[7047]);
     layer3_out[5760] <= layer2_out[5458];
     layer3_out[5761] <= ~(layer2_out[5355] ^ layer2_out[5356]);
     layer3_out[5762] <= layer2_out[9546];
     layer3_out[5763] <= layer2_out[11021];
     layer3_out[5764] <= ~layer2_out[2381];
     layer3_out[5765] <= ~layer2_out[9004] | layer2_out[9003];
     layer3_out[5766] <= layer2_out[7835] & ~layer2_out[7834];
     layer3_out[5767] <= ~(layer2_out[6233] | layer2_out[6234]);
     layer3_out[5768] <= layer2_out[5762] & ~layer2_out[5761];
     layer3_out[5769] <= layer2_out[3720] & ~layer2_out[3719];
     layer3_out[5770] <= layer2_out[9347] & layer2_out[9348];
     layer3_out[5771] <= ~(layer2_out[6789] ^ layer2_out[6790]);
     layer3_out[5772] <= layer2_out[305] & ~layer2_out[306];
     layer3_out[5773] <= ~layer2_out[7768];
     layer3_out[5774] <= layer2_out[7266] ^ layer2_out[7267];
     layer3_out[5775] <= ~layer2_out[9247];
     layer3_out[5776] <= layer2_out[9293];
     layer3_out[5777] <= layer2_out[3263];
     layer3_out[5778] <= layer2_out[1482] & ~layer2_out[1481];
     layer3_out[5779] <= layer2_out[7329];
     layer3_out[5780] <= layer2_out[5647] & layer2_out[5648];
     layer3_out[5781] <= ~(layer2_out[6865] | layer2_out[6866]);
     layer3_out[5782] <= ~layer2_out[2493];
     layer3_out[5783] <= layer2_out[4356];
     layer3_out[5784] <= ~layer2_out[3086];
     layer3_out[5785] <= layer2_out[7940];
     layer3_out[5786] <= layer2_out[6982] & ~layer2_out[6981];
     layer3_out[5787] <= layer2_out[1761];
     layer3_out[5788] <= layer2_out[5162] | layer2_out[5163];
     layer3_out[5789] <= ~layer2_out[7767];
     layer3_out[5790] <= layer2_out[8975];
     layer3_out[5791] <= layer2_out[2393] & layer2_out[2394];
     layer3_out[5792] <= layer2_out[6273] & layer2_out[6274];
     layer3_out[5793] <= layer2_out[2290] & ~layer2_out[2291];
     layer3_out[5794] <= ~(layer2_out[9147] | layer2_out[9148]);
     layer3_out[5795] <= layer2_out[3782];
     layer3_out[5796] <= ~layer2_out[2888];
     layer3_out[5797] <= layer2_out[6523] & ~layer2_out[6522];
     layer3_out[5798] <= ~layer2_out[5967];
     layer3_out[5799] <= ~(layer2_out[5169] | layer2_out[5170]);
     layer3_out[5800] <= ~(layer2_out[10193] | layer2_out[10194]);
     layer3_out[5801] <= ~layer2_out[5939] | layer2_out[5938];
     layer3_out[5802] <= ~(layer2_out[1842] | layer2_out[1843]);
     layer3_out[5803] <= layer2_out[5558];
     layer3_out[5804] <= ~(layer2_out[8797] | layer2_out[8798]);
     layer3_out[5805] <= ~(layer2_out[597] ^ layer2_out[598]);
     layer3_out[5806] <= layer2_out[1032] & ~layer2_out[1031];
     layer3_out[5807] <= ~(layer2_out[6079] | layer2_out[6080]);
     layer3_out[5808] <= layer2_out[1065] & ~layer2_out[1066];
     layer3_out[5809] <= ~layer2_out[3564];
     layer3_out[5810] <= layer2_out[4823];
     layer3_out[5811] <= layer2_out[2542] & ~layer2_out[2543];
     layer3_out[5812] <= ~layer2_out[11193];
     layer3_out[5813] <= ~(layer2_out[5422] | layer2_out[5423]);
     layer3_out[5814] <= layer2_out[10135] & layer2_out[10136];
     layer3_out[5815] <= layer2_out[10324];
     layer3_out[5816] <= layer2_out[6471];
     layer3_out[5817] <= ~layer2_out[6689] | layer2_out[6688];
     layer3_out[5818] <= layer2_out[2217];
     layer3_out[5819] <= ~layer2_out[8782];
     layer3_out[5820] <= layer2_out[1702] & ~layer2_out[1703];
     layer3_out[5821] <= ~layer2_out[706];
     layer3_out[5822] <= layer2_out[7079] & ~layer2_out[7080];
     layer3_out[5823] <= ~layer2_out[9839];
     layer3_out[5824] <= ~(layer2_out[10452] ^ layer2_out[10453]);
     layer3_out[5825] <= layer2_out[10579] & ~layer2_out[10580];
     layer3_out[5826] <= layer2_out[3245];
     layer3_out[5827] <= layer2_out[10418];
     layer3_out[5828] <= layer2_out[6607] & layer2_out[6608];
     layer3_out[5829] <= layer2_out[1267] & ~layer2_out[1268];
     layer3_out[5830] <= layer2_out[5393] ^ layer2_out[5394];
     layer3_out[5831] <= layer2_out[2994];
     layer3_out[5832] <= layer2_out[2229] ^ layer2_out[2230];
     layer3_out[5833] <= layer2_out[3149] | layer2_out[3150];
     layer3_out[5834] <= ~(layer2_out[6221] & layer2_out[6222]);
     layer3_out[5835] <= layer2_out[3016] & ~layer2_out[3015];
     layer3_out[5836] <= layer2_out[10264] & layer2_out[10265];
     layer3_out[5837] <= layer2_out[6657] & ~layer2_out[6656];
     layer3_out[5838] <= layer2_out[9829] & layer2_out[9830];
     layer3_out[5839] <= layer2_out[242] & ~layer2_out[241];
     layer3_out[5840] <= layer2_out[2079] & ~layer2_out[2078];
     layer3_out[5841] <= ~(layer2_out[10232] ^ layer2_out[10233]);
     layer3_out[5842] <= ~(layer2_out[8651] ^ layer2_out[8652]);
     layer3_out[5843] <= ~layer2_out[1579];
     layer3_out[5844] <= ~layer2_out[4814] | layer2_out[4813];
     layer3_out[5845] <= layer2_out[10334] & ~layer2_out[10335];
     layer3_out[5846] <= layer2_out[9966] & ~layer2_out[9965];
     layer3_out[5847] <= layer2_out[5306];
     layer3_out[5848] <= layer2_out[41] & layer2_out[42];
     layer3_out[5849] <= ~layer2_out[10278];
     layer3_out[5850] <= layer2_out[6964] & layer2_out[6965];
     layer3_out[5851] <= layer2_out[4344] ^ layer2_out[4345];
     layer3_out[5852] <= layer2_out[10829] ^ layer2_out[10830];
     layer3_out[5853] <= layer2_out[5259] & ~layer2_out[5258];
     layer3_out[5854] <= layer2_out[472] & layer2_out[473];
     layer3_out[5855] <= ~(layer2_out[900] ^ layer2_out[901]);
     layer3_out[5856] <= layer2_out[2787];
     layer3_out[5857] <= ~(layer2_out[11558] | layer2_out[11559]);
     layer3_out[5858] <= ~layer2_out[291];
     layer3_out[5859] <= layer2_out[9666] & ~layer2_out[9667];
     layer3_out[5860] <= ~layer2_out[2536];
     layer3_out[5861] <= layer2_out[4444] & ~layer2_out[4445];
     layer3_out[5862] <= ~layer2_out[10994];
     layer3_out[5863] <= ~(layer2_out[8305] ^ layer2_out[8306]);
     layer3_out[5864] <= layer2_out[4587] & ~layer2_out[4588];
     layer3_out[5865] <= ~layer2_out[11388];
     layer3_out[5866] <= ~(layer2_out[4768] | layer2_out[4769]);
     layer3_out[5867] <= layer2_out[9581] & ~layer2_out[9582];
     layer3_out[5868] <= ~layer2_out[3124];
     layer3_out[5869] <= layer2_out[3299];
     layer3_out[5870] <= layer2_out[6602] & layer2_out[6603];
     layer3_out[5871] <= ~(layer2_out[5374] ^ layer2_out[5375]);
     layer3_out[5872] <= ~(layer2_out[6555] & layer2_out[6556]);
     layer3_out[5873] <= ~layer2_out[8455];
     layer3_out[5874] <= ~layer2_out[2443];
     layer3_out[5875] <= layer2_out[5948] & layer2_out[5949];
     layer3_out[5876] <= ~layer2_out[2424];
     layer3_out[5877] <= layer2_out[11334] & ~layer2_out[11335];
     layer3_out[5878] <= layer2_out[9467] & ~layer2_out[9466];
     layer3_out[5879] <= ~layer2_out[10670];
     layer3_out[5880] <= layer2_out[6642] ^ layer2_out[6643];
     layer3_out[5881] <= layer2_out[5894] & ~layer2_out[5895];
     layer3_out[5882] <= layer2_out[1637] & ~layer2_out[1638];
     layer3_out[5883] <= ~layer2_out[9308];
     layer3_out[5884] <= ~(layer2_out[1827] | layer2_out[1828]);
     layer3_out[5885] <= layer2_out[2284] ^ layer2_out[2285];
     layer3_out[5886] <= ~layer2_out[1553];
     layer3_out[5887] <= layer2_out[9599] & ~layer2_out[9600];
     layer3_out[5888] <= ~(layer2_out[3548] & layer2_out[3549]);
     layer3_out[5889] <= ~layer2_out[3944] | layer2_out[3943];
     layer3_out[5890] <= layer2_out[2706] & ~layer2_out[2705];
     layer3_out[5891] <= ~(layer2_out[8959] ^ layer2_out[8960]);
     layer3_out[5892] <= ~(layer2_out[9919] ^ layer2_out[9920]);
     layer3_out[5893] <= layer2_out[10057];
     layer3_out[5894] <= layer2_out[5746];
     layer3_out[5895] <= ~layer2_out[10103];
     layer3_out[5896] <= ~(layer2_out[10435] | layer2_out[10436]);
     layer3_out[5897] <= ~layer2_out[9573];
     layer3_out[5898] <= ~layer2_out[3567];
     layer3_out[5899] <= layer2_out[4364] & ~layer2_out[4365];
     layer3_out[5900] <= layer2_out[11251];
     layer3_out[5901] <= layer2_out[144] & ~layer2_out[145];
     layer3_out[5902] <= layer2_out[4434];
     layer3_out[5903] <= ~layer2_out[9263];
     layer3_out[5904] <= layer2_out[372] & ~layer2_out[373];
     layer3_out[5905] <= layer2_out[4224] ^ layer2_out[4225];
     layer3_out[5906] <= layer2_out[5454];
     layer3_out[5907] <= layer2_out[8113] ^ layer2_out[8114];
     layer3_out[5908] <= ~(layer2_out[8160] | layer2_out[8161]);
     layer3_out[5909] <= ~layer2_out[7373];
     layer3_out[5910] <= ~(layer2_out[10373] | layer2_out[10374]);
     layer3_out[5911] <= layer2_out[9396] & layer2_out[9397];
     layer3_out[5912] <= ~layer2_out[5389];
     layer3_out[5913] <= ~(layer2_out[4087] & layer2_out[4088]);
     layer3_out[5914] <= layer2_out[7564] & layer2_out[7565];
     layer3_out[5915] <= ~layer2_out[1028];
     layer3_out[5916] <= ~layer2_out[3255];
     layer3_out[5917] <= layer2_out[787] & layer2_out[788];
     layer3_out[5918] <= ~(layer2_out[10763] | layer2_out[10764]);
     layer3_out[5919] <= layer2_out[8202] & layer2_out[8203];
     layer3_out[5920] <= layer2_out[5054] & ~layer2_out[5053];
     layer3_out[5921] <= layer2_out[2418] | layer2_out[2419];
     layer3_out[5922] <= layer2_out[4518] ^ layer2_out[4519];
     layer3_out[5923] <= ~(layer2_out[6179] & layer2_out[6180]);
     layer3_out[5924] <= ~(layer2_out[10063] | layer2_out[10064]);
     layer3_out[5925] <= layer2_out[7831] & ~layer2_out[7832];
     layer3_out[5926] <= ~(layer2_out[7872] ^ layer2_out[7873]);
     layer3_out[5927] <= ~(layer2_out[263] | layer2_out[264]);
     layer3_out[5928] <= layer2_out[8786] & ~layer2_out[8785];
     layer3_out[5929] <= layer2_out[9038] | layer2_out[9039];
     layer3_out[5930] <= layer2_out[9486];
     layer3_out[5931] <= ~layer2_out[1284] | layer2_out[1285];
     layer3_out[5932] <= ~(layer2_out[5070] ^ layer2_out[5071]);
     layer3_out[5933] <= ~(layer2_out[3797] ^ layer2_out[3798]);
     layer3_out[5934] <= layer2_out[9425];
     layer3_out[5935] <= layer2_out[9678] & layer2_out[9679];
     layer3_out[5936] <= ~(layer2_out[8524] | layer2_out[8525]);
     layer3_out[5937] <= ~layer2_out[5478];
     layer3_out[5938] <= layer2_out[7533] & ~layer2_out[7534];
     layer3_out[5939] <= ~(layer2_out[5133] | layer2_out[5134]);
     layer3_out[5940] <= layer2_out[2596] ^ layer2_out[2597];
     layer3_out[5941] <= layer2_out[10013] & layer2_out[10014];
     layer3_out[5942] <= layer2_out[3319] & ~layer2_out[3318];
     layer3_out[5943] <= ~layer2_out[11407];
     layer3_out[5944] <= ~layer2_out[3969];
     layer3_out[5945] <= ~layer2_out[2743] | layer2_out[2744];
     layer3_out[5946] <= layer2_out[1560] & layer2_out[1561];
     layer3_out[5947] <= ~layer2_out[250] | layer2_out[251];
     layer3_out[5948] <= layer2_out[8079] & layer2_out[8080];
     layer3_out[5949] <= ~(layer2_out[6962] | layer2_out[6963]);
     layer3_out[5950] <= ~layer2_out[7195];
     layer3_out[5951] <= ~(layer2_out[9461] ^ layer2_out[9462]);
     layer3_out[5952] <= layer2_out[10337] & ~layer2_out[10338];
     layer3_out[5953] <= ~layer2_out[11325];
     layer3_out[5954] <= ~layer2_out[10675];
     layer3_out[5955] <= ~(layer2_out[2642] | layer2_out[2643]);
     layer3_out[5956] <= ~layer2_out[9906];
     layer3_out[5957] <= ~layer2_out[9361] | layer2_out[9362];
     layer3_out[5958] <= layer2_out[11790] & layer2_out[11791];
     layer3_out[5959] <= ~(layer2_out[10922] ^ layer2_out[10923]);
     layer3_out[5960] <= layer2_out[5580] ^ layer2_out[5581];
     layer3_out[5961] <= layer2_out[1363] & ~layer2_out[1364];
     layer3_out[5962] <= ~(layer2_out[10367] | layer2_out[10368]);
     layer3_out[5963] <= layer2_out[7615];
     layer3_out[5964] <= ~(layer2_out[1098] & layer2_out[1099]);
     layer3_out[5965] <= layer2_out[2187] ^ layer2_out[2188];
     layer3_out[5966] <= ~layer2_out[4305];
     layer3_out[5967] <= layer2_out[10147];
     layer3_out[5968] <= layer2_out[10020];
     layer3_out[5969] <= ~(layer2_out[11610] | layer2_out[11611]);
     layer3_out[5970] <= layer2_out[1206] & ~layer2_out[1207];
     layer3_out[5971] <= ~(layer2_out[11228] & layer2_out[11229]);
     layer3_out[5972] <= layer2_out[7384];
     layer3_out[5973] <= ~layer2_out[5665];
     layer3_out[5974] <= layer2_out[6413] & layer2_out[6414];
     layer3_out[5975] <= ~layer2_out[2996];
     layer3_out[5976] <= layer2_out[9507];
     layer3_out[5977] <= layer2_out[9837] & layer2_out[9838];
     layer3_out[5978] <= ~layer2_out[10822];
     layer3_out[5979] <= ~layer2_out[4368];
     layer3_out[5980] <= layer2_out[8617] ^ layer2_out[8618];
     layer3_out[5981] <= ~layer2_out[8976];
     layer3_out[5982] <= layer2_out[9888];
     layer3_out[5983] <= ~layer2_out[11884];
     layer3_out[5984] <= ~layer2_out[9951];
     layer3_out[5985] <= layer2_out[11874];
     layer3_out[5986] <= 1'b0;
     layer3_out[5987] <= ~layer2_out[6042];
     layer3_out[5988] <= ~(layer2_out[11531] ^ layer2_out[11532]);
     layer3_out[5989] <= layer2_out[9158] & layer2_out[9159];
     layer3_out[5990] <= layer2_out[3691];
     layer3_out[5991] <= ~layer2_out[415];
     layer3_out[5992] <= layer2_out[11469];
     layer3_out[5993] <= ~(layer2_out[2289] ^ layer2_out[2290]);
     layer3_out[5994] <= ~layer2_out[9815];
     layer3_out[5995] <= layer2_out[2006] & ~layer2_out[2005];
     layer3_out[5996] <= ~layer2_out[4967];
     layer3_out[5997] <= layer2_out[6386] ^ layer2_out[6387];
     layer3_out[5998] <= layer2_out[3300] | layer2_out[3301];
     layer3_out[5999] <= layer2_out[920] & layer2_out[921];
     layer3_out[6000] <= ~(layer2_out[648] & layer2_out[649]);
     layer3_out[6001] <= ~(layer2_out[9542] ^ layer2_out[9543]);
     layer3_out[6002] <= layer2_out[7968] & layer2_out[7969];
     layer3_out[6003] <= layer2_out[9642] & ~layer2_out[9641];
     layer3_out[6004] <= ~layer2_out[2450];
     layer3_out[6005] <= layer2_out[7818] ^ layer2_out[7819];
     layer3_out[6006] <= ~layer2_out[2446];
     layer3_out[6007] <= ~layer2_out[2760];
     layer3_out[6008] <= ~layer2_out[3236];
     layer3_out[6009] <= layer2_out[8238] & layer2_out[8239];
     layer3_out[6010] <= ~layer2_out[5326];
     layer3_out[6011] <= ~layer2_out[7813] | layer2_out[7812];
     layer3_out[6012] <= layer2_out[9871];
     layer3_out[6013] <= ~layer2_out[4677] | layer2_out[4676];
     layer3_out[6014] <= ~layer2_out[11248];
     layer3_out[6015] <= layer2_out[7711];
     layer3_out[6016] <= layer2_out[11100];
     layer3_out[6017] <= ~layer2_out[7358];
     layer3_out[6018] <= ~(layer2_out[11105] & layer2_out[11106]);
     layer3_out[6019] <= layer2_out[6330];
     layer3_out[6020] <= ~layer2_out[6958];
     layer3_out[6021] <= layer2_out[7600] ^ layer2_out[7601];
     layer3_out[6022] <= ~(layer2_out[6911] & layer2_out[6912]);
     layer3_out[6023] <= ~(layer2_out[11637] & layer2_out[11638]);
     layer3_out[6024] <= ~layer2_out[19] | layer2_out[20];
     layer3_out[6025] <= layer2_out[9289];
     layer3_out[6026] <= layer2_out[5006] & layer2_out[5007];
     layer3_out[6027] <= ~layer2_out[3298] | layer2_out[3297];
     layer3_out[6028] <= ~(layer2_out[6541] ^ layer2_out[6542]);
     layer3_out[6029] <= layer2_out[313] & ~layer2_out[312];
     layer3_out[6030] <= layer2_out[6741];
     layer3_out[6031] <= ~(layer2_out[11277] ^ layer2_out[11278]);
     layer3_out[6032] <= layer2_out[1708] | layer2_out[1709];
     layer3_out[6033] <= ~layer2_out[10617];
     layer3_out[6034] <= layer2_out[11071] & ~layer2_out[11072];
     layer3_out[6035] <= layer2_out[3669];
     layer3_out[6036] <= layer2_out[7308] & ~layer2_out[7309];
     layer3_out[6037] <= ~(layer2_out[10771] ^ layer2_out[10772]);
     layer3_out[6038] <= ~layer2_out[10329] | layer2_out[10330];
     layer3_out[6039] <= layer2_out[5969] & ~layer2_out[5970];
     layer3_out[6040] <= layer2_out[8408] & ~layer2_out[8407];
     layer3_out[6041] <= layer2_out[3804] ^ layer2_out[3805];
     layer3_out[6042] <= layer2_out[1005];
     layer3_out[6043] <= ~layer2_out[7332] | layer2_out[7333];
     layer3_out[6044] <= ~layer2_out[3070];
     layer3_out[6045] <= layer2_out[10481] & layer2_out[10482];
     layer3_out[6046] <= ~layer2_out[1749];
     layer3_out[6047] <= layer2_out[11191];
     layer3_out[6048] <= ~(layer2_out[1806] ^ layer2_out[1807]);
     layer3_out[6049] <= layer2_out[9293] & ~layer2_out[9292];
     layer3_out[6050] <= layer2_out[11309];
     layer3_out[6051] <= ~layer2_out[8180];
     layer3_out[6052] <= layer2_out[5316];
     layer3_out[6053] <= layer2_out[5080];
     layer3_out[6054] <= layer2_out[1410] ^ layer2_out[1411];
     layer3_out[6055] <= ~layer2_out[8470];
     layer3_out[6056] <= ~(layer2_out[734] ^ layer2_out[735]);
     layer3_out[6057] <= ~layer2_out[1975] | layer2_out[1976];
     layer3_out[6058] <= ~layer2_out[2466] | layer2_out[2467];
     layer3_out[6059] <= layer2_out[655] & ~layer2_out[656];
     layer3_out[6060] <= ~(layer2_out[1510] | layer2_out[1511]);
     layer3_out[6061] <= ~(layer2_out[10653] ^ layer2_out[10654]);
     layer3_out[6062] <= ~(layer2_out[4486] ^ layer2_out[4487]);
     layer3_out[6063] <= ~(layer2_out[11604] ^ layer2_out[11605]);
     layer3_out[6064] <= layer2_out[827] & ~layer2_out[828];
     layer3_out[6065] <= layer2_out[409] ^ layer2_out[410];
     layer3_out[6066] <= layer2_out[7329] & ~layer2_out[7328];
     layer3_out[6067] <= ~(layer2_out[3582] & layer2_out[3583]);
     layer3_out[6068] <= layer2_out[7743];
     layer3_out[6069] <= layer2_out[3271];
     layer3_out[6070] <= ~(layer2_out[10307] & layer2_out[10308]);
     layer3_out[6071] <= ~layer2_out[697];
     layer3_out[6072] <= layer2_out[6739] & layer2_out[6740];
     layer3_out[6073] <= layer2_out[987];
     layer3_out[6074] <= ~layer2_out[6922];
     layer3_out[6075] <= ~(layer2_out[10836] | layer2_out[10837]);
     layer3_out[6076] <= layer2_out[11407] ^ layer2_out[11408];
     layer3_out[6077] <= layer2_out[944];
     layer3_out[6078] <= ~layer2_out[3696] | layer2_out[3697];
     layer3_out[6079] <= ~(layer2_out[7416] ^ layer2_out[7417]);
     layer3_out[6080] <= layer2_out[9542];
     layer3_out[6081] <= layer2_out[3114];
     layer3_out[6082] <= ~layer2_out[8711];
     layer3_out[6083] <= ~(layer2_out[1752] ^ layer2_out[1753]);
     layer3_out[6084] <= ~layer2_out[10914];
     layer3_out[6085] <= ~(layer2_out[11650] ^ layer2_out[11651]);
     layer3_out[6086] <= layer2_out[665] & layer2_out[666];
     layer3_out[6087] <= ~layer2_out[4874];
     layer3_out[6088] <= layer2_out[5889] ^ layer2_out[5890];
     layer3_out[6089] <= ~layer2_out[5133];
     layer3_out[6090] <= ~(layer2_out[3277] ^ layer2_out[3278]);
     layer3_out[6091] <= ~layer2_out[1368];
     layer3_out[6092] <= ~layer2_out[7160];
     layer3_out[6093] <= layer2_out[1866];
     layer3_out[6094] <= ~(layer2_out[2341] ^ layer2_out[2342]);
     layer3_out[6095] <= layer2_out[7825] ^ layer2_out[7826];
     layer3_out[6096] <= layer2_out[3951] ^ layer2_out[3952];
     layer3_out[6097] <= ~layer2_out[1041];
     layer3_out[6098] <= ~(layer2_out[836] ^ layer2_out[837]);
     layer3_out[6099] <= ~layer2_out[9422];
     layer3_out[6100] <= layer2_out[5419] & ~layer2_out[5420];
     layer3_out[6101] <= ~layer2_out[5008] | layer2_out[5007];
     layer3_out[6102] <= layer2_out[4959] ^ layer2_out[4960];
     layer3_out[6103] <= ~layer2_out[3843] | layer2_out[3842];
     layer3_out[6104] <= layer2_out[6640];
     layer3_out[6105] <= ~(layer2_out[7441] & layer2_out[7442]);
     layer3_out[6106] <= ~layer2_out[10322];
     layer3_out[6107] <= layer2_out[8125];
     layer3_out[6108] <= layer2_out[1788] & layer2_out[1789];
     layer3_out[6109] <= ~layer2_out[11895] | layer2_out[11894];
     layer3_out[6110] <= layer2_out[245];
     layer3_out[6111] <= layer2_out[882];
     layer3_out[6112] <= ~(layer2_out[9503] ^ layer2_out[9504]);
     layer3_out[6113] <= layer2_out[44];
     layer3_out[6114] <= ~layer2_out[1232] | layer2_out[1233];
     layer3_out[6115] <= ~layer2_out[6196];
     layer3_out[6116] <= layer2_out[1340] & ~layer2_out[1339];
     layer3_out[6117] <= ~layer2_out[4003];
     layer3_out[6118] <= layer2_out[4173] ^ layer2_out[4174];
     layer3_out[6119] <= ~layer2_out[33];
     layer3_out[6120] <= ~(layer2_out[5700] | layer2_out[5701]);
     layer3_out[6121] <= ~layer2_out[2907];
     layer3_out[6122] <= layer2_out[4680];
     layer3_out[6123] <= ~layer2_out[7677] | layer2_out[7676];
     layer3_out[6124] <= layer2_out[6952];
     layer3_out[6125] <= layer2_out[422] ^ layer2_out[423];
     layer3_out[6126] <= ~(layer2_out[2173] ^ layer2_out[2174]);
     layer3_out[6127] <= ~layer2_out[1513] | layer2_out[1514];
     layer3_out[6128] <= layer2_out[572] ^ layer2_out[573];
     layer3_out[6129] <= ~(layer2_out[6942] ^ layer2_out[6943]);
     layer3_out[6130] <= layer2_out[11494] | layer2_out[11495];
     layer3_out[6131] <= ~(layer2_out[3829] ^ layer2_out[3830]);
     layer3_out[6132] <= ~layer2_out[4012];
     layer3_out[6133] <= layer2_out[9481] ^ layer2_out[9482];
     layer3_out[6134] <= layer2_out[7325] & layer2_out[7326];
     layer3_out[6135] <= ~layer2_out[1317];
     layer3_out[6136] <= ~(layer2_out[8117] ^ layer2_out[8118]);
     layer3_out[6137] <= layer2_out[4038] ^ layer2_out[4039];
     layer3_out[6138] <= ~(layer2_out[10542] & layer2_out[10543]);
     layer3_out[6139] <= ~(layer2_out[2371] & layer2_out[2372]);
     layer3_out[6140] <= layer2_out[5891] ^ layer2_out[5892];
     layer3_out[6141] <= ~(layer2_out[4892] | layer2_out[4893]);
     layer3_out[6142] <= layer2_out[9549] & ~layer2_out[9548];
     layer3_out[6143] <= ~layer2_out[4012];
     layer3_out[6144] <= ~layer2_out[3230] | layer2_out[3231];
     layer3_out[6145] <= ~layer2_out[8822];
     layer3_out[6146] <= layer2_out[1561] & layer2_out[1562];
     layer3_out[6147] <= ~(layer2_out[6222] & layer2_out[6223]);
     layer3_out[6148] <= ~(layer2_out[7439] & layer2_out[7440]);
     layer3_out[6149] <= layer2_out[1864] | layer2_out[1865];
     layer3_out[6150] <= layer2_out[5599];
     layer3_out[6151] <= layer2_out[4019];
     layer3_out[6152] <= ~layer2_out[5624] | layer2_out[5623];
     layer3_out[6153] <= layer2_out[711] ^ layer2_out[712];
     layer3_out[6154] <= ~layer2_out[6484];
     layer3_out[6155] <= layer2_out[1154] & ~layer2_out[1155];
     layer3_out[6156] <= ~layer2_out[1199];
     layer3_out[6157] <= ~layer2_out[11728];
     layer3_out[6158] <= layer2_out[11495] ^ layer2_out[11496];
     layer3_out[6159] <= layer2_out[11301] & layer2_out[11302];
     layer3_out[6160] <= layer2_out[11339] ^ layer2_out[11340];
     layer3_out[6161] <= ~layer2_out[3200];
     layer3_out[6162] <= ~layer2_out[10961];
     layer3_out[6163] <= ~layer2_out[1365];
     layer3_out[6164] <= layer2_out[4145] ^ layer2_out[4146];
     layer3_out[6165] <= layer2_out[2890] & layer2_out[2891];
     layer3_out[6166] <= ~(layer2_out[7302] ^ layer2_out[7303]);
     layer3_out[6167] <= ~layer2_out[5963];
     layer3_out[6168] <= ~layer2_out[6852];
     layer3_out[6169] <= layer2_out[933] & ~layer2_out[932];
     layer3_out[6170] <= layer2_out[5708];
     layer3_out[6171] <= layer2_out[4057];
     layer3_out[6172] <= layer2_out[8296] | layer2_out[8297];
     layer3_out[6173] <= ~layer2_out[4149];
     layer3_out[6174] <= layer2_out[460];
     layer3_out[6175] <= ~(layer2_out[9847] | layer2_out[9848]);
     layer3_out[6176] <= layer2_out[7043] & layer2_out[7044];
     layer3_out[6177] <= layer2_out[11788] ^ layer2_out[11789];
     layer3_out[6178] <= ~(layer2_out[3538] | layer2_out[3539]);
     layer3_out[6179] <= layer2_out[2196];
     layer3_out[6180] <= layer2_out[2566];
     layer3_out[6181] <= layer2_out[3669] ^ layer2_out[3670];
     layer3_out[6182] <= ~layer2_out[10279] | layer2_out[10280];
     layer3_out[6183] <= ~layer2_out[8803];
     layer3_out[6184] <= layer2_out[5689];
     layer3_out[6185] <= ~(layer2_out[5903] | layer2_out[5904]);
     layer3_out[6186] <= layer2_out[1109];
     layer3_out[6187] <= ~layer2_out[10163] | layer2_out[10162];
     layer3_out[6188] <= layer2_out[11136] & ~layer2_out[11137];
     layer3_out[6189] <= ~layer2_out[6391] | layer2_out[6392];
     layer3_out[6190] <= layer2_out[5640];
     layer3_out[6191] <= layer2_out[10014] & layer2_out[10015];
     layer3_out[6192] <= layer2_out[2555] & layer2_out[2556];
     layer3_out[6193] <= ~(layer2_out[1023] ^ layer2_out[1024]);
     layer3_out[6194] <= ~layer2_out[2865];
     layer3_out[6195] <= layer2_out[5215];
     layer3_out[6196] <= ~layer2_out[9213];
     layer3_out[6197] <= layer2_out[2599];
     layer3_out[6198] <= layer2_out[4690] & ~layer2_out[4691];
     layer3_out[6199] <= layer2_out[5545];
     layer3_out[6200] <= ~layer2_out[3548] | layer2_out[3547];
     layer3_out[6201] <= layer2_out[627];
     layer3_out[6202] <= layer2_out[11661] ^ layer2_out[11662];
     layer3_out[6203] <= layer2_out[10952];
     layer3_out[6204] <= ~(layer2_out[338] ^ layer2_out[339]);
     layer3_out[6205] <= layer2_out[7333] & layer2_out[7334];
     layer3_out[6206] <= layer2_out[625];
     layer3_out[6207] <= layer2_out[1958] | layer2_out[1959];
     layer3_out[6208] <= ~layer2_out[5148];
     layer3_out[6209] <= ~layer2_out[8720];
     layer3_out[6210] <= ~layer2_out[36];
     layer3_out[6211] <= layer2_out[11557];
     layer3_out[6212] <= ~(layer2_out[1209] ^ layer2_out[1210]);
     layer3_out[6213] <= ~layer2_out[5607];
     layer3_out[6214] <= layer2_out[4460];
     layer3_out[6215] <= layer2_out[1438] & layer2_out[1439];
     layer3_out[6216] <= ~layer2_out[970];
     layer3_out[6217] <= ~(layer2_out[6996] | layer2_out[6997]);
     layer3_out[6218] <= layer2_out[7459] ^ layer2_out[7460];
     layer3_out[6219] <= ~(layer2_out[9008] ^ layer2_out[9009]);
     layer3_out[6220] <= layer2_out[4906] & ~layer2_out[4907];
     layer3_out[6221] <= layer2_out[346] ^ layer2_out[347];
     layer3_out[6222] <= ~(layer2_out[2541] & layer2_out[2542]);
     layer3_out[6223] <= ~layer2_out[5394];
     layer3_out[6224] <= layer2_out[2140] | layer2_out[2141];
     layer3_out[6225] <= ~layer2_out[4516];
     layer3_out[6226] <= layer2_out[690];
     layer3_out[6227] <= ~(layer2_out[5440] ^ layer2_out[5441]);
     layer3_out[6228] <= ~(layer2_out[8439] & layer2_out[8440]);
     layer3_out[6229] <= layer2_out[6348] & ~layer2_out[6347];
     layer3_out[6230] <= ~layer2_out[10131] | layer2_out[10132];
     layer3_out[6231] <= ~(layer2_out[8144] & layer2_out[8145]);
     layer3_out[6232] <= layer2_out[8912];
     layer3_out[6233] <= ~(layer2_out[4446] | layer2_out[4447]);
     layer3_out[6234] <= layer2_out[4456];
     layer3_out[6235] <= ~(layer2_out[5552] ^ layer2_out[5553]);
     layer3_out[6236] <= layer2_out[229] ^ layer2_out[230];
     layer3_out[6237] <= layer2_out[7877];
     layer3_out[6238] <= ~layer2_out[5401];
     layer3_out[6239] <= ~layer2_out[11652];
     layer3_out[6240] <= layer2_out[7817];
     layer3_out[6241] <= ~layer2_out[1380] | layer2_out[1381];
     layer3_out[6242] <= layer2_out[3604] & ~layer2_out[3603];
     layer3_out[6243] <= layer2_out[3812];
     layer3_out[6244] <= ~(layer2_out[5270] & layer2_out[5271]);
     layer3_out[6245] <= layer2_out[11074];
     layer3_out[6246] <= layer2_out[2315];
     layer3_out[6247] <= layer2_out[1174];
     layer3_out[6248] <= ~layer2_out[8259];
     layer3_out[6249] <= layer2_out[5594] ^ layer2_out[5595];
     layer3_out[6250] <= layer2_out[2492];
     layer3_out[6251] <= layer2_out[6285];
     layer3_out[6252] <= layer2_out[4896] ^ layer2_out[4897];
     layer3_out[6253] <= ~(layer2_out[11087] ^ layer2_out[11088]);
     layer3_out[6254] <= ~layer2_out[4787];
     layer3_out[6255] <= ~layer2_out[3246];
     layer3_out[6256] <= layer2_out[10796];
     layer3_out[6257] <= layer2_out[3663];
     layer3_out[6258] <= layer2_out[8372] & layer2_out[8373];
     layer3_out[6259] <= layer2_out[5010];
     layer3_out[6260] <= layer2_out[9420];
     layer3_out[6261] <= layer2_out[1768];
     layer3_out[6262] <= ~layer2_out[1743] | layer2_out[1744];
     layer3_out[6263] <= ~(layer2_out[1192] | layer2_out[1193]);
     layer3_out[6264] <= layer2_out[5683] & ~layer2_out[5684];
     layer3_out[6265] <= layer2_out[704] & layer2_out[705];
     layer3_out[6266] <= layer2_out[6838] ^ layer2_out[6839];
     layer3_out[6267] <= ~layer2_out[11518];
     layer3_out[6268] <= ~(layer2_out[797] ^ layer2_out[798]);
     layer3_out[6269] <= ~(layer2_out[4778] ^ layer2_out[4779]);
     layer3_out[6270] <= layer2_out[616] & ~layer2_out[615];
     layer3_out[6271] <= layer2_out[10204] & ~layer2_out[10205];
     layer3_out[6272] <= layer2_out[7963];
     layer3_out[6273] <= ~(layer2_out[7233] ^ layer2_out[7234]);
     layer3_out[6274] <= ~layer2_out[10191] | layer2_out[10190];
     layer3_out[6275] <= ~layer2_out[6002];
     layer3_out[6276] <= layer2_out[4703] & ~layer2_out[4702];
     layer3_out[6277] <= layer2_out[6231] ^ layer2_out[6232];
     layer3_out[6278] <= layer2_out[5930];
     layer3_out[6279] <= ~(layer2_out[9979] & layer2_out[9980]);
     layer3_out[6280] <= layer2_out[2098] | layer2_out[2099];
     layer3_out[6281] <= layer2_out[2326];
     layer3_out[6282] <= layer2_out[11353] & layer2_out[11354];
     layer3_out[6283] <= layer2_out[10817];
     layer3_out[6284] <= ~layer2_out[499];
     layer3_out[6285] <= layer2_out[11908];
     layer3_out[6286] <= ~(layer2_out[5785] ^ layer2_out[5786]);
     layer3_out[6287] <= ~(layer2_out[9485] ^ layer2_out[9486]);
     layer3_out[6288] <= ~(layer2_out[2632] & layer2_out[2633]);
     layer3_out[6289] <= ~layer2_out[3672];
     layer3_out[6290] <= ~layer2_out[6970];
     layer3_out[6291] <= layer2_out[11107] & ~layer2_out[11108];
     layer3_out[6292] <= layer2_out[8420];
     layer3_out[6293] <= layer2_out[6151] ^ layer2_out[6152];
     layer3_out[6294] <= layer2_out[8658] & layer2_out[8659];
     layer3_out[6295] <= ~layer2_out[7674];
     layer3_out[6296] <= layer2_out[5484] & ~layer2_out[5483];
     layer3_out[6297] <= ~layer2_out[6775];
     layer3_out[6298] <= ~layer2_out[4200];
     layer3_out[6299] <= ~layer2_out[6178];
     layer3_out[6300] <= ~layer2_out[11222];
     layer3_out[6301] <= layer2_out[6575];
     layer3_out[6302] <= layer2_out[5512] ^ layer2_out[5513];
     layer3_out[6303] <= ~layer2_out[920];
     layer3_out[6304] <= ~layer2_out[261];
     layer3_out[6305] <= layer2_out[9750] | layer2_out[9751];
     layer3_out[6306] <= ~layer2_out[1765];
     layer3_out[6307] <= layer2_out[4039] | layer2_out[4040];
     layer3_out[6308] <= layer2_out[6934];
     layer3_out[6309] <= layer2_out[9050];
     layer3_out[6310] <= layer2_out[6943];
     layer3_out[6311] <= ~(layer2_out[11876] ^ layer2_out[11877]);
     layer3_out[6312] <= layer2_out[805];
     layer3_out[6313] <= layer2_out[3552] ^ layer2_out[3553];
     layer3_out[6314] <= layer2_out[11675] & ~layer2_out[11674];
     layer3_out[6315] <= ~(layer2_out[6346] | layer2_out[6347]);
     layer3_out[6316] <= layer2_out[5849] | layer2_out[5850];
     layer3_out[6317] <= ~layer2_out[8815];
     layer3_out[6318] <= layer2_out[3512];
     layer3_out[6319] <= layer2_out[1796];
     layer3_out[6320] <= layer2_out[4679] | layer2_out[4680];
     layer3_out[6321] <= layer2_out[1652] ^ layer2_out[1653];
     layer3_out[6322] <= layer2_out[11260];
     layer3_out[6323] <= ~layer2_out[92];
     layer3_out[6324] <= layer2_out[8850] ^ layer2_out[8851];
     layer3_out[6325] <= ~(layer2_out[2846] & layer2_out[2847]);
     layer3_out[6326] <= ~layer2_out[9639];
     layer3_out[6327] <= layer2_out[5807] & ~layer2_out[5808];
     layer3_out[6328] <= ~layer2_out[9220];
     layer3_out[6329] <= ~(layer2_out[6675] ^ layer2_out[6676]);
     layer3_out[6330] <= ~layer2_out[9402] | layer2_out[9403];
     layer3_out[6331] <= ~(layer2_out[9726] ^ layer2_out[9727]);
     layer3_out[6332] <= layer2_out[10686] ^ layer2_out[10687];
     layer3_out[6333] <= ~layer2_out[3188];
     layer3_out[6334] <= ~(layer2_out[9587] ^ layer2_out[9588]);
     layer3_out[6335] <= layer2_out[6927];
     layer3_out[6336] <= layer2_out[327] ^ layer2_out[328];
     layer3_out[6337] <= layer2_out[5649] ^ layer2_out[5650];
     layer3_out[6338] <= ~(layer2_out[9727] & layer2_out[9728]);
     layer3_out[6339] <= 1'b1;
     layer3_out[6340] <= ~(layer2_out[11285] ^ layer2_out[11286]);
     layer3_out[6341] <= layer2_out[1063] & ~layer2_out[1062];
     layer3_out[6342] <= ~(layer2_out[5954] ^ layer2_out[5955]);
     layer3_out[6343] <= ~layer2_out[9978];
     layer3_out[6344] <= ~layer2_out[3392] | layer2_out[3391];
     layer3_out[6345] <= layer2_out[966] & layer2_out[967];
     layer3_out[6346] <= ~layer2_out[6679];
     layer3_out[6347] <= layer2_out[7181] ^ layer2_out[7182];
     layer3_out[6348] <= layer2_out[11298];
     layer3_out[6349] <= layer2_out[6534] | layer2_out[6535];
     layer3_out[6350] <= ~(layer2_out[4691] | layer2_out[4692]);
     layer3_out[6351] <= layer2_out[11056] | layer2_out[11057];
     layer3_out[6352] <= ~layer2_out[1731];
     layer3_out[6353] <= layer2_out[715];
     layer3_out[6354] <= ~layer2_out[11605];
     layer3_out[6355] <= layer2_out[4344];
     layer3_out[6356] <= layer2_out[555];
     layer3_out[6357] <= ~layer2_out[10778];
     layer3_out[6358] <= ~layer2_out[4188];
     layer3_out[6359] <= layer2_out[11858] & ~layer2_out[11857];
     layer3_out[6360] <= ~layer2_out[9837];
     layer3_out[6361] <= ~(layer2_out[7568] | layer2_out[7569]);
     layer3_out[6362] <= ~layer2_out[10272];
     layer3_out[6363] <= layer2_out[775] & ~layer2_out[774];
     layer3_out[6364] <= ~(layer2_out[1877] | layer2_out[1878]);
     layer3_out[6365] <= ~layer2_out[8379];
     layer3_out[6366] <= layer2_out[9701] & layer2_out[9702];
     layer3_out[6367] <= ~layer2_out[681];
     layer3_out[6368] <= layer2_out[7992] | layer2_out[7993];
     layer3_out[6369] <= layer2_out[5225] ^ layer2_out[5226];
     layer3_out[6370] <= layer2_out[5788];
     layer3_out[6371] <= ~(layer2_out[4623] ^ layer2_out[4624]);
     layer3_out[6372] <= layer2_out[9228] | layer2_out[9229];
     layer3_out[6373] <= layer2_out[9299];
     layer3_out[6374] <= layer2_out[2567];
     layer3_out[6375] <= ~layer2_out[7835];
     layer3_out[6376] <= layer2_out[5953] ^ layer2_out[5954];
     layer3_out[6377] <= ~(layer2_out[5019] ^ layer2_out[5020]);
     layer3_out[6378] <= layer2_out[8719] & ~layer2_out[8720];
     layer3_out[6379] <= layer2_out[1000];
     layer3_out[6380] <= ~layer2_out[389] | layer2_out[390];
     layer3_out[6381] <= layer2_out[10318];
     layer3_out[6382] <= layer2_out[5719] | layer2_out[5720];
     layer3_out[6383] <= ~(layer2_out[10570] & layer2_out[10571]);
     layer3_out[6384] <= ~(layer2_out[6034] ^ layer2_out[6035]);
     layer3_out[6385] <= ~(layer2_out[11816] | layer2_out[11817]);
     layer3_out[6386] <= ~layer2_out[6444];
     layer3_out[6387] <= layer2_out[9208];
     layer3_out[6388] <= ~layer2_out[10677] | layer2_out[10676];
     layer3_out[6389] <= ~(layer2_out[576] | layer2_out[577]);
     layer3_out[6390] <= layer2_out[11355] ^ layer2_out[11356];
     layer3_out[6391] <= layer2_out[1295] & ~layer2_out[1294];
     layer3_out[6392] <= ~layer2_out[4910];
     layer3_out[6393] <= layer2_out[3125] ^ layer2_out[3126];
     layer3_out[6394] <= ~(layer2_out[1906] ^ layer2_out[1907]);
     layer3_out[6395] <= ~(layer2_out[11218] ^ layer2_out[11219]);
     layer3_out[6396] <= ~(layer2_out[9535] & layer2_out[9536]);
     layer3_out[6397] <= layer2_out[7827] ^ layer2_out[7828];
     layer3_out[6398] <= layer2_out[9861];
     layer3_out[6399] <= layer2_out[238] & ~layer2_out[237];
     layer3_out[6400] <= layer2_out[6723] ^ layer2_out[6724];
     layer3_out[6401] <= layer2_out[8094];
     layer3_out[6402] <= ~layer2_out[5916];
     layer3_out[6403] <= ~(layer2_out[6464] ^ layer2_out[6465]);
     layer3_out[6404] <= ~(layer2_out[11428] ^ layer2_out[11429]);
     layer3_out[6405] <= ~(layer2_out[10560] ^ layer2_out[10561]);
     layer3_out[6406] <= ~layer2_out[8692] | layer2_out[8693];
     layer3_out[6407] <= layer2_out[1671] | layer2_out[1672];
     layer3_out[6408] <= ~(layer2_out[7976] ^ layer2_out[7977]);
     layer3_out[6409] <= ~layer2_out[3693];
     layer3_out[6410] <= ~layer2_out[5421];
     layer3_out[6411] <= ~(layer2_out[7320] ^ layer2_out[7321]);
     layer3_out[6412] <= layer2_out[1056] ^ layer2_out[1057];
     layer3_out[6413] <= layer2_out[8093] | layer2_out[8094];
     layer3_out[6414] <= layer2_out[7646];
     layer3_out[6415] <= layer2_out[9893];
     layer3_out[6416] <= layer2_out[4090] & layer2_out[4091];
     layer3_out[6417] <= ~(layer2_out[1217] ^ layer2_out[1218]);
     layer3_out[6418] <= ~layer2_out[896] | layer2_out[897];
     layer3_out[6419] <= layer2_out[10000];
     layer3_out[6420] <= layer2_out[1614] ^ layer2_out[1615];
     layer3_out[6421] <= layer2_out[11148];
     layer3_out[6422] <= layer2_out[6171];
     layer3_out[6423] <= layer2_out[2699] & ~layer2_out[2700];
     layer3_out[6424] <= layer2_out[9393] | layer2_out[9394];
     layer3_out[6425] <= ~layer2_out[5963];
     layer3_out[6426] <= layer2_out[7664] & ~layer2_out[7663];
     layer3_out[6427] <= ~(layer2_out[4732] ^ layer2_out[4733]);
     layer3_out[6428] <= layer2_out[9751] | layer2_out[9752];
     layer3_out[6429] <= ~layer2_out[8283];
     layer3_out[6430] <= layer2_out[3964] & layer2_out[3965];
     layer3_out[6431] <= ~layer2_out[1757];
     layer3_out[6432] <= ~layer2_out[5364] | layer2_out[5363];
     layer3_out[6433] <= ~(layer2_out[6756] ^ layer2_out[6757]);
     layer3_out[6434] <= ~(layer2_out[3845] | layer2_out[3846]);
     layer3_out[6435] <= layer2_out[4042] & layer2_out[4043];
     layer3_out[6436] <= layer2_out[7611] | layer2_out[7612];
     layer3_out[6437] <= layer2_out[11116] ^ layer2_out[11117];
     layer3_out[6438] <= layer2_out[4504] ^ layer2_out[4505];
     layer3_out[6439] <= ~layer2_out[7359];
     layer3_out[6440] <= ~(layer2_out[3777] ^ layer2_out[3778]);
     layer3_out[6441] <= ~layer2_out[6484];
     layer3_out[6442] <= ~layer2_out[5802];
     layer3_out[6443] <= layer2_out[10647] & ~layer2_out[10648];
     layer3_out[6444] <= layer2_out[10081] | layer2_out[10082];
     layer3_out[6445] <= ~(layer2_out[8806] & layer2_out[8807]);
     layer3_out[6446] <= ~(layer2_out[3330] & layer2_out[3331]);
     layer3_out[6447] <= ~layer2_out[9268];
     layer3_out[6448] <= ~layer2_out[1810];
     layer3_out[6449] <= layer2_out[3507];
     layer3_out[6450] <= ~(layer2_out[1566] ^ layer2_out[1567]);
     layer3_out[6451] <= ~(layer2_out[9398] ^ layer2_out[9399]);
     layer3_out[6452] <= layer2_out[9655] ^ layer2_out[9656];
     layer3_out[6453] <= layer2_out[4761] ^ layer2_out[4762];
     layer3_out[6454] <= layer2_out[3096] | layer2_out[3097];
     layer3_out[6455] <= ~(layer2_out[4427] ^ layer2_out[4428]);
     layer3_out[6456] <= ~layer2_out[6940];
     layer3_out[6457] <= ~(layer2_out[3721] ^ layer2_out[3722]);
     layer3_out[6458] <= layer2_out[3109] & ~layer2_out[3110];
     layer3_out[6459] <= layer2_out[1996] | layer2_out[1997];
     layer3_out[6460] <= ~(layer2_out[3518] | layer2_out[3519]);
     layer3_out[6461] <= ~layer2_out[638];
     layer3_out[6462] <= layer2_out[7293] | layer2_out[7294];
     layer3_out[6463] <= layer2_out[4539];
     layer3_out[6464] <= ~layer2_out[6970];
     layer3_out[6465] <= ~(layer2_out[7423] & layer2_out[7424]);
     layer3_out[6466] <= ~(layer2_out[9978] & layer2_out[9979]);
     layer3_out[6467] <= layer2_out[10258] & layer2_out[10259];
     layer3_out[6468] <= ~(layer2_out[1251] ^ layer2_out[1252]);
     layer3_out[6469] <= ~layer2_out[1222];
     layer3_out[6470] <= ~layer2_out[9740];
     layer3_out[6471] <= ~(layer2_out[289] ^ layer2_out[290]);
     layer3_out[6472] <= layer2_out[4729] | layer2_out[4730];
     layer3_out[6473] <= layer2_out[7824];
     layer3_out[6474] <= ~(layer2_out[5075] ^ layer2_out[5076]);
     layer3_out[6475] <= layer2_out[11103] ^ layer2_out[11104];
     layer3_out[6476] <= layer2_out[6441];
     layer3_out[6477] <= ~(layer2_out[3550] ^ layer2_out[3551]);
     layer3_out[6478] <= layer2_out[9146] & ~layer2_out[9145];
     layer3_out[6479] <= layer2_out[1082] ^ layer2_out[1083];
     layer3_out[6480] <= ~layer2_out[7444];
     layer3_out[6481] <= layer2_out[3598];
     layer3_out[6482] <= layer2_out[7635];
     layer3_out[6483] <= layer2_out[1579];
     layer3_out[6484] <= ~(layer2_out[1368] | layer2_out[1369]);
     layer3_out[6485] <= layer2_out[4643];
     layer3_out[6486] <= layer2_out[10841];
     layer3_out[6487] <= layer2_out[4183] ^ layer2_out[4184];
     layer3_out[6488] <= ~layer2_out[3713];
     layer3_out[6489] <= layer2_out[6216];
     layer3_out[6490] <= ~(layer2_out[1083] ^ layer2_out[1084]);
     layer3_out[6491] <= ~layer2_out[2527];
     layer3_out[6492] <= ~(layer2_out[782] ^ layer2_out[783]);
     layer3_out[6493] <= layer2_out[4482];
     layer3_out[6494] <= layer2_out[7566];
     layer3_out[6495] <= ~(layer2_out[3448] & layer2_out[3449]);
     layer3_out[6496] <= ~(layer2_out[6359] ^ layer2_out[6360]);
     layer3_out[6497] <= layer2_out[3608] & ~layer2_out[3607];
     layer3_out[6498] <= layer2_out[3102];
     layer3_out[6499] <= ~layer2_out[4736];
     layer3_out[6500] <= layer2_out[11374];
     layer3_out[6501] <= ~(layer2_out[3875] & layer2_out[3876]);
     layer3_out[6502] <= ~layer2_out[11409];
     layer3_out[6503] <= layer2_out[4831] ^ layer2_out[4832];
     layer3_out[6504] <= ~layer2_out[444] | layer2_out[445];
     layer3_out[6505] <= ~layer2_out[2804] | layer2_out[2803];
     layer3_out[6506] <= layer2_out[2510] ^ layer2_out[2511];
     layer3_out[6507] <= ~layer2_out[10871];
     layer3_out[6508] <= layer2_out[3272] | layer2_out[3273];
     layer3_out[6509] <= layer2_out[8770] & ~layer2_out[8769];
     layer3_out[6510] <= layer2_out[7048] & layer2_out[7049];
     layer3_out[6511] <= layer2_out[1830] & layer2_out[1831];
     layer3_out[6512] <= ~(layer2_out[3409] | layer2_out[3410]);
     layer3_out[6513] <= layer2_out[6100] ^ layer2_out[6101];
     layer3_out[6514] <= layer2_out[11358];
     layer3_out[6515] <= ~layer2_out[2791];
     layer3_out[6516] <= layer2_out[3500] ^ layer2_out[3501];
     layer3_out[6517] <= layer2_out[2327] ^ layer2_out[2328];
     layer3_out[6518] <= ~layer2_out[4544];
     layer3_out[6519] <= ~(layer2_out[11710] & layer2_out[11711]);
     layer3_out[6520] <= layer2_out[609] ^ layer2_out[610];
     layer3_out[6521] <= ~(layer2_out[9889] ^ layer2_out[9890]);
     layer3_out[6522] <= layer2_out[2631];
     layer3_out[6523] <= layer2_out[2227];
     layer3_out[6524] <= ~layer2_out[8745];
     layer3_out[6525] <= layer2_out[4410];
     layer3_out[6526] <= ~(layer2_out[9198] ^ layer2_out[9199]);
     layer3_out[6527] <= layer2_out[9694] | layer2_out[9695];
     layer3_out[6528] <= layer2_out[1692] | layer2_out[1693];
     layer3_out[6529] <= layer2_out[5475] | layer2_out[5476];
     layer3_out[6530] <= ~layer2_out[11317];
     layer3_out[6531] <= layer2_out[341] ^ layer2_out[342];
     layer3_out[6532] <= layer2_out[10844];
     layer3_out[6533] <= layer2_out[1486];
     layer3_out[6534] <= ~(layer2_out[4140] ^ layer2_out[4141]);
     layer3_out[6535] <= ~layer2_out[1426];
     layer3_out[6536] <= ~layer2_out[1352] | layer2_out[1353];
     layer3_out[6537] <= ~(layer2_out[9011] & layer2_out[9012]);
     layer3_out[6538] <= layer2_out[8733] & ~layer2_out[8732];
     layer3_out[6539] <= ~(layer2_out[11290] | layer2_out[11291]);
     layer3_out[6540] <= ~(layer2_out[9052] ^ layer2_out[9053]);
     layer3_out[6541] <= layer2_out[6267] & layer2_out[6268];
     layer3_out[6542] <= layer2_out[7644] & ~layer2_out[7643];
     layer3_out[6543] <= layer2_out[1888];
     layer3_out[6544] <= layer2_out[6204];
     layer3_out[6545] <= ~layer2_out[9876] | layer2_out[9875];
     layer3_out[6546] <= layer2_out[3555];
     layer3_out[6547] <= layer2_out[3343];
     layer3_out[6548] <= ~(layer2_out[6936] & layer2_out[6937]);
     layer3_out[6549] <= layer2_out[5609] ^ layer2_out[5610];
     layer3_out[6550] <= layer2_out[8211];
     layer3_out[6551] <= ~layer2_out[11702];
     layer3_out[6552] <= layer2_out[1919] & ~layer2_out[1920];
     layer3_out[6553] <= layer2_out[447];
     layer3_out[6554] <= layer2_out[1050] ^ layer2_out[1051];
     layer3_out[6555] <= layer2_out[10122] & layer2_out[10123];
     layer3_out[6556] <= layer2_out[10154] ^ layer2_out[10155];
     layer3_out[6557] <= ~layer2_out[3255];
     layer3_out[6558] <= layer2_out[2775] | layer2_out[2776];
     layer3_out[6559] <= ~layer2_out[455];
     layer3_out[6560] <= ~layer2_out[8175] | layer2_out[8176];
     layer3_out[6561] <= ~layer2_out[11732] | layer2_out[11731];
     layer3_out[6562] <= layer2_out[2189] & ~layer2_out[2190];
     layer3_out[6563] <= ~layer2_out[9363] | layer2_out[9362];
     layer3_out[6564] <= ~layer2_out[739] | layer2_out[738];
     layer3_out[6565] <= ~layer2_out[726];
     layer3_out[6566] <= layer2_out[737] ^ layer2_out[738];
     layer3_out[6567] <= layer2_out[5602] & layer2_out[5603];
     layer3_out[6568] <= ~layer2_out[11939] | layer2_out[11940];
     layer3_out[6569] <= ~layer2_out[10213] | layer2_out[10212];
     layer3_out[6570] <= layer2_out[7900];
     layer3_out[6571] <= layer2_out[2617] | layer2_out[2618];
     layer3_out[6572] <= ~(layer2_out[1574] ^ layer2_out[1575]);
     layer3_out[6573] <= layer2_out[4155] & layer2_out[4156];
     layer3_out[6574] <= layer2_out[6636] ^ layer2_out[6637];
     layer3_out[6575] <= layer2_out[11687] | layer2_out[11688];
     layer3_out[6576] <= layer2_out[10043];
     layer3_out[6577] <= layer2_out[5587] & ~layer2_out[5588];
     layer3_out[6578] <= ~(layer2_out[7248] & layer2_out[7249]);
     layer3_out[6579] <= layer2_out[2979] & layer2_out[2980];
     layer3_out[6580] <= ~layer2_out[10627];
     layer3_out[6581] <= layer2_out[46];
     layer3_out[6582] <= layer2_out[7] | layer2_out[8];
     layer3_out[6583] <= layer2_out[122];
     layer3_out[6584] <= layer2_out[5436];
     layer3_out[6585] <= ~(layer2_out[11758] & layer2_out[11759]);
     layer3_out[6586] <= ~(layer2_out[164] ^ layer2_out[165]);
     layer3_out[6587] <= ~layer2_out[4742];
     layer3_out[6588] <= ~(layer2_out[579] ^ layer2_out[580]);
     layer3_out[6589] <= ~(layer2_out[9430] & layer2_out[9431]);
     layer3_out[6590] <= ~layer2_out[7099];
     layer3_out[6591] <= ~(layer2_out[11870] ^ layer2_out[11871]);
     layer3_out[6592] <= ~layer2_out[8370];
     layer3_out[6593] <= ~(layer2_out[3700] & layer2_out[3701]);
     layer3_out[6594] <= layer2_out[9504] & layer2_out[9505];
     layer3_out[6595] <= ~(layer2_out[8359] & layer2_out[8360]);
     layer3_out[6596] <= ~layer2_out[11202] | layer2_out[11203];
     layer3_out[6597] <= ~layer2_out[6438];
     layer3_out[6598] <= layer2_out[4126] ^ layer2_out[4127];
     layer3_out[6599] <= ~(layer2_out[9500] | layer2_out[9501]);
     layer3_out[6600] <= layer2_out[6397];
     layer3_out[6601] <= layer2_out[8778] | layer2_out[8779];
     layer3_out[6602] <= ~layer2_out[5626] | layer2_out[5625];
     layer3_out[6603] <= ~layer2_out[2802] | layer2_out[2803];
     layer3_out[6604] <= layer2_out[10645] | layer2_out[10646];
     layer3_out[6605] <= ~layer2_out[823] | layer2_out[824];
     layer3_out[6606] <= ~layer2_out[7160];
     layer3_out[6607] <= ~(layer2_out[1093] ^ layer2_out[1094]);
     layer3_out[6608] <= ~layer2_out[11750];
     layer3_out[6609] <= layer2_out[11544];
     layer3_out[6610] <= layer2_out[4719] | layer2_out[4720];
     layer3_out[6611] <= layer2_out[8965];
     layer3_out[6612] <= ~(layer2_out[7601] ^ layer2_out[7602]);
     layer3_out[6613] <= layer2_out[6023] ^ layer2_out[6024];
     layer3_out[6614] <= layer2_out[10699];
     layer3_out[6615] <= layer2_out[9602] & ~layer2_out[9603];
     layer3_out[6616] <= ~(layer2_out[4004] ^ layer2_out[4005]);
     layer3_out[6617] <= layer2_out[4552];
     layer3_out[6618] <= layer2_out[1784] ^ layer2_out[1785];
     layer3_out[6619] <= layer2_out[4372] | layer2_out[4373];
     layer3_out[6620] <= ~(layer2_out[5619] & layer2_out[5620]);
     layer3_out[6621] <= layer2_out[902] ^ layer2_out[903];
     layer3_out[6622] <= ~layer2_out[7931] | layer2_out[7930];
     layer3_out[6623] <= layer2_out[5678] & ~layer2_out[5679];
     layer3_out[6624] <= layer2_out[5320] ^ layer2_out[5321];
     layer3_out[6625] <= layer2_out[5439] & ~layer2_out[5438];
     layer3_out[6626] <= ~layer2_out[9769];
     layer3_out[6627] <= layer2_out[2349];
     layer3_out[6628] <= ~layer2_out[6000];
     layer3_out[6629] <= layer2_out[8699] & layer2_out[8700];
     layer3_out[6630] <= ~layer2_out[411];
     layer3_out[6631] <= layer2_out[3853];
     layer3_out[6632] <= ~(layer2_out[6828] ^ layer2_out[6829]);
     layer3_out[6633] <= layer2_out[10056];
     layer3_out[6634] <= ~layer2_out[7449];
     layer3_out[6635] <= ~layer2_out[2818] | layer2_out[2817];
     layer3_out[6636] <= layer2_out[11321] ^ layer2_out[11322];
     layer3_out[6637] <= ~layer2_out[8902];
     layer3_out[6638] <= ~(layer2_out[1340] ^ layer2_out[1341]);
     layer3_out[6639] <= ~(layer2_out[503] ^ layer2_out[504]);
     layer3_out[6640] <= layer2_out[8415] ^ layer2_out[8416];
     layer3_out[6641] <= layer2_out[1655] & ~layer2_out[1656];
     layer3_out[6642] <= layer2_out[9450] & ~layer2_out[9449];
     layer3_out[6643] <= layer2_out[6054] & ~layer2_out[6055];
     layer3_out[6644] <= ~layer2_out[9992];
     layer3_out[6645] <= layer2_out[3154];
     layer3_out[6646] <= ~(layer2_out[4968] | layer2_out[4969]);
     layer3_out[6647] <= layer2_out[9557] & ~layer2_out[9558];
     layer3_out[6648] <= ~layer2_out[11816];
     layer3_out[6649] <= layer2_out[1857] & layer2_out[1858];
     layer3_out[6650] <= ~(layer2_out[5373] ^ layer2_out[5374]);
     layer3_out[6651] <= layer2_out[9457];
     layer3_out[6652] <= layer2_out[4249] & layer2_out[4250];
     layer3_out[6653] <= ~layer2_out[6628];
     layer3_out[6654] <= ~layer2_out[9145];
     layer3_out[6655] <= ~(layer2_out[8052] ^ layer2_out[8053]);
     layer3_out[6656] <= layer2_out[6566] ^ layer2_out[6567];
     layer3_out[6657] <= ~layer2_out[9472] | layer2_out[9473];
     layer3_out[6658] <= layer2_out[8563];
     layer3_out[6659] <= layer2_out[136];
     layer3_out[6660] <= ~layer2_out[2665];
     layer3_out[6661] <= layer2_out[4054] | layer2_out[4055];
     layer3_out[6662] <= layer2_out[9698];
     layer3_out[6663] <= layer2_out[6995];
     layer3_out[6664] <= ~layer2_out[2163];
     layer3_out[6665] <= ~(layer2_out[7203] ^ layer2_out[7204]);
     layer3_out[6666] <= layer2_out[10149];
     layer3_out[6667] <= layer2_out[1781] & layer2_out[1782];
     layer3_out[6668] <= ~(layer2_out[6677] ^ layer2_out[6678]);
     layer3_out[6669] <= layer2_out[7800] & ~layer2_out[7799];
     layer3_out[6670] <= layer2_out[4116] & ~layer2_out[4117];
     layer3_out[6671] <= layer2_out[5549];
     layer3_out[6672] <= ~(layer2_out[356] & layer2_out[357]);
     layer3_out[6673] <= ~layer2_out[1395];
     layer3_out[6674] <= ~layer2_out[6638];
     layer3_out[6675] <= layer2_out[7817];
     layer3_out[6676] <= layer2_out[5131];
     layer3_out[6677] <= layer2_out[11119] | layer2_out[11120];
     layer3_out[6678] <= ~(layer2_out[11551] | layer2_out[11552]);
     layer3_out[6679] <= ~(layer2_out[3880] | layer2_out[3881]);
     layer3_out[6680] <= layer2_out[922] & ~layer2_out[923];
     layer3_out[6681] <= ~layer2_out[8254];
     layer3_out[6682] <= ~layer2_out[10329] | layer2_out[10328];
     layer3_out[6683] <= ~layer2_out[5795] | layer2_out[5794];
     layer3_out[6684] <= layer2_out[7307] & layer2_out[7308];
     layer3_out[6685] <= ~(layer2_out[7456] & layer2_out[7457]);
     layer3_out[6686] <= layer2_out[441];
     layer3_out[6687] <= ~(layer2_out[11741] | layer2_out[11742]);
     layer3_out[6688] <= ~layer2_out[9828];
     layer3_out[6689] <= ~layer2_out[6922] | layer2_out[6921];
     layer3_out[6690] <= ~(layer2_out[10220] | layer2_out[10221]);
     layer3_out[6691] <= ~(layer2_out[11756] | layer2_out[11757]);
     layer3_out[6692] <= layer2_out[3353] ^ layer2_out[3354];
     layer3_out[6693] <= ~(layer2_out[1227] ^ layer2_out[1228]);
     layer3_out[6694] <= layer2_out[6646];
     layer3_out[6695] <= ~layer2_out[11904];
     layer3_out[6696] <= layer2_out[1203] & ~layer2_out[1204];
     layer3_out[6697] <= layer2_out[2752];
     layer3_out[6698] <= layer2_out[2185] & ~layer2_out[2186];
     layer3_out[6699] <= layer2_out[6976] & ~layer2_out[6977];
     layer3_out[6700] <= ~layer2_out[833];
     layer3_out[6701] <= layer2_out[834] ^ layer2_out[835];
     layer3_out[6702] <= layer2_out[6689] & layer2_out[6690];
     layer3_out[6703] <= ~(layer2_out[7994] & layer2_out[7995]);
     layer3_out[6704] <= layer2_out[933];
     layer3_out[6705] <= layer2_out[5478] & layer2_out[5479];
     layer3_out[6706] <= ~layer2_out[3788];
     layer3_out[6707] <= ~layer2_out[340] | layer2_out[339];
     layer3_out[6708] <= ~layer2_out[8656];
     layer3_out[6709] <= ~(layer2_out[4114] & layer2_out[4115]);
     layer3_out[6710] <= ~layer2_out[10226];
     layer3_out[6711] <= layer2_out[4069] ^ layer2_out[4070];
     layer3_out[6712] <= ~(layer2_out[634] | layer2_out[635]);
     layer3_out[6713] <= layer2_out[2444] & layer2_out[2445];
     layer3_out[6714] <= layer2_out[1698] ^ layer2_out[1699];
     layer3_out[6715] <= layer2_out[2278] ^ layer2_out[2279];
     layer3_out[6716] <= layer2_out[5793];
     layer3_out[6717] <= layer2_out[11780] ^ layer2_out[11781];
     layer3_out[6718] <= layer2_out[11299] ^ layer2_out[11300];
     layer3_out[6719] <= ~layer2_out[2774] | layer2_out[2775];
     layer3_out[6720] <= layer2_out[866] & layer2_out[867];
     layer3_out[6721] <= layer2_out[775] ^ layer2_out[776];
     layer3_out[6722] <= layer2_out[2694] & ~layer2_out[2695];
     layer3_out[6723] <= layer2_out[9930] & layer2_out[9931];
     layer3_out[6724] <= ~(layer2_out[7175] & layer2_out[7176]);
     layer3_out[6725] <= ~layer2_out[5253] | layer2_out[5252];
     layer3_out[6726] <= ~(layer2_out[4124] ^ layer2_out[4125]);
     layer3_out[6727] <= ~(layer2_out[5333] & layer2_out[5334]);
     layer3_out[6728] <= ~layer2_out[5523];
     layer3_out[6729] <= layer2_out[1699] ^ layer2_out[1700];
     layer3_out[6730] <= layer2_out[8506] & ~layer2_out[8505];
     layer3_out[6731] <= layer2_out[6975];
     layer3_out[6732] <= layer2_out[391];
     layer3_out[6733] <= layer2_out[6786];
     layer3_out[6734] <= ~layer2_out[6409];
     layer3_out[6735] <= layer2_out[1909];
     layer3_out[6736] <= layer2_out[8641];
     layer3_out[6737] <= ~layer2_out[3098] | layer2_out[3099];
     layer3_out[6738] <= ~layer2_out[11160];
     layer3_out[6739] <= ~layer2_out[4347];
     layer3_out[6740] <= layer2_out[11398] & ~layer2_out[11397];
     layer3_out[6741] <= ~(layer2_out[11340] ^ layer2_out[11341]);
     layer3_out[6742] <= ~(layer2_out[10101] ^ layer2_out[10102]);
     layer3_out[6743] <= ~(layer2_out[9564] | layer2_out[9565]);
     layer3_out[6744] <= ~layer2_out[5843] | layer2_out[5844];
     layer3_out[6745] <= layer2_out[7158] & ~layer2_out[7159];
     layer3_out[6746] <= layer2_out[7743] & ~layer2_out[7744];
     layer3_out[6747] <= ~layer2_out[6909];
     layer3_out[6748] <= ~(layer2_out[4649] | layer2_out[4650]);
     layer3_out[6749] <= ~layer2_out[7012];
     layer3_out[6750] <= layer2_out[4350] ^ layer2_out[4351];
     layer3_out[6751] <= layer2_out[8727] | layer2_out[8728];
     layer3_out[6752] <= layer2_out[2237] & ~layer2_out[2238];
     layer3_out[6753] <= ~layer2_out[9000];
     layer3_out[6754] <= layer2_out[5210];
     layer3_out[6755] <= ~(layer2_out[4048] & layer2_out[4049]);
     layer3_out[6756] <= ~layer2_out[158];
     layer3_out[6757] <= ~(layer2_out[2530] & layer2_out[2531]);
     layer3_out[6758] <= layer2_out[4211];
     layer3_out[6759] <= layer2_out[8335] | layer2_out[8336];
     layer3_out[6760] <= layer2_out[4701];
     layer3_out[6761] <= layer2_out[11033] & ~layer2_out[11034];
     layer3_out[6762] <= layer2_out[3984] | layer2_out[3985];
     layer3_out[6763] <= layer2_out[4330];
     layer3_out[6764] <= ~(layer2_out[526] & layer2_out[527]);
     layer3_out[6765] <= ~layer2_out[6236] | layer2_out[6235];
     layer3_out[6766] <= layer2_out[3812] & layer2_out[3813];
     layer3_out[6767] <= ~layer2_out[2882];
     layer3_out[6768] <= layer2_out[6048];
     layer3_out[6769] <= layer2_out[1404] & layer2_out[1405];
     layer3_out[6770] <= ~layer2_out[2229] | layer2_out[2228];
     layer3_out[6771] <= layer2_out[5630];
     layer3_out[6772] <= ~(layer2_out[6638] | layer2_out[6639]);
     layer3_out[6773] <= layer2_out[1974];
     layer3_out[6774] <= layer2_out[11436];
     layer3_out[6775] <= layer2_out[5807] & ~layer2_out[5806];
     layer3_out[6776] <= layer2_out[6931];
     layer3_out[6777] <= ~layer2_out[2372] | layer2_out[2373];
     layer3_out[6778] <= layer2_out[1030] & ~layer2_out[1031];
     layer3_out[6779] <= layer2_out[4271];
     layer3_out[6780] <= layer2_out[8514] ^ layer2_out[8515];
     layer3_out[6781] <= ~layer2_out[5450];
     layer3_out[6782] <= layer2_out[5443];
     layer3_out[6783] <= layer2_out[9024];
     layer3_out[6784] <= layer2_out[2915] & layer2_out[2916];
     layer3_out[6785] <= ~layer2_out[6870] | layer2_out[6871];
     layer3_out[6786] <= ~layer2_out[3308];
     layer3_out[6787] <= ~(layer2_out[8970] | layer2_out[8971]);
     layer3_out[6788] <= layer2_out[11496] | layer2_out[11497];
     layer3_out[6789] <= layer2_out[588];
     layer3_out[6790] <= layer2_out[1483];
     layer3_out[6791] <= layer2_out[5208] & ~layer2_out[5209];
     layer3_out[6792] <= ~(layer2_out[10614] & layer2_out[10615]);
     layer3_out[6793] <= layer2_out[5702] & layer2_out[5703];
     layer3_out[6794] <= layer2_out[11445];
     layer3_out[6795] <= layer2_out[9918];
     layer3_out[6796] <= ~(layer2_out[2250] & layer2_out[2251]);
     layer3_out[6797] <= layer2_out[7214];
     layer3_out[6798] <= ~layer2_out[9958];
     layer3_out[6799] <= layer2_out[3466] ^ layer2_out[3467];
     layer3_out[6800] <= ~(layer2_out[5705] ^ layer2_out[5706]);
     layer3_out[6801] <= ~layer2_out[8815] | layer2_out[8814];
     layer3_out[6802] <= ~(layer2_out[6107] | layer2_out[6108]);
     layer3_out[6803] <= ~(layer2_out[6903] ^ layer2_out[6904]);
     layer3_out[6804] <= ~(layer2_out[10629] | layer2_out[10630]);
     layer3_out[6805] <= ~(layer2_out[5667] ^ layer2_out[5668]);
     layer3_out[6806] <= layer2_out[512];
     layer3_out[6807] <= ~(layer2_out[4812] | layer2_out[4813]);
     layer3_out[6808] <= layer2_out[10041];
     layer3_out[6809] <= ~layer2_out[4357];
     layer3_out[6810] <= ~layer2_out[1523];
     layer3_out[6811] <= layer2_out[6211] ^ layer2_out[6212];
     layer3_out[6812] <= ~layer2_out[5412];
     layer3_out[6813] <= ~layer2_out[4031];
     layer3_out[6814] <= ~layer2_out[2558];
     layer3_out[6815] <= layer2_out[5016];
     layer3_out[6816] <= ~layer2_out[1581];
     layer3_out[6817] <= ~(layer2_out[2552] ^ layer2_out[2553]);
     layer3_out[6818] <= layer2_out[10297];
     layer3_out[6819] <= ~layer2_out[8178] | layer2_out[8177];
     layer3_out[6820] <= layer2_out[9688];
     layer3_out[6821] <= layer2_out[11984] & ~layer2_out[11983];
     layer3_out[6822] <= layer2_out[8754] | layer2_out[8755];
     layer3_out[6823] <= ~(layer2_out[7956] ^ layer2_out[7957]);
     layer3_out[6824] <= layer2_out[296] & layer2_out[297];
     layer3_out[6825] <= ~(layer2_out[2725] & layer2_out[2726]);
     layer3_out[6826] <= layer2_out[400] | layer2_out[401];
     layer3_out[6827] <= ~(layer2_out[8800] & layer2_out[8801]);
     layer3_out[6828] <= ~layer2_out[10271] | layer2_out[10270];
     layer3_out[6829] <= ~layer2_out[10309];
     layer3_out[6830] <= ~layer2_out[8646];
     layer3_out[6831] <= ~(layer2_out[6799] & layer2_out[6800]);
     layer3_out[6832] <= layer2_out[8599] ^ layer2_out[8600];
     layer3_out[6833] <= layer2_out[8500] & ~layer2_out[8499];
     layer3_out[6834] <= layer2_out[4373];
     layer3_out[6835] <= ~layer2_out[1150];
     layer3_out[6836] <= layer2_out[2406];
     layer3_out[6837] <= ~(layer2_out[1243] | layer2_out[1244]);
     layer3_out[6838] <= layer2_out[8571];
     layer3_out[6839] <= layer2_out[5618];
     layer3_out[6840] <= ~layer2_out[7006];
     layer3_out[6841] <= layer2_out[2316] ^ layer2_out[2317];
     layer3_out[6842] <= ~layer2_out[8452];
     layer3_out[6843] <= ~layer2_out[11706] | layer2_out[11705];
     layer3_out[6844] <= layer2_out[4064] & ~layer2_out[4063];
     layer3_out[6845] <= layer2_out[2365] & layer2_out[2366];
     layer3_out[6846] <= ~(layer2_out[11722] ^ layer2_out[11723]);
     layer3_out[6847] <= ~(layer2_out[6007] | layer2_out[6008]);
     layer3_out[6848] <= ~(layer2_out[68] ^ layer2_out[69]);
     layer3_out[6849] <= ~layer2_out[642];
     layer3_out[6850] <= layer2_out[11676];
     layer3_out[6851] <= ~(layer2_out[477] | layer2_out[478]);
     layer3_out[6852] <= layer2_out[7598];
     layer3_out[6853] <= layer2_out[989];
     layer3_out[6854] <= ~(layer2_out[7703] | layer2_out[7704]);
     layer3_out[6855] <= ~layer2_out[8984];
     layer3_out[6856] <= layer2_out[8658];
     layer3_out[6857] <= ~layer2_out[11602];
     layer3_out[6858] <= ~layer2_out[615] | layer2_out[614];
     layer3_out[6859] <= layer2_out[8275] ^ layer2_out[8276];
     layer3_out[6860] <= layer2_out[7859] ^ layer2_out[7860];
     layer3_out[6861] <= ~(layer2_out[2470] ^ layer2_out[2471]);
     layer3_out[6862] <= layer2_out[6658];
     layer3_out[6863] <= layer2_out[5910];
     layer3_out[6864] <= layer2_out[645] ^ layer2_out[646];
     layer3_out[6865] <= ~layer2_out[4129];
     layer3_out[6866] <= layer2_out[10215];
     layer3_out[6867] <= ~layer2_out[2007];
     layer3_out[6868] <= ~layer2_out[8186] | layer2_out[8185];
     layer3_out[6869] <= layer2_out[4414] & ~layer2_out[4413];
     layer3_out[6870] <= layer2_out[6370];
     layer3_out[6871] <= layer2_out[10330] & layer2_out[10331];
     layer3_out[6872] <= ~layer2_out[446] | layer2_out[447];
     layer3_out[6873] <= layer2_out[1896] ^ layer2_out[1897];
     layer3_out[6874] <= layer2_out[3716] & ~layer2_out[3717];
     layer3_out[6875] <= ~layer2_out[9932] | layer2_out[9933];
     layer3_out[6876] <= ~layer2_out[3787];
     layer3_out[6877] <= layer2_out[2418];
     layer3_out[6878] <= layer2_out[1116];
     layer3_out[6879] <= layer2_out[2246] ^ layer2_out[2247];
     layer3_out[6880] <= ~(layer2_out[6612] & layer2_out[6613]);
     layer3_out[6881] <= ~layer2_out[9647] | layer2_out[9646];
     layer3_out[6882] <= ~(layer2_out[9596] & layer2_out[9597]);
     layer3_out[6883] <= layer2_out[6845];
     layer3_out[6884] <= layer2_out[11336] ^ layer2_out[11337];
     layer3_out[6885] <= layer2_out[5650];
     layer3_out[6886] <= ~layer2_out[10736];
     layer3_out[6887] <= layer2_out[8056] ^ layer2_out[8057];
     layer3_out[6888] <= ~(layer2_out[1910] ^ layer2_out[1911]);
     layer3_out[6889] <= ~layer2_out[4715];
     layer3_out[6890] <= layer2_out[10749];
     layer3_out[6891] <= layer2_out[11656];
     layer3_out[6892] <= layer2_out[6712] & ~layer2_out[6713];
     layer3_out[6893] <= ~layer2_out[4989] | layer2_out[4990];
     layer3_out[6894] <= ~(layer2_out[11732] & layer2_out[11733]);
     layer3_out[6895] <= layer2_out[5353] & ~layer2_out[5354];
     layer3_out[6896] <= layer2_out[8635] & layer2_out[8636];
     layer3_out[6897] <= ~layer2_out[7939];
     layer3_out[6898] <= layer2_out[9945];
     layer3_out[6899] <= layer2_out[7393] ^ layer2_out[7394];
     layer3_out[6900] <= ~(layer2_out[9108] ^ layer2_out[9109]);
     layer3_out[6901] <= layer2_out[4386] ^ layer2_out[4387];
     layer3_out[6902] <= ~(layer2_out[3933] ^ layer2_out[3934]);
     layer3_out[6903] <= layer2_out[186] & layer2_out[187];
     layer3_out[6904] <= ~(layer2_out[2991] | layer2_out[2992]);
     layer3_out[6905] <= ~(layer2_out[3408] & layer2_out[3409]);
     layer3_out[6906] <= layer2_out[6900] ^ layer2_out[6901];
     layer3_out[6907] <= layer2_out[5989] & ~layer2_out[5990];
     layer3_out[6908] <= layer2_out[1341] | layer2_out[1342];
     layer3_out[6909] <= ~layer2_out[3779];
     layer3_out[6910] <= layer2_out[6619] & ~layer2_out[6618];
     layer3_out[6911] <= ~(layer2_out[7894] ^ layer2_out[7895]);
     layer3_out[6912] <= ~(layer2_out[5278] & layer2_out[5279]);
     layer3_out[6913] <= ~layer2_out[9357];
     layer3_out[6914] <= ~layer2_out[68] | layer2_out[67];
     layer3_out[6915] <= ~(layer2_out[2584] | layer2_out[2585]);
     layer3_out[6916] <= layer2_out[10266] ^ layer2_out[10267];
     layer3_out[6917] <= layer2_out[1445] & layer2_out[1446];
     layer3_out[6918] <= ~layer2_out[11846] | layer2_out[11845];
     layer3_out[6919] <= layer2_out[326] & ~layer2_out[325];
     layer3_out[6920] <= ~layer2_out[8330];
     layer3_out[6921] <= ~(layer2_out[1874] ^ layer2_out[1875]);
     layer3_out[6922] <= layer2_out[2459] & ~layer2_out[2460];
     layer3_out[6923] <= layer2_out[2376] ^ layer2_out[2377];
     layer3_out[6924] <= ~layer2_out[2806] | layer2_out[2805];
     layer3_out[6925] <= layer2_out[4939];
     layer3_out[6926] <= ~(layer2_out[1018] ^ layer2_out[1019]);
     layer3_out[6927] <= ~(layer2_out[5143] ^ layer2_out[5144]);
     layer3_out[6928] <= ~(layer2_out[9155] & layer2_out[9156]);
     layer3_out[6929] <= ~layer2_out[4377] | layer2_out[4376];
     layer3_out[6930] <= ~layer2_out[4842] | layer2_out[4843];
     layer3_out[6931] <= ~(layer2_out[8] ^ layer2_out[9]);
     layer3_out[6932] <= ~(layer2_out[879] ^ layer2_out[880]);
     layer3_out[6933] <= layer2_out[5839];
     layer3_out[6934] <= layer2_out[1495] & ~layer2_out[1496];
     layer3_out[6935] <= ~(layer2_out[4179] & layer2_out[4180]);
     layer3_out[6936] <= ~layer2_out[4898];
     layer3_out[6937] <= ~layer2_out[2605];
     layer3_out[6938] <= ~layer2_out[1986];
     layer3_out[6939] <= ~layer2_out[1574] | layer2_out[1573];
     layer3_out[6940] <= ~layer2_out[4115] | layer2_out[4116];
     layer3_out[6941] <= ~layer2_out[3418] | layer2_out[3417];
     layer3_out[6942] <= ~layer2_out[6403] | layer2_out[6402];
     layer3_out[6943] <= layer2_out[236] ^ layer2_out[237];
     layer3_out[6944] <= layer2_out[2555];
     layer3_out[6945] <= layer2_out[6314];
     layer3_out[6946] <= ~layer2_out[5924];
     layer3_out[6947] <= ~(layer2_out[1881] & layer2_out[1882]);
     layer3_out[6948] <= ~layer2_out[4924] | layer2_out[4925];
     layer3_out[6949] <= layer2_out[10853] & layer2_out[10854];
     layer3_out[6950] <= ~(layer2_out[4765] ^ layer2_out[4766]);
     layer3_out[6951] <= layer2_out[7029];
     layer3_out[6952] <= ~(layer2_out[8615] ^ layer2_out[8616]);
     layer3_out[6953] <= layer2_out[11642];
     layer3_out[6954] <= ~layer2_out[5892];
     layer3_out[6955] <= layer2_out[3404] & ~layer2_out[3403];
     layer3_out[6956] <= ~(layer2_out[9844] ^ layer2_out[9845]);
     layer3_out[6957] <= ~layer2_out[10668];
     layer3_out[6958] <= layer2_out[7570] | layer2_out[7571];
     layer3_out[6959] <= layer2_out[2518];
     layer3_out[6960] <= ~(layer2_out[359] ^ layer2_out[360]);
     layer3_out[6961] <= layer2_out[6897];
     layer3_out[6962] <= layer2_out[6640];
     layer3_out[6963] <= ~(layer2_out[3632] & layer2_out[3633]);
     layer3_out[6964] <= layer2_out[11885];
     layer3_out[6965] <= ~layer2_out[8444] | layer2_out[8445];
     layer3_out[6966] <= layer2_out[5463] & ~layer2_out[5462];
     layer3_out[6967] <= ~(layer2_out[1978] ^ layer2_out[1979]);
     layer3_out[6968] <= ~layer2_out[1961];
     layer3_out[6969] <= ~(layer2_out[6730] ^ layer2_out[6731]);
     layer3_out[6970] <= layer2_out[735];
     layer3_out[6971] <= layer2_out[6342] | layer2_out[6343];
     layer3_out[6972] <= ~(layer2_out[4322] | layer2_out[4323]);
     layer3_out[6973] <= ~(layer2_out[3005] ^ layer2_out[3006]);
     layer3_out[6974] <= ~layer2_out[3182];
     layer3_out[6975] <= ~layer2_out[2032] | layer2_out[2033];
     layer3_out[6976] <= layer2_out[10866];
     layer3_out[6977] <= layer2_out[3789] ^ layer2_out[3790];
     layer3_out[6978] <= ~layer2_out[7287] | layer2_out[7288];
     layer3_out[6979] <= ~(layer2_out[358] | layer2_out[359]);
     layer3_out[6980] <= layer2_out[11734] ^ layer2_out[11735];
     layer3_out[6981] <= layer2_out[1444];
     layer3_out[6982] <= layer2_out[10264];
     layer3_out[6983] <= ~layer2_out[6391] | layer2_out[6390];
     layer3_out[6984] <= ~layer2_out[5194];
     layer3_out[6985] <= ~(layer2_out[6406] ^ layer2_out[6407]);
     layer3_out[6986] <= layer2_out[1926];
     layer3_out[6987] <= ~layer2_out[8835] | layer2_out[8834];
     layer3_out[6988] <= layer2_out[11669];
     layer3_out[6989] <= layer2_out[11049] ^ layer2_out[11050];
     layer3_out[6990] <= ~layer2_out[4406];
     layer3_out[6991] <= layer2_out[10684] ^ layer2_out[10685];
     layer3_out[6992] <= ~(layer2_out[10058] & layer2_out[10059]);
     layer3_out[6993] <= ~(layer2_out[8831] & layer2_out[8832]);
     layer3_out[6994] <= ~(layer2_out[5812] ^ layer2_out[5813]);
     layer3_out[6995] <= ~layer2_out[4197] | layer2_out[4196];
     layer3_out[6996] <= ~layer2_out[5712] | layer2_out[5711];
     layer3_out[6997] <= layer2_out[2093];
     layer3_out[6998] <= layer2_out[4415];
     layer3_out[6999] <= ~layer2_out[8298];
     layer3_out[7000] <= layer2_out[3061] | layer2_out[3062];
     layer3_out[7001] <= layer2_out[1213] | layer2_out[1214];
     layer3_out[7002] <= layer2_out[3657] ^ layer2_out[3658];
     layer3_out[7003] <= ~(layer2_out[5831] ^ layer2_out[5832]);
     layer3_out[7004] <= ~(layer2_out[10766] ^ layer2_out[10767]);
     layer3_out[7005] <= layer2_out[3621];
     layer3_out[7006] <= layer2_out[8309];
     layer3_out[7007] <= ~layer2_out[5236];
     layer3_out[7008] <= layer2_out[7419] & layer2_out[7420];
     layer3_out[7009] <= layer2_out[259] & layer2_out[260];
     layer3_out[7010] <= ~layer2_out[2345] | layer2_out[2346];
     layer3_out[7011] <= layer2_out[1351];
     layer3_out[7012] <= ~layer2_out[7297];
     layer3_out[7013] <= layer2_out[2752];
     layer3_out[7014] <= ~layer2_out[8404];
     layer3_out[7015] <= layer2_out[9101] & ~layer2_out[9100];
     layer3_out[7016] <= ~(layer2_out[6187] ^ layer2_out[6188]);
     layer3_out[7017] <= ~layer2_out[11711];
     layer3_out[7018] <= ~(layer2_out[7513] ^ layer2_out[7514]);
     layer3_out[7019] <= ~layer2_out[4185];
     layer3_out[7020] <= ~layer2_out[11215];
     layer3_out[7021] <= ~layer2_out[8075] | layer2_out[8074];
     layer3_out[7022] <= ~layer2_out[9803];
     layer3_out[7023] <= ~(layer2_out[3455] | layer2_out[3456]);
     layer3_out[7024] <= layer2_out[3244];
     layer3_out[7025] <= layer2_out[11911];
     layer3_out[7026] <= layer2_out[6424];
     layer3_out[7027] <= ~(layer2_out[8638] ^ layer2_out[8639]);
     layer3_out[7028] <= ~layer2_out[4890] | layer2_out[4891];
     layer3_out[7029] <= ~(layer2_out[11920] ^ layer2_out[11921]);
     layer3_out[7030] <= layer2_out[8694] & layer2_out[8695];
     layer3_out[7031] <= ~layer2_out[11782] | layer2_out[11781];
     layer3_out[7032] <= layer2_out[4955] & ~layer2_out[4954];
     layer3_out[7033] <= layer2_out[8026] & layer2_out[8027];
     layer3_out[7034] <= layer2_out[4195] | layer2_out[4196];
     layer3_out[7035] <= ~(layer2_out[2380] ^ layer2_out[2381]);
     layer3_out[7036] <= layer2_out[11212] & ~layer2_out[11211];
     layer3_out[7037] <= ~layer2_out[5922] | layer2_out[5923];
     layer3_out[7038] <= layer2_out[10252] & ~layer2_out[10253];
     layer3_out[7039] <= layer2_out[10198];
     layer3_out[7040] <= ~layer2_out[3031];
     layer3_out[7041] <= ~layer2_out[5686] | layer2_out[5687];
     layer3_out[7042] <= layer2_out[4628] | layer2_out[4629];
     layer3_out[7043] <= layer2_out[8017];
     layer3_out[7044] <= layer2_out[1811] ^ layer2_out[1812];
     layer3_out[7045] <= layer2_out[10439] | layer2_out[10440];
     layer3_out[7046] <= ~layer2_out[4165];
     layer3_out[7047] <= layer2_out[8234];
     layer3_out[7048] <= ~layer2_out[5077];
     layer3_out[7049] <= layer2_out[2123] & ~layer2_out[2124];
     layer3_out[7050] <= layer2_out[8576] | layer2_out[8577];
     layer3_out[7051] <= ~layer2_out[9867];
     layer3_out[7052] <= layer2_out[9713] ^ layer2_out[9714];
     layer3_out[7053] <= layer2_out[290] & ~layer2_out[291];
     layer3_out[7054] <= ~layer2_out[5997];
     layer3_out[7055] <= ~(layer2_out[11601] | layer2_out[11602]);
     layer3_out[7056] <= ~layer2_out[9812] | layer2_out[9811];
     layer3_out[7057] <= ~layer2_out[357];
     layer3_out[7058] <= layer2_out[1852];
     layer3_out[7059] <= ~(layer2_out[10188] ^ layer2_out[10189]);
     layer3_out[7060] <= layer2_out[6963] ^ layer2_out[6964];
     layer3_out[7061] <= layer2_out[4265] & layer2_out[4266];
     layer3_out[7062] <= layer2_out[5434];
     layer3_out[7063] <= ~(layer2_out[5204] ^ layer2_out[5205]);
     layer3_out[7064] <= layer2_out[4246] | layer2_out[4247];
     layer3_out[7065] <= layer2_out[3381] ^ layer2_out[3382];
     layer3_out[7066] <= layer2_out[2020];
     layer3_out[7067] <= ~(layer2_out[5248] ^ layer2_out[5249]);
     layer3_out[7068] <= layer2_out[3743];
     layer3_out[7069] <= layer2_out[2688];
     layer3_out[7070] <= layer2_out[9620] ^ layer2_out[9621];
     layer3_out[7071] <= layer2_out[6183];
     layer3_out[7072] <= ~(layer2_out[10177] | layer2_out[10178]);
     layer3_out[7073] <= ~layer2_out[2573] | layer2_out[2574];
     layer3_out[7074] <= layer2_out[7702] ^ layer2_out[7703];
     layer3_out[7075] <= ~layer2_out[10908];
     layer3_out[7076] <= layer2_out[8031] & layer2_out[8032];
     layer3_out[7077] <= ~(layer2_out[8104] ^ layer2_out[8105]);
     layer3_out[7078] <= layer2_out[4376] & ~layer2_out[4375];
     layer3_out[7079] <= layer2_out[6843];
     layer3_out[7080] <= layer2_out[11337];
     layer3_out[7081] <= ~layer2_out[1373] | layer2_out[1372];
     layer3_out[7082] <= layer2_out[1412] & layer2_out[1413];
     layer3_out[7083] <= layer2_out[5809] & layer2_out[5810];
     layer3_out[7084] <= layer2_out[465];
     layer3_out[7085] <= layer2_out[8868] ^ layer2_out[8869];
     layer3_out[7086] <= ~layer2_out[7444];
     layer3_out[7087] <= ~(layer2_out[2310] ^ layer2_out[2311]);
     layer3_out[7088] <= ~layer2_out[9037];
     layer3_out[7089] <= layer2_out[2034];
     layer3_out[7090] <= ~layer2_out[7659];
     layer3_out[7091] <= ~(layer2_out[8971] & layer2_out[8972]);
     layer3_out[7092] <= layer2_out[11126];
     layer3_out[7093] <= ~layer2_out[100];
     layer3_out[7094] <= ~(layer2_out[9465] ^ layer2_out[9466]);
     layer3_out[7095] <= layer2_out[6700] & ~layer2_out[6701];
     layer3_out[7096] <= ~layer2_out[4708] | layer2_out[4707];
     layer3_out[7097] <= layer2_out[10035];
     layer3_out[7098] <= layer2_out[1233];
     layer3_out[7099] <= ~(layer2_out[9925] & layer2_out[9926]);
     layer3_out[7100] <= ~layer2_out[6403];
     layer3_out[7101] <= ~layer2_out[6857];
     layer3_out[7102] <= ~layer2_out[9093];
     layer3_out[7103] <= layer2_out[7924];
     layer3_out[7104] <= ~(layer2_out[4144] ^ layer2_out[4145]);
     layer3_out[7105] <= ~(layer2_out[9163] ^ layer2_out[9164]);
     layer3_out[7106] <= layer2_out[1710] | layer2_out[1711];
     layer3_out[7107] <= layer2_out[3435] ^ layer2_out[3436];
     layer3_out[7108] <= layer2_out[6771] & ~layer2_out[6770];
     layer3_out[7109] <= layer2_out[11823];
     layer3_out[7110] <= layer2_out[407] ^ layer2_out[408];
     layer3_out[7111] <= layer2_out[10345];
     layer3_out[7112] <= ~(layer2_out[8019] | layer2_out[8020]);
     layer3_out[7113] <= ~layer2_out[537];
     layer3_out[7114] <= ~layer2_out[10810];
     layer3_out[7115] <= ~layer2_out[11473] | layer2_out[11474];
     layer3_out[7116] <= ~layer2_out[11135] | layer2_out[11136];
     layer3_out[7117] <= layer2_out[5774] & ~layer2_out[5773];
     layer3_out[7118] <= ~layer2_out[9516];
     layer3_out[7119] <= ~(layer2_out[10067] ^ layer2_out[10068]);
     layer3_out[7120] <= ~layer2_out[10973];
     layer3_out[7121] <= ~layer2_out[11025];
     layer3_out[7122] <= layer2_out[10413];
     layer3_out[7123] <= ~layer2_out[10511] | layer2_out[10512];
     layer3_out[7124] <= ~layer2_out[1860];
     layer3_out[7125] <= ~layer2_out[8142] | layer2_out[8141];
     layer3_out[7126] <= ~layer2_out[4741];
     layer3_out[7127] <= ~(layer2_out[11975] ^ layer2_out[11976]);
     layer3_out[7128] <= layer2_out[4763];
     layer3_out[7129] <= layer2_out[6003] | layer2_out[6004];
     layer3_out[7130] <= ~(layer2_out[1317] & layer2_out[1318]);
     layer3_out[7131] <= layer2_out[3190];
     layer3_out[7132] <= layer2_out[11718];
     layer3_out[7133] <= ~(layer2_out[5234] ^ layer2_out[5235]);
     layer3_out[7134] <= ~layer2_out[4301];
     layer3_out[7135] <= ~(layer2_out[5865] | layer2_out[5866]);
     layer3_out[7136] <= ~layer2_out[6580];
     layer3_out[7137] <= ~(layer2_out[2414] | layer2_out[2415]);
     layer3_out[7138] <= layer2_out[3965] | layer2_out[3966];
     layer3_out[7139] <= layer2_out[3752] & ~layer2_out[3751];
     layer3_out[7140] <= layer2_out[4957];
     layer3_out[7141] <= layer2_out[5605] & ~layer2_out[5604];
     layer3_out[7142] <= layer2_out[1517] & layer2_out[1518];
     layer3_out[7143] <= layer2_out[10385] & ~layer2_out[10386];
     layer3_out[7144] <= ~(layer2_out[3558] ^ layer2_out[3559]);
     layer3_out[7145] <= ~(layer2_out[6418] ^ layer2_out[6419]);
     layer3_out[7146] <= ~(layer2_out[5098] | layer2_out[5099]);
     layer3_out[7147] <= ~layer2_out[3004];
     layer3_out[7148] <= ~layer2_out[9759];
     layer3_out[7149] <= ~(layer2_out[10725] ^ layer2_out[10726]);
     layer3_out[7150] <= ~layer2_out[1535];
     layer3_out[7151] <= layer2_out[8138];
     layer3_out[7152] <= ~layer2_out[424];
     layer3_out[7153] <= layer2_out[10985] & ~layer2_out[10986];
     layer3_out[7154] <= ~layer2_out[1279];
     layer3_out[7155] <= ~layer2_out[1304];
     layer3_out[7156] <= ~(layer2_out[2082] | layer2_out[2083]);
     layer3_out[7157] <= layer2_out[4974];
     layer3_out[7158] <= ~layer2_out[3066] | layer2_out[3067];
     layer3_out[7159] <= ~layer2_out[4995];
     layer3_out[7160] <= ~(layer2_out[10069] & layer2_out[10070]);
     layer3_out[7161] <= ~layer2_out[7659];
     layer3_out[7162] <= layer2_out[7319] ^ layer2_out[7320];
     layer3_out[7163] <= layer2_out[3621];
     layer3_out[7164] <= layer2_out[10718];
     layer3_out[7165] <= ~layer2_out[10139];
     layer3_out[7166] <= layer2_out[3431] & layer2_out[3432];
     layer3_out[7167] <= layer2_out[3907];
     layer3_out[7168] <= layer2_out[2337] ^ layer2_out[2338];
     layer3_out[7169] <= ~layer2_out[4574];
     layer3_out[7170] <= layer2_out[4671];
     layer3_out[7171] <= ~layer2_out[2665];
     layer3_out[7172] <= ~layer2_out[6827];
     layer3_out[7173] <= ~layer2_out[4449];
     layer3_out[7174] <= layer2_out[3052] ^ layer2_out[3053];
     layer3_out[7175] <= layer2_out[9674] & ~layer2_out[9673];
     layer3_out[7176] <= ~layer2_out[1050] | layer2_out[1049];
     layer3_out[7177] <= ~(layer2_out[3559] | layer2_out[3560]);
     layer3_out[7178] <= ~layer2_out[8046];
     layer3_out[7179] <= layer2_out[7969] | layer2_out[7970];
     layer3_out[7180] <= layer2_out[4914];
     layer3_out[7181] <= ~(layer2_out[1820] | layer2_out[1821]);
     layer3_out[7182] <= ~layer2_out[9982];
     layer3_out[7183] <= layer2_out[7861];
     layer3_out[7184] <= layer2_out[2287];
     layer3_out[7185] <= layer2_out[9562] ^ layer2_out[9563];
     layer3_out[7186] <= ~(layer2_out[4727] & layer2_out[4728]);
     layer3_out[7187] <= layer2_out[10888] | layer2_out[10889];
     layer3_out[7188] <= layer2_out[1775] & layer2_out[1776];
     layer3_out[7189] <= layer2_out[8369] & ~layer2_out[8368];
     layer3_out[7190] <= layer2_out[9528] | layer2_out[9529];
     layer3_out[7191] <= layer2_out[1947];
     layer3_out[7192] <= layer2_out[3926] & ~layer2_out[3927];
     layer3_out[7193] <= ~layer2_out[603];
     layer3_out[7194] <= ~layer2_out[1892] | layer2_out[1893];
     layer3_out[7195] <= layer2_out[8666] & layer2_out[8667];
     layer3_out[7196] <= ~layer2_out[11733];
     layer3_out[7197] <= ~layer2_out[11143];
     layer3_out[7198] <= ~layer2_out[9578] | layer2_out[9579];
     layer3_out[7199] <= layer2_out[10332] ^ layer2_out[10333];
     layer3_out[7200] <= ~layer2_out[5629];
     layer3_out[7201] <= ~layer2_out[11406];
     layer3_out[7202] <= ~layer2_out[3317];
     layer3_out[7203] <= layer2_out[11159] & ~layer2_out[11158];
     layer3_out[7204] <= layer2_out[8317];
     layer3_out[7205] <= ~layer2_out[240];
     layer3_out[7206] <= ~layer2_out[3776];
     layer3_out[7207] <= layer2_out[3058];
     layer3_out[7208] <= ~(layer2_out[4197] | layer2_out[4198]);
     layer3_out[7209] <= ~(layer2_out[11953] | layer2_out[11954]);
     layer3_out[7210] <= ~layer2_out[2331];
     layer3_out[7211] <= layer2_out[11206] ^ layer2_out[11207];
     layer3_out[7212] <= layer2_out[11503] | layer2_out[11504];
     layer3_out[7213] <= layer2_out[1349] ^ layer2_out[1350];
     layer3_out[7214] <= layer2_out[11997] & ~layer2_out[11998];
     layer3_out[7215] <= layer2_out[10592];
     layer3_out[7216] <= ~layer2_out[4459];
     layer3_out[7217] <= ~layer2_out[10032];
     layer3_out[7218] <= layer2_out[2011];
     layer3_out[7219] <= layer2_out[7971] & ~layer2_out[7970];
     layer3_out[7220] <= ~layer2_out[3217];
     layer3_out[7221] <= layer2_out[10488] & layer2_out[10489];
     layer3_out[7222] <= layer2_out[10763];
     layer3_out[7223] <= ~layer2_out[3144];
     layer3_out[7224] <= layer2_out[4709];
     layer3_out[7225] <= layer2_out[1496] & ~layer2_out[1497];
     layer3_out[7226] <= ~(layer2_out[2531] ^ layer2_out[2532]);
     layer3_out[7227] <= ~(layer2_out[4445] | layer2_out[4446]);
     layer3_out[7228] <= layer2_out[6988] ^ layer2_out[6989];
     layer3_out[7229] <= ~layer2_out[6040];
     layer3_out[7230] <= layer2_out[2] & layer2_out[3];
     layer3_out[7231] <= ~layer2_out[9583];
     layer3_out[7232] <= ~(layer2_out[3953] | layer2_out[3954]);
     layer3_out[7233] <= layer2_out[3738];
     layer3_out[7234] <= layer2_out[2604] & ~layer2_out[2603];
     layer3_out[7235] <= ~(layer2_out[4379] ^ layer2_out[4380]);
     layer3_out[7236] <= layer2_out[10445];
     layer3_out[7237] <= layer2_out[9496] ^ layer2_out[9497];
     layer3_out[7238] <= ~layer2_out[4363];
     layer3_out[7239] <= ~layer2_out[6331];
     layer3_out[7240] <= ~layer2_out[2478];
     layer3_out[7241] <= layer2_out[158] & ~layer2_out[157];
     layer3_out[7242] <= layer2_out[3542] & layer2_out[3543];
     layer3_out[7243] <= layer2_out[4256] & layer2_out[4257];
     layer3_out[7244] <= layer2_out[5779];
     layer3_out[7245] <= ~layer2_out[394];
     layer3_out[7246] <= layer2_out[9319];
     layer3_out[7247] <= layer2_out[6704];
     layer3_out[7248] <= ~(layer2_out[4772] & layer2_out[4773]);
     layer3_out[7249] <= layer2_out[113] ^ layer2_out[114];
     layer3_out[7250] <= ~layer2_out[566];
     layer3_out[7251] <= ~(layer2_out[3604] ^ layer2_out[3605]);
     layer3_out[7252] <= ~(layer2_out[4667] | layer2_out[4668]);
     layer3_out[7253] <= layer2_out[6505];
     layer3_out[7254] <= layer2_out[72];
     layer3_out[7255] <= layer2_out[10752] & ~layer2_out[10751];
     layer3_out[7256] <= layer2_out[9495];
     layer3_out[7257] <= layer2_out[6577] & ~layer2_out[6576];
     layer3_out[7258] <= layer2_out[699] & ~layer2_out[698];
     layer3_out[7259] <= ~layer2_out[7089];
     layer3_out[7260] <= layer2_out[10581] ^ layer2_out[10582];
     layer3_out[7261] <= layer2_out[7739] & ~layer2_out[7740];
     layer3_out[7262] <= ~layer2_out[4200];
     layer3_out[7263] <= layer2_out[11718];
     layer3_out[7264] <= layer2_out[5806] & ~layer2_out[5805];
     layer3_out[7265] <= layer2_out[2806];
     layer3_out[7266] <= layer2_out[1691] & layer2_out[1692];
     layer3_out[7267] <= layer2_out[9231] & ~layer2_out[9230];
     layer3_out[7268] <= ~(layer2_out[4750] ^ layer2_out[4751]);
     layer3_out[7269] <= layer2_out[676];
     layer3_out[7270] <= ~layer2_out[2111];
     layer3_out[7271] <= layer2_out[4583] & ~layer2_out[4582];
     layer3_out[7272] <= layer2_out[8598] & ~layer2_out[8599];
     layer3_out[7273] <= layer2_out[6769] & ~layer2_out[6770];
     layer3_out[7274] <= ~layer2_out[3588];
     layer3_out[7275] <= layer2_out[6504];
     layer3_out[7276] <= layer2_out[7725] ^ layer2_out[7726];
     layer3_out[7277] <= layer2_out[6030] & ~layer2_out[6029];
     layer3_out[7278] <= ~layer2_out[3884];
     layer3_out[7279] <= ~layer2_out[6340];
     layer3_out[7280] <= layer2_out[4632] & layer2_out[4633];
     layer3_out[7281] <= layer2_out[1292];
     layer3_out[7282] <= ~layer2_out[2118];
     layer3_out[7283] <= ~(layer2_out[9686] & layer2_out[9687]);
     layer3_out[7284] <= layer2_out[3802] & ~layer2_out[3803];
     layer3_out[7285] <= ~layer2_out[7346];
     layer3_out[7286] <= ~(layer2_out[2968] ^ layer2_out[2969]);
     layer3_out[7287] <= ~(layer2_out[3224] & layer2_out[3225]);
     layer3_out[7288] <= ~layer2_out[2329];
     layer3_out[7289] <= layer2_out[9237] & ~layer2_out[9238];
     layer3_out[7290] <= layer2_out[9397] & ~layer2_out[9398];
     layer3_out[7291] <= layer2_out[4654] & layer2_out[4655];
     layer3_out[7292] <= layer2_out[3291] & ~layer2_out[3290];
     layer3_out[7293] <= layer2_out[6220] & ~layer2_out[6219];
     layer3_out[7294] <= ~(layer2_out[8295] | layer2_out[8296]);
     layer3_out[7295] <= ~(layer2_out[11326] ^ layer2_out[11327]);
     layer3_out[7296] <= layer2_out[3154] & layer2_out[3155];
     layer3_out[7297] <= layer2_out[386];
     layer3_out[7298] <= layer2_out[4279] & layer2_out[4280];
     layer3_out[7299] <= layer2_out[10708];
     layer3_out[7300] <= layer2_out[2674] & ~layer2_out[2673];
     layer3_out[7301] <= layer2_out[10111] & ~layer2_out[10110];
     layer3_out[7302] <= layer2_out[8540] ^ layer2_out[8541];
     layer3_out[7303] <= layer2_out[9392];
     layer3_out[7304] <= layer2_out[5880] & ~layer2_out[5881];
     layer3_out[7305] <= ~(layer2_out[10983] ^ layer2_out[10984]);
     layer3_out[7306] <= layer2_out[7729];
     layer3_out[7307] <= ~layer2_out[1715] | layer2_out[1716];
     layer3_out[7308] <= layer2_out[10455];
     layer3_out[7309] <= layer2_out[9113];
     layer3_out[7310] <= layer2_out[8340] | layer2_out[8341];
     layer3_out[7311] <= layer2_out[11109];
     layer3_out[7312] <= ~layer2_out[4668];
     layer3_out[7313] <= layer2_out[4075] ^ layer2_out[4076];
     layer3_out[7314] <= layer2_out[4830];
     layer3_out[7315] <= ~(layer2_out[419] | layer2_out[420]);
     layer3_out[7316] <= layer2_out[4339] & ~layer2_out[4338];
     layer3_out[7317] <= layer2_out[9543] & ~layer2_out[9544];
     layer3_out[7318] <= layer2_out[8198] & layer2_out[8199];
     layer3_out[7319] <= ~layer2_out[7327];
     layer3_out[7320] <= ~layer2_out[2967];
     layer3_out[7321] <= layer2_out[4268] & layer2_out[4269];
     layer3_out[7322] <= layer2_out[3270];
     layer3_out[7323] <= ~layer2_out[5842];
     layer3_out[7324] <= ~layer2_out[3935];
     layer3_out[7325] <= layer2_out[802];
     layer3_out[7326] <= ~(layer2_out[6868] | layer2_out[6869]);
     layer3_out[7327] <= layer2_out[5427] & ~layer2_out[5428];
     layer3_out[7328] <= layer2_out[8520];
     layer3_out[7329] <= layer2_out[2402];
     layer3_out[7330] <= layer2_out[3309] | layer2_out[3310];
     layer3_out[7331] <= layer2_out[11134];
     layer3_out[7332] <= layer2_out[2348] | layer2_out[2349];
     layer3_out[7333] <= ~(layer2_out[4996] | layer2_out[4997]);
     layer3_out[7334] <= ~layer2_out[4217] | layer2_out[4216];
     layer3_out[7335] <= ~layer2_out[11066] | layer2_out[11067];
     layer3_out[7336] <= ~layer2_out[11181] | layer2_out[11180];
     layer3_out[7337] <= layer2_out[11434];
     layer3_out[7338] <= ~layer2_out[7436];
     layer3_out[7339] <= layer2_out[6453] & layer2_out[6454];
     layer3_out[7340] <= layer2_out[495];
     layer3_out[7341] <= ~layer2_out[6292];
     layer3_out[7342] <= layer2_out[1869] ^ layer2_out[1870];
     layer3_out[7343] <= ~(layer2_out[5556] | layer2_out[5557]);
     layer3_out[7344] <= ~(layer2_out[3571] ^ layer2_out[3572]);
     layer3_out[7345] <= layer2_out[1769] & ~layer2_out[1768];
     layer3_out[7346] <= layer2_out[1511];
     layer3_out[7347] <= layer2_out[5923];
     layer3_out[7348] <= layer2_out[11361] & ~layer2_out[11362];
     layer3_out[7349] <= layer2_out[4225] & layer2_out[4226];
     layer3_out[7350] <= layer2_out[8848] & layer2_out[8849];
     layer3_out[7351] <= ~layer2_out[8552];
     layer3_out[7352] <= layer2_out[695] & layer2_out[696];
     layer3_out[7353] <= layer2_out[5061];
     layer3_out[7354] <= layer2_out[3710];
     layer3_out[7355] <= ~(layer2_out[7260] | layer2_out[7261]);
     layer3_out[7356] <= ~layer2_out[9809];
     layer3_out[7357] <= layer2_out[3649] ^ layer2_out[3650];
     layer3_out[7358] <= layer2_out[2845];
     layer3_out[7359] <= layer2_out[9729];
     layer3_out[7360] <= layer2_out[6862];
     layer3_out[7361] <= ~(layer2_out[3648] | layer2_out[3649]);
     layer3_out[7362] <= layer2_out[9197];
     layer3_out[7363] <= layer2_out[10343];
     layer3_out[7364] <= layer2_out[1281] & ~layer2_out[1282];
     layer3_out[7365] <= layer2_out[4182] | layer2_out[4183];
     layer3_out[7366] <= ~layer2_out[2905];
     layer3_out[7367] <= layer2_out[5209] & ~layer2_out[5210];
     layer3_out[7368] <= layer2_out[7455] & layer2_out[7456];
     layer3_out[7369] <= layer2_out[9018];
     layer3_out[7370] <= layer2_out[9804] & layer2_out[9805];
     layer3_out[7371] <= layer2_out[3084] & ~layer2_out[3085];
     layer3_out[7372] <= ~(layer2_out[2999] | layer2_out[3000]);
     layer3_out[7373] <= ~layer2_out[9400];
     layer3_out[7374] <= ~layer2_out[1900];
     layer3_out[7375] <= layer2_out[5616];
     layer3_out[7376] <= ~layer2_out[8299];
     layer3_out[7377] <= ~layer2_out[1850];
     layer3_out[7378] <= layer2_out[6812] & layer2_out[6813];
     layer3_out[7379] <= layer2_out[7865] ^ layer2_out[7866];
     layer3_out[7380] <= layer2_out[5899];
     layer3_out[7381] <= layer2_out[5736] & layer2_out[5737];
     layer3_out[7382] <= ~(layer2_out[5926] | layer2_out[5927]);
     layer3_out[7383] <= layer2_out[786];
     layer3_out[7384] <= layer2_out[1570] ^ layer2_out[1571];
     layer3_out[7385] <= layer2_out[11597] & layer2_out[11598];
     layer3_out[7386] <= layer2_out[6908];
     layer3_out[7387] <= layer2_out[5212];
     layer3_out[7388] <= layer2_out[11624] & ~layer2_out[11623];
     layer3_out[7389] <= ~(layer2_out[9306] | layer2_out[9307]);
     layer3_out[7390] <= ~layer2_out[6615] | layer2_out[6614];
     layer3_out[7391] <= layer2_out[6284];
     layer3_out[7392] <= ~layer2_out[6092];
     layer3_out[7393] <= layer2_out[2358] & layer2_out[2359];
     layer3_out[7394] <= layer2_out[8323] & layer2_out[8324];
     layer3_out[7395] <= layer2_out[1803];
     layer3_out[7396] <= layer2_out[10531];
     layer3_out[7397] <= ~layer2_out[8823] | layer2_out[8824];
     layer3_out[7398] <= ~layer2_out[7524];
     layer3_out[7399] <= layer2_out[2138];
     layer3_out[7400] <= layer2_out[731];
     layer3_out[7401] <= layer2_out[7388];
     layer3_out[7402] <= layer2_out[9297];
     layer3_out[7403] <= layer2_out[3221] | layer2_out[3222];
     layer3_out[7404] <= ~layer2_out[9864];
     layer3_out[7405] <= layer2_out[10565] & ~layer2_out[10566];
     layer3_out[7406] <= ~(layer2_out[1521] | layer2_out[1522]);
     layer3_out[7407] <= layer2_out[5051] & layer2_out[5052];
     layer3_out[7408] <= layer2_out[1602];
     layer3_out[7409] <= layer2_out[9041] & layer2_out[9042];
     layer3_out[7410] <= layer2_out[8388] ^ layer2_out[8389];
     layer3_out[7411] <= ~(layer2_out[680] | layer2_out[681]);
     layer3_out[7412] <= layer2_out[11351];
     layer3_out[7413] <= layer2_out[4245];
     layer3_out[7414] <= ~layer2_out[5352];
     layer3_out[7415] <= ~layer2_out[1999];
     layer3_out[7416] <= layer2_out[5531] & ~layer2_out[5530];
     layer3_out[7417] <= layer2_out[4697] & layer2_out[4698];
     layer3_out[7418] <= ~layer2_out[3592];
     layer3_out[7419] <= layer2_out[7996] & layer2_out[7997];
     layer3_out[7420] <= layer2_out[9920] & layer2_out[9921];
     layer3_out[7421] <= ~layer2_out[5038];
     layer3_out[7422] <= layer2_out[4367];
     layer3_out[7423] <= ~(layer2_out[11166] | layer2_out[11167]);
     layer3_out[7424] <= layer2_out[6487];
     layer3_out[7425] <= layer2_out[9904] & ~layer2_out[9905];
     layer3_out[7426] <= layer2_out[5620] ^ layer2_out[5621];
     layer3_out[7427] <= layer2_out[11986];
     layer3_out[7428] <= layer2_out[2793] & ~layer2_out[2792];
     layer3_out[7429] <= layer2_out[6388];
     layer3_out[7430] <= layer2_out[9782] & layer2_out[9783];
     layer3_out[7431] <= layer2_out[1516] & layer2_out[1517];
     layer3_out[7432] <= ~(layer2_out[8261] | layer2_out[8262]);
     layer3_out[7433] <= ~layer2_out[9206];
     layer3_out[7434] <= layer2_out[7180];
     layer3_out[7435] <= layer2_out[1650] & ~layer2_out[1649];
     layer3_out[7436] <= ~layer2_out[6206];
     layer3_out[7437] <= layer2_out[5565] & ~layer2_out[5564];
     layer3_out[7438] <= ~(layer2_out[10814] | layer2_out[10815]);
     layer3_out[7439] <= ~layer2_out[7791];
     layer3_out[7440] <= layer2_out[11746];
     layer3_out[7441] <= layer2_out[2868];
     layer3_out[7442] <= ~layer2_out[5230];
     layer3_out[7443] <= layer2_out[4504];
     layer3_out[7444] <= ~layer2_out[3340];
     layer3_out[7445] <= layer2_out[4137] ^ layer2_out[4138];
     layer3_out[7446] <= layer2_out[4889];
     layer3_out[7447] <= layer2_out[6953];
     layer3_out[7448] <= ~(layer2_out[6622] | layer2_out[6623]);
     layer3_out[7449] <= ~layer2_out[7883];
     layer3_out[7450] <= layer2_out[5048] ^ layer2_out[5049];
     layer3_out[7451] <= ~layer2_out[236];
     layer3_out[7452] <= ~layer2_out[442];
     layer3_out[7453] <= ~layer2_out[7479];
     layer3_out[7454] <= ~(layer2_out[416] ^ layer2_out[417]);
     layer3_out[7455] <= layer2_out[7990] & ~layer2_out[7991];
     layer3_out[7456] <= layer2_out[4893] | layer2_out[4894];
     layer3_out[7457] <= layer2_out[392] ^ layer2_out[393];
     layer3_out[7458] <= ~layer2_out[4136];
     layer3_out[7459] <= ~layer2_out[5655];
     layer3_out[7460] <= layer2_out[4133];
     layer3_out[7461] <= ~(layer2_out[4651] ^ layer2_out[4652]);
     layer3_out[7462] <= ~(layer2_out[6056] | layer2_out[6057]);
     layer3_out[7463] <= layer2_out[7231];
     layer3_out[7464] <= layer2_out[11237];
     layer3_out[7465] <= ~(layer2_out[10128] ^ layer2_out[10129]);
     layer3_out[7466] <= layer2_out[10590] | layer2_out[10591];
     layer3_out[7467] <= ~layer2_out[3961];
     layer3_out[7468] <= ~(layer2_out[3941] | layer2_out[3942]);
     layer3_out[7469] <= ~(layer2_out[450] | layer2_out[451]);
     layer3_out[7470] <= layer2_out[10026] & ~layer2_out[10025];
     layer3_out[7471] <= layer2_out[7015];
     layer3_out[7472] <= layer2_out[6695];
     layer3_out[7473] <= layer2_out[11446] & layer2_out[11447];
     layer3_out[7474] <= ~layer2_out[364];
     layer3_out[7475] <= ~layer2_out[11227] | layer2_out[11226];
     layer3_out[7476] <= ~(layer2_out[7849] | layer2_out[7850]);
     layer3_out[7477] <= layer2_out[6385] ^ layer2_out[6386];
     layer3_out[7478] <= ~(layer2_out[5219] | layer2_out[5220]);
     layer3_out[7479] <= ~layer2_out[1333];
     layer3_out[7480] <= layer2_out[10364];
     layer3_out[7481] <= layer2_out[6661];
     layer3_out[7482] <= ~layer2_out[7819];
     layer3_out[7483] <= ~layer2_out[3191];
     layer3_out[7484] <= ~layer2_out[1744];
     layer3_out[7485] <= layer2_out[1777] & ~layer2_out[1778];
     layer3_out[7486] <= layer2_out[6950];
     layer3_out[7487] <= layer2_out[11577] & ~layer2_out[11578];
     layer3_out[7488] <= layer2_out[2681] & ~layer2_out[2682];
     layer3_out[7489] <= ~layer2_out[1727];
     layer3_out[7490] <= ~(layer2_out[6513] ^ layer2_out[6514]);
     layer3_out[7491] <= layer2_out[1878] & layer2_out[1879];
     layer3_out[7492] <= layer2_out[5783] & ~layer2_out[5784];
     layer3_out[7493] <= ~(layer2_out[10217] ^ layer2_out[10218]);
     layer3_out[7494] <= ~(layer2_out[6004] ^ layer2_out[6005]);
     layer3_out[7495] <= layer2_out[2887] & ~layer2_out[2888];
     layer3_out[7496] <= ~layer2_out[11150];
     layer3_out[7497] <= layer2_out[554] & ~layer2_out[553];
     layer3_out[7498] <= layer2_out[10511] & ~layer2_out[10510];
     layer3_out[7499] <= ~(layer2_out[4822] | layer2_out[4823]);
     layer3_out[7500] <= layer2_out[2138];
     layer3_out[7501] <= layer2_out[10541] & layer2_out[10542];
     layer3_out[7502] <= ~(layer2_out[3846] ^ layer2_out[3847]);
     layer3_out[7503] <= ~layer2_out[3212];
     layer3_out[7504] <= ~(layer2_out[9454] ^ layer2_out[9455]);
     layer3_out[7505] <= ~layer2_out[6630];
     layer3_out[7506] <= layer2_out[7461];
     layer3_out[7507] <= ~layer2_out[7277] | layer2_out[7278];
     layer3_out[7508] <= ~layer2_out[599] | layer2_out[598];
     layer3_out[7509] <= ~(layer2_out[11161] | layer2_out[11162]);
     layer3_out[7510] <= ~(layer2_out[205] | layer2_out[206]);
     layer3_out[7511] <= layer2_out[8288];
     layer3_out[7512] <= layer2_out[620] & ~layer2_out[619];
     layer3_out[7513] <= layer2_out[4835] | layer2_out[4836];
     layer3_out[7514] <= layer2_out[2401] & layer2_out[2402];
     layer3_out[7515] <= layer2_out[11177] & ~layer2_out[11176];
     layer3_out[7516] <= layer2_out[9570];
     layer3_out[7517] <= layer2_out[5715] & ~layer2_out[5716];
     layer3_out[7518] <= ~layer2_out[1330];
     layer3_out[7519] <= ~(layer2_out[7112] ^ layer2_out[7113]);
     layer3_out[7520] <= ~(layer2_out[10267] | layer2_out[10268]);
     layer3_out[7521] <= layer2_out[2183];
     layer3_out[7522] <= ~layer2_out[539];
     layer3_out[7523] <= layer2_out[917] & layer2_out[918];
     layer3_out[7524] <= ~(layer2_out[4576] ^ layer2_out[4577]);
     layer3_out[7525] <= ~layer2_out[11937];
     layer3_out[7526] <= layer2_out[11994] & ~layer2_out[11993];
     layer3_out[7527] <= layer2_out[10138];
     layer3_out[7528] <= layer2_out[5812];
     layer3_out[7529] <= layer2_out[352] | layer2_out[353];
     layer3_out[7530] <= layer2_out[7453] & ~layer2_out[7454];
     layer3_out[7531] <= layer2_out[8534];
     layer3_out[7532] <= ~(layer2_out[4009] & layer2_out[4010]);
     layer3_out[7533] <= layer2_out[1757] & ~layer2_out[1756];
     layer3_out[7534] <= layer2_out[8321] & ~layer2_out[8320];
     layer3_out[7535] <= layer2_out[5060] & layer2_out[5061];
     layer3_out[7536] <= layer2_out[5185] ^ layer2_out[5186];
     layer3_out[7537] <= ~layer2_out[5521];
     layer3_out[7538] <= layer2_out[8667] & ~layer2_out[8668];
     layer3_out[7539] <= layer2_out[1993] ^ layer2_out[1994];
     layer3_out[7540] <= ~layer2_out[4767];
     layer3_out[7541] <= ~layer2_out[5021] | layer2_out[5022];
     layer3_out[7542] <= layer2_out[895];
     layer3_out[7543] <= layer2_out[7001] & layer2_out[7002];
     layer3_out[7544] <= layer2_out[5332] & layer2_out[5333];
     layer3_out[7545] <= ~layer2_out[11460];
     layer3_out[7546] <= ~layer2_out[5967];
     layer3_out[7547] <= layer2_out[10384];
     layer3_out[7548] <= layer2_out[318] & ~layer2_out[319];
     layer3_out[7549] <= layer2_out[8362] & layer2_out[8363];
     layer3_out[7550] <= ~layer2_out[6247];
     layer3_out[7551] <= layer2_out[2408] & ~layer2_out[2409];
     layer3_out[7552] <= layer2_out[6011] & ~layer2_out[6012];
     layer3_out[7553] <= layer2_out[2560] & ~layer2_out[2559];
     layer3_out[7554] <= ~layer2_out[982] | layer2_out[983];
     layer3_out[7555] <= layer2_out[10361] & ~layer2_out[10362];
     layer3_out[7556] <= ~layer2_out[7252] | layer2_out[7251];
     layer3_out[7557] <= ~(layer2_out[8866] | layer2_out[8867]);
     layer3_out[7558] <= ~(layer2_out[4482] | layer2_out[4483]);
     layer3_out[7559] <= layer2_out[1161] & ~layer2_out[1162];
     layer3_out[7560] <= layer2_out[6588] ^ layer2_out[6589];
     layer3_out[7561] <= layer2_out[7521] & layer2_out[7522];
     layer3_out[7562] <= ~layer2_out[2355];
     layer3_out[7563] <= ~(layer2_out[11254] | layer2_out[11255]);
     layer3_out[7564] <= ~layer2_out[7107];
     layer3_out[7565] <= layer2_out[3780] & layer2_out[3781];
     layer3_out[7566] <= ~layer2_out[9795];
     layer3_out[7567] <= layer2_out[3305];
     layer3_out[7568] <= layer2_out[6255] ^ layer2_out[6256];
     layer3_out[7569] <= layer2_out[487];
     layer3_out[7570] <= layer2_out[3857] & layer2_out[3858];
     layer3_out[7571] <= ~layer2_out[253];
     layer3_out[7572] <= layer2_out[5397];
     layer3_out[7573] <= layer2_out[10803];
     layer3_out[7574] <= ~(layer2_out[8767] | layer2_out[8768]);
     layer3_out[7575] <= layer2_out[11751] ^ layer2_out[11752];
     layer3_out[7576] <= layer2_out[2872] & layer2_out[2873];
     layer3_out[7577] <= layer2_out[5882];
     layer3_out[7578] <= layer2_out[7240] & layer2_out[7241];
     layer3_out[7579] <= ~(layer2_out[1045] | layer2_out[1046]);
     layer3_out[7580] <= layer2_out[5751];
     layer3_out[7581] <= layer2_out[6481] & layer2_out[6482];
     layer3_out[7582] <= layer2_out[1568];
     layer3_out[7583] <= layer2_out[11620];
     layer3_out[7584] <= layer2_out[7475] & layer2_out[7476];
     layer3_out[7585] <= layer2_out[3839] & ~layer2_out[3840];
     layer3_out[7586] <= layer2_out[7788] ^ layer2_out[7789];
     layer3_out[7587] <= ~(layer2_out[4767] | layer2_out[4768]);
     layer3_out[7588] <= ~layer2_out[3209];
     layer3_out[7589] <= ~(layer2_out[9684] ^ layer2_out[9685]);
     layer3_out[7590] <= ~layer2_out[1969];
     layer3_out[7591] <= layer2_out[1916] & ~layer2_out[1917];
     layer3_out[7592] <= layer2_out[5150] & layer2_out[5151];
     layer3_out[7593] <= layer2_out[1832] ^ layer2_out[1833];
     layer3_out[7594] <= ~(layer2_out[3473] | layer2_out[3474]);
     layer3_out[7595] <= layer2_out[11778] & ~layer2_out[11777];
     layer3_out[7596] <= layer2_out[4984];
     layer3_out[7597] <= layer2_out[5178];
     layer3_out[7598] <= layer2_out[4835];
     layer3_out[7599] <= layer2_out[4894] & layer2_out[4895];
     layer3_out[7600] <= ~(layer2_out[451] | layer2_out[452]);
     layer3_out[7601] <= layer2_out[11396] | layer2_out[11397];
     layer3_out[7602] <= ~layer2_out[3000];
     layer3_out[7603] <= layer2_out[8896];
     layer3_out[7604] <= layer2_out[554] & layer2_out[555];
     layer3_out[7605] <= layer2_out[1734] | layer2_out[1735];
     layer3_out[7606] <= layer2_out[11754] & layer2_out[11755];
     layer3_out[7607] <= ~(layer2_out[8242] | layer2_out[8243]);
     layer3_out[7608] <= layer2_out[3811] & ~layer2_out[3810];
     layer3_out[7609] <= layer2_out[4580];
     layer3_out[7610] <= ~(layer2_out[8594] ^ layer2_out[8595]);
     layer3_out[7611] <= layer2_out[9600] & layer2_out[9601];
     layer3_out[7612] <= ~layer2_out[2995];
     layer3_out[7613] <= layer2_out[10023] & ~layer2_out[10022];
     layer3_out[7614] <= ~layer2_out[1407];
     layer3_out[7615] <= ~layer2_out[335];
     layer3_out[7616] <= ~layer2_out[1008] | layer2_out[1009];
     layer3_out[7617] <= ~layer2_out[4441] | layer2_out[4440];
     layer3_out[7618] <= layer2_out[9781] & ~layer2_out[9780];
     layer3_out[7619] <= layer2_out[5490];
     layer3_out[7620] <= ~layer2_out[10441] | layer2_out[10440];
     layer3_out[7621] <= layer2_out[11546] & ~layer2_out[11547];
     layer3_out[7622] <= layer2_out[5931];
     layer3_out[7623] <= layer2_out[11056];
     layer3_out[7624] <= ~layer2_out[2730];
     layer3_out[7625] <= layer2_out[11226];
     layer3_out[7626] <= layer2_out[8955] & ~layer2_out[8956];
     layer3_out[7627] <= layer2_out[276];
     layer3_out[7628] <= ~layer2_out[2690];
     layer3_out[7629] <= ~layer2_out[4936];
     layer3_out[7630] <= layer2_out[6667] | layer2_out[6668];
     layer3_out[7631] <= ~(layer2_out[492] | layer2_out[493]);
     layer3_out[7632] <= ~layer2_out[1478];
     layer3_out[7633] <= layer2_out[9455] & layer2_out[9456];
     layer3_out[7634] <= layer2_out[7263];
     layer3_out[7635] <= layer2_out[2587];
     layer3_out[7636] <= layer2_out[5482];
     layer3_out[7637] <= ~layer2_out[10472];
     layer3_out[7638] <= ~layer2_out[511];
     layer3_out[7639] <= ~layer2_out[10667];
     layer3_out[7640] <= layer2_out[11145];
     layer3_out[7641] <= ~layer2_out[7206];
     layer3_out[7642] <= layer2_out[1048];
     layer3_out[7643] <= layer2_out[6338];
     layer3_out[7644] <= ~(layer2_out[3513] ^ layer2_out[3514]);
     layer3_out[7645] <= layer2_out[3440];
     layer3_out[7646] <= layer2_out[10349] & ~layer2_out[10348];
     layer3_out[7647] <= ~layer2_out[10432];
     layer3_out[7648] <= layer2_out[10740] | layer2_out[10741];
     layer3_out[7649] <= ~layer2_out[11626];
     layer3_out[7650] <= ~(layer2_out[7991] | layer2_out[7992]);
     layer3_out[7651] <= ~layer2_out[10237];
     layer3_out[7652] <= ~(layer2_out[3416] | layer2_out[3417]);
     layer3_out[7653] <= layer2_out[6311];
     layer3_out[7654] <= ~layer2_out[1825];
     layer3_out[7655] <= layer2_out[739] & ~layer2_out[740];
     layer3_out[7656] <= ~layer2_out[134] | layer2_out[133];
     layer3_out[7657] <= layer2_out[6817] & layer2_out[6818];
     layer3_out[7658] <= layer2_out[8187];
     layer3_out[7659] <= layer2_out[10211] & ~layer2_out[10212];
     layer3_out[7660] <= ~layer2_out[10206];
     layer3_out[7661] <= ~layer2_out[6405] | layer2_out[6404];
     layer3_out[7662] <= layer2_out[2488] & ~layer2_out[2489];
     layer3_out[7663] <= ~layer2_out[4612];
     layer3_out[7664] <= ~(layer2_out[551] ^ layer2_out[552]);
     layer3_out[7665] <= ~(layer2_out[8285] | layer2_out[8286]);
     layer3_out[7666] <= layer2_out[6889] & ~layer2_out[6888];
     layer3_out[7667] <= layer2_out[942];
     layer3_out[7668] <= ~(layer2_out[8538] | layer2_out[8539]);
     layer3_out[7669] <= layer2_out[960];
     layer3_out[7670] <= ~layer2_out[6836];
     layer3_out[7671] <= layer2_out[2887] & ~layer2_out[2886];
     layer3_out[7672] <= ~layer2_out[5744];
     layer3_out[7673] <= ~(layer2_out[11547] | layer2_out[11548]);
     layer3_out[7674] <= layer2_out[8817];
     layer3_out[7675] <= layer2_out[583] & ~layer2_out[584];
     layer3_out[7676] <= ~layer2_out[9643];
     layer3_out[7677] <= layer2_out[960] & ~layer2_out[959];
     layer3_out[7678] <= ~layer2_out[9770] | layer2_out[9769];
     layer3_out[7679] <= layer2_out[3311];
     layer3_out[7680] <= ~layer2_out[7021] | layer2_out[7020];
     layer3_out[7681] <= ~(layer2_out[5318] | layer2_out[5319]);
     layer3_out[7682] <= ~layer2_out[9852];
     layer3_out[7683] <= layer2_out[954];
     layer3_out[7684] <= layer2_out[7360] & ~layer2_out[7361];
     layer3_out[7685] <= layer2_out[6220];
     layer3_out[7686] <= layer2_out[8820] & layer2_out[8821];
     layer3_out[7687] <= layer2_out[8018] | layer2_out[8019];
     layer3_out[7688] <= layer2_out[10644];
     layer3_out[7689] <= ~(layer2_out[6998] | layer2_out[6999]);
     layer3_out[7690] <= ~layer2_out[7821];
     layer3_out[7691] <= ~layer2_out[8474];
     layer3_out[7692] <= layer2_out[200];
     layer3_out[7693] <= layer2_out[8691];
     layer3_out[7694] <= layer2_out[4788] ^ layer2_out[4789];
     layer3_out[7695] <= layer2_out[3863];
     layer3_out[7696] <= layer2_out[5888];
     layer3_out[7697] <= layer2_out[9173];
     layer3_out[7698] <= ~layer2_out[8410] | layer2_out[8411];
     layer3_out[7699] <= ~layer2_out[2466];
     layer3_out[7700] <= layer2_out[605];
     layer3_out[7701] <= ~layer2_out[9696];
     layer3_out[7702] <= layer2_out[7595];
     layer3_out[7703] <= ~(layer2_out[6066] | layer2_out[6067]);
     layer3_out[7704] <= layer2_out[875] ^ layer2_out[876];
     layer3_out[7705] <= ~layer2_out[1163];
     layer3_out[7706] <= ~layer2_out[2824];
     layer3_out[7707] <= ~(layer2_out[4403] & layer2_out[4404]);
     layer3_out[7708] <= ~(layer2_out[1630] ^ layer2_out[1631]);
     layer3_out[7709] <= layer2_out[11302] & ~layer2_out[11303];
     layer3_out[7710] <= layer2_out[137] | layer2_out[138];
     layer3_out[7711] <= layer2_out[5800] ^ layer2_out[5801];
     layer3_out[7712] <= layer2_out[71] & ~layer2_out[70];
     layer3_out[7713] <= ~(layer2_out[5659] ^ layer2_out[5660]);
     layer3_out[7714] <= ~(layer2_out[11940] ^ layer2_out[11941]);
     layer3_out[7715] <= ~(layer2_out[10223] & layer2_out[10224]);
     layer3_out[7716] <= ~(layer2_out[5254] | layer2_out[5255]);
     layer3_out[7717] <= layer2_out[2154] ^ layer2_out[2155];
     layer3_out[7718] <= ~(layer2_out[3740] ^ layer2_out[3741]);
     layer3_out[7719] <= ~layer2_out[5348];
     layer3_out[7720] <= layer2_out[6777] & layer2_out[6778];
     layer3_out[7721] <= layer2_out[8304] & ~layer2_out[8303];
     layer3_out[7722] <= ~layer2_out[4027];
     layer3_out[7723] <= ~(layer2_out[4015] | layer2_out[4016]);
     layer3_out[7724] <= ~layer2_out[2260];
     layer3_out[7725] <= layer2_out[3088] & layer2_out[3089];
     layer3_out[7726] <= layer2_out[10265] & layer2_out[10266];
     layer3_out[7727] <= ~layer2_out[8843];
     layer3_out[7728] <= layer2_out[8106];
     layer3_out[7729] <= ~layer2_out[2350];
     layer3_out[7730] <= ~layer2_out[4977];
     layer3_out[7731] <= ~layer2_out[8998] | layer2_out[8999];
     layer3_out[7732] <= layer2_out[3928] & ~layer2_out[3927];
     layer3_out[7733] <= ~(layer2_out[3451] ^ layer2_out[3452]);
     layer3_out[7734] <= layer2_out[8535];
     layer3_out[7735] <= layer2_out[5094] & ~layer2_out[5095];
     layer3_out[7736] <= layer2_out[8448] & ~layer2_out[8447];
     layer3_out[7737] <= layer2_out[7536];
     layer3_out[7738] <= ~(layer2_out[2355] | layer2_out[2356]);
     layer3_out[7739] <= ~layer2_out[4594] | layer2_out[4595];
     layer3_out[7740] <= ~layer2_out[7759];
     layer3_out[7741] <= ~(layer2_out[3828] & layer2_out[3829]);
     layer3_out[7742] <= layer2_out[10948] & ~layer2_out[10947];
     layer3_out[7743] <= ~layer2_out[9798] | layer2_out[9799];
     layer3_out[7744] <= ~layer2_out[106];
     layer3_out[7745] <= layer2_out[11476] & layer2_out[11477];
     layer3_out[7746] <= ~layer2_out[470];
     layer3_out[7747] <= layer2_out[8014] & ~layer2_out[8013];
     layer3_out[7748] <= layer2_out[2815] & ~layer2_out[2814];
     layer3_out[7749] <= layer2_out[11617] ^ layer2_out[11618];
     layer3_out[7750] <= ~(layer2_out[4277] | layer2_out[4278]);
     layer3_out[7751] <= ~layer2_out[5206];
     layer3_out[7752] <= ~layer2_out[9259];
     layer3_out[7753] <= ~layer2_out[1939];
     layer3_out[7754] <= layer2_out[7642];
     layer3_out[7755] <= layer2_out[11595] & ~layer2_out[11596];
     layer3_out[7756] <= ~(layer2_out[9367] ^ layer2_out[9368]);
     layer3_out[7757] <= ~(layer2_out[418] | layer2_out[419]);
     layer3_out[7758] <= layer2_out[605] & ~layer2_out[604];
     layer3_out[7759] <= ~layer2_out[5851] | layer2_out[5852];
     layer3_out[7760] <= ~(layer2_out[9277] | layer2_out[9278]);
     layer3_out[7761] <= layer2_out[4320] & ~layer2_out[4319];
     layer3_out[7762] <= ~(layer2_out[4479] | layer2_out[4480]);
     layer3_out[7763] <= ~(layer2_out[9717] ^ layer2_out[9718]);
     layer3_out[7764] <= layer2_out[3714] & ~layer2_out[3713];
     layer3_out[7765] <= layer2_out[7528] & ~layer2_out[7527];
     layer3_out[7766] <= layer2_out[7060];
     layer3_out[7767] <= layer2_out[8341] & ~layer2_out[8342];
     layer3_out[7768] <= layer2_out[3654];
     layer3_out[7769] <= layer2_out[914] & ~layer2_out[913];
     layer3_out[7770] <= layer2_out[9805] & ~layer2_out[9806];
     layer3_out[7771] <= layer2_out[4616] & layer2_out[4617];
     layer3_out[7772] <= layer2_out[6941] & ~layer2_out[6940];
     layer3_out[7773] <= ~layer2_out[10291];
     layer3_out[7774] <= layer2_out[9291] & ~layer2_out[9292];
     layer3_out[7775] <= layer2_out[5561] ^ layer2_out[5562];
     layer3_out[7776] <= layer2_out[4317];
     layer3_out[7777] <= layer2_out[5560];
     layer3_out[7778] <= ~layer2_out[11917];
     layer3_out[7779] <= ~(layer2_out[2749] | layer2_out[2750]);
     layer3_out[7780] <= ~layer2_out[10934] | layer2_out[10935];
     layer3_out[7781] <= layer2_out[7239] & layer2_out[7240];
     layer3_out[7782] <= layer2_out[2644] & layer2_out[2645];
     layer3_out[7783] <= layer2_out[10494] & ~layer2_out[10495];
     layer3_out[7784] <= layer2_out[4558] & ~layer2_out[4557];
     layer3_out[7785] <= ~layer2_out[1815] | layer2_out[1814];
     layer3_out[7786] <= ~layer2_out[1085];
     layer3_out[7787] <= ~(layer2_out[9611] & layer2_out[9612]);
     layer3_out[7788] <= layer2_out[8580] ^ layer2_out[8581];
     layer3_out[7789] <= layer2_out[10404] ^ layer2_out[10405];
     layer3_out[7790] <= layer2_out[7246] ^ layer2_out[7247];
     layer3_out[7791] <= layer2_out[1123];
     layer3_out[7792] <= ~layer2_out[2796];
     layer3_out[7793] <= layer2_out[1587] ^ layer2_out[1588];
     layer3_out[7794] <= layer2_out[8367] & ~layer2_out[8368];
     layer3_out[7795] <= ~layer2_out[4352];
     layer3_out[7796] <= layer2_out[2494];
     layer3_out[7797] <= layer2_out[6226];
     layer3_out[7798] <= layer2_out[5581] & layer2_out[5582];
     layer3_out[7799] <= layer2_out[11901];
     layer3_out[7800] <= ~layer2_out[7484];
     layer3_out[7801] <= layer2_out[1967] & ~layer2_out[1966];
     layer3_out[7802] <= ~(layer2_out[1884] | layer2_out[1885]);
     layer3_out[7803] <= layer2_out[8942];
     layer3_out[7804] <= layer2_out[9661];
     layer3_out[7805] <= layer2_out[2374];
     layer3_out[7806] <= ~layer2_out[984];
     layer3_out[7807] <= layer2_out[5183] & layer2_out[5184];
     layer3_out[7808] <= ~layer2_out[5561] | layer2_out[5560];
     layer3_out[7809] <= ~(layer2_out[8267] | layer2_out[8268]);
     layer3_out[7810] <= layer2_out[10210] ^ layer2_out[10211];
     layer3_out[7811] <= layer2_out[747];
     layer3_out[7812] <= ~layer2_out[5629];
     layer3_out[7813] <= ~layer2_out[10652];
     layer3_out[7814] <= layer2_out[722] & ~layer2_out[721];
     layer3_out[7815] <= ~layer2_out[6065];
     layer3_out[7816] <= ~layer2_out[6742];
     layer3_out[7817] <= ~(layer2_out[4721] | layer2_out[4722]);
     layer3_out[7818] <= layer2_out[8011] & ~layer2_out[8012];
     layer3_out[7819] <= layer2_out[6965];
     layer3_out[7820] <= layer2_out[1754];
     layer3_out[7821] <= layer2_out[9813] & ~layer2_out[9814];
     layer3_out[7822] <= layer2_out[2685];
     layer3_out[7823] <= layer2_out[8885];
     layer3_out[7824] <= ~(layer2_out[11534] ^ layer2_out[11535]);
     layer3_out[7825] <= layer2_out[6024] & ~layer2_out[6025];
     layer3_out[7826] <= layer2_out[1157] & ~layer2_out[1158];
     layer3_out[7827] <= layer2_out[8489];
     layer3_out[7828] <= layer2_out[6684];
     layer3_out[7829] <= layer2_out[3206] & ~layer2_out[3207];
     layer3_out[7830] <= ~(layer2_out[3889] | layer2_out[3890]);
     layer3_out[7831] <= layer2_out[5616];
     layer3_out[7832] <= layer2_out[11606];
     layer3_out[7833] <= ~layer2_out[835];
     layer3_out[7834] <= layer2_out[1733];
     layer3_out[7835] <= ~(layer2_out[4204] ^ layer2_out[4205]);
     layer3_out[7836] <= ~(layer2_out[4598] | layer2_out[4599]);
     layer3_out[7837] <= layer2_out[4022] ^ layer2_out[4023];
     layer3_out[7838] <= ~layer2_out[4755];
     layer3_out[7839] <= ~layer2_out[2474];
     layer3_out[7840] <= layer2_out[7378];
     layer3_out[7841] <= ~layer2_out[8866];
     layer3_out[7842] <= ~layer2_out[7849];
     layer3_out[7843] <= layer2_out[2057];
     layer3_out[7844] <= layer2_out[2176] & ~layer2_out[2177];
     layer3_out[7845] <= layer2_out[10133];
     layer3_out[7846] <= layer2_out[8848] & ~layer2_out[8847];
     layer3_out[7847] <= ~(layer2_out[9104] | layer2_out[9105]);
     layer3_out[7848] <= ~(layer2_out[10767] | layer2_out[10768]);
     layer3_out[7849] <= ~layer2_out[5851];
     layer3_out[7850] <= layer2_out[11514] | layer2_out[11515];
     layer3_out[7851] <= layer2_out[5978] & ~layer2_out[5979];
     layer3_out[7852] <= layer2_out[4639] ^ layer2_out[4640];
     layer3_out[7853] <= layer2_out[2738];
     layer3_out[7854] <= layer2_out[7657] & layer2_out[7658];
     layer3_out[7855] <= layer2_out[2022] & ~layer2_out[2021];
     layer3_out[7856] <= layer2_out[8934] | layer2_out[8935];
     layer3_out[7857] <= layer2_out[11335] ^ layer2_out[11336];
     layer3_out[7858] <= ~layer2_out[6318];
     layer3_out[7859] <= layer2_out[7342] | layer2_out[7343];
     layer3_out[7860] <= ~(layer2_out[10490] & layer2_out[10491]);
     layer3_out[7861] <= layer2_out[10383] & ~layer2_out[10382];
     layer3_out[7862] <= ~layer2_out[2109];
     layer3_out[7863] <= layer2_out[10605];
     layer3_out[7864] <= layer2_out[2233];
     layer3_out[7865] <= ~(layer2_out[11768] | layer2_out[11769]);
     layer3_out[7866] <= layer2_out[5155];
     layer3_out[7867] <= ~layer2_out[7189];
     layer3_out[7868] <= ~(layer2_out[2981] & layer2_out[2982]);
     layer3_out[7869] <= ~layer2_out[3708];
     layer3_out[7870] <= layer2_out[10671];
     layer3_out[7871] <= layer2_out[6987];
     layer3_out[7872] <= layer2_out[9209];
     layer3_out[7873] <= ~layer2_out[11166];
     layer3_out[7874] <= ~layer2_out[4629] | layer2_out[4630];
     layer3_out[7875] <= ~layer2_out[7874];
     layer3_out[7876] <= ~(layer2_out[1091] ^ layer2_out[1092]);
     layer3_out[7877] <= ~layer2_out[9007];
     layer3_out[7878] <= layer2_out[810] ^ layer2_out[811];
     layer3_out[7879] <= ~(layer2_out[4370] & layer2_out[4371]);
     layer3_out[7880] <= layer2_out[11955];
     layer3_out[7881] <= layer2_out[5096] ^ layer2_out[5097];
     layer3_out[7882] <= layer2_out[7717] & ~layer2_out[7716];
     layer3_out[7883] <= layer2_out[7042] & layer2_out[7043];
     layer3_out[7884] <= ~layer2_out[4022];
     layer3_out[7885] <= ~layer2_out[3659];
     layer3_out[7886] <= ~layer2_out[6905];
     layer3_out[7887] <= layer2_out[407];
     layer3_out[7888] <= layer2_out[11831] & ~layer2_out[11830];
     layer3_out[7889] <= ~layer2_out[10659];
     layer3_out[7890] <= ~(layer2_out[4030] | layer2_out[4031]);
     layer3_out[7891] <= layer2_out[1912] & ~layer2_out[1913];
     layer3_out[7892] <= layer2_out[4511] & ~layer2_out[4510];
     layer3_out[7893] <= ~(layer2_out[7715] | layer2_out[7716]);
     layer3_out[7894] <= ~layer2_out[5662];
     layer3_out[7895] <= layer2_out[1785];
     layer3_out[7896] <= layer2_out[9033];
     layer3_out[7897] <= ~(layer2_out[1936] ^ layer2_out[1937]);
     layer3_out[7898] <= ~layer2_out[9192];
     layer3_out[7899] <= layer2_out[8042];
     layer3_out[7900] <= layer2_out[6421] & ~layer2_out[6420];
     layer3_out[7901] <= ~(layer2_out[1799] ^ layer2_out[1800]);
     layer3_out[7902] <= layer2_out[3395] & layer2_out[3396];
     layer3_out[7903] <= layer2_out[3838] & layer2_out[3839];
     layer3_out[7904] <= ~layer2_out[3501] | layer2_out[3502];
     layer3_out[7905] <= ~(layer2_out[5138] | layer2_out[5139]);
     layer3_out[7906] <= layer2_out[6771] & ~layer2_out[6772];
     layer3_out[7907] <= ~layer2_out[9556];
     layer3_out[7908] <= layer2_out[10012] & ~layer2_out[10011];
     layer3_out[7909] <= layer2_out[4217] ^ layer2_out[4218];
     layer3_out[7910] <= layer2_out[4112] & ~layer2_out[4111];
     layer3_out[7911] <= ~layer2_out[8588] | layer2_out[8589];
     layer3_out[7912] <= layer2_out[5430];
     layer3_out[7913] <= ~(layer2_out[3064] | layer2_out[3065]);
     layer3_out[7914] <= layer2_out[1344];
     layer3_out[7915] <= ~(layer2_out[4016] | layer2_out[4017]);
     layer3_out[7916] <= layer2_out[10806] & ~layer2_out[10807];
     layer3_out[7917] <= layer2_out[3580] & ~layer2_out[3579];
     layer3_out[7918] <= ~(layer2_out[7283] | layer2_out[7284]);
     layer3_out[7919] <= layer2_out[2397];
     layer3_out[7920] <= layer2_out[11546];
     layer3_out[7921] <= layer2_out[2691];
     layer3_out[7922] <= ~layer2_out[2946];
     layer3_out[7923] <= layer2_out[3082] & ~layer2_out[3083];
     layer3_out[7924] <= layer2_out[7476];
     layer3_out[7925] <= ~layer2_out[11432];
     layer3_out[7926] <= layer2_out[3009] & ~layer2_out[3008];
     layer3_out[7927] <= ~layer2_out[7892];
     layer3_out[7928] <= layer2_out[9550];
     layer3_out[7929] <= layer2_out[8132] ^ layer2_out[8133];
     layer3_out[7930] <= layer2_out[10246];
     layer3_out[7931] <= ~layer2_out[5733];
     layer3_out[7932] <= layer2_out[11131] & ~layer2_out[11130];
     layer3_out[7933] <= ~(layer2_out[9099] | layer2_out[9100]);
     layer3_out[7934] <= layer2_out[7650] ^ layer2_out[7651];
     layer3_out[7935] <= layer2_out[10536] ^ layer2_out[10537];
     layer3_out[7936] <= layer2_out[10553] & ~layer2_out[10552];
     layer3_out[7937] <= layer2_out[11832] & ~layer2_out[11833];
     layer3_out[7938] <= ~layer2_out[8460];
     layer3_out[7939] <= layer2_out[6719];
     layer3_out[7940] <= layer2_out[1376];
     layer3_out[7941] <= ~(layer2_out[2134] ^ layer2_out[2135]);
     layer3_out[7942] <= ~layer2_out[3199];
     layer3_out[7943] <= ~(layer2_out[10224] & layer2_out[10225]);
     layer3_out[7944] <= ~(layer2_out[3103] | layer2_out[3104]);
     layer3_out[7945] <= ~layer2_out[2442];
     layer3_out[7946] <= layer2_out[4786] & ~layer2_out[4787];
     layer3_out[7947] <= layer2_out[830] | layer2_out[831];
     layer3_out[7948] <= ~(layer2_out[1591] | layer2_out[1592]);
     layer3_out[7949] <= layer2_out[6819] | layer2_out[6820];
     layer3_out[7950] <= layer2_out[9424];
     layer3_out[7951] <= ~(layer2_out[10092] & layer2_out[10093]);
     layer3_out[7952] <= layer2_out[2744] & layer2_out[2745];
     layer3_out[7953] <= ~layer2_out[10459];
     layer3_out[7954] <= ~layer2_out[1088];
     layer3_out[7955] <= layer2_out[5400];
     layer3_out[7956] <= layer2_out[4963] & ~layer2_out[4962];
     layer3_out[7957] <= ~layer2_out[3034];
     layer3_out[7958] <= layer2_out[5436];
     layer3_out[7959] <= ~layer2_out[9279];
     layer3_out[7960] <= layer2_out[2433];
     layer3_out[7961] <= layer2_out[4476];
     layer3_out[7962] <= layer2_out[5151];
     layer3_out[7963] <= ~layer2_out[3756];
     layer3_out[7964] <= ~layer2_out[11187];
     layer3_out[7965] <= ~layer2_out[1023] | layer2_out[1022];
     layer3_out[7966] <= layer2_out[10062] & ~layer2_out[10063];
     layer3_out[7967] <= layer2_out[2158] & ~layer2_out[2159];
     layer3_out[7968] <= ~layer2_out[2515];
     layer3_out[7969] <= layer2_out[3428];
     layer3_out[7970] <= layer2_out[7790] & ~layer2_out[7791];
     layer3_out[7971] <= ~(layer2_out[5870] | layer2_out[5871]);
     layer3_out[7972] <= layer2_out[448];
     layer3_out[7973] <= layer2_out[4915];
     layer3_out[7974] <= layer2_out[7413] | layer2_out[7414];
     layer3_out[7975] <= ~(layer2_out[2941] ^ layer2_out[2942]);
     layer3_out[7976] <= layer2_out[5279] & layer2_out[5280];
     layer3_out[7977] <= ~layer2_out[781];
     layer3_out[7978] <= layer2_out[105] & ~layer2_out[106];
     layer3_out[7979] <= ~layer2_out[5642] | layer2_out[5643];
     layer3_out[7980] <= layer2_out[3156] & layer2_out[3157];
     layer3_out[7981] <= ~layer2_out[1532];
     layer3_out[7982] <= layer2_out[3419] & ~layer2_out[3418];
     layer3_out[7983] <= layer2_out[6129] & ~layer2_out[6130];
     layer3_out[7984] <= layer2_out[11202];
     layer3_out[7985] <= ~(layer2_out[9256] & layer2_out[9257]);
     layer3_out[7986] <= ~(layer2_out[5856] ^ layer2_out[5857]);
     layer3_out[7987] <= layer2_out[8558];
     layer3_out[7988] <= layer2_out[7150];
     layer3_out[7989] <= layer2_out[2162] & ~layer2_out[2161];
     layer3_out[7990] <= layer2_out[6494] ^ layer2_out[6495];
     layer3_out[7991] <= layer2_out[5902];
     layer3_out[7992] <= ~(layer2_out[414] ^ layer2_out[415]);
     layer3_out[7993] <= layer2_out[10703] & ~layer2_out[10704];
     layer3_out[7994] <= layer2_out[11278] & ~layer2_out[11279];
     layer3_out[7995] <= layer2_out[10905] & ~layer2_out[10904];
     layer3_out[7996] <= layer2_out[7295] & ~layer2_out[7294];
     layer3_out[7997] <= layer2_out[1400] | layer2_out[1401];
     layer3_out[7998] <= layer2_out[9619] ^ layer2_out[9620];
     layer3_out[7999] <= layer2_out[11681] ^ layer2_out[11682];
     layer3_out[8000] <= ~(layer2_out[6138] | layer2_out[6139]);
     layer3_out[8001] <= layer2_out[11182];
     layer3_out[8002] <= ~layer2_out[537];
     layer3_out[8003] <= layer2_out[4991];
     layer3_out[8004] <= ~layer2_out[4941];
     layer3_out[8005] <= layer2_out[2576] ^ layer2_out[2577];
     layer3_out[8006] <= ~layer2_out[6581];
     layer3_out[8007] <= layer2_out[6555];
     layer3_out[8008] <= layer2_out[11430];
     layer3_out[8009] <= layer2_out[4083] ^ layer2_out[4084];
     layer3_out[8010] <= ~layer2_out[4283];
     layer3_out[8011] <= ~layer2_out[4949];
     layer3_out[8012] <= layer2_out[11031] & ~layer2_out[11030];
     layer3_out[8013] <= layer2_out[992] & ~layer2_out[991];
     layer3_out[8014] <= ~layer2_out[3570];
     layer3_out[8015] <= layer2_out[3377] ^ layer2_out[3378];
     layer3_out[8016] <= layer2_out[5010] & ~layer2_out[5009];
     layer3_out[8017] <= ~(layer2_out[5145] & layer2_out[5146]);
     layer3_out[8018] <= layer2_out[4883];
     layer3_out[8019] <= layer2_out[204] & ~layer2_out[205];
     layer3_out[8020] <= layer2_out[9753] | layer2_out[9754];
     layer3_out[8021] <= layer2_out[2413] & layer2_out[2414];
     layer3_out[8022] <= layer2_out[3054] & ~layer2_out[3053];
     layer3_out[8023] <= ~(layer2_out[822] & layer2_out[823]);
     layer3_out[8024] <= ~layer2_out[4009];
     layer3_out[8025] <= layer2_out[1460];
     layer3_out[8026] <= layer2_out[7778] & layer2_out[7779];
     layer3_out[8027] <= layer2_out[1297] & ~layer2_out[1298];
     layer3_out[8028] <= ~layer2_out[859];
     layer3_out[8029] <= layer2_out[9121];
     layer3_out[8030] <= ~layer2_out[9524];
     layer3_out[8031] <= ~(layer2_out[189] ^ layer2_out[190]);
     layer3_out[8032] <= layer2_out[10529] & ~layer2_out[10528];
     layer3_out[8033] <= ~(layer2_out[5243] & layer2_out[5244]);
     layer3_out[8034] <= layer2_out[5515] ^ layer2_out[5516];
     layer3_out[8035] <= layer2_out[11792];
     layer3_out[8036] <= layer2_out[3407];
     layer3_out[8037] <= layer2_out[11095] & ~layer2_out[11096];
     layer3_out[8038] <= layer2_out[7972] & ~layer2_out[7973];
     layer3_out[8039] <= ~layer2_out[10258];
     layer3_out[8040] <= ~layer2_out[7575];
     layer3_out[8041] <= layer2_out[5846] ^ layer2_out[5847];
     layer3_out[8042] <= layer2_out[609];
     layer3_out[8043] <= layer2_out[7668] & ~layer2_out[7669];
     layer3_out[8044] <= ~(layer2_out[8081] | layer2_out[8082]);
     layer3_out[8045] <= ~(layer2_out[3614] | layer2_out[3615]);
     layer3_out[8046] <= layer2_out[7036];
     layer3_out[8047] <= layer2_out[6659];
     layer3_out[8048] <= layer2_out[10583] & ~layer2_out[10584];
     layer3_out[8049] <= ~(layer2_out[363] | layer2_out[364]);
     layer3_out[8050] <= layer2_out[2544] & ~layer2_out[2543];
     layer3_out[8051] <= ~(layer2_out[11663] | layer2_out[11664]);
     layer3_out[8052] <= ~layer2_out[4728];
     layer3_out[8053] <= ~(layer2_out[55] ^ layer2_out[56]);
     layer3_out[8054] <= ~layer2_out[3572];
     layer3_out[8055] <= layer2_out[367];
     layer3_out[8056] <= layer2_out[11638] & ~layer2_out[11639];
     layer3_out[8057] <= ~(layer2_out[2148] | layer2_out[2149]);
     layer3_out[8058] <= ~(layer2_out[6871] & layer2_out[6872]);
     layer3_out[8059] <= layer2_out[1811] & ~layer2_out[1810];
     layer3_out[8060] <= ~(layer2_out[5682] | layer2_out[5683]);
     layer3_out[8061] <= layer2_out[8440] & layer2_out[8441];
     layer3_out[8062] <= ~(layer2_out[4493] ^ layer2_out[4494]);
     layer3_out[8063] <= layer2_out[6849] & layer2_out[6850];
     layer3_out[8064] <= layer2_out[4867] & ~layer2_out[4866];
     layer3_out[8065] <= layer2_out[4158] & layer2_out[4159];
     layer3_out[8066] <= layer2_out[7615] ^ layer2_out[7616];
     layer3_out[8067] <= ~(layer2_out[10149] | layer2_out[10150]);
     layer3_out[8068] <= layer2_out[4720] & ~layer2_out[4721];
     layer3_out[8069] <= layer2_out[4138] ^ layer2_out[4139];
     layer3_out[8070] <= layer2_out[7235] & ~layer2_out[7236];
     layer3_out[8071] <= layer2_out[1249] & layer2_out[1250];
     layer3_out[8072] <= ~layer2_out[3118];
     layer3_out[8073] <= ~layer2_out[4045];
     layer3_out[8074] <= layer2_out[4578] | layer2_out[4579];
     layer3_out[8075] <= layer2_out[1916] & ~layer2_out[1915];
     layer3_out[8076] <= layer2_out[8650] & layer2_out[8651];
     layer3_out[8077] <= layer2_out[10689] & ~layer2_out[10688];
     layer3_out[8078] <= layer2_out[11977] ^ layer2_out[11978];
     layer3_out[8079] <= ~(layer2_out[5294] | layer2_out[5295]);
     layer3_out[8080] <= ~layer2_out[8410];
     layer3_out[8081] <= layer2_out[6040] ^ layer2_out[6041];
     layer3_out[8082] <= layer2_out[5488] & layer2_out[5489];
     layer3_out[8083] <= layer2_out[4231] ^ layer2_out[4232];
     layer3_out[8084] <= ~layer2_out[5264];
     layer3_out[8085] <= layer2_out[2203];
     layer3_out[8086] <= layer2_out[1452] & ~layer2_out[1453];
     layer3_out[8087] <= layer2_out[578];
     layer3_out[8088] <= ~layer2_out[1104];
     layer3_out[8089] <= layer2_out[2834] & ~layer2_out[2833];
     layer3_out[8090] <= layer2_out[1830] & ~layer2_out[1829];
     layer3_out[8091] <= ~(layer2_out[9223] | layer2_out[9224]);
     layer3_out[8092] <= layer2_out[6780];
     layer3_out[8093] <= layer2_out[1876] & ~layer2_out[1875];
     layer3_out[8094] <= ~(layer2_out[3854] | layer2_out[3855]);
     layer3_out[8095] <= ~layer2_out[4561];
     layer3_out[8096] <= ~layer2_out[1030];
     layer3_out[8097] <= ~layer2_out[6737];
     layer3_out[8098] <= layer2_out[1132];
     layer3_out[8099] <= ~layer2_out[7386];
     layer3_out[8100] <= layer2_out[1582] | layer2_out[1583];
     layer3_out[8101] <= ~layer2_out[9241];
     layer3_out[8102] <= layer2_out[1495];
     layer3_out[8103] <= layer2_out[2843];
     layer3_out[8104] <= layer2_out[6086] & ~layer2_out[6087];
     layer3_out[8105] <= layer2_out[4730] & layer2_out[4731];
     layer3_out[8106] <= layer2_out[1258];
     layer3_out[8107] <= layer2_out[6854] & layer2_out[6855];
     layer3_out[8108] <= layer2_out[3433] & ~layer2_out[3432];
     layer3_out[8109] <= layer2_out[710];
     layer3_out[8110] <= ~(layer2_out[7645] | layer2_out[7646]);
     layer3_out[8111] <= ~layer2_out[3415];
     layer3_out[8112] <= layer2_out[2992];
     layer3_out[8113] <= ~(layer2_out[140] | layer2_out[141]);
     layer3_out[8114] <= ~layer2_out[6868];
     layer3_out[8115] <= ~layer2_out[11420];
     layer3_out[8116] <= layer2_out[7940];
     layer3_out[8117] <= layer2_out[1807] & layer2_out[1808];
     layer3_out[8118] <= layer2_out[11849] & layer2_out[11850];
     layer3_out[8119] <= ~layer2_out[1885];
     layer3_out[8120] <= layer2_out[2668] | layer2_out[2669];
     layer3_out[8121] <= layer2_out[3522];
     layer3_out[8122] <= layer2_out[8422];
     layer3_out[8123] <= layer2_out[8665] & ~layer2_out[8666];
     layer3_out[8124] <= layer2_out[11356] ^ layer2_out[11357];
     layer3_out[8125] <= layer2_out[9754] & ~layer2_out[9755];
     layer3_out[8126] <= layer2_out[8076] & layer2_out[8077];
     layer3_out[8127] <= layer2_out[6170] & layer2_out[6171];
     layer3_out[8128] <= ~layer2_out[1628];
     layer3_out[8129] <= layer2_out[722] ^ layer2_out[723];
     layer3_out[8130] <= ~(layer2_out[10075] | layer2_out[10076]);
     layer3_out[8131] <= layer2_out[11591] & ~layer2_out[11592];
     layer3_out[8132] <= layer2_out[7736];
     layer3_out[8133] <= ~(layer2_out[9337] | layer2_out[9338]);
     layer3_out[8134] <= layer2_out[7205];
     layer3_out[8135] <= layer2_out[3486];
     layer3_out[8136] <= layer2_out[2234];
     layer3_out[8137] <= layer2_out[75] & layer2_out[76];
     layer3_out[8138] <= ~layer2_out[9277];
     layer3_out[8139] <= ~(layer2_out[6424] | layer2_out[6425]);
     layer3_out[8140] <= ~layer2_out[4422];
     layer3_out[8141] <= ~layer2_out[7028];
     layer3_out[8142] <= ~(layer2_out[4844] | layer2_out[4845]);
     layer3_out[8143] <= ~layer2_out[11890] | layer2_out[11891];
     layer3_out[8144] <= layer2_out[842] & ~layer2_out[843];
     layer3_out[8145] <= ~layer2_out[2813];
     layer3_out[8146] <= ~layer2_out[3562];
     layer3_out[8147] <= layer2_out[8878];
     layer3_out[8148] <= ~layer2_out[2583];
     layer3_out[8149] <= ~(layer2_out[8486] ^ layer2_out[8487]);
     layer3_out[8150] <= layer2_out[9468] & ~layer2_out[9469];
     layer3_out[8151] <= layer2_out[2430];
     layer3_out[8152] <= layer2_out[3242];
     layer3_out[8153] <= ~(layer2_out[23] & layer2_out[24]);
     layer3_out[8154] <= ~layer2_out[6128] | layer2_out[6129];
     layer3_out[8155] <= ~(layer2_out[3389] | layer2_out[3390]);
     layer3_out[8156] <= layer2_out[2859];
     layer3_out[8157] <= ~layer2_out[8256] | layer2_out[8257];
     layer3_out[8158] <= ~layer2_out[6297];
     layer3_out[8159] <= ~(layer2_out[2974] | layer2_out[2975]);
     layer3_out[8160] <= layer2_out[8059];
     layer3_out[8161] <= ~(layer2_out[1136] | layer2_out[1137]);
     layer3_out[8162] <= ~(layer2_out[11868] ^ layer2_out[11869]);
     layer3_out[8163] <= ~(layer2_out[10970] | layer2_out[10971]);
     layer3_out[8164] <= layer2_out[7455] & ~layer2_out[7454];
     layer3_out[8165] <= ~layer2_out[1240];
     layer3_out[8166] <= layer2_out[7547] | layer2_out[7548];
     layer3_out[8167] <= ~(layer2_out[6847] | layer2_out[6848]);
     layer3_out[8168] <= ~layer2_out[8128];
     layer3_out[8169] <= ~(layer2_out[13] ^ layer2_out[14]);
     layer3_out[8170] <= layer2_out[11422];
     layer3_out[8171] <= layer2_out[9073];
     layer3_out[8172] <= ~layer2_out[8491];
     layer3_out[8173] <= layer2_out[10881] & ~layer2_out[10882];
     layer3_out[8174] <= layer2_out[10081] & ~layer2_out[10080];
     layer3_out[8175] <= layer2_out[895];
     layer3_out[8176] <= layer2_out[2390] & layer2_out[2391];
     layer3_out[8177] <= layer2_out[9960];
     layer3_out[8178] <= layer2_out[11980] & ~layer2_out[11979];
     layer3_out[8179] <= layer2_out[9266] & layer2_out[9267];
     layer3_out[8180] <= ~layer2_out[9075];
     layer3_out[8181] <= ~layer2_out[6798];
     layer3_out[8182] <= layer2_out[10047];
     layer3_out[8183] <= layer2_out[5641] & ~layer2_out[5642];
     layer3_out[8184] <= ~(layer2_out[6906] | layer2_out[6907]);
     layer3_out[8185] <= layer2_out[10447] & layer2_out[10448];
     layer3_out[8186] <= layer2_out[9533] & layer2_out[9534];
     layer3_out[8187] <= layer2_out[2630];
     layer3_out[8188] <= ~(layer2_out[3073] | layer2_out[3074]);
     layer3_out[8189] <= layer2_out[2538] & ~layer2_out[2539];
     layer3_out[8190] <= ~layer2_out[6620];
     layer3_out[8191] <= ~(layer2_out[5172] ^ layer2_out[5173]);
     layer3_out[8192] <= layer2_out[11524] & ~layer2_out[11523];
     layer3_out[8193] <= layer2_out[7916] & layer2_out[7917];
     layer3_out[8194] <= ~(layer2_out[1923] | layer2_out[1924]);
     layer3_out[8195] <= ~layer2_out[181];
     layer3_out[8196] <= layer2_out[11714];
     layer3_out[8197] <= ~(layer2_out[3939] ^ layer2_out[3940]);
     layer3_out[8198] <= ~layer2_out[4463];
     layer3_out[8199] <= layer2_out[1474] & ~layer2_out[1475];
     layer3_out[8200] <= ~(layer2_out[5742] ^ layer2_out[5743]);
     layer3_out[8201] <= layer2_out[1154] & ~layer2_out[1153];
     layer3_out[8202] <= ~layer2_out[4514];
     layer3_out[8203] <= ~layer2_out[5066];
     layer3_out[8204] <= layer2_out[3782] & layer2_out[3783];
     layer3_out[8205] <= ~(layer2_out[7202] | layer2_out[7203]);
     layer3_out[8206] <= ~layer2_out[9043];
     layer3_out[8207] <= layer2_out[2277] & layer2_out[2278];
     layer3_out[8208] <= layer2_out[234] & ~layer2_out[233];
     layer3_out[8209] <= layer2_out[4554] & layer2_out[4555];
     layer3_out[8210] <= ~(layer2_out[9747] | layer2_out[9748]);
     layer3_out[8211] <= ~layer2_out[1145] | layer2_out[1144];
     layer3_out[8212] <= ~layer2_out[6533] | layer2_out[6532];
     layer3_out[8213] <= layer2_out[5980];
     layer3_out[8214] <= layer2_out[7975] ^ layer2_out[7976];
     layer3_out[8215] <= layer2_out[6887];
     layer3_out[8216] <= layer2_out[6489];
     layer3_out[8217] <= ~(layer2_out[7370] | layer2_out[7371]);
     layer3_out[8218] <= layer2_out[7733] & ~layer2_out[7734];
     layer3_out[8219] <= ~layer2_out[3695];
     layer3_out[8220] <= ~(layer2_out[2288] ^ layer2_out[2289]);
     layer3_out[8221] <= ~layer2_out[7735] | layer2_out[7736];
     layer3_out[8222] <= ~layer2_out[5826];
     layer3_out[8223] <= ~layer2_out[6496];
     layer3_out[8224] <= layer2_out[10860] & layer2_out[10861];
     layer3_out[8225] <= ~(layer2_out[9241] | layer2_out[9242]);
     layer3_out[8226] <= layer2_out[5384];
     layer3_out[8227] <= layer2_out[10518];
     layer3_out[8228] <= layer2_out[11957] & ~layer2_out[11956];
     layer3_out[8229] <= ~(layer2_out[9229] | layer2_out[9230]);
     layer3_out[8230] <= ~layer2_out[558] | layer2_out[557];
     layer3_out[8231] <= ~(layer2_out[3868] | layer2_out[3869]);
     layer3_out[8232] <= layer2_out[1035];
     layer3_out[8233] <= layer2_out[6059] & ~layer2_out[6060];
     layer3_out[8234] <= layer2_out[10297];
     layer3_out[8235] <= layer2_out[7713] & ~layer2_out[7714];
     layer3_out[8236] <= layer2_out[1912] & ~layer2_out[1911];
     layer3_out[8237] <= ~(layer2_out[11813] | layer2_out[11814]);
     layer3_out[8238] <= ~layer2_out[108] | layer2_out[109];
     layer3_out[8239] <= layer2_out[6201];
     layer3_out[8240] <= ~layer2_out[10992];
     layer3_out[8241] <= ~layer2_out[3947];
     layer3_out[8242] <= layer2_out[6547] & ~layer2_out[6548];
     layer3_out[8243] <= layer2_out[9079] & layer2_out[9080];
     layer3_out[8244] <= ~layer2_out[5945];
     layer3_out[8245] <= layer2_out[7922];
     layer3_out[8246] <= layer2_out[5928];
     layer3_out[8247] <= layer2_out[1619];
     layer3_out[8248] <= layer2_out[6276] & ~layer2_out[6275];
     layer3_out[8249] <= layer2_out[11425] & layer2_out[11426];
     layer3_out[8250] <= layer2_out[4492] & layer2_out[4493];
     layer3_out[8251] <= layer2_out[6098];
     layer3_out[8252] <= ~(layer2_out[9856] | layer2_out[9857]);
     layer3_out[8253] <= layer2_out[3928] & ~layer2_out[3929];
     layer3_out[8254] <= layer2_out[10903] & ~layer2_out[10904];
     layer3_out[8255] <= ~(layer2_out[9825] ^ layer2_out[9826]);
     layer3_out[8256] <= layer2_out[5755] & ~layer2_out[5754];
     layer3_out[8257] <= ~layer2_out[6884];
     layer3_out[8258] <= layer2_out[3850] & ~layer2_out[3851];
     layer3_out[8259] <= ~layer2_out[7628] | layer2_out[7629];
     layer3_out[8260] <= layer2_out[10655];
     layer3_out[8261] <= layer2_out[6919] & ~layer2_out[6920];
     layer3_out[8262] <= ~(layer2_out[6278] | layer2_out[6279]);
     layer3_out[8263] <= ~(layer2_out[1746] & layer2_out[1747]);
     layer3_out[8264] <= ~layer2_out[149];
     layer3_out[8265] <= ~(layer2_out[3482] & layer2_out[3483]);
     layer3_out[8266] <= layer2_out[9877] ^ layer2_out[9878];
     layer3_out[8267] <= layer2_out[10780] & ~layer2_out[10779];
     layer3_out[8268] <= layer2_out[530];
     layer3_out[8269] <= ~layer2_out[9647];
     layer3_out[8270] <= layer2_out[11945];
     layer3_out[8271] <= ~(layer2_out[7734] | layer2_out[7735]);
     layer3_out[8272] <= ~(layer2_out[4465] | layer2_out[4466]);
     layer3_out[8273] <= layer2_out[8563] & layer2_out[8564];
     layer3_out[8274] <= ~(layer2_out[9831] ^ layer2_out[9832]);
     layer3_out[8275] <= ~layer2_out[930];
     layer3_out[8276] <= ~layer2_out[10874];
     layer3_out[8277] <= layer2_out[2841];
     layer3_out[8278] <= ~layer2_out[3941] | layer2_out[3940];
     layer3_out[8279] <= ~(layer2_out[7950] | layer2_out[7951]);
     layer3_out[8280] <= layer2_out[8647] | layer2_out[8648];
     layer3_out[8281] <= layer2_out[8758] & ~layer2_out[8759];
     layer3_out[8282] <= ~(layer2_out[10088] ^ layer2_out[10089]);
     layer3_out[8283] <= ~layer2_out[3269] | layer2_out[3268];
     layer3_out[8284] <= ~(layer2_out[3647] | layer2_out[3648]);
     layer3_out[8285] <= layer2_out[6930];
     layer3_out[8286] <= layer2_out[10152] & ~layer2_out[10151];
     layer3_out[8287] <= layer2_out[7262];
     layer3_out[8288] <= layer2_out[3376];
     layer3_out[8289] <= layer2_out[6157] & layer2_out[6158];
     layer3_out[8290] <= layer2_out[49];
     layer3_out[8291] <= ~layer2_out[1635];
     layer3_out[8292] <= ~layer2_out[4771];
     layer3_out[8293] <= ~layer2_out[10840];
     layer3_out[8294] <= ~layer2_out[548];
     layer3_out[8295] <= layer2_out[404] & layer2_out[405];
     layer3_out[8296] <= layer2_out[3974];
     layer3_out[8297] <= layer2_out[3274];
     layer3_out[8298] <= layer2_out[5228];
     layer3_out[8299] <= ~(layer2_out[6168] ^ layer2_out[6169]);
     layer3_out[8300] <= layer2_out[4194] & ~layer2_out[4195];
     layer3_out[8301] <= ~layer2_out[4599];
     layer3_out[8302] <= layer2_out[320] & layer2_out[321];
     layer3_out[8303] <= ~layer2_out[7422];
     layer3_out[8304] <= ~layer2_out[11587];
     layer3_out[8305] <= layer2_out[1621] & ~layer2_out[1622];
     layer3_out[8306] <= layer2_out[1290] & layer2_out[1291];
     layer3_out[8307] <= ~layer2_out[8741];
     layer3_out[8308] <= layer2_out[4125] & layer2_out[4126];
     layer3_out[8309] <= ~layer2_out[10734];
     layer3_out[8310] <= ~layer2_out[4096];
     layer3_out[8311] <= ~(layer2_out[5803] & layer2_out[5804]);
     layer3_out[8312] <= ~(layer2_out[5854] | layer2_out[5855]);
     layer3_out[8313] <= ~layer2_out[8991];
     layer3_out[8314] <= layer2_out[4452];
     layer3_out[8315] <= layer2_out[9369];
     layer3_out[8316] <= layer2_out[891];
     layer3_out[8317] <= ~layer2_out[1315];
     layer3_out[8318] <= layer2_out[813];
     layer3_out[8319] <= layer2_out[8148];
     layer3_out[8320] <= layer2_out[10941] & ~layer2_out[10942];
     layer3_out[8321] <= ~layer2_out[2654];
     layer3_out[8322] <= ~(layer2_out[4917] | layer2_out[4918]);
     layer3_out[8323] <= layer2_out[8753] & ~layer2_out[8754];
     layer3_out[8324] <= layer2_out[4804];
     layer3_out[8325] <= layer2_out[673];
     layer3_out[8326] <= ~layer2_out[3611];
     layer3_out[8327] <= layer2_out[172] & ~layer2_out[171];
     layer3_out[8328] <= layer2_out[485] & layer2_out[486];
     layer3_out[8329] <= layer2_out[331] & layer2_out[332];
     layer3_out[8330] <= layer2_out[6821];
     layer3_out[8331] <= layer2_out[221];
     layer3_out[8332] <= ~layer2_out[10891];
     layer3_out[8333] <= layer2_out[1650];
     layer3_out[8334] <= layer2_out[1632];
     layer3_out[8335] <= ~layer2_out[10130];
     layer3_out[8336] <= layer2_out[7823] & ~layer2_out[7822];
     layer3_out[8337] <= layer2_out[11699];
     layer3_out[8338] <= layer2_out[7368] & ~layer2_out[7369];
     layer3_out[8339] <= ~layer2_out[7127];
     layer3_out[8340] <= ~(layer2_out[4276] | layer2_out[4277]);
     layer3_out[8341] <= layer2_out[2150] & ~layer2_out[2151];
     layer3_out[8342] <= layer2_out[6080];
     layer3_out[8343] <= ~(layer2_out[10180] | layer2_out[10181]);
     layer3_out[8344] <= layer2_out[4098] & ~layer2_out[4097];
     layer3_out[8345] <= layer2_out[10770] & ~layer2_out[10769];
     layer3_out[8346] <= ~layer2_out[10663];
     layer3_out[8347] <= layer2_out[2848];
     layer3_out[8348] <= ~(layer2_out[3622] ^ layer2_out[3623]);
     layer3_out[8349] <= layer2_out[37];
     layer3_out[8350] <= layer2_out[3688] & ~layer2_out[3689];
     layer3_out[8351] <= ~layer2_out[8629];
     layer3_out[8352] <= ~(layer2_out[2122] ^ layer2_out[2123]);
     layer3_out[8353] <= ~layer2_out[9894];
     layer3_out[8354] <= ~layer2_out[8953];
     layer3_out[8355] <= layer2_out[6725] & ~layer2_out[6726];
     layer3_out[8356] <= layer2_out[7227] & ~layer2_out[7226];
     layer3_out[8357] <= ~layer2_out[6292];
     layer3_out[8358] <= layer2_out[986];
     layer3_out[8359] <= ~layer2_out[2696];
     layer3_out[8360] <= layer2_out[1817] & layer2_out[1818];
     layer3_out[8361] <= layer2_out[3283] ^ layer2_out[3284];
     layer3_out[8362] <= layer2_out[1808] & layer2_out[1809];
     layer3_out[8363] <= ~layer2_out[4816];
     layer3_out[8364] <= layer2_out[5738] & layer2_out[5739];
     layer3_out[8365] <= ~(layer2_out[4908] ^ layer2_out[4909]);
     layer3_out[8366] <= layer2_out[939] & layer2_out[940];
     layer3_out[8367] <= ~layer2_out[1999];
     layer3_out[8368] <= layer2_out[3866] & ~layer2_out[3867];
     layer3_out[8369] <= layer2_out[3296] & ~layer2_out[3295];
     layer3_out[8370] <= ~(layer2_out[3093] | layer2_out[3094]);
     layer3_out[8371] <= ~(layer2_out[2894] | layer2_out[2895]);
     layer3_out[8372] <= ~(layer2_out[4919] ^ layer2_out[4920]);
     layer3_out[8373] <= layer2_out[11853] & ~layer2_out[11854];
     layer3_out[8374] <= layer2_out[4804];
     layer3_out[8375] <= layer2_out[3264] ^ layer2_out[3265];
     layer3_out[8376] <= layer2_out[8154] & ~layer2_out[8155];
     layer3_out[8377] <= ~layer2_out[6134];
     layer3_out[8378] <= layer2_out[3618];
     layer3_out[8379] <= layer2_out[1063] ^ layer2_out[1064];
     layer3_out[8380] <= ~(layer2_out[1037] | layer2_out[1038]);
     layer3_out[8381] <= layer2_out[11093] ^ layer2_out[11094];
     layer3_out[8382] <= layer2_out[11445] | layer2_out[11446];
     layer3_out[8383] <= layer2_out[4032] | layer2_out[4033];
     layer3_out[8384] <= layer2_out[312];
     layer3_out[8385] <= ~(layer2_out[7450] ^ layer2_out[7451]);
     layer3_out[8386] <= ~layer2_out[5088];
     layer3_out[8387] <= layer2_out[5454] & ~layer2_out[5453];
     layer3_out[8388] <= layer2_out[5323];
     layer3_out[8389] <= layer2_out[7234];
     layer3_out[8390] <= ~layer2_out[9045] | layer2_out[9046];
     layer3_out[8391] <= ~layer2_out[1313];
     layer3_out[8392] <= layer2_out[2319] & layer2_out[2320];
     layer3_out[8393] <= layer2_out[1974] & layer2_out[1975];
     layer3_out[8394] <= layer2_out[9458] & ~layer2_out[9459];
     layer3_out[8395] <= ~(layer2_out[9756] & layer2_out[9757]);
     layer3_out[8396] <= ~layer2_out[7167];
     layer3_out[8397] <= layer2_out[1348] & layer2_out[1349];
     layer3_out[8398] <= layer2_out[973];
     layer3_out[8399] <= ~(layer2_out[7889] ^ layer2_out[7890]);
     layer3_out[8400] <= layer2_out[11780];
     layer3_out[8401] <= layer2_out[3933];
     layer3_out[8402] <= layer2_out[8763];
     layer3_out[8403] <= layer2_out[11500];
     layer3_out[8404] <= ~layer2_out[9112];
     layer3_out[8405] <= ~layer2_out[10554];
     layer3_out[8406] <= ~layer2_out[4122];
     layer3_out[8407] <= ~layer2_out[9610];
     layer3_out[8408] <= ~(layer2_out[6727] & layer2_out[6728]);
     layer3_out[8409] <= ~layer2_out[1499];
     layer3_out[8410] <= ~layer2_out[11832];
     layer3_out[8411] <= layer2_out[4247] | layer2_out[4248];
     layer3_out[8412] <= ~layer2_out[10066];
     layer3_out[8413] <= layer2_out[97];
     layer3_out[8414] <= layer2_out[11740] ^ layer2_out[11741];
     layer3_out[8415] <= layer2_out[7833] & layer2_out[7834];
     layer3_out[8416] <= layer2_out[2205] ^ layer2_out[2206];
     layer3_out[8417] <= layer2_out[1196] ^ layer2_out[1197];
     layer3_out[8418] <= ~layer2_out[10285] | layer2_out[10284];
     layer3_out[8419] <= ~layer2_out[4957];
     layer3_out[8420] <= layer2_out[3013] | layer2_out[3014];
     layer3_out[8421] <= ~(layer2_out[10335] | layer2_out[10336]);
     layer3_out[8422] <= ~layer2_out[6647];
     layer3_out[8423] <= layer2_out[4606] & ~layer2_out[4605];
     layer3_out[8424] <= ~layer2_out[826];
     layer3_out[8425] <= ~layer2_out[4499] | layer2_out[4498];
     layer3_out[8426] <= ~(layer2_out[7959] ^ layer2_out[7960]);
     layer3_out[8427] <= layer2_out[2375];
     layer3_out[8428] <= ~layer2_out[4297];
     layer3_out[8429] <= layer2_out[6051] ^ layer2_out[6052];
     layer3_out[8430] <= ~layer2_out[3279];
     layer3_out[8431] <= ~layer2_out[5396] | layer2_out[5395];
     layer3_out[8432] <= layer2_out[4731] ^ layer2_out[4732];
     layer3_out[8433] <= ~(layer2_out[10176] ^ layer2_out[10177]);
     layer3_out[8434] <= ~layer2_out[6459] | layer2_out[6460];
     layer3_out[8435] <= layer2_out[7649] & ~layer2_out[7650];
     layer3_out[8436] <= ~(layer2_out[232] ^ layer2_out[233]);
     layer3_out[8437] <= ~layer2_out[10914];
     layer3_out[8438] <= layer2_out[103] | layer2_out[104];
     layer3_out[8439] <= ~(layer2_out[8168] ^ layer2_out[8169]);
     layer3_out[8440] <= layer2_out[11090] & layer2_out[11091];
     layer3_out[8441] <= ~layer2_out[4949] | layer2_out[4948];
     layer3_out[8442] <= layer2_out[4897] & layer2_out[4898];
     layer3_out[8443] <= ~(layer2_out[5573] ^ layer2_out[5574]);
     layer3_out[8444] <= layer2_out[4872] ^ layer2_out[4873];
     layer3_out[8445] <= layer2_out[5381];
     layer3_out[8446] <= ~layer2_out[5680] | layer2_out[5681];
     layer3_out[8447] <= layer2_out[4467];
     layer3_out[8448] <= layer2_out[3799] & ~layer2_out[3798];
     layer3_out[8449] <= ~(layer2_out[6793] | layer2_out[6794]);
     layer3_out[8450] <= layer2_out[9973];
     layer3_out[8451] <= ~layer2_out[6437];
     layer3_out[8452] <= layer2_out[8596] & layer2_out[8597];
     layer3_out[8453] <= layer2_out[508];
     layer3_out[8454] <= layer2_out[758];
     layer3_out[8455] <= ~(layer2_out[8457] | layer2_out[8458]);
     layer3_out[8456] <= ~layer2_out[2504];
     layer3_out[8457] <= layer2_out[10594];
     layer3_out[8458] <= ~layer2_out[7951];
     layer3_out[8459] <= layer2_out[1064] & layer2_out[1065];
     layer3_out[8460] <= ~layer2_out[1308];
     layer3_out[8461] <= layer2_out[524];
     layer3_out[8462] <= ~layer2_out[9435];
     layer3_out[8463] <= ~layer2_out[11301];
     layer3_out[8464] <= ~layer2_out[8832] | layer2_out[8833];
     layer3_out[8465] <= layer2_out[4675] | layer2_out[4676];
     layer3_out[8466] <= layer2_out[1618];
     layer3_out[8467] <= layer2_out[8707] & ~layer2_out[8708];
     layer3_out[8468] <= ~(layer2_out[1374] | layer2_out[1375]);
     layer3_out[8469] <= ~layer2_out[6528];
     layer3_out[8470] <= layer2_out[7692];
     layer3_out[8471] <= layer2_out[6837] ^ layer2_out[6838];
     layer3_out[8472] <= ~(layer2_out[1501] ^ layer2_out[1502]);
     layer3_out[8473] <= ~(layer2_out[2964] ^ layer2_out[2965]);
     layer3_out[8474] <= ~layer2_out[11976] | layer2_out[11977];
     layer3_out[8475] <= ~(layer2_out[5888] ^ layer2_out[5889]);
     layer3_out[8476] <= layer2_out[10827] ^ layer2_out[10828];
     layer3_out[8477] <= layer2_out[6515];
     layer3_out[8478] <= ~layer2_out[5203] | layer2_out[5202];
     layer3_out[8479] <= layer2_out[1876] ^ layer2_out[1877];
     layer3_out[8480] <= ~layer2_out[11123];
     layer3_out[8481] <= layer2_out[11230];
     layer3_out[8482] <= layer2_out[3382] & layer2_out[3383];
     layer3_out[8483] <= layer2_out[9243] ^ layer2_out[9244];
     layer3_out[8484] <= ~(layer2_out[11065] ^ layer2_out[11066]);
     layer3_out[8485] <= layer2_out[1366] ^ layer2_out[1367];
     layer3_out[8486] <= ~layer2_out[8726];
     layer3_out[8487] <= layer2_out[10074] & ~layer2_out[10073];
     layer3_out[8488] <= layer2_out[2147];
     layer3_out[8489] <= layer2_out[223] ^ layer2_out[224];
     layer3_out[8490] <= ~(layer2_out[9] & layer2_out[10]);
     layer3_out[8491] <= layer2_out[9862];
     layer3_out[8492] <= ~layer2_out[4306];
     layer3_out[8493] <= layer2_out[9176];
     layer3_out[8494] <= layer2_out[776];
     layer3_out[8495] <= layer2_out[3895];
     layer3_out[8496] <= ~(layer2_out[11567] | layer2_out[11568]);
     layer3_out[8497] <= ~layer2_out[7042] | layer2_out[7041];
     layer3_out[8498] <= layer2_out[11223] | layer2_out[11224];
     layer3_out[8499] <= layer2_out[9097] & ~layer2_out[9096];
     layer3_out[8500] <= layer2_out[9616] ^ layer2_out[9617];
     layer3_out[8501] <= ~(layer2_out[9116] ^ layer2_out[9117]);
     layer3_out[8502] <= ~layer2_out[10518] | layer2_out[10517];
     layer3_out[8503] <= layer2_out[2270] & ~layer2_out[2269];
     layer3_out[8504] <= layer2_out[7575] ^ layer2_out[7576];
     layer3_out[8505] <= layer2_out[9595];
     layer3_out[8506] <= layer2_out[9840] | layer2_out[9841];
     layer3_out[8507] <= layer2_out[11582];
     layer3_out[8508] <= ~layer2_out[3619] | layer2_out[3620];
     layer3_out[8509] <= ~layer2_out[9151] | layer2_out[9150];
     layer3_out[8510] <= ~(layer2_out[238] | layer2_out[239]);
     layer3_out[8511] <= ~(layer2_out[4060] ^ layer2_out[4061]);
     layer3_out[8512] <= layer2_out[8001];
     layer3_out[8513] <= layer2_out[8195] ^ layer2_out[8196];
     layer3_out[8514] <= layer2_out[1445];
     layer3_out[8515] <= layer2_out[9915] & ~layer2_out[9914];
     layer3_out[8516] <= layer2_out[4356];
     layer3_out[8517] <= layer2_out[6327];
     layer3_out[8518] <= ~layer2_out[771] | layer2_out[772];
     layer3_out[8519] <= ~layer2_out[11931];
     layer3_out[8520] <= layer2_out[65];
     layer3_out[8521] <= layer2_out[1027] & ~layer2_out[1026];
     layer3_out[8522] <= layer2_out[5124] & ~layer2_out[5123];
     layer3_out[8523] <= layer2_out[1302] & layer2_out[1303];
     layer3_out[8524] <= layer2_out[2629];
     layer3_out[8525] <= ~layer2_out[6463];
     layer3_out[8526] <= ~layer2_out[9127] | layer2_out[9128];
     layer3_out[8527] <= ~(layer2_out[514] ^ layer2_out[515]);
     layer3_out[8528] <= layer2_out[8767];
     layer3_out[8529] <= ~(layer2_out[11271] ^ layer2_out[11272]);
     layer3_out[8530] <= layer2_out[8426];
     layer3_out[8531] <= ~(layer2_out[1371] ^ layer2_out[1372]);
     layer3_out[8532] <= ~layer2_out[3993];
     layer3_out[8533] <= layer2_out[818];
     layer3_out[8534] <= ~(layer2_out[1214] ^ layer2_out[1215]);
     layer3_out[8535] <= ~(layer2_out[7903] & layer2_out[7904]);
     layer3_out[8536] <= ~layer2_out[2338] | layer2_out[2339];
     layer3_out[8537] <= ~layer2_out[2602];
     layer3_out[8538] <= layer2_out[10480] & ~layer2_out[10481];
     layer3_out[8539] <= layer2_out[10717];
     layer3_out[8540] <= ~layer2_out[8312];
     layer3_out[8541] <= ~(layer2_out[4921] & layer2_out[4922]);
     layer3_out[8542] <= layer2_out[8014] ^ layer2_out[8015];
     layer3_out[8543] <= layer2_out[7501] & layer2_out[7502];
     layer3_out[8544] <= layer2_out[8801] & layer2_out[8802];
     layer3_out[8545] <= ~(layer2_out[11671] & layer2_out[11672]);
     layer3_out[8546] <= ~layer2_out[2422] | layer2_out[2423];
     layer3_out[8547] <= ~(layer2_out[4387] ^ layer2_out[4388]);
     layer3_out[8548] <= ~(layer2_out[7119] | layer2_out[7120]);
     layer3_out[8549] <= ~(layer2_out[1487] | layer2_out[1488]);
     layer3_out[8550] <= layer2_out[3028];
     layer3_out[8551] <= ~layer2_out[3447] | layer2_out[3448];
     layer3_out[8552] <= layer2_out[9491] & ~layer2_out[9492];
     layer3_out[8553] <= ~(layer2_out[279] & layer2_out[280]);
     layer3_out[8554] <= ~layer2_out[6457];
     layer3_out[8555] <= ~layer2_out[6055];
     layer3_out[8556] <= layer2_out[8680] & ~layer2_out[8679];
     layer3_out[8557] <= layer2_out[701] & ~layer2_out[702];
     layer3_out[8558] <= layer2_out[97] & ~layer2_out[96];
     layer3_out[8559] <= layer2_out[7895] & layer2_out[7896];
     layer3_out[8560] <= layer2_out[11080];
     layer3_out[8561] <= ~layer2_out[278];
     layer3_out[8562] <= ~layer2_out[2190];
     layer3_out[8563] <= layer2_out[10721] & ~layer2_out[10722];
     layer3_out[8564] <= layer2_out[4253] & layer2_out[4254];
     layer3_out[8565] <= ~layer2_out[10] | layer2_out[11];
     layer3_out[8566] <= layer2_out[11354] & ~layer2_out[11355];
     layer3_out[8567] <= ~layer2_out[3946];
     layer3_out[8568] <= layer2_out[9766];
     layer3_out[8569] <= layer2_out[2581];
     layer3_out[8570] <= layer2_out[1128] & layer2_out[1129];
     layer3_out[8571] <= ~(layer2_out[6121] | layer2_out[6122]);
     layer3_out[8572] <= layer2_out[6433] ^ layer2_out[6434];
     layer3_out[8573] <= layer2_out[8374] | layer2_out[8375];
     layer3_out[8574] <= ~(layer2_out[10389] & layer2_out[10390]);
     layer3_out[8575] <= ~(layer2_out[246] ^ layer2_out[247]);
     layer3_out[8576] <= ~layer2_out[704];
     layer3_out[8577] <= ~(layer2_out[3730] & layer2_out[3731]);
     layer3_out[8578] <= ~(layer2_out[3321] | layer2_out[3322]);
     layer3_out[8579] <= layer2_out[719] | layer2_out[720];
     layer3_out[8580] <= ~layer2_out[4249] | layer2_out[4248];
     layer3_out[8581] <= layer2_out[1300] ^ layer2_out[1301];
     layer3_out[8582] <= layer2_out[10721];
     layer3_out[8583] <= layer2_out[647];
     layer3_out[8584] <= layer2_out[4847] ^ layer2_out[4848];
     layer3_out[8585] <= ~(layer2_out[617] ^ layer2_out[618]);
     layer3_out[8586] <= layer2_out[636];
     layer3_out[8587] <= ~(layer2_out[2096] ^ layer2_out[2097]);
     layer3_out[8588] <= ~layer2_out[2807];
     layer3_out[8589] <= layer2_out[10386] | layer2_out[10387];
     layer3_out[8590] <= ~layer2_out[3139];
     layer3_out[8591] <= layer2_out[3784];
     layer3_out[8592] <= ~(layer2_out[5239] & layer2_out[5240]);
     layer3_out[8593] <= ~layer2_out[5080];
     layer3_out[8594] <= layer2_out[292];
     layer3_out[8595] <= ~layer2_out[3065];
     layer3_out[8596] <= layer2_out[10466] ^ layer2_out[10467];
     layer3_out[8597] <= layer2_out[4518];
     layer3_out[8598] <= ~layer2_out[9513] | layer2_out[9514];
     layer3_out[8599] <= layer2_out[8382] & layer2_out[8383];
     layer3_out[8600] <= ~(layer2_out[11215] | layer2_out[11216]);
     layer3_out[8601] <= layer2_out[2658] ^ layer2_out[2659];
     layer3_out[8602] <= layer2_out[2499] & ~layer2_out[2498];
     layer3_out[8603] <= ~layer2_out[4980];
     layer3_out[8604] <= layer2_out[8127] & ~layer2_out[8126];
     layer3_out[8605] <= layer2_out[1968] ^ layer2_out[1969];
     layer3_out[8606] <= ~layer2_out[8436];
     layer3_out[8607] <= layer2_out[6925] | layer2_out[6926];
     layer3_out[8608] <= ~layer2_out[5411];
     layer3_out[8609] <= layer2_out[9345] & ~layer2_out[9344];
     layer3_out[8610] <= layer2_out[11208];
     layer3_out[8611] <= layer2_out[4521] & ~layer2_out[4520];
     layer3_out[8612] <= layer2_out[4136];
     layer3_out[8613] <= layer2_out[3010] ^ layer2_out[3011];
     layer3_out[8614] <= ~layer2_out[6491] | layer2_out[6490];
     layer3_out[8615] <= layer2_out[900];
     layer3_out[8616] <= layer2_out[7093] & ~layer2_out[7094];
     layer3_out[8617] <= ~(layer2_out[11310] | layer2_out[11311]);
     layer3_out[8618] <= layer2_out[11721] | layer2_out[11722];
     layer3_out[8619] <= layer2_out[9531] | layer2_out[9532];
     layer3_out[8620] <= layer2_out[231];
     layer3_out[8621] <= layer2_out[143] & layer2_out[144];
     layer3_out[8622] <= ~layer2_out[10181] | layer2_out[10182];
     layer3_out[8623] <= layer2_out[11839];
     layer3_out[8624] <= layer2_out[8973];
     layer3_out[8625] <= ~(layer2_out[10462] | layer2_out[10463]);
     layer3_out[8626] <= layer2_out[10376] ^ layer2_out[10377];
     layer3_out[8627] <= layer2_out[7516] ^ layer2_out[7517];
     layer3_out[8628] <= ~(layer2_out[10189] & layer2_out[10190]);
     layer3_out[8629] <= layer2_out[5713];
     layer3_out[8630] <= layer2_out[7221];
     layer3_out[8631] <= ~layer2_out[8401];
     layer3_out[8632] <= layer2_out[8244];
     layer3_out[8633] <= ~(layer2_out[3606] | layer2_out[3607]);
     layer3_out[8634] <= ~layer2_out[11823];
     layer3_out[8635] <= layer2_out[5253];
     layer3_out[8636] <= layer2_out[2079];
     layer3_out[8637] <= ~layer2_out[9253] | layer2_out[9254];
     layer3_out[8638] <= ~(layer2_out[226] & layer2_out[227]);
     layer3_out[8639] <= ~(layer2_out[437] | layer2_out[438]);
     layer3_out[8640] <= layer2_out[6526];
     layer3_out[8641] <= layer2_out[1681];
     layer3_out[8642] <= layer2_out[8564] | layer2_out[8565];
     layer3_out[8643] <= layer2_out[6844];
     layer3_out[8644] <= layer2_out[2447] & layer2_out[2448];
     layer3_out[8645] <= ~layer2_out[2262] | layer2_out[2263];
     layer3_out[8646] <= layer2_out[5195];
     layer3_out[8647] <= layer2_out[5369] & ~layer2_out[5370];
     layer3_out[8648] <= layer2_out[6321] & layer2_out[6322];
     layer3_out[8649] <= layer2_out[10916] & ~layer2_out[10917];
     layer3_out[8650] <= layer2_out[5464] ^ layer2_out[5465];
     layer3_out[8651] <= ~layer2_out[9108];
     layer3_out[8652] <= layer2_out[11508] & ~layer2_out[11507];
     layer3_out[8653] <= ~(layer2_out[2097] | layer2_out[2098]);
     layer3_out[8654] <= layer2_out[9656] ^ layer2_out[9657];
     layer3_out[8655] <= ~layer2_out[10826] | layer2_out[10825];
     layer3_out[8656] <= layer2_out[8601] | layer2_out[8602];
     layer3_out[8657] <= layer2_out[4007] | layer2_out[4008];
     layer3_out[8658] <= layer2_out[5217] ^ layer2_out[5218];
     layer3_out[8659] <= ~layer2_out[11156];
     layer3_out[8660] <= layer2_out[4933] & layer2_out[4934];
     layer3_out[8661] <= ~layer2_out[6914] | layer2_out[6915];
     layer3_out[8662] <= layer2_out[10588];
     layer3_out[8663] <= ~layer2_out[1234] | layer2_out[1235];
     layer3_out[8664] <= ~layer2_out[5053] | layer2_out[5052];
     layer3_out[8665] <= layer2_out[2409];
     layer3_out[8666] <= ~layer2_out[7272] | layer2_out[7271];
     layer3_out[8667] <= layer2_out[9474];
     layer3_out[8668] <= layer2_out[6394] ^ layer2_out[6395];
     layer3_out[8669] <= ~(layer2_out[10394] & layer2_out[10395]);
     layer3_out[8670] <= ~layer2_out[10933];
     layer3_out[8671] <= layer2_out[2639] ^ layer2_out[2640];
     layer3_out[8672] <= layer2_out[8250];
     layer3_out[8673] <= ~layer2_out[6037] | layer2_out[6036];
     layer3_out[8674] <= ~layer2_out[11352] | layer2_out[11351];
     layer3_out[8675] <= layer2_out[11016] & layer2_out[11017];
     layer3_out[8676] <= ~layer2_out[8938] | layer2_out[8939];
     layer3_out[8677] <= layer2_out[2985];
     layer3_out[8678] <= ~layer2_out[1170];
     layer3_out[8679] <= ~layer2_out[9711];
     layer3_out[8680] <= ~layer2_out[9068];
     layer3_out[8681] <= ~layer2_out[1046];
     layer3_out[8682] <= ~layer2_out[3048];
     layer3_out[8683] <= layer2_out[5191] & ~layer2_out[5192];
     layer3_out[8684] <= ~layer2_out[10935];
     layer3_out[8685] <= ~layer2_out[6823];
     layer3_out[8686] <= ~layer2_out[1718];
     layer3_out[8687] <= ~(layer2_out[11314] & layer2_out[11315]);
     layer3_out[8688] <= ~(layer2_out[7163] ^ layer2_out[7164]);
     layer3_out[8689] <= layer2_out[462];
     layer3_out[8690] <= layer2_out[3401] & layer2_out[3402];
     layer3_out[8691] <= ~layer2_out[1623] | layer2_out[1624];
     layer3_out[8692] <= layer2_out[2561] ^ layer2_out[2562];
     layer3_out[8693] <= ~layer2_out[855];
     layer3_out[8694] <= layer2_out[10949] & ~layer2_out[10948];
     layer3_out[8695] <= layer2_out[7514] ^ layer2_out[7515];
     layer3_out[8696] <= ~layer2_out[9075];
     layer3_out[8697] <= layer2_out[3260] ^ layer2_out[3261];
     layer3_out[8698] <= layer2_out[6120] & ~layer2_out[6121];
     layer3_out[8699] <= layer2_out[3267];
     layer3_out[8700] <= layer2_out[10469];
     layer3_out[8701] <= ~layer2_out[3824];
     layer3_out[8702] <= layer2_out[7942];
     layer3_out[8703] <= layer2_out[2475];
     layer3_out[8704] <= ~(layer2_out[11114] | layer2_out[11115]);
     layer3_out[8705] <= ~layer2_out[833];
     layer3_out[8706] <= layer2_out[5774] & ~layer2_out[5775];
     layer3_out[8707] <= layer2_out[8818] ^ layer2_out[8819];
     layer3_out[8708] <= ~layer2_out[1646];
     layer3_out[8709] <= ~(layer2_out[5307] & layer2_out[5308]);
     layer3_out[8710] <= layer2_out[2544] & ~layer2_out[2545];
     layer3_out[8711] <= layer2_out[1898];
     layer3_out[8712] <= ~(layer2_out[7946] | layer2_out[7947]);
     layer3_out[8713] <= layer2_out[9882] & ~layer2_out[9881];
     layer3_out[8714] <= ~layer2_out[1322];
     layer3_out[8715] <= layer2_out[11143];
     layer3_out[8716] <= layer2_out[2299];
     layer3_out[8717] <= ~(layer2_out[5346] & layer2_out[5347]);
     layer3_out[8718] <= layer2_out[8636];
     layer3_out[8719] <= layer2_out[510];
     layer3_out[8720] <= layer2_out[11641];
     layer3_out[8721] <= ~layer2_out[306];
     layer3_out[8722] <= ~(layer2_out[1126] & layer2_out[1127]);
     layer3_out[8723] <= layer2_out[4193];
     layer3_out[8724] <= layer2_out[6492] & layer2_out[6493];
     layer3_out[8725] <= layer2_out[1533] ^ layer2_out[1534];
     layer3_out[8726] <= layer2_out[1703];
     layer3_out[8727] <= layer2_out[5861] & ~layer2_out[5860];
     layer3_out[8728] <= layer2_out[1486] & ~layer2_out[1485];
     layer3_out[8729] <= layer2_out[11743] & ~layer2_out[11744];
     layer3_out[8730] <= ~(layer2_out[4494] ^ layer2_out[4495]);
     layer3_out[8731] <= layer2_out[9974];
     layer3_out[8732] <= layer2_out[10289] & layer2_out[10290];
     layer3_out[8733] <= ~layer2_out[533] | layer2_out[532];
     layer3_out[8734] <= ~(layer2_out[4272] | layer2_out[4273]);
     layer3_out[8735] <= ~(layer2_out[3095] ^ layer2_out[3096]);
     layer3_out[8736] <= ~layer2_out[687];
     layer3_out[8737] <= ~(layer2_out[4930] ^ layer2_out[4931]);
     layer3_out[8738] <= layer2_out[7038] & ~layer2_out[7037];
     layer3_out[8739] <= layer2_out[6249] ^ layer2_out[6250];
     layer3_out[8740] <= ~(layer2_out[11188] ^ layer2_out[11189]);
     layer3_out[8741] <= layer2_out[3419] ^ layer2_out[3420];
     layer3_out[8742] <= layer2_out[9203];
     layer3_out[8743] <= ~(layer2_out[2715] | layer2_out[2716]);
     layer3_out[8744] <= layer2_out[1145] & ~layer2_out[1146];
     layer3_out[8745] <= layer2_out[1853] & layer2_out[1854];
     layer3_out[8746] <= ~layer2_out[7964];
     layer3_out[8747] <= layer2_out[9401];
     layer3_out[8748] <= ~layer2_out[9865];
     layer3_out[8749] <= layer2_out[1954];
     layer3_out[8750] <= layer2_out[362] ^ layer2_out[363];
     layer3_out[8751] <= ~(layer2_out[11054] ^ layer2_out[11055]);
     layer3_out[8752] <= ~(layer2_out[4091] ^ layer2_out[4092]);
     layer3_out[8753] <= ~layer2_out[11072];
     layer3_out[8754] <= ~(layer2_out[6800] | layer2_out[6801]);
     layer3_out[8755] <= layer2_out[9218] | layer2_out[9219];
     layer3_out[8756] <= layer2_out[4937];
     layer3_out[8757] <= layer2_out[621];
     layer3_out[8758] <= ~layer2_out[10906] | layer2_out[10907];
     layer3_out[8759] <= ~layer2_out[2181];
     layer3_out[8760] <= layer2_out[4926] & ~layer2_out[4925];
     layer3_out[8761] <= ~layer2_out[5431];
     layer3_out[8762] <= layer2_out[4062] | layer2_out[4063];
     layer3_out[8763] <= ~(layer2_out[11611] | layer2_out[11612]);
     layer3_out[8764] <= ~(layer2_out[1684] | layer2_out[1685]);
     layer3_out[8765] <= ~layer2_out[1863];
     layer3_out[8766] <= layer2_out[9423] ^ layer2_out[9424];
     layer3_out[8767] <= ~layer2_out[3362] | layer2_out[3361];
     layer3_out[8768] <= layer2_out[2647];
     layer3_out[8769] <= ~layer2_out[7206];
     layer3_out[8770] <= layer2_out[11950] & ~layer2_out[11949];
     layer3_out[8771] <= layer2_out[360] | layer2_out[361];
     layer3_out[8772] <= ~layer2_out[8543];
     layer3_out[8773] <= layer2_out[2178] ^ layer2_out[2179];
     layer3_out[8774] <= layer2_out[2214];
     layer3_out[8775] <= layer2_out[90] & ~layer2_out[91];
     layer3_out[8776] <= layer2_out[6500] & ~layer2_out[6501];
     layer3_out[8777] <= ~(layer2_out[8788] & layer2_out[8789]);
     layer3_out[8778] <= ~(layer2_out[11315] & layer2_out[11316]);
     layer3_out[8779] <= ~layer2_out[3390];
     layer3_out[8780] <= layer2_out[8148];
     layer3_out[8781] <= ~layer2_out[9509] | layer2_out[9508];
     layer3_out[8782] <= ~layer2_out[3918] | layer2_out[3919];
     layer3_out[8783] <= ~layer2_out[80];
     layer3_out[8784] <= layer2_out[10585];
     layer3_out[8785] <= ~layer2_out[1994];
     layer3_out[8786] <= layer2_out[10491] ^ layer2_out[10492];
     layer3_out[8787] <= ~layer2_out[762];
     layer3_out[8788] <= ~layer2_out[5471];
     layer3_out[8789] <= ~layer2_out[336] | layer2_out[335];
     layer3_out[8790] <= layer2_out[9059] & layer2_out[9060];
     layer3_out[8791] <= layer2_out[9142] ^ layer2_out[9143];
     layer3_out[8792] <= ~(layer2_out[10526] & layer2_out[10527]);
     layer3_out[8793] <= ~(layer2_out[7399] & layer2_out[7400]);
     layer3_out[8794] <= layer2_out[6099];
     layer3_out[8795] <= layer2_out[8205] & ~layer2_out[8206];
     layer3_out[8796] <= layer2_out[8306] | layer2_out[8307];
     layer3_out[8797] <= layer2_out[2095] ^ layer2_out[2096];
     layer3_out[8798] <= layer2_out[11147];
     layer3_out[8799] <= ~layer2_out[6398] | layer2_out[6399];
     layer3_out[8800] <= ~(layer2_out[8899] & layer2_out[8900]);
     layer3_out[8801] <= layer2_out[3396] ^ layer2_out[3397];
     layer3_out[8802] <= ~layer2_out[8192];
     layer3_out[8803] <= layer2_out[3706];
     layer3_out[8804] <= layer2_out[3375] & ~layer2_out[3374];
     layer3_out[8805] <= ~layer2_out[11956];
     layer3_out[8806] <= layer2_out[990];
     layer3_out[8807] <= layer2_out[9882];
     layer3_out[8808] <= ~layer2_out[8644];
     layer3_out[8809] <= layer2_out[6752];
     layer3_out[8810] <= layer2_out[5187];
     layer3_out[8811] <= layer2_out[9899] & ~layer2_out[9898];
     layer3_out[8812] <= ~(layer2_out[7690] ^ layer2_out[7691]);
     layer3_out[8813] <= ~(layer2_out[2221] ^ layer2_out[2222]);
     layer3_out[8814] <= layer2_out[10700] & layer2_out[10701];
     layer3_out[8815] <= layer2_out[2637] & ~layer2_out[2638];
     layer3_out[8816] <= ~layer2_out[11847];
     layer3_out[8817] <= ~(layer2_out[7720] | layer2_out[7721]);
     layer3_out[8818] <= ~layer2_out[11077];
     layer3_out[8819] <= ~(layer2_out[10589] ^ layer2_out[10590]);
     layer3_out[8820] <= ~layer2_out[11530];
     layer3_out[8821] <= layer2_out[2496];
     layer3_out[8822] <= layer2_out[3934];
     layer3_out[8823] <= layer2_out[3675];
     layer3_out[8824] <= layer2_out[176];
     layer3_out[8825] <= layer2_out[7955];
     layer3_out[8826] <= layer2_out[3651];
     layer3_out[8827] <= layer2_out[11972];
     layer3_out[8828] <= layer2_out[8557] ^ layer2_out[8558];
     layer3_out[8829] <= layer2_out[7288] | layer2_out[7289];
     layer3_out[8830] <= ~layer2_out[1719] | layer2_out[1720];
     layer3_out[8831] <= layer2_out[8914] | layer2_out[8915];
     layer3_out[8832] <= layer2_out[9225];
     layer3_out[8833] <= layer2_out[670];
     layer3_out[8834] <= layer2_out[9476] & layer2_out[9477];
     layer3_out[8835] <= layer2_out[3591];
     layer3_out[8836] <= layer2_out[3990];
     layer3_out[8837] <= ~(layer2_out[8096] & layer2_out[8097]);
     layer3_out[8838] <= ~(layer2_out[10520] ^ layer2_out[10521]);
     layer3_out[8839] <= ~layer2_out[9048] | layer2_out[9047];
     layer3_out[8840] <= layer2_out[6778] ^ layer2_out[6779];
     layer3_out[8841] <= layer2_out[10910] & layer2_out[10911];
     layer3_out[8842] <= layer2_out[7165];
     layer3_out[8843] <= layer2_out[11805];
     layer3_out[8844] <= ~layer2_out[4072];
     layer3_out[8845] <= layer2_out[7929] & ~layer2_out[7930];
     layer3_out[8846] <= ~layer2_out[5473];
     layer3_out[8847] <= layer2_out[109] | layer2_out[110];
     layer3_out[8848] <= layer2_out[1717];
     layer3_out[8849] <= ~layer2_out[8151];
     layer3_out[8850] <= ~layer2_out[8303];
     layer3_out[8851] <= layer2_out[6308] ^ layer2_out[6309];
     layer3_out[8852] <= layer2_out[7245] & ~layer2_out[7246];
     layer3_out[8853] <= layer2_out[892];
     layer3_out[8854] <= layer2_out[406] & ~layer2_out[405];
     layer3_out[8855] <= layer2_out[1149] ^ layer2_out[1150];
     layer3_out[8856] <= ~layer2_out[9184];
     layer3_out[8857] <= ~layer2_out[6642];
     layer3_out[8858] <= ~layer2_out[3289];
     layer3_out[8859] <= layer2_out[1584] ^ layer2_out[1585];
     layer3_out[8860] <= ~layer2_out[2827];
     layer3_out[8861] <= ~layer2_out[9549];
     layer3_out[8862] <= ~layer2_out[1230];
     layer3_out[8863] <= layer2_out[4597] & ~layer2_out[4598];
     layer3_out[8864] <= layer2_out[1061] & ~layer2_out[1062];
     layer3_out[8865] <= ~layer2_out[2286];
     layer3_out[8866] <= layer2_out[6565] & ~layer2_out[6566];
     layer3_out[8867] <= layer2_out[1937] | layer2_out[1938];
     layer3_out[8868] <= ~(layer2_out[3503] & layer2_out[3504]);
     layer3_out[8869] <= ~layer2_out[11342] | layer2_out[11343];
     layer3_out[8870] <= ~layer2_out[10508] | layer2_out[10507];
     layer3_out[8871] <= layer2_out[8244];
     layer3_out[8872] <= ~layer2_out[4267];
     layer3_out[8873] <= layer2_out[11441] & ~layer2_out[11442];
     layer3_out[8874] <= ~(layer2_out[1755] & layer2_out[1756]);
     layer3_out[8875] <= layer2_out[8888] & ~layer2_out[8889];
     layer3_out[8876] <= layer2_out[6898] & ~layer2_out[6897];
     layer3_out[8877] <= layer2_out[10879] & ~layer2_out[10880];
     layer3_out[8878] <= ~layer2_out[10772] | layer2_out[10773];
     layer3_out[8879] <= layer2_out[5233] & ~layer2_out[5234];
     layer3_out[8880] <= ~(layer2_out[1790] | layer2_out[1791]);
     layer3_out[8881] <= ~layer2_out[7312] | layer2_out[7311];
     layer3_out[8882] <= layer2_out[5377] & ~layer2_out[5376];
     layer3_out[8883] <= layer2_out[11208] & layer2_out[11209];
     layer3_out[8884] <= ~(layer2_out[7463] & layer2_out[7464]);
     layer3_out[8885] <= layer2_out[6217] | layer2_out[6218];
     layer3_out[8886] <= layer2_out[9932];
     layer3_out[8887] <= ~(layer2_out[11513] ^ layer2_out[11514]);
     layer3_out[8888] <= layer2_out[7396] & ~layer2_out[7395];
     layer3_out[8889] <= ~layer2_out[3827] | layer2_out[3826];
     layer3_out[8890] <= layer2_out[11461] | layer2_out[11462];
     layer3_out[8891] <= layer2_out[2838] ^ layer2_out[2839];
     layer3_out[8892] <= layer2_out[9530] | layer2_out[9531];
     layer3_out[8893] <= layer2_out[9190] & ~layer2_out[9189];
     layer3_out[8894] <= layer2_out[1116] | layer2_out[1117];
     layer3_out[8895] <= layer2_out[8007] & ~layer2_out[8008];
     layer3_out[8896] <= layer2_out[5414] & ~layer2_out[5415];
     layer3_out[8897] <= layer2_out[8539] & layer2_out[8540];
     layer3_out[8898] <= layer2_out[11270] & ~layer2_out[11269];
     layer3_out[8899] <= layer2_out[1360] & layer2_out[1361];
     layer3_out[8900] <= layer2_out[3714];
     layer3_out[8901] <= layer2_out[1465] | layer2_out[1466];
     layer3_out[8902] <= layer2_out[1280];
     layer3_out[8903] <= ~layer2_out[8387];
     layer3_out[8904] <= layer2_out[8639] ^ layer2_out[8640];
     layer3_out[8905] <= layer2_out[3296] & ~layer2_out[3297];
     layer3_out[8906] <= ~(layer2_out[5361] ^ layer2_out[5362]);
     layer3_out[8907] <= layer2_out[5222] | layer2_out[5223];
     layer3_out[8908] <= ~(layer2_out[7721] & layer2_out[7722]);
     layer3_out[8909] <= layer2_out[10909] | layer2_out[10910];
     layer3_out[8910] <= ~(layer2_out[1674] | layer2_out[1675]);
     layer3_out[8911] <= ~layer2_out[7803];
     layer3_out[8912] <= layer2_out[11034] ^ layer2_out[11035];
     layer3_out[8913] <= layer2_out[6326] | layer2_out[6327];
     layer3_out[8914] <= layer2_out[5757];
     layer3_out[8915] <= layer2_out[8428] & layer2_out[8429];
     layer3_out[8916] <= ~layer2_out[10125];
     layer3_out[8917] <= ~layer2_out[7403];
     layer3_out[8918] <= layer2_out[4262];
     layer3_out[8919] <= layer2_out[11706];
     layer3_out[8920] <= layer2_out[329] | layer2_out[330];
     layer3_out[8921] <= layer2_out[271] & ~layer2_out[270];
     layer3_out[8922] <= ~(layer2_out[9439] & layer2_out[9440]);
     layer3_out[8923] <= layer2_out[6884] & layer2_out[6885];
     layer3_out[8924] <= ~(layer2_out[4609] | layer2_out[4610]);
     layer3_out[8925] <= layer2_out[9278] | layer2_out[9279];
     layer3_out[8926] <= ~layer2_out[6833] | layer2_out[6832];
     layer3_out[8927] <= ~(layer2_out[11817] & layer2_out[11818]);
     layer3_out[8928] <= ~(layer2_out[2084] | layer2_out[2085]);
     layer3_out[8929] <= ~layer2_out[8028];
     layer3_out[8930] <= ~layer2_out[962];
     layer3_out[8931] <= layer2_out[3718] & ~layer2_out[3719];
     layer3_out[8932] <= ~(layer2_out[5086] | layer2_out[5087]);
     layer3_out[8933] <= layer2_out[6553];
     layer3_out[8934] <= layer2_out[9700] ^ layer2_out[9701];
     layer3_out[8935] <= layer2_out[2334];
     layer3_out[8936] <= ~(layer2_out[2546] ^ layer2_out[2547]);
     layer3_out[8937] <= ~(layer2_out[3022] ^ layer2_out[3023]);
     layer3_out[8938] <= ~(layer2_out[5231] ^ layer2_out[5232]);
     layer3_out[8939] <= layer2_out[1421] & layer2_out[1422];
     layer3_out[8940] <= layer2_out[4566];
     layer3_out[8941] <= layer2_out[7798] | layer2_out[7799];
     layer3_out[8942] <= layer2_out[143] & ~layer2_out[142];
     layer3_out[8943] <= layer2_out[2823] & layer2_out[2824];
     layer3_out[8944] <= layer2_out[10594];
     layer3_out[8945] <= layer2_out[4281];
     layer3_out[8946] <= ~(layer2_out[2200] & layer2_out[2201]);
     layer3_out[8947] <= ~(layer2_out[4624] | layer2_out[4625]);
     layer3_out[8948] <= ~layer2_out[9495] | layer2_out[9494];
     layer3_out[8949] <= ~layer2_out[322];
     layer3_out[8950] <= layer2_out[10819] & ~layer2_out[10818];
     layer3_out[8951] <= layer2_out[4269] ^ layer2_out[4270];
     layer3_out[8952] <= layer2_out[11197] | layer2_out[11198];
     layer3_out[8953] <= layer2_out[11601];
     layer3_out[8954] <= layer2_out[9452];
     layer3_out[8955] <= layer2_out[7928] & layer2_out[7929];
     layer3_out[8956] <= ~layer2_out[935] | layer2_out[936];
     layer3_out[8957] <= ~layer2_out[874];
     layer3_out[8958] <= ~layer2_out[130];
     layer3_out[8959] <= layer2_out[9815] | layer2_out[9816];
     layer3_out[8960] <= ~layer2_out[9407];
     layer3_out[8961] <= ~(layer2_out[5524] & layer2_out[5525]);
     layer3_out[8962] <= layer2_out[1724] & ~layer2_out[1723];
     layer3_out[8963] <= layer2_out[5796] ^ layer2_out[5797];
     layer3_out[8964] <= ~(layer2_out[1193] & layer2_out[1194]);
     layer3_out[8965] <= layer2_out[2967] | layer2_out[2968];
     layer3_out[8966] <= layer2_out[9413];
     layer3_out[8967] <= layer2_out[1856] ^ layer2_out[1857];
     layer3_out[8968] <= layer2_out[8416] ^ layer2_out[8417];
     layer3_out[8969] <= ~(layer2_out[1721] | layer2_out[1722]);
     layer3_out[8970] <= layer2_out[8962] & ~layer2_out[8963];
     layer3_out[8971] <= layer2_out[7052];
     layer3_out[8972] <= ~layer2_out[11292];
     layer3_out[8973] <= layer2_out[8723];
     layer3_out[8974] <= ~layer2_out[8642];
     layer3_out[8975] <= layer2_out[11440] ^ layer2_out[11441];
     layer3_out[8976] <= layer2_out[10098] ^ layer2_out[10099];
     layer3_out[8977] <= layer2_out[11966] & layer2_out[11967];
     layer3_out[8978] <= layer2_out[1839];
     layer3_out[8979] <= ~layer2_out[7362];
     layer3_out[8980] <= ~(layer2_out[6715] | layer2_out[6716]);
     layer3_out[8981] <= layer2_out[3134] | layer2_out[3135];
     layer3_out[8982] <= layer2_out[6173] & layer2_out[6174];
     layer3_out[8983] <= ~(layer2_out[8583] | layer2_out[8584]);
     layer3_out[8984] <= ~layer2_out[9101];
     layer3_out[8985] <= ~(layer2_out[11449] | layer2_out[11450]);
     layer3_out[8986] <= layer2_out[4569] & ~layer2_out[4568];
     layer3_out[8987] <= ~layer2_out[9776];
     layer3_out[8988] <= ~(layer2_out[1017] ^ layer2_out[1018]);
     layer3_out[8989] <= ~(layer2_out[2804] | layer2_out[2805]);
     layer3_out[8990] <= layer2_out[5488];
     layer3_out[8991] <= layer2_out[3400];
     layer3_out[8992] <= ~layer2_out[6801];
     layer3_out[8993] <= ~(layer2_out[3562] ^ layer2_out[3563]);
     layer3_out[8994] <= ~(layer2_out[10048] ^ layer2_out[10049]);
     layer3_out[8995] <= ~layer2_out[2707];
     layer3_out[8996] <= layer2_out[4312] & layer2_out[4313];
     layer3_out[8997] <= ~layer2_out[11869];
     layer3_out[8998] <= layer2_out[6932];
     layer3_out[8999] <= layer2_out[5189];
     layer3_out[9000] <= layer2_out[8997];
     layer3_out[9001] <= layer2_out[2058] | layer2_out[2059];
     layer3_out[9002] <= layer2_out[2629] ^ layer2_out[2630];
     layer3_out[9003] <= layer2_out[8685] ^ layer2_out[8686];
     layer3_out[9004] <= layer2_out[5440];
     layer3_out[9005] <= ~(layer2_out[8443] ^ layer2_out[8444]);
     layer3_out[9006] <= ~(layer2_out[4024] | layer2_out[4025]);
     layer3_out[9007] <= layer2_out[20];
     layer3_out[9008] <= layer2_out[11582] & ~layer2_out[11583];
     layer3_out[9009] <= layer2_out[11705];
     layer3_out[9010] <= layer2_out[4531] ^ layer2_out[4532];
     layer3_out[9011] <= ~(layer2_out[5197] ^ layer2_out[5198]);
     layer3_out[9012] <= layer2_out[2590];
     layer3_out[9013] <= layer2_out[436] & ~layer2_out[437];
     layer3_out[9014] <= layer2_out[9283];
     layer3_out[9015] <= ~(layer2_out[6673] & layer2_out[6674]);
     layer3_out[9016] <= ~layer2_out[4694];
     layer3_out[9017] <= layer2_out[5348];
     layer3_out[9018] <= ~(layer2_out[6795] | layer2_out[6796]);
     layer3_out[9019] <= ~(layer2_out[1379] & layer2_out[1380]);
     layer3_out[9020] <= ~(layer2_out[2622] | layer2_out[2623]);
     layer3_out[9021] <= layer2_out[2950] | layer2_out[2951];
     layer3_out[9022] <= layer2_out[6164] & ~layer2_out[6163];
     layer3_out[9023] <= ~layer2_out[2900];
     layer3_out[9024] <= layer2_out[11091] | layer2_out[11092];
     layer3_out[9025] <= layer2_out[3293] & layer2_out[3294];
     layer3_out[9026] <= layer2_out[7543] & ~layer2_out[7544];
     layer3_out[9027] <= ~layer2_out[2139];
     layer3_out[9028] <= ~layer2_out[11618];
     layer3_out[9029] <= ~layer2_out[5877];
     layer3_out[9030] <= ~layer2_out[53];
     layer3_out[9031] <= ~(layer2_out[11882] | layer2_out[11883]);
     layer3_out[9032] <= layer2_out[1076];
     layer3_out[9033] <= ~layer2_out[1559];
     layer3_out[9034] <= ~(layer2_out[1451] | layer2_out[1452]);
     layer3_out[9035] <= ~layer2_out[7620] | layer2_out[7621];
     layer3_out[9036] <= ~(layer2_out[6232] ^ layer2_out[6233]);
     layer3_out[9037] <= ~layer2_out[2192];
     layer3_out[9038] <= layer2_out[5177] & layer2_out[5178];
     layer3_out[9039] <= ~(layer2_out[10136] ^ layer2_out[10137]);
     layer3_out[9040] <= ~layer2_out[1796];
     layer3_out[9041] <= ~layer2_out[9796] | layer2_out[9797];
     layer3_out[9042] <= layer2_out[7447] ^ layer2_out[7448];
     layer3_out[9043] <= layer2_out[5447];
     layer3_out[9044] <= layer2_out[9892];
     layer3_out[9045] <= ~layer2_out[3690];
     layer3_out[9046] <= ~(layer2_out[7623] ^ layer2_out[7624]);
     layer3_out[9047] <= layer2_out[8763];
     layer3_out[9048] <= layer2_out[11633] & ~layer2_out[11634];
     layer3_out[9049] <= ~layer2_out[2152] | layer2_out[2151];
     layer3_out[9050] <= layer2_out[2891] & layer2_out[2892];
     layer3_out[9051] <= ~(layer2_out[7866] ^ layer2_out[7867]);
     layer3_out[9052] <= layer2_out[1987];
     layer3_out[9053] <= ~(layer2_out[5567] | layer2_out[5568]);
     layer3_out[9054] <= ~layer2_out[10085];
     layer3_out[9055] <= ~(layer2_out[4453] ^ layer2_out[4454]);
     layer3_out[9056] <= ~(layer2_out[4584] ^ layer2_out[4585]);
     layer3_out[9057] <= ~layer2_out[2678];
     layer3_out[9058] <= layer2_out[8418];
     layer3_out[9059] <= layer2_out[9286] & ~layer2_out[9285];
     layer3_out[9060] <= layer2_out[7881];
     layer3_out[9061] <= layer2_out[1260];
     layer3_out[9062] <= layer2_out[9444] & layer2_out[9445];
     layer3_out[9063] <= layer2_out[1921] & ~layer2_out[1920];
     layer3_out[9064] <= layer2_out[2636] ^ layer2_out[2637];
     layer3_out[9065] <= layer2_out[2863] & ~layer2_out[2864];
     layer3_out[9066] <= ~layer2_out[10162] | layer2_out[10161];
     layer3_out[9067] <= ~layer2_out[1964];
     layer3_out[9068] <= ~layer2_out[11824] | layer2_out[11825];
     layer3_out[9069] <= layer2_out[2054] ^ layer2_out[2055];
     layer3_out[9070] <= ~layer2_out[1213];
     layer3_out[9071] <= layer2_out[6575];
     layer3_out[9072] <= ~layer2_out[7264];
     layer3_out[9073] <= ~layer2_out[1593];
     layer3_out[9074] <= layer2_out[7268] ^ layer2_out[7269];
     layer3_out[9075] <= layer2_out[1236];
     layer3_out[9076] <= ~(layer2_out[910] ^ layer2_out[911]);
     layer3_out[9077] <= ~layer2_out[3530];
     layer3_out[9078] <= layer2_out[8060];
     layer3_out[9079] <= layer2_out[7334] ^ layer2_out[7335];
     layer3_out[9080] <= layer2_out[3626] | layer2_out[3627];
     layer3_out[9081] <= ~layer2_out[5498];
     layer3_out[9082] <= ~layer2_out[10397];
     layer3_out[9083] <= layer2_out[2811] ^ layer2_out[2812];
     layer3_out[9084] <= layer2_out[1705] & layer2_out[1706];
     layer3_out[9085] <= layer2_out[754] & layer2_out[755];
     layer3_out[9086] <= ~(layer2_out[1576] ^ layer2_out[1577]);
     layer3_out[9087] <= ~layer2_out[6673] | layer2_out[6672];
     layer3_out[9088] <= layer2_out[3668];
     layer3_out[9089] <= ~layer2_out[8136];
     layer3_out[9090] <= layer2_out[5531] & layer2_out[5532];
     layer3_out[9091] <= ~layer2_out[7535];
     layer3_out[9092] <= ~(layer2_out[3380] ^ layer2_out[3381]);
     layer3_out[9093] <= ~(layer2_out[8434] & layer2_out[8435]);
     layer3_out[9094] <= layer2_out[6898] & ~layer2_out[6899];
     layer3_out[9095] <= layer2_out[8352];
     layer3_out[9096] <= layer2_out[544];
     layer3_out[9097] <= ~layer2_out[3873];
     layer3_out[9098] <= layer2_out[5690];
     layer3_out[9099] <= ~(layer2_out[10105] | layer2_out[10106]);
     layer3_out[9100] <= ~layer2_out[1354] | layer2_out[1353];
     layer3_out[9101] <= layer2_out[1128] & ~layer2_out[1127];
     layer3_out[9102] <= layer2_out[5555] ^ layer2_out[5556];
     layer3_out[9103] <= ~(layer2_out[10739] | layer2_out[10740]);
     layer3_out[9104] <= ~layer2_out[1362] | layer2_out[1363];
     layer3_out[9105] <= layer2_out[5735];
     layer3_out[9106] <= layer2_out[5015] ^ layer2_out[5016];
     layer3_out[9107] <= layer2_out[4592] & layer2_out[4593];
     layer3_out[9108] <= layer2_out[780] & ~layer2_out[781];
     layer3_out[9109] <= layer2_out[5268] | layer2_out[5269];
     layer3_out[9110] <= ~layer2_out[262] | layer2_out[263];
     layer3_out[9111] <= ~(layer2_out[2041] ^ layer2_out[2042]);
     layer3_out[9112] <= ~layer2_out[2437];
     layer3_out[9113] <= ~layer2_out[8787];
     layer3_out[9114] <= layer2_out[272];
     layer3_out[9115] <= layer2_out[4171] & layer2_out[4172];
     layer3_out[9116] <= layer2_out[175] & layer2_out[176];
     layer3_out[9117] <= layer2_out[10641] & ~layer2_out[10640];
     layer3_out[9118] <= layer2_out[4556];
     layer3_out[9119] <= layer2_out[10883] & ~layer2_out[10882];
     layer3_out[9120] <= ~(layer2_out[9854] | layer2_out[9855]);
     layer3_out[9121] <= ~(layer2_out[8625] | layer2_out[8626]);
     layer3_out[9122] <= layer2_out[7567] & layer2_out[7568];
     layer3_out[9123] <= layer2_out[10230];
     layer3_out[9124] <= layer2_out[4035] & layer2_out[4036];
     layer3_out[9125] <= ~layer2_out[6502];
     layer3_out[9126] <= ~(layer2_out[3443] ^ layer2_out[3444]);
     layer3_out[9127] <= ~(layer2_out[5768] & layer2_out[5769]);
     layer3_out[9128] <= ~layer2_out[6728] | layer2_out[6729];
     layer3_out[9129] <= ~layer2_out[1593];
     layer3_out[9130] <= ~layer2_out[11438];
     layer3_out[9131] <= ~layer2_out[1347];
     layer3_out[9132] <= ~layer2_out[7783];
     layer3_out[9133] <= ~layer2_out[7290];
     layer3_out[9134] <= layer2_out[7299];
     layer3_out[9135] <= layer2_out[11298] & ~layer2_out[11299];
     layer3_out[9136] <= ~(layer2_out[10005] & layer2_out[10006]);
     layer3_out[9137] <= layer2_out[8428];
     layer3_out[9138] <= ~(layer2_out[6621] ^ layer2_out[6622]);
     layer3_out[9139] <= layer2_out[3893];
     layer3_out[9140] <= ~layer2_out[8463];
     layer3_out[9141] <= layer2_out[5050];
     layer3_out[9142] <= ~(layer2_out[2361] & layer2_out[2362]);
     layer3_out[9143] <= layer2_out[6319] & ~layer2_out[6318];
     layer3_out[9144] <= ~(layer2_out[8121] | layer2_out[8122]);
     layer3_out[9145] <= ~layer2_out[6428];
     layer3_out[9146] <= ~layer2_out[10099] | layer2_out[10100];
     layer3_out[9147] <= ~(layer2_out[6131] & layer2_out[6132]);
     layer3_out[9148] <= layer2_out[3173];
     layer3_out[9149] <= ~(layer2_out[5389] & layer2_out[5390]);
     layer3_out[9150] <= ~layer2_out[9137];
     layer3_out[9151] <= layer2_out[4703] & layer2_out[4704];
     layer3_out[9152] <= layer2_out[7879] & ~layer2_out[7880];
     layer3_out[9153] <= layer2_out[9421];
     layer3_out[9154] <= layer2_out[5285];
     layer3_out[9155] <= ~layer2_out[9555];
     layer3_out[9156] <= layer2_out[3896] | layer2_out[3897];
     layer3_out[9157] <= layer2_out[8345] & layer2_out[8346];
     layer3_out[9158] <= layer2_out[7605];
     layer3_out[9159] <= layer2_out[7585] & layer2_out[7586];
     layer3_out[9160] <= layer2_out[10979] ^ layer2_out[10980];
     layer3_out[9161] <= layer2_out[3122] & layer2_out[3123];
     layer3_out[9162] <= layer2_out[4218] & layer2_out[4219];
     layer3_out[9163] <= layer2_out[3537];
     layer3_out[9164] <= layer2_out[4383];
     layer3_out[9165] <= layer2_out[11099];
     layer3_out[9166] <= ~(layer2_out[11559] ^ layer2_out[11560]);
     layer3_out[9167] <= layer2_out[957];
     layer3_out[9168] <= layer2_out[3212];
     layer3_out[9169] <= ~layer2_out[11883];
     layer3_out[9170] <= ~layer2_out[5663];
     layer3_out[9171] <= layer2_out[2198] | layer2_out[2199];
     layer3_out[9172] <= layer2_out[500];
     layer3_out[9173] <= layer2_out[5782];
     layer3_out[9174] <= layer2_out[40];
     layer3_out[9175] <= layer2_out[3500];
     layer3_out[9176] <= ~layer2_out[11485];
     layer3_out[9177] <= layer2_out[6251] ^ layer2_out[6252];
     layer3_out[9178] <= ~(layer2_out[8393] | layer2_out[8394]);
     layer3_out[9179] <= ~layer2_out[6276] | layer2_out[6277];
     layer3_out[9180] <= layer2_out[3222] ^ layer2_out[3223];
     layer3_out[9181] <= layer2_out[1400] & ~layer2_out[1399];
     layer3_out[9182] <= ~layer2_out[5608];
     layer3_out[9183] <= layer2_out[5969] & ~layer2_out[5968];
     layer3_out[9184] <= ~layer2_out[6692];
     layer3_out[9185] <= layer2_out[3765] & ~layer2_out[3766];
     layer3_out[9186] <= ~(layer2_out[7036] & layer2_out[7037]);
     layer3_out[9187] <= ~layer2_out[9639];
     layer3_out[9188] <= ~layer2_out[8438];
     layer3_out[9189] <= layer2_out[9433];
     layer3_out[9190] <= layer2_out[1545];
     layer3_out[9191] <= layer2_out[9703] | layer2_out[9704];
     layer3_out[9192] <= ~layer2_out[5628] | layer2_out[5627];
     layer3_out[9193] <= layer2_out[3079];
     layer3_out[9194] <= layer2_out[10864] & layer2_out[10865];
     layer3_out[9195] <= ~layer2_out[10438] | layer2_out[10437];
     layer3_out[9196] <= layer2_out[6445] & ~layer2_out[6446];
     layer3_out[9197] <= ~layer2_out[11399];
     layer3_out[9198] <= ~layer2_out[757];
     layer3_out[9199] <= ~(layer2_out[3033] & layer2_out[3034]);
     layer3_out[9200] <= ~(layer2_out[98] ^ layer2_out[99]);
     layer3_out[9201] <= ~layer2_out[2672];
     layer3_out[9202] <= ~(layer2_out[1569] | layer2_out[1570]);
     layer3_out[9203] <= layer2_out[4076];
     layer3_out[9204] <= ~layer2_out[4756] | layer2_out[4755];
     layer3_out[9205] <= ~(layer2_out[11463] ^ layer2_out[11464]);
     layer3_out[9206] <= ~layer2_out[1186];
     layer3_out[9207] <= ~layer2_out[9036] | layer2_out[9035];
     layer3_out[9208] <= ~layer2_out[4503];
     layer3_out[9209] <= layer2_out[1052];
     layer3_out[9210] <= layer2_out[7925];
     layer3_out[9211] <= ~(layer2_out[10884] ^ layer2_out[10885]);
     layer3_out[9212] <= layer2_out[4006];
     layer3_out[9213] <= layer2_out[3777] & ~layer2_out[3776];
     layer3_out[9214] <= layer2_out[2090];
     layer3_out[9215] <= ~layer2_out[1629];
     layer3_out[9216] <= ~(layer2_out[11695] ^ layer2_out[11696]);
     layer3_out[9217] <= ~(layer2_out[5741] & layer2_out[5742]);
     layer3_out[9218] <= ~(layer2_out[4064] | layer2_out[4065]);
     layer3_out[9219] <= ~(layer2_out[1502] | layer2_out[1503]);
     layer3_out[9220] <= layer2_out[7458];
     layer3_out[9221] <= ~layer2_out[6062];
     layer3_out[9222] <= ~layer2_out[9912] | layer2_out[9911];
     layer3_out[9223] <= ~layer2_out[2955];
     layer3_out[9224] <= ~(layer2_out[10175] & layer2_out[10176]);
     layer3_out[9225] <= ~(layer2_out[1882] ^ layer2_out[1883]);
     layer3_out[9226] <= ~layer2_out[565];
     layer3_out[9227] <= layer2_out[7560];
     layer3_out[9228] <= layer2_out[7813] & ~layer2_out[7814];
     layer3_out[9229] <= ~layer2_out[9407];
     layer3_out[9230] <= layer2_out[1535] & ~layer2_out[1534];
     layer3_out[9231] <= ~layer2_out[3949];
     layer3_out[9232] <= ~layer2_out[37];
     layer3_out[9233] <= layer2_out[4623];
     layer3_out[9234] <= layer2_out[2204];
     layer3_out[9235] <= ~(layer2_out[10745] ^ layer2_out[10746]);
     layer3_out[9236] <= layer2_out[6570];
     layer3_out[9237] <= ~layer2_out[256];
     layer3_out[9238] <= layer2_out[8672] & ~layer2_out[8673];
     layer3_out[9239] <= ~(layer2_out[4174] | layer2_out[4175]);
     layer3_out[9240] <= layer2_out[10585];
     layer3_out[9241] <= layer2_out[11632] & layer2_out[11633];
     layer3_out[9242] <= layer2_out[5767] & ~layer2_out[5766];
     layer3_out[9243] <= ~layer2_out[10826];
     layer3_out[9244] <= ~layer2_out[9232];
     layer3_out[9245] <= ~(layer2_out[10929] & layer2_out[10930]);
     layer3_out[9246] <= layer2_out[2276];
     layer3_out[9247] <= layer2_out[733];
     layer3_out[9248] <= layer2_out[8715];
     layer3_out[9249] <= ~layer2_out[6867];
     layer3_out[9250] <= layer2_out[8814];
     layer3_out[9251] <= ~(layer2_out[4758] & layer2_out[4759]);
     layer3_out[9252] <= layer2_out[8208];
     layer3_out[9253] <= ~layer2_out[7671];
     layer3_out[9254] <= layer2_out[8377] | layer2_out[8378];
     layer3_out[9255] <= layer2_out[4750];
     layer3_out[9256] <= layer2_out[1338] & ~layer2_out[1337];
     layer3_out[9257] <= ~layer2_out[11392] | layer2_out[11391];
     layer3_out[9258] <= layer2_out[4487];
     layer3_out[9259] <= ~layer2_out[4740];
     layer3_out[9260] <= layer2_out[6028];
     layer3_out[9261] <= ~layer2_out[1114];
     layer3_out[9262] <= layer2_out[6244];
     layer3_out[9263] <= ~layer2_out[3070] | layer2_out[3071];
     layer3_out[9264] <= ~layer2_out[8135];
     layer3_out[9265] <= ~layer2_out[9858];
     layer3_out[9266] <= ~(layer2_out[11518] | layer2_out[11519]);
     layer3_out[9267] <= ~layer2_out[2064];
     layer3_out[9268] <= layer2_out[7757];
     layer3_out[9269] <= ~layer2_out[2065] | layer2_out[2066];
     layer3_out[9270] <= layer2_out[8932] & layer2_out[8933];
     layer3_out[9271] <= layer2_out[8738];
     layer3_out[9272] <= layer2_out[213] & layer2_out[214];
     layer3_out[9273] <= ~(layer2_out[8105] | layer2_out[8106]);
     layer3_out[9274] <= layer2_out[3007];
     layer3_out[9275] <= layer2_out[3990];
     layer3_out[9276] <= layer2_out[840] ^ layer2_out[841];
     layer3_out[9277] <= ~layer2_out[9955];
     layer3_out[9278] <= ~(layer2_out[2238] ^ layer2_out[2239]);
     layer3_out[9279] <= ~layer2_out[5548];
     layer3_out[9280] <= layer2_out[2718] | layer2_out[2719];
     layer3_out[9281] <= ~layer2_out[11401];
     layer3_out[9282] <= layer2_out[7422] ^ layer2_out[7423];
     layer3_out[9283] <= ~layer2_out[10465];
     layer3_out[9284] <= layer2_out[11720];
     layer3_out[9285] <= ~(layer2_out[10461] | layer2_out[10462]);
     layer3_out[9286] <= layer2_out[4838] & ~layer2_out[4837];
     layer3_out[9287] <= layer2_out[5527] & ~layer2_out[5528];
     layer3_out[9288] <= layer2_out[10712];
     layer3_out[9289] <= ~layer2_out[4400] | layer2_out[4401];
     layer3_out[9290] <= ~(layer2_out[2351] ^ layer2_out[2352]);
     layer3_out[9291] <= layer2_out[8396];
     layer3_out[9292] <= layer2_out[387] | layer2_out[388];
     layer3_out[9293] <= ~layer2_out[10959];
     layer3_out[9294] <= ~layer2_out[8807] | layer2_out[8808];
     layer3_out[9295] <= ~layer2_out[582];
     layer3_out[9296] <= layer2_out[7472] ^ layer2_out[7473];
     layer3_out[9297] <= layer2_out[5540] & ~layer2_out[5541];
     layer3_out[9298] <= layer2_out[2746] ^ layer2_out[2747];
     layer3_out[9299] <= layer2_out[10097] ^ layer2_out[10098];
     layer3_out[9300] <= ~(layer2_out[1286] & layer2_out[1287]);
     layer3_out[9301] <= layer2_out[9862];
     layer3_out[9302] <= ~layer2_out[9970] | layer2_out[9971];
     layer3_out[9303] <= layer2_out[11871] | layer2_out[11872];
     layer3_out[9304] <= layer2_out[10116] & layer2_out[10117];
     layer3_out[9305] <= layer2_out[9876] ^ layer2_out[9877];
     layer3_out[9306] <= ~(layer2_out[11814] | layer2_out[11815]);
     layer3_out[9307] <= ~(layer2_out[8067] ^ layer2_out[8068]);
     layer3_out[9308] <= ~(layer2_out[2471] | layer2_out[2472]);
     layer3_out[9309] <= layer2_out[3753] ^ layer2_out[3754];
     layer3_out[9310] <= layer2_out[8048];
     layer3_out[9311] <= layer2_out[9270] & ~layer2_out[9271];
     layer3_out[9312] <= layer2_out[396];
     layer3_out[9313] <= ~layer2_out[3148] | layer2_out[3149];
     layer3_out[9314] <= layer2_out[10402] & layer2_out[10403];
     layer3_out[9315] <= layer2_out[7469] & ~layer2_out[7468];
     layer3_out[9316] <= ~layer2_out[10370] | layer2_out[10371];
     layer3_out[9317] <= layer2_out[6139] & layer2_out[6140];
     layer3_out[9318] <= layer2_out[4596] & ~layer2_out[4595];
     layer3_out[9319] <= layer2_out[6602];
     layer3_out[9320] <= ~layer2_out[2577] | layer2_out[2578];
     layer3_out[9321] <= layer2_out[7081] & layer2_out[7082];
     layer3_out[9322] <= ~(layer2_out[1456] ^ layer2_out[1457]);
     layer3_out[9323] <= layer2_out[2600] & ~layer2_out[2599];
     layer3_out[9324] <= ~layer2_out[5830];
     layer3_out[9325] <= ~(layer2_out[1891] ^ layer2_out[1892]);
     layer3_out[9326] <= layer2_out[6536] & ~layer2_out[6537];
     layer3_out[9327] <= layer2_out[3575] & layer2_out[3576];
     layer3_out[9328] <= layer2_out[9216] & ~layer2_out[9217];
     layer3_out[9329] <= ~(layer2_out[3609] | layer2_out[3610]);
     layer3_out[9330] <= ~layer2_out[6361] | layer2_out[6360];
     layer3_out[9331] <= ~(layer2_out[5632] ^ layer2_out[5633]);
     layer3_out[9332] <= ~(layer2_out[5280] & layer2_out[5281]);
     layer3_out[9333] <= ~layer2_out[11785] | layer2_out[11786];
     layer3_out[9334] <= ~layer2_out[6692];
     layer3_out[9335] <= layer2_out[10472] | layer2_out[10473];
     layer3_out[9336] <= ~(layer2_out[7101] & layer2_out[7102]);
     layer3_out[9337] <= ~layer2_out[10933];
     layer3_out[9338] <= ~layer2_out[11265];
     layer3_out[9339] <= ~(layer2_out[1929] & layer2_out[1930]);
     layer3_out[9340] <= layer2_out[1291] ^ layer2_out[1292];
     layer3_out[9341] <= ~layer2_out[8169] | layer2_out[8170];
     layer3_out[9342] <= layer2_out[3490] & ~layer2_out[3491];
     layer3_out[9343] <= ~(layer2_out[4215] | layer2_out[4216]);
     layer3_out[9344] <= ~layer2_out[11964];
     layer3_out[9345] <= ~layer2_out[5731] | layer2_out[5730];
     layer3_out[9346] <= layer2_out[8882] | layer2_out[8883];
     layer3_out[9347] <= layer2_out[2621];
     layer3_out[9348] <= layer2_out[6870];
     layer3_out[9349] <= ~(layer2_out[6523] | layer2_out[6524]);
     layer3_out[9350] <= layer2_out[972];
     layer3_out[9351] <= ~layer2_out[6694];
     layer3_out[9352] <= layer2_out[9885] ^ layer2_out[9886];
     layer3_out[9353] <= layer2_out[8986];
     layer3_out[9354] <= layer2_out[7115] & ~layer2_out[7116];
     layer3_out[9355] <= ~(layer2_out[10531] | layer2_out[10532]);
     layer3_out[9356] <= ~layer2_out[7481];
     layer3_out[9357] <= ~layer2_out[3749];
     layer3_out[9358] <= ~layer2_out[5091];
     layer3_out[9359] <= ~(layer2_out[1356] | layer2_out[1357]);
     layer3_out[9360] <= layer2_out[11982];
     layer3_out[9361] <= ~(layer2_out[6768] ^ layer2_out[6769]);
     layer3_out[9362] <= ~(layer2_out[6610] | layer2_out[6611]);
     layer3_out[9363] <= ~(layer2_out[11659] | layer2_out[11660]);
     layer3_out[9364] <= ~layer2_out[10397];
     layer3_out[9365] <= ~layer2_out[3820] | layer2_out[3819];
     layer3_out[9366] <= ~(layer2_out[9791] | layer2_out[9792]);
     layer3_out[9367] <= layer2_out[6239];
     layer3_out[9368] <= layer2_out[5256] & ~layer2_out[5255];
     layer3_out[9369] <= layer2_out[11404] & ~layer2_out[11405];
     layer3_out[9370] <= layer2_out[7238];
     layer3_out[9371] <= layer2_out[7317];
     layer3_out[9372] <= layer2_out[9723];
     layer3_out[9373] <= layer2_out[9405] | layer2_out[9406];
     layer3_out[9374] <= ~layer2_out[5402] | layer2_out[5403];
     layer3_out[9375] <= layer2_out[2114] & ~layer2_out[2115];
     layer3_out[9376] <= ~layer2_out[10708] | layer2_out[10709];
     layer3_out[9377] <= ~layer2_out[9132] | layer2_out[9133];
     layer3_out[9378] <= ~layer2_out[8858] | layer2_out[8857];
     layer3_out[9379] <= ~(layer2_out[8020] & layer2_out[8021]);
     layer3_out[9380] <= ~layer2_out[2528];
     layer3_out[9381] <= ~layer2_out[9732] | layer2_out[9731];
     layer3_out[9382] <= ~(layer2_out[5572] ^ layer2_out[5573]);
     layer3_out[9383] <= layer2_out[5735];
     layer3_out[9384] <= layer2_out[5153];
     layer3_out[9385] <= ~(layer2_out[9923] | layer2_out[9924]);
     layer3_out[9386] <= layer2_out[1226] & ~layer2_out[1225];
     layer3_out[9387] <= layer2_out[11263] & ~layer2_out[11264];
     layer3_out[9388] <= ~layer2_out[5445] | layer2_out[5444];
     layer3_out[9389] <= ~layer2_out[5533];
     layer3_out[9390] <= layer2_out[8252];
     layer3_out[9391] <= ~layer2_out[7724];
     layer3_out[9392] <= ~layer2_out[11284];
     layer3_out[9393] <= layer2_out[3187] | layer2_out[3188];
     layer3_out[9394] <= layer2_out[682];
     layer3_out[9395] <= ~(layer2_out[59] | layer2_out[60]);
     layer3_out[9396] <= ~layer2_out[10077];
     layer3_out[9397] <= ~(layer2_out[1125] & layer2_out[1126]);
     layer3_out[9398] <= ~layer2_out[170];
     layer3_out[9399] <= layer2_out[10950];
     layer3_out[9400] <= ~layer2_out[8166] | layer2_out[8165];
     layer3_out[9401] <= ~layer2_out[11708];
     layer3_out[9402] <= layer2_out[7091] ^ layer2_out[7092];
     layer3_out[9403] <= layer2_out[7999];
     layer3_out[9404] <= ~layer2_out[7854] | layer2_out[7855];
     layer3_out[9405] <= ~(layer2_out[2884] & layer2_out[2885]);
     layer3_out[9406] <= layer2_out[1521];
     layer3_out[9407] <= layer2_out[2761];
     layer3_out[9408] <= layer2_out[10457] & ~layer2_out[10456];
     layer3_out[9409] <= layer2_out[9758] & ~layer2_out[9757];
     layer3_out[9410] <= layer2_out[2518] ^ layer2_out[2519];
     layer3_out[9411] <= ~layer2_out[7583];
     layer3_out[9412] <= layer2_out[11982] & ~layer2_out[11983];
     layer3_out[9413] <= layer2_out[8347] ^ layer2_out[8348];
     layer3_out[9414] <= ~layer2_out[3982] | layer2_out[3983];
     layer3_out[9415] <= layer2_out[4105] & layer2_out[4106];
     layer3_out[9416] <= ~(layer2_out[9088] & layer2_out[9089]);
     layer3_out[9417] <= layer2_out[2415] & ~layer2_out[2416];
     layer3_out[9418] <= layer2_out[707] & ~layer2_out[706];
     layer3_out[9419] <= layer2_out[1319];
     layer3_out[9420] <= ~layer2_out[10433];
     layer3_out[9421] <= ~(layer2_out[8982] ^ layer2_out[8983]);
     layer3_out[9422] <= layer2_out[9481] & ~layer2_out[9480];
     layer3_out[9423] <= ~layer2_out[4339];
     layer3_out[9424] <= layer2_out[5449];
     layer3_out[9425] <= layer2_out[8157];
     layer3_out[9426] <= layer2_out[10259] & ~layer2_out[10260];
     layer3_out[9427] <= layer2_out[3915];
     layer3_out[9428] <= layer2_out[7419] & ~layer2_out[7418];
     layer3_out[9429] <= layer2_out[1183] & layer2_out[1184];
     layer3_out[9430] <= layer2_out[2954] & ~layer2_out[2953];
     layer3_out[9431] <= layer2_out[2756];
     layer3_out[9432] <= ~layer2_out[9369] | layer2_out[9370];
     layer3_out[9433] <= ~layer2_out[5913];
     layer3_out[9434] <= ~layer2_out[9872] | layer2_out[9873];
     layer3_out[9435] <= ~layer2_out[1203];
     layer3_out[9436] <= ~(layer2_out[1636] & layer2_out[1637]);
     layer3_out[9437] <= ~(layer2_out[9183] ^ layer2_out[9184]);
     layer3_out[9438] <= layer2_out[7452];
     layer3_out[9439] <= ~layer2_out[4102];
     layer3_out[9440] <= ~(layer2_out[5362] ^ layer2_out[5363]);
     layer3_out[9441] <= layer2_out[10513] & ~layer2_out[10512];
     layer3_out[9442] <= layer2_out[7005];
     layer3_out[9443] <= ~(layer2_out[8149] | layer2_out[8150]);
     layer3_out[9444] <= layer2_out[4036] | layer2_out[4037];
     layer3_out[9445] <= layer2_out[5095];
     layer3_out[9446] <= layer2_out[811] & ~layer2_out[812];
     layer3_out[9447] <= ~layer2_out[9975];
     layer3_out[9448] <= layer2_out[120] ^ layer2_out[121];
     layer3_out[9449] <= ~layer2_out[8846] | layer2_out[8847];
     layer3_out[9450] <= layer2_out[5287] & layer2_out[5288];
     layer3_out[9451] <= layer2_out[7283];
     layer3_out[9452] <= layer2_out[2737] & ~layer2_out[2738];
     layer3_out[9453] <= layer2_out[901] ^ layer2_out[902];
     layer3_out[9454] <= layer2_out[5409];
     layer3_out[9455] <= layer2_out[5140] ^ layer2_out[5141];
     layer3_out[9456] <= layer2_out[848] & layer2_out[849];
     layer3_out[9457] <= ~layer2_out[6466];
     layer3_out[9458] <= ~layer2_out[1199];
     layer3_out[9459] <= layer2_out[2932] | layer2_out[2933];
     layer3_out[9460] <= ~(layer2_out[3936] & layer2_out[3937]);
     layer3_out[9461] <= layer2_out[6615] & ~layer2_out[6616];
     layer3_out[9462] <= layer2_out[11992];
     layer3_out[9463] <= layer2_out[8968] & layer2_out[8969];
     layer3_out[9464] <= ~layer2_out[1385];
     layer3_out[9465] <= layer2_out[8356] & layer2_out[8357];
     layer3_out[9466] <= layer2_out[9014];
     layer3_out[9467] <= layer2_out[7104] & ~layer2_out[7103];
     layer3_out[9468] <= ~layer2_out[10550] | layer2_out[10549];
     layer3_out[9469] <= layer2_out[1360];
     layer3_out[9470] <= ~layer2_out[7003];
     layer3_out[9471] <= layer2_out[66] | layer2_out[67];
     layer3_out[9472] <= ~layer2_out[1792];
     layer3_out[9473] <= ~layer2_out[10347];
     layer3_out[9474] <= ~(layer2_out[6049] ^ layer2_out[6050]);
     layer3_out[9475] <= layer2_out[11524] | layer2_out[11525];
     layer3_out[9476] <= layer2_out[685] | layer2_out[686];
     layer3_out[9477] <= layer2_out[5199];
     layer3_out[9478] <= ~layer2_out[2232] | layer2_out[2231];
     layer3_out[9479] <= layer2_out[9957] ^ layer2_out[9958];
     layer3_out[9480] <= layer2_out[11251];
     layer3_out[9481] <= layer2_out[2688] ^ layer2_out[2689];
     layer3_out[9482] <= layer2_out[8820];
     layer3_out[9483] <= ~(layer2_out[11585] ^ layer2_out[11586]);
     layer3_out[9484] <= ~layer2_out[10563] | layer2_out[10564];
     layer3_out[9485] <= layer2_out[11103];
     layer3_out[9486] <= layer2_out[6111] ^ layer2_out[6112];
     layer3_out[9487] <= ~layer2_out[2174] | layer2_out[2175];
     layer3_out[9488] <= layer2_out[7786] ^ layer2_out[7787];
     layer3_out[9489] <= layer2_out[770] & ~layer2_out[771];
     layer3_out[9490] <= ~layer2_out[6531] | layer2_out[6532];
     layer3_out[9491] <= ~layer2_out[6420];
     layer3_out[9492] <= ~layer2_out[10119];
     layer3_out[9493] <= ~layer2_out[2548];
     layer3_out[9494] <= ~layer2_out[2973];
     layer3_out[9495] <= ~layer2_out[1834];
     layer3_out[9496] <= ~(layer2_out[3322] | layer2_out[3323]);
     layer3_out[9497] <= ~layer2_out[6755];
     layer3_out[9498] <= layer2_out[8951] ^ layer2_out[8952];
     layer3_out[9499] <= layer2_out[1481];
     layer3_out[9500] <= layer2_out[7007] ^ layer2_out[7008];
     layer3_out[9501] <= ~(layer2_out[9113] | layer2_out[9114]);
     layer3_out[9502] <= layer2_out[8234];
     layer3_out[9503] <= ~layer2_out[283];
     layer3_out[9504] <= ~(layer2_out[5972] | layer2_out[5973]);
     layer3_out[9505] <= layer2_out[11878] ^ layer2_out[11879];
     layer3_out[9506] <= ~layer2_out[7851];
     layer3_out[9507] <= ~(layer2_out[7338] | layer2_out[7339]);
     layer3_out[9508] <= ~layer2_out[17] | layer2_out[18];
     layer3_out[9509] <= layer2_out[11673] & layer2_out[11674];
     layer3_out[9510] <= ~layer2_out[10446] | layer2_out[10447];
     layer3_out[9511] <= layer2_out[228] ^ layer2_out[229];
     layer3_out[9512] <= layer2_out[6208] | layer2_out[6209];
     layer3_out[9513] <= ~layer2_out[5675] | layer2_out[5674];
     layer3_out[9514] <= layer2_out[8230];
     layer3_out[9515] <= ~layer2_out[2011];
     layer3_out[9516] <= layer2_out[1437] | layer2_out[1438];
     layer3_out[9517] <= layer2_out[2753] ^ layer2_out[2754];
     layer3_out[9518] <= ~layer2_out[8442];
     layer3_out[9519] <= layer2_out[240];
     layer3_out[9520] <= ~layer2_out[7781];
     layer3_out[9521] <= layer2_out[1037];
     layer3_out[9522] <= layer2_out[10657] & ~layer2_out[10658];
     layer3_out[9523] <= layer2_out[10015];
     layer3_out[9524] <= ~(layer2_out[5769] & layer2_out[5770]);
     layer3_out[9525] <= ~layer2_out[8923];
     layer3_out[9526] <= ~(layer2_out[7569] | layer2_out[7570]);
     layer3_out[9527] <= layer2_out[5100];
     layer3_out[9528] <= layer2_out[32] & ~layer2_out[31];
     layer3_out[9529] <= ~(layer2_out[7664] ^ layer2_out[7665]);
     layer3_out[9530] <= ~layer2_out[10213] | layer2_out[10214];
     layer3_out[9531] <= layer2_out[9171];
     layer3_out[9532] <= layer2_out[11443] & ~layer2_out[11444];
     layer3_out[9533] <= ~(layer2_out[9012] | layer2_out[9013]);
     layer3_out[9534] <= layer2_out[1707];
     layer3_out[9535] <= ~layer2_out[8594];
     layer3_out[9536] <= ~layer2_out[3428];
     layer3_out[9537] <= ~(layer2_out[11029] | layer2_out[11030]);
     layer3_out[9538] <= layer2_out[5800];
     layer3_out[9539] <= ~layer2_out[493] | layer2_out[494];
     layer3_out[9540] <= ~(layer2_out[3186] ^ layer2_out[3187]);
     layer3_out[9541] <= ~layer2_out[10939];
     layer3_out[9542] <= ~layer2_out[5458] | layer2_out[5459];
     layer3_out[9543] <= ~layer2_out[10987] | layer2_out[10988];
     layer3_out[9544] <= ~(layer2_out[7096] | layer2_out[7097]);
     layer3_out[9545] <= layer2_out[7151];
     layer3_out[9546] <= ~layer2_out[10053] | layer2_out[10054];
     layer3_out[9547] <= ~layer2_out[8323];
     layer3_out[9548] <= layer2_out[11068];
     layer3_out[9549] <= layer2_out[32];
     layer3_out[9550] <= ~layer2_out[7675] | layer2_out[7676];
     layer3_out[9551] <= ~layer2_out[11667];
     layer3_out[9552] <= layer2_out[2927] & layer2_out[2928];
     layer3_out[9553] <= ~layer2_out[11472];
     layer3_out[9554] <= ~(layer2_out[9509] & layer2_out[9510]);
     layer3_out[9555] <= layer2_out[8939] & layer2_out[8940];
     layer3_out[9556] <= ~layer2_out[2223];
     layer3_out[9557] <= ~layer2_out[1687];
     layer3_out[9558] <= ~(layer2_out[7464] | layer2_out[7465]);
     layer3_out[9559] <= layer2_out[7292] ^ layer2_out[7293];
     layer3_out[9560] <= ~layer2_out[1927];
     layer3_out[9561] <= layer2_out[10167];
     layer3_out[9562] <= ~layer2_out[7648];
     layer3_out[9563] <= ~layer2_out[10800] | layer2_out[10801];
     layer3_out[9564] <= ~layer2_out[11922];
     layer3_out[9565] <= ~layer2_out[2369];
     layer3_out[9566] <= layer2_out[4944] ^ layer2_out[4945];
     layer3_out[9567] <= ~(layer2_out[7110] | layer2_out[7111]);
     layer3_out[9568] <= ~layer2_out[2703];
     layer3_out[9569] <= layer2_out[8544] & layer2_out[8545];
     layer3_out[9570] <= ~(layer2_out[10414] ^ layer2_out[10415]);
     layer3_out[9571] <= ~(layer2_out[5739] ^ layer2_out[5740]);
     layer3_out[9572] <= layer2_out[8011];
     layer3_out[9573] <= layer2_out[3161] & ~layer2_out[3160];
     layer3_out[9574] <= ~layer2_out[4958];
     layer3_out[9575] <= ~(layer2_out[7027] ^ layer2_out[7028]);
     layer3_out[9576] <= layer2_out[6664] | layer2_out[6665];
     layer3_out[9577] <= layer2_out[4461] | layer2_out[4462];
     layer3_out[9578] <= ~layer2_out[325] | layer2_out[324];
     layer3_out[9579] <= ~layer2_out[1625] | layer2_out[1624];
     layer3_out[9580] <= ~layer2_out[2882];
     layer3_out[9581] <= ~(layer2_out[8482] ^ layer2_out[8483]);
     layer3_out[9582] <= layer2_out[10109];
     layer3_out[9583] <= ~layer2_out[506] | layer2_out[505];
     layer3_out[9584] <= layer2_out[6913] ^ layer2_out[6914];
     layer3_out[9585] <= ~(layer2_out[8799] ^ layer2_out[8800]);
     layer3_out[9586] <= layer2_out[3657] & ~layer2_out[3656];
     layer3_out[9587] <= layer2_out[10325] & layer2_out[10326];
     layer3_out[9588] <= layer2_out[5896] & layer2_out[5897];
     layer3_out[9589] <= layer2_out[8036] | layer2_out[8037];
     layer3_out[9590] <= ~layer2_out[1562];
     layer3_out[9591] <= layer2_out[10877];
     layer3_out[9592] <= ~layer2_out[3045];
     layer3_out[9593] <= ~layer2_out[2530];
     layer3_out[9594] <= ~layer2_out[4481];
     layer3_out[9595] <= layer2_out[6454] ^ layer2_out[6455];
     layer3_out[9596] <= layer2_out[7808] & ~layer2_out[7809];
     layer3_out[9597] <= ~layer2_out[10838] | layer2_out[10837];
     layer3_out[9598] <= layer2_out[9880] & ~layer2_out[9881];
     layer3_out[9599] <= layer2_out[6112] ^ layer2_out[6113];
     layer3_out[9600] <= layer2_out[10737];
     layer3_out[9601] <= ~layer2_out[6812] | layer2_out[6811];
     layer3_out[9602] <= layer2_out[6959] ^ layer2_out[6960];
     layer3_out[9603] <= layer2_out[1383] & ~layer2_out[1382];
     layer3_out[9604] <= ~layer2_out[1054];
     layer3_out[9605] <= layer2_out[8466] & layer2_out[8467];
     layer3_out[9606] <= layer2_out[4412] | layer2_out[4413];
     layer3_out[9607] <= ~layer2_out[11184];
     layer3_out[9608] <= layer2_out[10170] ^ layer2_out[10171];
     layer3_out[9609] <= layer2_out[6158] & layer2_out[6159];
     layer3_out[9610] <= layer2_out[3688];
     layer3_out[9611] <= ~(layer2_out[7425] & layer2_out[7426]);
     layer3_out[9612] <= ~(layer2_out[8876] | layer2_out[8877]);
     layer3_out[9613] <= layer2_out[7352] & ~layer2_out[7351];
     layer3_out[9614] <= ~layer2_out[612] | layer2_out[611];
     layer3_out[9615] <= layer2_out[3083] & layer2_out[3084];
     layer3_out[9616] <= ~(layer2_out[11168] | layer2_out[11169]);
     layer3_out[9617] <= ~(layer2_out[1066] | layer2_out[1067]);
     layer3_out[9618] <= ~layer2_out[3590];
     layer3_out[9619] <= layer2_out[3184];
     layer3_out[9620] <= ~(layer2_out[6236] ^ layer2_out[6237]);
     layer3_out[9621] <= layer2_out[10795] & ~layer2_out[10794];
     layer3_out[9622] <= layer2_out[11652];
     layer3_out[9623] <= ~(layer2_out[929] | layer2_out[930]);
     layer3_out[9624] <= layer2_out[10318] ^ layer2_out[10319];
     layer3_out[9625] <= ~layer2_out[8330] | layer2_out[8331];
     layer3_out[9626] <= ~layer2_out[8701];
     layer3_out[9627] <= layer2_out[11658] ^ layer2_out[11659];
     layer3_out[9628] <= ~(layer2_out[5467] | layer2_out[5468]);
     layer3_out[9629] <= ~layer2_out[5261];
     layer3_out[9630] <= ~(layer2_out[8609] | layer2_out[8610]);
     layer3_out[9631] <= layer2_out[8049] & layer2_out[8050];
     layer3_out[9632] <= ~(layer2_out[8550] ^ layer2_out[8551]);
     layer3_out[9633] <= layer2_out[7050] & ~layer2_out[7049];
     layer3_out[9634] <= ~(layer2_out[5506] ^ layer2_out[5507]);
     layer3_out[9635] <= ~(layer2_out[988] | layer2_out[989]);
     layer3_out[9636] <= ~layer2_out[876];
     layer3_out[9637] <= ~layer2_out[7893];
     layer3_out[9638] <= layer2_out[11412];
     layer3_out[9639] <= ~layer2_out[11242];
     layer3_out[9640] <= ~(layer2_out[7838] ^ layer2_out[7839]);
     layer3_out[9641] <= layer2_out[11621] & ~layer2_out[11620];
     layer3_out[9642] <= layer2_out[7280] & ~layer2_out[7279];
     layer3_out[9643] <= layer2_out[4646] & layer2_out[4647];
     layer3_out[9644] <= layer2_out[353] ^ layer2_out[354];
     layer3_out[9645] <= layer2_out[3837];
     layer3_out[9646] <= ~layer2_out[5695];
     layer3_out[9647] <= layer2_out[2865] & ~layer2_out[2866];
     layer3_out[9648] <= layer2_out[3514];
     layer3_out[9649] <= layer2_out[4448] & layer2_out[4449];
     layer3_out[9650] <= layer2_out[9249] ^ layer2_out[9250];
     layer3_out[9651] <= layer2_out[2383] | layer2_out[2384];
     layer3_out[9652] <= ~layer2_out[3913];
     layer3_out[9653] <= layer2_out[5783] & ~layer2_out[5782];
     layer3_out[9654] <= layer2_out[8281] ^ layer2_out[8282];
     layer3_out[9655] <= ~layer2_out[155];
     layer3_out[9656] <= ~layer2_out[793] | layer2_out[792];
     layer3_out[9657] <= layer2_out[4520] & ~layer2_out[4519];
     layer3_out[9658] <= layer2_out[3011];
     layer3_out[9659] <= ~(layer2_out[10183] | layer2_out[10184]);
     layer3_out[9660] <= layer2_out[7687] | layer2_out[7688];
     layer3_out[9661] <= ~layer2_out[3540];
     layer3_out[9662] <= layer2_out[6085];
     layer3_out[9663] <= ~(layer2_out[4545] | layer2_out[4546]);
     layer3_out[9664] <= layer2_out[10895] & ~layer2_out[10896];
     layer3_out[9665] <= ~layer2_out[6442] | layer2_out[6443];
     layer3_out[9666] <= layer2_out[9693] | layer2_out[9694];
     layer3_out[9667] <= layer2_out[5855];
     layer3_out[9668] <= layer2_out[2772] | layer2_out[2773];
     layer3_out[9669] <= layer2_out[10983];
     layer3_out[9670] <= ~(layer2_out[5071] ^ layer2_out[5072]);
     layer3_out[9671] <= layer2_out[1627];
     layer3_out[9672] <= ~layer2_out[8935];
     layer3_out[9673] <= layer2_out[3682] ^ layer2_out[3683];
     layer3_out[9674] <= ~layer2_out[2378] | layer2_out[2379];
     layer3_out[9675] <= layer2_out[8917];
     layer3_out[9676] <= layer2_out[1780];
     layer3_out[9677] <= layer2_out[9703];
     layer3_out[9678] <= layer2_out[7632];
     layer3_out[9679] <= ~layer2_out[11961] | layer2_out[11960];
     layer3_out[9680] <= layer2_out[11749];
     layer3_out[9681] <= ~(layer2_out[3194] | layer2_out[3195]);
     layer3_out[9682] <= ~layer2_out[10122] | layer2_out[10121];
     layer3_out[9683] <= layer2_out[6667] & ~layer2_out[6666];
     layer3_out[9684] <= layer2_out[3446] & layer2_out[3447];
     layer3_out[9685] <= ~(layer2_out[8714] & layer2_out[8715]);
     layer3_out[9686] <= layer2_out[2610];
     layer3_out[9687] <= ~layer2_out[8367] | layer2_out[8366];
     layer3_out[9688] <= layer2_out[1463];
     layer3_out[9689] <= ~(layer2_out[851] | layer2_out[852]);
     layer3_out[9690] <= ~layer2_out[5625];
     layer3_out[9691] <= layer2_out[10514] & layer2_out[10515];
     layer3_out[9692] <= layer2_out[4056] & ~layer2_out[4055];
     layer3_out[9693] <= layer2_out[9770] & layer2_out[9771];
     layer3_out[9694] <= layer2_out[3047];
     layer3_out[9695] <= ~layer2_out[9737];
     layer3_out[9696] <= layer2_out[10920] & layer2_out[10921];
     layer3_out[9697] <= layer2_out[9607];
     layer3_out[9698] <= layer2_out[5809];
     layer3_out[9699] <= layer2_out[5337];
     layer3_out[9700] <= layer2_out[2318] & ~layer2_out[2319];
     layer3_out[9701] <= layer2_out[2109] & layer2_out[2110];
     layer3_out[9702] <= layer2_out[6568] & ~layer2_out[6567];
     layer3_out[9703] <= layer2_out[11715] ^ layer2_out[11716];
     layer3_out[9704] <= ~layer2_out[8628] | layer2_out[8627];
     layer3_out[9705] <= layer2_out[2929] & ~layer2_out[2930];
     layer3_out[9706] <= ~layer2_out[8752];
     layer3_out[9707] <= ~(layer2_out[4242] | layer2_out[4243]);
     layer3_out[9708] <= layer2_out[5726] & ~layer2_out[5725];
     layer3_out[9709] <= layer2_out[2271];
     layer3_out[9710] <= ~layer2_out[3784];
     layer3_out[9711] <= layer2_out[5826] & ~layer2_out[5825];
     layer3_out[9712] <= layer2_out[4309] & ~layer2_out[4310];
     layer3_out[9713] <= ~(layer2_out[4426] ^ layer2_out[4427]);
     layer3_out[9714] <= layer2_out[11281];
     layer3_out[9715] <= ~layer2_out[8034] | layer2_out[8035];
     layer3_out[9716] <= layer2_out[10682] ^ layer2_out[10683];
     layer3_out[9717] <= layer2_out[5748];
     layer3_out[9718] <= ~layer2_out[2926];
     layer3_out[9719] <= ~layer2_out[132];
     layer3_out[9720] <= layer2_out[3248] ^ layer2_out[3249];
     layer3_out[9721] <= ~(layer2_out[8017] | layer2_out[8018]);
     layer3_out[9722] <= layer2_out[7744] ^ layer2_out[7745];
     layer3_out[9723] <= layer2_out[8728] & layer2_out[8729];
     layer3_out[9724] <= layer2_out[9916];
     layer3_out[9725] <= ~layer2_out[3464];
     layer3_out[9726] <= layer2_out[9321] ^ layer2_out[9322];
     layer3_out[9727] <= layer2_out[1459] & ~layer2_out[1460];
     layer3_out[9728] <= layer2_out[3316] | layer2_out[3317];
     layer3_out[9729] <= layer2_out[7864] ^ layer2_out[7865];
     layer3_out[9730] <= layer2_out[1954] & layer2_out[1955];
     layer3_out[9731] <= layer2_out[2302];
     layer3_out[9732] <= layer2_out[4236] & ~layer2_out[4237];
     layer3_out[9733] <= ~(layer2_out[1370] ^ layer2_out[1371]);
     layer3_out[9734] <= layer2_out[10781] & ~layer2_out[10780];
     layer3_out[9735] <= layer2_out[2264];
     layer3_out[9736] <= layer2_out[1921] & layer2_out[1922];
     layer3_out[9737] <= layer2_out[1440] & layer2_out[1441];
     layer3_out[9738] <= layer2_out[6961];
     layer3_out[9739] <= ~layer2_out[10045];
     layer3_out[9740] <= ~(layer2_out[8139] | layer2_out[8140]);
     layer3_out[9741] <= layer2_out[2293] & ~layer2_out[2294];
     layer3_out[9742] <= layer2_out[6804] & ~layer2_out[6805];
     layer3_out[9743] <= ~layer2_out[2312] | layer2_out[2313];
     layer3_out[9744] <= layer2_out[8726] & ~layer2_out[8727];
     layer3_out[9745] <= layer2_out[8653];
     layer3_out[9746] <= ~(layer2_out[7025] | layer2_out[7026]);
     layer3_out[9747] <= ~(layer2_out[1323] & layer2_out[1324]);
     layer3_out[9748] <= ~layer2_out[8655];
     layer3_out[9749] <= layer2_out[1614] & ~layer2_out[1613];
     layer3_out[9750] <= ~layer2_out[1705] | layer2_out[1704];
     layer3_out[9751] <= layer2_out[1653] & layer2_out[1654];
     layer3_out[9752] <= ~layer2_out[9122];
     layer3_out[9753] <= layer2_out[7122] & ~layer2_out[7123];
     layer3_out[9754] <= ~(layer2_out[5030] | layer2_out[5031]);
     layer3_out[9755] <= layer2_out[7535];
     layer3_out[9756] <= layer2_out[7297];
     layer3_out[9757] <= layer2_out[9843] ^ layer2_out[9844];
     layer3_out[9758] <= layer2_out[10971] & ~layer2_out[10972];
     layer3_out[9759] <= layer2_out[1834] & ~layer2_out[1833];
     layer3_out[9760] <= ~layer2_out[3051] | layer2_out[3052];
     layer3_out[9761] <= layer2_out[1332];
     layer3_out[9762] <= ~layer2_out[10356];
     layer3_out[9763] <= layer2_out[9034] & ~layer2_out[9035];
     layer3_out[9764] <= ~layer2_out[3464] | layer2_out[3465];
     layer3_out[9765] <= layer2_out[9095];
     layer3_out[9766] <= ~layer2_out[26];
     layer3_out[9767] <= layer2_out[8574] & layer2_out[8575];
     layer3_out[9768] <= ~layer2_out[5590];
     layer3_out[9769] <= layer2_out[5403] ^ layer2_out[5404];
     layer3_out[9770] <= ~layer2_out[2340];
     layer3_out[9771] <= ~layer2_out[11257];
     layer3_out[9772] <= ~layer2_out[3349];
     layer3_out[9773] <= layer2_out[1087];
     layer3_out[9774] <= ~(layer2_out[1689] | layer2_out[1690]);
     layer3_out[9775] <= layer2_out[8529] | layer2_out[8530];
     layer3_out[9776] <= layer2_out[2615];
     layer3_out[9777] <= ~(layer2_out[1427] | layer2_out[1428]);
     layer3_out[9778] <= ~(layer2_out[1508] ^ layer2_out[1509]);
     layer3_out[9779] <= layer2_out[7431] & ~layer2_out[7430];
     layer3_out[9780] <= layer2_out[7949] & ~layer2_out[7948];
     layer3_out[9781] <= layer2_out[10981] & layer2_out[10982];
     layer3_out[9782] <= layer2_out[11803];
     layer3_out[9783] <= layer2_out[7844] & ~layer2_out[7843];
     layer3_out[9784] <= layer2_out[1493] & layer2_out[1494];
     layer3_out[9785] <= layer2_out[5768] & ~layer2_out[5767];
     layer3_out[9786] <= ~(layer2_out[6125] ^ layer2_out[6126]);
     layer3_out[9787] <= layer2_out[1678] & ~layer2_out[1679];
     layer3_out[9788] <= layer2_out[8101] & layer2_out[8102];
     layer3_out[9789] <= layer2_out[11707] & layer2_out[11708];
     layer3_out[9790] <= layer2_out[4631];
     layer3_out[9791] <= ~(layer2_out[679] ^ layer2_out[680]);
     layer3_out[9792] <= ~(layer2_out[1269] ^ layer2_out[1270]);
     layer3_out[9793] <= layer2_out[4143] & ~layer2_out[4144];
     layer3_out[9794] <= ~(layer2_out[9124] | layer2_out[9125]);
     layer3_out[9795] <= layer2_out[10537];
     layer3_out[9796] <= layer2_out[6031] & ~layer2_out[6030];
     layer3_out[9797] <= layer2_out[3126] ^ layer2_out[3127];
     layer3_out[9798] <= layer2_out[10502] & layer2_out[10503];
     layer3_out[9799] <= ~layer2_out[9460] | layer2_out[9461];
     layer3_out[9800] <= layer2_out[9207] & ~layer2_out[9208];
     layer3_out[9801] <= layer2_out[10691];
     layer3_out[9802] <= ~layer2_out[1138];
     layer3_out[9803] <= layer2_out[10299];
     layer3_out[9804] <= ~layer2_out[5640];
     layer3_out[9805] <= ~(layer2_out[3831] ^ layer2_out[3832]);
     layer3_out[9806] <= ~layer2_out[3876] | layer2_out[3877];
     layer3_out[9807] <= layer2_out[4760];
     layer3_out[9808] <= ~(layer2_out[7694] ^ layer2_out[7695]);
     layer3_out[9809] <= layer2_out[9676] & layer2_out[9677];
     layer3_out[9810] <= ~(layer2_out[6572] & layer2_out[6573]);
     layer3_out[9811] <= ~(layer2_out[6136] ^ layer2_out[6137]);
     layer3_out[9812] <= ~layer2_out[4540];
     layer3_out[9813] <= ~(layer2_out[73] | layer2_out[74]);
     layer3_out[9814] <= ~(layer2_out[998] | layer2_out[999]);
     layer3_out[9815] <= ~layer2_out[11987] | layer2_out[11988];
     layer3_out[9816] <= layer2_out[5899] ^ layer2_out[5900];
     layer3_out[9817] <= layer2_out[1525];
     layer3_out[9818] <= ~layer2_out[4336];
     layer3_out[9819] <= layer2_out[4869];
     layer3_out[9820] <= layer2_out[5701];
     layer3_out[9821] <= layer2_out[4523];
     layer3_out[9822] <= ~(layer2_out[4877] | layer2_out[4878]);
     layer3_out[9823] <= ~(layer2_out[2924] | layer2_out[2925]);
     layer3_out[9824] <= layer2_out[11533] & layer2_out[11534];
     layer3_out[9825] <= ~(layer2_out[2429] & layer2_out[2430]);
     layer3_out[9826] <= ~layer2_out[5] | layer2_out[6];
     layer3_out[9827] <= layer2_out[8578] & ~layer2_out[8579];
     layer3_out[9828] <= layer2_out[9366] & layer2_out[9367];
     layer3_out[9829] <= ~layer2_out[5329];
     layer3_out[9830] <= ~layer2_out[5484];
     layer3_out[9831] <= ~layer2_out[10437];
     layer3_out[9832] <= ~(layer2_out[10290] ^ layer2_out[10291]);
     layer3_out[9833] <= ~(layer2_out[3778] | layer2_out[3779]);
     layer3_out[9834] <= layer2_out[3086];
     layer3_out[9835] <= ~layer2_out[1376];
     layer3_out[9836] <= layer2_out[7065] & ~layer2_out[7064];
     layer3_out[9837] <= ~(layer2_out[6257] | layer2_out[6258]);
     layer3_out[9838] <= ~layer2_out[3894];
     layer3_out[9839] <= layer2_out[11205] & ~layer2_out[11204];
     layer3_out[9840] <= layer2_out[7084];
     layer3_out[9841] <= layer2_out[9968];
     layer3_out[9842] <= ~(layer2_out[11628] & layer2_out[11629]);
     layer3_out[9843] <= ~layer2_out[1320];
     layer3_out[9844] <= layer2_out[6355] & ~layer2_out[6356];
     layer3_out[9845] <= layer2_out[6794] ^ layer2_out[6795];
     layer3_out[9846] <= layer2_out[10155] | layer2_out[10156];
     layer3_out[9847] <= ~layer2_out[4437];
     layer3_out[9848] <= ~layer2_out[7416];
     layer3_out[9849] <= layer2_out[8397] & layer2_out[8398];
     layer3_out[9850] <= layer2_out[10486] & ~layer2_out[10487];
     layer3_out[9851] <= ~layer2_out[10179];
     layer3_out[9852] <= ~(layer2_out[3738] | layer2_out[3739]);
     layer3_out[9853] <= ~(layer2_out[9289] | layer2_out[9290]);
     layer3_out[9854] <= layer2_out[8855] & ~layer2_out[8856];
     layer3_out[9855] <= ~layer2_out[8617];
     layer3_out[9856] <= ~(layer2_out[10002] | layer2_out[10003]);
     layer3_out[9857] <= ~layer2_out[600];
     layer3_out[9858] <= layer2_out[6852] ^ layer2_out[6853];
     layer3_out[9859] <= ~layer2_out[267] | layer2_out[268];
     layer3_out[9860] <= layer2_out[1113] & ~layer2_out[1112];
     layer3_out[9861] <= layer2_out[7944] & ~layer2_out[7943];
     layer3_out[9862] <= layer2_out[2257] & layer2_out[2258];
     layer3_out[9863] <= layer2_out[11076];
     layer3_out[9864] <= layer2_out[1081];
     layer3_out[9865] <= layer2_out[9853];
     layer3_out[9866] <= ~layer2_out[7212];
     layer3_out[9867] <= ~(layer2_out[5212] ^ layer2_out[5213]);
     layer3_out[9868] <= ~layer2_out[7161] | layer2_out[7162];
     layer3_out[9869] <= layer2_out[482] & layer2_out[483];
     layer3_out[9870] <= ~layer2_out[4938];
     layer3_out[9871] <= layer2_out[3727];
     layer3_out[9872] <= layer2_out[11266] & layer2_out[11267];
     layer3_out[9873] <= layer2_out[79];
     layer3_out[9874] <= ~layer2_out[10315];
     layer3_out[9875] <= layer2_out[8229] ^ layer2_out[8230];
     layer3_out[9876] <= layer2_out[9874] & layer2_out[9875];
     layer3_out[9877] <= layer2_out[5588] ^ layer2_out[5589];
     layer3_out[9878] <= layer2_out[11241];
     layer3_out[9879] <= ~layer2_out[4635];
     layer3_out[9880] <= layer2_out[8611] & ~layer2_out[8612];
     layer3_out[9881] <= layer2_out[3147];
     layer3_out[9882] <= ~layer2_out[6210];
     layer3_out[9883] <= layer2_out[11058];
     layer3_out[9884] <= ~layer2_out[11424];
     layer3_out[9885] <= layer2_out[6339];
     layer3_out[9886] <= ~layer2_out[10565];
     layer3_out[9887] <= layer2_out[2220] & layer2_out[2221];
     layer3_out[9888] <= ~layer2_out[4867];
     layer3_out[9889] <= ~layer2_out[11482];
     layer3_out[9890] <= layer2_out[7209] | layer2_out[7210];
     layer3_out[9891] <= ~layer2_out[9314];
     layer3_out[9892] <= layer2_out[3534] & ~layer2_out[3535];
     layer3_out[9893] <= ~layer2_out[3395];
     layer3_out[9894] <= ~(layer2_out[2873] | layer2_out[2874]);
     layer3_out[9895] <= layer2_out[9233] & layer2_out[9234];
     layer3_out[9896] <= layer2_out[5365];
     layer3_out[9897] <= ~layer2_out[10635];
     layer3_out[9898] <= ~(layer2_out[8039] & layer2_out[8040]);
     layer3_out[9899] <= ~layer2_out[10052];
     layer3_out[9900] <= layer2_out[7771] | layer2_out[7772];
     layer3_out[9901] <= layer2_out[5580];
     layer3_out[9902] <= layer2_out[3468] & layer2_out[3469];
     layer3_out[9903] <= ~layer2_out[10451];
     layer3_out[9904] <= layer2_out[5951];
     layer3_out[9905] <= ~(layer2_out[132] | layer2_out[133]);
     layer3_out[9906] <= layer2_out[4574] & layer2_out[4575];
     layer3_out[9907] <= ~(layer2_out[5131] | layer2_out[5132]);
     layer3_out[9908] <= ~layer2_out[6718];
     layer3_out[9909] <= layer2_out[7593];
     layer3_out[9910] <= layer2_out[4065];
     layer3_out[9911] <= layer2_out[11195] | layer2_out[11196];
     layer3_out[9912] <= layer2_out[5243] & ~layer2_out[5242];
     layer3_out[9913] <= layer2_out[11465];
     layer3_out[9914] <= layer2_out[10569];
     layer3_out[9915] <= layer2_out[6750] ^ layer2_out[6751];
     layer3_out[9916] <= layer2_out[778];
     layer3_out[9917] <= layer2_out[10920];
     layer3_out[9918] <= ~(layer2_out[6117] ^ layer2_out[6118]);
     layer3_out[9919] <= layer2_out[9157] & ~layer2_out[9158];
     layer3_out[9920] <= ~layer2_out[7885];
     layer3_out[9921] <= layer2_out[11025];
     layer3_out[9922] <= ~(layer2_out[10697] ^ layer2_out[10698]);
     layer3_out[9923] <= layer2_out[1762] & layer2_out[1763];
     layer3_out[9924] <= layer2_out[10650] ^ layer2_out[10651];
     layer3_out[9925] <= layer2_out[8783] & ~layer2_out[8784];
     layer3_out[9926] <= ~layer2_out[6417];
     layer3_out[9927] <= ~layer2_out[8714];
     layer3_out[9928] <= layer2_out[3498] ^ layer2_out[3499];
     layer3_out[9929] <= ~layer2_out[6722];
     layer3_out[9930] <= ~(layer2_out[6496] | layer2_out[6497]);
     layer3_out[9931] <= layer2_out[11155] & ~layer2_out[11156];
     layer3_out[9932] <= ~layer2_out[5918];
     layer3_out[9933] <= layer2_out[9561];
     layer3_out[9934] <= ~layer2_out[7533];
     layer3_out[9935] <= layer2_out[11797] & ~layer2_out[11796];
     layer3_out[9936] <= ~(layer2_out[9521] ^ layer2_out[9522]);
     layer3_out[9937] <= ~layer2_out[8894];
     layer3_out[9938] <= ~layer2_out[11471] | layer2_out[11470];
     layer3_out[9939] <= ~(layer2_out[7540] & layer2_out[7541]);
     layer3_out[9940] <= ~(layer2_out[4295] | layer2_out[4296]);
     layer3_out[9941] <= layer2_out[1873] ^ layer2_out[1874];
     layer3_out[9942] <= layer2_out[7352];
     layer3_out[9943] <= ~(layer2_out[6682] & layer2_out[6683]);
     layer3_out[9944] <= ~layer2_out[6984];
     layer3_out[9945] <= layer2_out[3874] ^ layer2_out[3875];
     layer3_out[9946] <= layer2_out[7606] & layer2_out[7607];
     layer3_out[9947] <= layer2_out[10193] & ~layer2_out[10192];
     layer3_out[9948] <= layer2_out[9520] & ~layer2_out[9519];
     layer3_out[9949] <= ~(layer2_out[10354] ^ layer2_out[10355]);
     layer3_out[9950] <= layer2_out[8097];
     layer3_out[9951] <= ~layer2_out[3285];
     layer3_out[9952] <= layer2_out[2025];
     layer3_out[9953] <= layer2_out[5496] & layer2_out[5497];
     layer3_out[9954] <= layer2_out[11723];
     layer3_out[9955] <= ~layer2_out[8308];
     layer3_out[9956] <= layer2_out[8716];
     layer3_out[9957] <= ~(layer2_out[5310] & layer2_out[5311]);
     layer3_out[9958] <= ~(layer2_out[10588] & layer2_out[10589]);
     layer3_out[9959] <= layer2_out[2709] ^ layer2_out[2710];
     layer3_out[9960] <= layer2_out[8103] & layer2_out[8104];
     layer3_out[9961] <= layer2_out[8907];
     layer3_out[9962] <= layer2_out[7050];
     layer3_out[9963] <= layer2_out[7170];
     layer3_out[9964] <= layer2_out[11000] & ~layer2_out[10999];
     layer3_out[9965] <= ~layer2_out[801];
     layer3_out[9966] <= layer2_out[5893];
     layer3_out[9967] <= layer2_out[6633] ^ layer2_out[6634];
     layer3_out[9968] <= ~layer2_out[657];
     layer3_out[9969] <= ~layer2_out[5158];
     layer3_out[9970] <= layer2_out[8861] & ~layer2_out[8860];
     layer3_out[9971] <= layer2_out[4826];
     layer3_out[9972] <= layer2_out[11049];
     layer3_out[9973] <= ~layer2_out[2429];
     layer3_out[9974] <= ~layer2_out[3365] | layer2_out[3366];
     layer3_out[9975] <= layer2_out[8963] | layer2_out[8964];
     layer3_out[9976] <= layer2_out[8228] & layer2_out[8229];
     layer3_out[9977] <= ~layer2_out[7763];
     layer3_out[9978] <= ~layer2_out[886];
     layer3_out[9979] <= layer2_out[3670] | layer2_out[3671];
     layer3_out[9980] <= ~layer2_out[9445];
     layer3_out[9981] <= ~(layer2_out[9265] & layer2_out[9266]);
     layer3_out[9982] <= ~layer2_out[3203];
     layer3_out[9983] <= ~(layer2_out[2936] | layer2_out[2937]);
     layer3_out[9984] <= ~(layer2_out[6449] ^ layer2_out[6450]);
     layer3_out[9985] <= layer2_out[8389] & ~layer2_out[8390];
     layer3_out[9986] <= layer2_out[11877] & layer2_out[11878];
     layer3_out[9987] <= ~layer2_out[2721];
     layer3_out[9988] <= ~(layer2_out[11911] | layer2_out[11912]);
     layer3_out[9989] <= layer2_out[1899] & layer2_out[1900];
     layer3_out[9990] <= layer2_out[2553];
     layer3_out[9991] <= ~layer2_out[7370];
     layer3_out[9992] <= layer2_out[9527] & ~layer2_out[9526];
     layer3_out[9993] <= ~layer2_out[5544];
     layer3_out[9994] <= layer2_out[2480];
     layer3_out[9995] <= ~layer2_out[6651];
     layer3_out[9996] <= ~layer2_out[2476] | layer2_out[2477];
     layer3_out[9997] <= layer2_out[3038];
     layer3_out[9998] <= layer2_out[9162] & ~layer2_out[9163];
     layer3_out[9999] <= layer2_out[1463];
     layer3_out[10000] <= ~layer2_out[3343];
     layer3_out[10001] <= layer2_out[4035] & ~layer2_out[4034];
     layer3_out[10002] <= ~layer2_out[4913];
     layer3_out[10003] <= layer2_out[8334] & ~layer2_out[8333];
     layer3_out[10004] <= ~layer2_out[8947];
     layer3_out[10005] <= layer2_out[11880] & layer2_out[11881];
     layer3_out[10006] <= layer2_out[9585] & ~layer2_out[9584];
     layer3_out[10007] <= ~layer2_out[6312];
     layer3_out[10008] <= layer2_out[10134] & ~layer2_out[10133];
     layer3_out[10009] <= ~layer2_out[4689];
     layer3_out[10010] <= ~layer2_out[2296];
     layer3_out[10011] <= layer2_out[7699] & layer2_out[7700];
     layer3_out[10012] <= layer2_out[2648];
     layer3_out[10013] <= ~layer2_out[5977];
     layer3_out[10014] <= ~layer2_out[4192];
     layer3_out[10015] <= layer2_out[7807];
     layer3_out[10016] <= ~layer2_out[7738];
     layer3_out[10017] <= ~layer2_out[5120] | layer2_out[5119];
     layer3_out[10018] <= ~layer2_out[10996] | layer2_out[10995];
     layer3_out[10019] <= ~(layer2_out[4416] | layer2_out[4417]);
     layer3_out[10020] <= layer2_out[4323];
     layer3_out[10021] <= layer2_out[8236] ^ layer2_out[8237];
     layer3_out[10022] <= ~(layer2_out[7584] | layer2_out[7585]);
     layer3_out[10023] <= ~layer2_out[4028];
     layer3_out[10024] <= layer2_out[11081];
     layer3_out[10025] <= layer2_out[6393] ^ layer2_out[6394];
     layer3_out[10026] <= ~layer2_out[6900] | layer2_out[6899];
     layer3_out[10027] <= ~(layer2_out[4780] ^ layer2_out[4781]);
     layer3_out[10028] <= layer2_out[1546];
     layer3_out[10029] <= ~layer2_out[6979];
     layer3_out[10030] <= ~layer2_out[3710];
     layer3_out[10031] <= layer2_out[7511] & ~layer2_out[7510];
     layer3_out[10032] <= layer2_out[8460];
     layer3_out[10033] <= layer2_out[6137] ^ layer2_out[6138];
     layer3_out[10034] <= ~layer2_out[3763];
     layer3_out[10035] <= ~layer2_out[7667] | layer2_out[7666];
     layer3_out[10036] <= ~(layer2_out[8003] | layer2_out[8004]);
     layer3_out[10037] <= layer2_out[2915];
     layer3_out[10038] <= ~(layer2_out[8348] & layer2_out[8349]);
     layer3_out[10039] <= ~layer2_out[11588];
     layer3_out[10040] <= layer2_out[8830] ^ layer2_out[8831];
     layer3_out[10041] <= layer2_out[11848];
     layer3_out[10042] <= ~(layer2_out[2043] | layer2_out[2044]);
     layer3_out[10043] <= ~layer2_out[4168] | layer2_out[4169];
     layer3_out[10044] <= layer2_out[2240] & ~layer2_out[2241];
     layer3_out[10045] <= layer2_out[5568];
     layer3_out[10046] <= layer2_out[4614] & ~layer2_out[4615];
     layer3_out[10047] <= layer2_out[7605] & layer2_out[7606];
     layer3_out[10048] <= layer2_out[1279] | layer2_out[1280];
     layer3_out[10049] <= ~layer2_out[10358];
     layer3_out[10050] <= ~(layer2_out[1619] | layer2_out[1620]);
     layer3_out[10051] <= ~layer2_out[2627];
     layer3_out[10052] <= ~(layer2_out[8706] | layer2_out[8707]);
     layer3_out[10053] <= layer2_out[9771] & layer2_out[9772];
     layer3_out[10054] <= ~layer2_out[9149];
     layer3_out[10055] <= layer2_out[2212] & ~layer2_out[2213];
     layer3_out[10056] <= ~(layer2_out[4175] ^ layer2_out[4176]);
     layer3_out[10057] <= ~(layer2_out[4792] & layer2_out[4793]);
     layer3_out[10058] <= layer2_out[7258] & ~layer2_out[7259];
     layer3_out[10059] <= ~(layer2_out[7797] | layer2_out[7798]);
     layer3_out[10060] <= ~layer2_out[11234];
     layer3_out[10061] <= layer2_out[7722] & ~layer2_out[7723];
     layer3_out[10062] <= layer2_out[4679];
     layer3_out[10063] <= layer2_out[10095];
     layer3_out[10064] <= layer2_out[9261];
     layer3_out[10065] <= layer2_out[3138] & ~layer2_out[3137];
     layer3_out[10066] <= layer2_out[2947] & layer2_out[2948];
     layer3_out[10067] <= ~layer2_out[6048];
     layer3_out[10068] <= ~(layer2_out[535] ^ layer2_out[536]);
     layer3_out[10069] <= ~(layer2_out[7432] ^ layer2_out[7433]);
     layer3_out[10070] <= ~layer2_out[1175];
     layer3_out[10071] <= ~layer2_out[1814] | layer2_out[1813];
     layer3_out[10072] <= layer2_out[10624] ^ layer2_out[10625];
     layer3_out[10073] <= layer2_out[9025];
     layer3_out[10074] <= layer2_out[9615] & layer2_out[9616];
     layer3_out[10075] <= ~layer2_out[753];
     layer3_out[10076] <= layer2_out[10617] & layer2_out[10618];
     layer3_out[10077] <= layer2_out[4080] & ~layer2_out[4081];
     layer3_out[10078] <= layer2_out[1615] & ~layer2_out[1616];
     layer3_out[10079] <= ~layer2_out[6579];
     layer3_out[10080] <= layer2_out[3225] & ~layer2_out[3226];
     layer3_out[10081] <= layer2_out[5231];
     layer3_out[10082] <= ~layer2_out[2680];
     layer3_out[10083] <= layer2_out[6164] ^ layer2_out[6165];
     layer3_out[10084] <= ~layer2_out[8906];
     layer3_out[10085] <= layer2_out[11000] & ~layer2_out[11001];
     layer3_out[10086] <= ~layer2_out[3999];
     layer3_out[10087] <= layer2_out[4129];
     layer3_out[10088] <= ~layer2_out[4173] | layer2_out[4172];
     layer3_out[10089] <= ~(layer2_out[136] | layer2_out[137]);
     layer3_out[10090] <= layer2_out[4590];
     layer3_out[10091] <= ~(layer2_out[10245] | layer2_out[10246]);
     layer3_out[10092] <= ~layer2_out[7364];
     layer3_out[10093] <= layer2_out[8412];
     layer3_out[10094] <= layer2_out[8305];
     layer3_out[10095] <= layer2_out[3655];
     layer3_out[10096] <= ~(layer2_out[527] ^ layer2_out[528]);
     layer3_out[10097] <= layer2_out[11543] ^ layer2_out[11544];
     layer3_out[10098] <= ~layer2_out[10675];
     layer3_out[10099] <= layer2_out[2067];
     layer3_out[10100] <= ~layer2_out[1681];
     layer3_out[10101] <= ~(layer2_out[4450] & layer2_out[4451]);
     layer3_out[10102] <= ~(layer2_out[162] ^ layer2_out[163]);
     layer3_out[10103] <= ~layer2_out[6831] | layer2_out[6832];
     layer3_out[10104] <= ~(layer2_out[7557] | layer2_out[7558]);
     layer3_out[10105] <= layer2_out[4697];
     layer3_out[10106] <= ~layer2_out[10292];
     layer3_out[10107] <= ~layer2_out[7466] | layer2_out[7465];
     layer3_out[10108] <= layer2_out[6931] & ~layer2_out[6932];
     layer3_out[10109] <= ~(layer2_out[193] | layer2_out[194]);
     layer3_out[10110] <= layer2_out[1718];
     layer3_out[10111] <= layer2_out[8671];
     layer3_out[10112] <= ~layer2_out[9986];
     layer3_out[10113] <= ~layer2_out[6926];
     layer3_out[10114] <= ~layer2_out[10896];
     layer3_out[10115] <= layer2_out[6996] & ~layer2_out[6995];
     layer3_out[10116] <= layer2_out[11701] & layer2_out[11702];
     layer3_out[10117] <= layer2_out[3167] & layer2_out[3168];
     layer3_out[10118] <= ~layer2_out[8613];
     layer3_out[10119] <= ~layer2_out[3088];
     layer3_out[10120] <= ~(layer2_out[9758] & layer2_out[9759]);
     layer3_out[10121] <= layer2_out[3677] & layer2_out[3678];
     layer3_out[10122] <= layer2_out[11968] & layer2_out[11969];
     layer3_out[10123] <= layer2_out[7490];
     layer3_out[10124] <= ~layer2_out[10858];
     layer3_out[10125] <= layer2_out[10169] ^ layer2_out[10170];
     layer3_out[10126] <= ~layer2_out[9295];
     layer3_out[10127] <= ~layer2_out[983];
     layer3_out[10128] <= ~layer2_out[6072];
     layer3_out[10129] <= layer2_out[5200];
     layer3_out[10130] <= ~layer2_out[11935];
     layer3_out[10131] <= layer2_out[8885] ^ layer2_out[8886];
     layer3_out[10132] <= layer2_out[5944] | layer2_out[5945];
     layer3_out[10133] <= layer2_out[2083] | layer2_out[2084];
     layer3_out[10134] <= layer2_out[6670] & ~layer2_out[6669];
     layer3_out[10135] <= layer2_out[7683] & ~layer2_out[7684];
     layer3_out[10136] <= ~(layer2_out[3736] | layer2_out[3737]);
     layer3_out[10137] <= ~layer2_out[6551];
     layer3_out[10138] <= ~layer2_out[4004];
     layer3_out[10139] <= ~layer2_out[8678];
     layer3_out[10140] <= ~(layer2_out[3683] ^ layer2_out[3684]);
     layer3_out[10141] <= layer2_out[3378] & ~layer2_out[3379];
     layer3_out[10142] <= layer2_out[11660] | layer2_out[11661];
     layer3_out[10143] <= layer2_out[1780];
     layer3_out[10144] <= ~(layer2_out[9833] ^ layer2_out[9834]);
     layer3_out[10145] <= ~layer2_out[3951];
     layer3_out[10146] <= layer2_out[4280] & layer2_out[4281];
     layer3_out[10147] <= layer2_out[6985] & ~layer2_out[6984];
     layer3_out[10148] <= layer2_out[8964] | layer2_out[8965];
     layer3_out[10149] <= layer2_out[4161] & ~layer2_out[4160];
     layer3_out[10150] <= layer2_out[11479] & ~layer2_out[11478];
     layer3_out[10151] <= ~layer2_out[11191] | layer2_out[11190];
     layer3_out[10152] <= ~layer2_out[8138] | layer2_out[8137];
     layer3_out[10153] <= layer2_out[9390];
     layer3_out[10154] <= layer2_out[6606];
     layer3_out[10155] <= layer2_out[10637];
     layer3_out[10156] <= ~(layer2_out[9963] ^ layer2_out[9964]);
     layer3_out[10157] <= layer2_out[7891];
     layer3_out[10158] <= layer2_out[4444] & ~layer2_out[4443];
     layer3_out[10159] <= ~(layer2_out[5955] & layer2_out[5956]);
     layer3_out[10160] <= ~layer2_out[9275] | layer2_out[9276];
     layer3_out[10161] <= layer2_out[3151];
     layer3_out[10162] <= ~(layer2_out[366] | layer2_out[367]);
     layer3_out[10163] <= layer2_out[10004];
     layer3_out[10164] <= layer2_out[6648] & layer2_out[6649];
     layer3_out[10165] <= ~layer2_out[10966] | layer2_out[10965];
     layer3_out[10166] <= ~layer2_out[4846] | layer2_out[4845];
     layer3_out[10167] <= ~layer2_out[6556] | layer2_out[6557];
     layer3_out[10168] <= layer2_out[1013] | layer2_out[1014];
     layer3_out[10169] <= layer2_out[10820] ^ layer2_out[10821];
     layer3_out[10170] <= layer2_out[11386];
     layer3_out[10171] <= layer2_out[10867] ^ layer2_out[10868];
     layer3_out[10172] <= ~(layer2_out[6345] | layer2_out[6346]);
     layer3_out[10173] <= ~layer2_out[4818];
     layer3_out[10174] <= ~layer2_out[3241] | layer2_out[3240];
     layer3_out[10175] <= layer2_out[11458] & layer2_out[11459];
     layer3_out[10176] <= layer2_out[6436];
     layer3_out[10177] <= ~(layer2_out[5638] & layer2_out[5639]);
     layer3_out[10178] <= layer2_out[7517];
     layer3_out[10179] <= layer2_out[161] & ~layer2_out[162];
     layer3_out[10180] <= layer2_out[8477] & layer2_out[8478];
     layer3_out[10181] <= ~layer2_out[11172] | layer2_out[11171];
     layer3_out[10182] <= layer2_out[2981];
     layer3_out[10183] <= ~layer2_out[9684];
     layer3_out[10184] <= layer2_out[11900] & ~layer2_out[11901];
     layer3_out[10185] <= layer2_out[9755] & layer2_out[9756];
     layer3_out[10186] <= layer2_out[5396];
     layer3_out[10187] <= layer2_out[1430] & layer2_out[1431];
     layer3_out[10188] <= layer2_out[5772];
     layer3_out[10189] <= layer2_out[8841];
     layer3_out[10190] <= ~layer2_out[6877];
     layer3_out[10191] <= layer2_out[6181];
     layer3_out[10192] <= layer2_out[330];
     layer3_out[10193] <= ~layer2_out[3267];
     layer3_out[10194] <= ~layer2_out[6448];
     layer3_out[10195] <= layer2_out[201];
     layer3_out[10196] <= layer2_out[10689] & ~layer2_out[10690];
     layer3_out[10197] <= ~(layer2_out[7034] & layer2_out[7035]);
     layer3_out[10198] <= ~layer2_out[5975] | layer2_out[5974];
     layer3_out[10199] <= layer2_out[4658];
     layer3_out[10200] <= layer2_out[300] ^ layer2_out[301];
     layer3_out[10201] <= layer2_out[6269] | layer2_out[6270];
     layer3_out[10202] <= layer2_out[9633];
     layer3_out[10203] <= ~(layer2_out[8498] ^ layer2_out[8499]);
     layer3_out[10204] <= ~(layer2_out[3717] ^ layer2_out[3718]);
     layer3_out[10205] <= ~(layer2_out[5358] | layer2_out[5359]);
     layer3_out[10206] <= ~(layer2_out[11980] & layer2_out[11981]);
     layer3_out[10207] <= ~layer2_out[7192];
     layer3_out[10208] <= layer2_out[8152];
     layer3_out[10209] <= layer2_out[11325] & layer2_out[11326];
     layer3_out[10210] <= layer2_out[7604] & ~layer2_out[7603];
     layer3_out[10211] <= ~(layer2_out[639] | layer2_out[640]);
     layer3_out[10212] <= layer2_out[11039] | layer2_out[11040];
     layer3_out[10213] <= layer2_out[6546];
     layer3_out[10214] <= ~layer2_out[8481];
     layer3_out[10215] <= ~(layer2_out[5592] & layer2_out[5593]);
     layer3_out[10216] <= ~layer2_out[2868];
     layer3_out[10217] <= layer2_out[6920];
     layer3_out[10218] <= ~layer2_out[2287];
     layer3_out[10219] <= ~layer2_out[11287];
     layer3_out[10220] <= layer2_out[4986];
     layer3_out[10221] <= layer2_out[2389];
     layer3_out[10222] <= ~layer2_out[265];
     layer3_out[10223] <= layer2_out[2766] | layer2_out[2767];
     layer3_out[10224] <= ~(layer2_out[9433] | layer2_out[9434]);
     layer3_out[10225] <= ~layer2_out[6483];
     layer3_out[10226] <= layer2_out[10787];
     layer3_out[10227] <= ~layer2_out[5723];
     layer3_out[10228] <= layer2_out[10260] & layer2_out[10261];
     layer3_out[10229] <= ~layer2_out[5791];
     layer3_out[10230] <= layer2_out[11763] & ~layer2_out[11764];
     layer3_out[10231] <= layer2_out[1070] ^ layer2_out[1071];
     layer3_out[10232] <= layer2_out[11586];
     layer3_out[10233] <= layer2_out[817] & ~layer2_out[816];
     layer3_out[10234] <= layer2_out[869];
     layer3_out[10235] <= ~(layer2_out[11052] ^ layer2_out[11053]);
     layer3_out[10236] <= layer2_out[7781] & layer2_out[7782];
     layer3_out[10237] <= layer2_out[9789] & ~layer2_out[9790];
     layer3_out[10238] <= ~(layer2_out[8634] ^ layer2_out[8635]);
     layer3_out[10239] <= layer2_out[10391] & ~layer2_out[10392];
     layer3_out[10240] <= layer2_out[8682] & ~layer2_out[8683];
     layer3_out[10241] <= layer2_out[1484];
     layer3_out[10242] <= ~(layer2_out[9097] ^ layer2_out[9098]);
     layer3_out[10243] <= layer2_out[2648] & layer2_out[2649];
     layer3_out[10244] <= layer2_out[2240];
     layer3_out[10245] <= layer2_out[1004] & layer2_out[1005];
     layer3_out[10246] <= layer2_out[3461];
     layer3_out[10247] <= layer2_out[2502] & ~layer2_out[2503];
     layer3_out[10248] <= layer2_out[4924];
     layer3_out[10249] <= layer2_out[5093];
     layer3_out[10250] <= ~layer2_out[3426];
     layer3_out[10251] <= ~(layer2_out[5875] | layer2_out[5876]);
     layer3_out[10252] <= ~layer2_out[8987] | layer2_out[8988];
     layer3_out[10253] <= layer2_out[86] & layer2_out[87];
     layer3_out[10254] <= layer2_out[10006] | layer2_out[10007];
     layer3_out[10255] <= layer2_out[5378] ^ layer2_out[5379];
     layer3_out[10256] <= ~(layer2_out[5226] & layer2_out[5227]);
     layer3_out[10257] <= layer2_out[10151] & ~layer2_out[10150];
     layer3_out[10258] <= layer2_out[11383] & layer2_out[11384];
     layer3_out[10259] <= ~layer2_out[7937];
     layer3_out[10260] <= layer2_out[6039];
     layer3_out[10261] <= layer2_out[6577] ^ layer2_out[6578];
     layer3_out[10262] <= layer2_out[8834];
     layer3_out[10263] <= layer2_out[3306] ^ layer2_out[3307];
     layer3_out[10264] <= ~(layer2_out[8688] ^ layer2_out[8689]);
     layer3_out[10265] <= ~(layer2_out[2320] ^ layer2_out[2321]);
     layer3_out[10266] <= ~(layer2_out[11243] ^ layer2_out[11244]);
     layer3_out[10267] <= ~layer2_out[8319];
     layer3_out[10268] <= layer2_out[5775];
     layer3_out[10269] <= ~(layer2_out[6148] ^ layer2_out[6149]);
     layer3_out[10270] <= layer2_out[6749] & ~layer2_out[6750];
     layer3_out[10271] <= ~(layer2_out[7777] ^ layer2_out[7778]);
     layer3_out[10272] <= ~(layer2_out[9679] | layer2_out[9680]);
     layer3_out[10273] <= layer2_out[7661];
     layer3_out[10274] <= layer2_out[9511];
     layer3_out[10275] <= layer2_out[10758];
     layer3_out[10276] <= layer2_out[5764] & ~layer2_out[5765];
     layer3_out[10277] <= ~layer2_out[1338] | layer2_out[1339];
     layer3_out[10278] <= layer2_out[8790];
     layer3_out[10279] <= ~layer2_out[5367];
     layer3_out[10280] <= layer2_out[4666] & layer2_out[4667];
     layer3_out[10281] <= layer2_out[2609] & layer2_out[2610];
     layer3_out[10282] <= ~layer2_out[7174] | layer2_out[7175];
     layer3_out[10283] <= ~layer2_out[7937];
     layer3_out[10284] <= ~(layer2_out[10405] | layer2_out[10406]);
     layer3_out[10285] <= layer2_out[8044] | layer2_out[8045];
     layer3_out[10286] <= layer2_out[288] & ~layer2_out[289];
     layer3_out[10287] <= layer2_out[6045] & ~layer2_out[6044];
     layer3_out[10288] <= layer2_out[9870] ^ layer2_out[9871];
     layer3_out[10289] <= layer2_out[2849];
     layer3_out[10290] <= ~layer2_out[11131] | layer2_out[11132];
     layer3_out[10291] <= ~layer2_out[9995] | layer2_out[9996];
     layer3_out[10292] <= ~(layer2_out[6594] ^ layer2_out[6595]);
     layer3_out[10293] <= layer2_out[3793];
     layer3_out[10294] <= layer2_out[3168];
     layer3_out[10295] <= layer2_out[5276];
     layer3_out[10296] <= ~layer2_out[11134];
     layer3_out[10297] <= ~(layer2_out[3412] | layer2_out[3413]);
     layer3_out[10298] <= layer2_out[1299];
     layer3_out[10299] <= layer2_out[10422];
     layer3_out[10300] <= layer2_out[5474] ^ layer2_out[5475];
     layer3_out[10301] <= ~layer2_out[11770];
     layer3_out[10302] <= layer2_out[2048] & layer2_out[2049];
     layer3_out[10303] <= ~layer2_out[1851];
     layer3_out[10304] <= layer2_out[10785] ^ layer2_out[10786];
     layer3_out[10305] <= ~(layer2_out[6224] | layer2_out[6225]);
     layer3_out[10306] <= layer2_out[6142];
     layer3_out[10307] <= layer2_out[11892];
     layer3_out[10308] <= layer2_out[285];
     layer3_out[10309] <= ~(layer2_out[10506] ^ layer2_out[10507]);
     layer3_out[10310] <= ~layer2_out[1879];
     layer3_out[10311] <= ~(layer2_out[9507] | layer2_out[9508]);
     layer3_out[10312] <= ~(layer2_out[8693] | layer2_out[8694]);
     layer3_out[10313] <= ~layer2_out[2248];
     layer3_out[10314] <= layer2_out[10678];
     layer3_out[10315] <= layer2_out[5021] & ~layer2_out[5020];
     layer3_out[10316] <= ~layer2_out[7506];
     layer3_out[10317] <= ~(layer2_out[293] & layer2_out[294]);
     layer3_out[10318] <= layer2_out[7488];
     layer3_out[10319] <= ~layer2_out[8735];
     layer3_out[10320] <= ~layer2_out[11113];
     layer3_out[10321] <= layer2_out[6109];
     layer3_out[10322] <= ~(layer2_out[11676] | layer2_out[11677]);
     layer3_out[10323] <= layer2_out[7583] & ~layer2_out[7584];
     layer3_out[10324] <= ~(layer2_out[49] ^ layer2_out[50]);
     layer3_out[10325] <= layer2_out[8900] & ~layer2_out[8901];
     layer3_out[10326] <= layer2_out[10430] & ~layer2_out[10429];
     layer3_out[10327] <= layer2_out[7176] & ~layer2_out[7177];
     layer3_out[10328] <= layer2_out[11803];
     layer3_out[10329] <= layer2_out[1628];
     layer3_out[10330] <= ~layer2_out[4548];
     layer3_out[10331] <= layer2_out[3258] ^ layer2_out[3259];
     layer3_out[10332] <= ~(layer2_out[9372] | layer2_out[9373]);
     layer3_out[10333] <= layer2_out[8886] & ~layer2_out[8887];
     layer3_out[10334] <= ~layer2_out[2207];
     layer3_out[10335] <= ~layer2_out[11991];
     layer3_out[10336] <= ~layer2_out[9053];
     layer3_out[10337] <= layer2_out[8089];
     layer3_out[10338] <= layer2_out[10461];
     layer3_out[10339] <= ~layer2_out[1442];
     layer3_out[10340] <= ~layer2_out[9903];
     layer3_out[10341] <= ~(layer2_out[6017] | layer2_out[6018]);
     layer3_out[10342] <= layer2_out[11271];
     layer3_out[10343] <= layer2_out[7871] | layer2_out[7872];
     layer3_out[10344] <= layer2_out[845];
     layer3_out[10345] <= layer2_out[7417] & ~layer2_out[7418];
     layer3_out[10346] <= layer2_out[2538];
     layer3_out[10347] <= ~layer2_out[11755];
     layer3_out[10348] <= layer2_out[4700];
     layer3_out[10349] <= layer2_out[9900] & ~layer2_out[9901];
     layer3_out[10350] <= layer2_out[59];
     layer3_out[10351] <= ~layer2_out[5691];
     layer3_out[10352] <= ~layer2_out[7257];
     layer3_out[10353] <= layer2_out[9794] & layer2_out[9795];
     layer3_out[10354] <= ~layer2_out[3675];
     layer3_out[10355] <= layer2_out[1356];
     layer3_out[10356] <= layer2_out[10174];
     layer3_out[10357] <= layer2_out[9004];
     layer3_out[10358] <= layer2_out[10474];
     layer3_out[10359] <= layer2_out[60];
     layer3_out[10360] <= layer2_out[7032] ^ layer2_out[7033];
     layer3_out[10361] <= ~(layer2_out[6657] & layer2_out[6658]);
     layer3_out[10362] <= ~layer2_out[6124];
     layer3_out[10363] <= ~(layer2_out[2906] | layer2_out[2907]);
     layer3_out[10364] <= layer2_out[478] ^ layer2_out[479];
     layer3_out[10365] <= ~layer2_out[3180] | layer2_out[3179];
     layer3_out[10366] <= layer2_out[784];
     layer3_out[10367] <= layer2_out[744];
     layer3_out[10368] <= layer2_out[2070];
     layer3_out[10369] <= layer2_out[481];
     layer3_out[10370] <= ~layer2_out[9917] | layer2_out[9918];
     layer3_out[10371] <= ~(layer2_out[6826] & layer2_out[6827]);
     layer3_out[10372] <= layer2_out[7724];
     layer3_out[10373] <= ~layer2_out[7775] | layer2_out[7776];
     layer3_out[10374] <= ~layer2_out[2582];
     layer3_out[10375] <= ~layer2_out[7406];
     layer3_out[10376] <= layer2_out[11479] & layer2_out[11480];
     layer3_out[10377] <= ~(layer2_out[8291] & layer2_out[8292]);
     layer3_out[10378] <= ~(layer2_out[10612] ^ layer2_out[10613]);
     layer3_out[10379] <= ~(layer2_out[11466] & layer2_out[11467]);
     layer3_out[10380] <= layer2_out[3258] & ~layer2_out[3257];
     layer3_out[10381] <= layer2_out[5424] & ~layer2_out[5423];
     layer3_out[10382] <= layer2_out[1421] & ~layer2_out[1420];
     layer3_out[10383] <= ~layer2_out[3285];
     layer3_out[10384] <= layer2_out[2623] & ~layer2_out[2624];
     layer3_out[10385] <= ~layer2_out[10117] | layer2_out[10118];
     layer3_out[10386] <= ~layer2_out[6813] | layer2_out[6814];
     layer3_out[10387] <= layer2_out[3445] | layer2_out[3446];
     layer3_out[10388] <= layer2_out[8503] ^ layer2_out[8504];
     layer3_out[10389] <= layer2_out[249];
     layer3_out[10390] <= ~layer2_out[9723] | layer2_out[9724];
     layer3_out[10391] <= ~(layer2_out[6245] | layer2_out[6246]);
     layer3_out[10392] <= layer2_out[9607] & ~layer2_out[9608];
     layer3_out[10393] <= layer2_out[11502] & ~layer2_out[11503];
     layer3_out[10394] <= ~layer2_out[2944] | layer2_out[2943];
     layer3_out[10395] <= layer2_out[13];
     layer3_out[10396] <= ~layer2_out[1394] | layer2_out[1393];
     layer3_out[10397] <= layer2_out[2978] & ~layer2_out[2977];
     layer3_out[10398] <= ~(layer2_out[6096] | layer2_out[6097]);
     layer3_out[10399] <= layer2_out[8290] & ~layer2_out[8291];
     layer3_out[10400] <= ~layer2_out[6825];
     layer3_out[10401] <= ~layer2_out[9628];
     layer3_out[10402] <= ~layer2_out[3923];
     layer3_out[10403] <= layer2_out[4764] & ~layer2_out[4765];
     layer3_out[10404] <= ~(layer2_out[7893] ^ layer2_out[7894]);
     layer3_out[10405] <= ~(layer2_out[3858] | layer2_out[3859]);
     layer3_out[10406] <= layer2_out[4610];
     layer3_out[10407] <= ~layer2_out[9988];
     layer3_out[10408] <= ~layer2_out[6702];
     layer3_out[10409] <= layer2_out[11194];
     layer3_out[10410] <= ~layer2_out[8170];
     layer3_out[10411] <= ~(layer2_out[7858] ^ layer2_out[7859]);
     layer3_out[10412] <= ~(layer2_out[8394] | layer2_out[8395]);
     layer3_out[10413] <= layer2_out[5681] ^ layer2_out[5682];
     layer3_out[10414] <= ~layer2_out[11511];
     layer3_out[10415] <= layer2_out[4478];
     layer3_out[10416] <= ~layer2_out[3492];
     layer3_out[10417] <= ~layer2_out[865];
     layer3_out[10418] <= layer2_out[2851];
     layer3_out[10419] <= ~(layer2_out[8070] | layer2_out[8071]);
     layer3_out[10420] <= layer2_out[1504] & layer2_out[1505];
     layer3_out[10421] <= ~layer2_out[6102];
     layer3_out[10422] <= ~(layer2_out[10023] | layer2_out[10024]);
     layer3_out[10423] <= layer2_out[6515];
     layer3_out[10424] <= layer2_out[1607] & ~layer2_out[1608];
     layer3_out[10425] <= ~layer2_out[967];
     layer3_out[10426] <= layer2_out[2318] & ~layer2_out[2317];
     layer3_out[10427] <= layer2_out[4169];
     layer3_out[10428] <= layer2_out[11840];
     layer3_out[10429] <= ~(layer2_out[2728] | layer2_out[2729]);
     layer3_out[10430] <= ~layer2_out[9117];
     layer3_out[10431] <= layer2_out[6185];
     layer3_out[10432] <= ~layer2_out[3687];
     layer3_out[10433] <= ~layer2_out[6591];
     layer3_out[10434] <= ~(layer2_out[6512] ^ layer2_out[6513]);
     layer3_out[10435] <= ~layer2_out[4889];
     layer3_out[10436] <= layer2_out[1528] & ~layer2_out[1527];
     layer3_out[10437] <= layer2_out[6254] & ~layer2_out[6253];
     layer3_out[10438] <= ~(layer2_out[4363] & layer2_out[4364]);
     layer3_out[10439] <= ~layer2_out[3968];
     layer3_out[10440] <= layer2_out[3437] ^ layer2_out[3438];
     layer3_out[10441] <= ~layer2_out[8839];
     layer3_out[10442] <= layer2_out[934] & layer2_out[935];
     layer3_out[10443] <= layer2_out[10575] & ~layer2_out[10574];
     layer3_out[10444] <= layer2_out[10578] & ~layer2_out[10577];
     layer3_out[10445] <= ~(layer2_out[5417] | layer2_out[5418]);
     layer3_out[10446] <= ~(layer2_out[8858] & layer2_out[8859]);
     layer3_out[10447] <= ~layer2_out[429] | layer2_out[430];
     layer3_out[10448] <= layer2_out[10004] & layer2_out[10005];
     layer3_out[10449] <= layer2_out[1333] ^ layer2_out[1334];
     layer3_out[10450] <= layer2_out[4077] & ~layer2_out[4078];
     layer3_out[10451] <= layer2_out[6289];
     layer3_out[10452] <= ~(layer2_out[11275] ^ layer2_out[11276]);
     layer3_out[10453] <= ~layer2_out[2986];
     layer3_out[10454] <= layer2_out[8028];
     layer3_out[10455] <= ~layer2_out[8898];
     layer3_out[10456] <= layer2_out[6758] & ~layer2_out[6757];
     layer3_out[10457] <= layer2_out[149] & ~layer2_out[148];
     layer3_out[10458] <= ~layer2_out[221];
     layer3_out[10459] <= layer2_out[6485] & layer2_out[6486];
     layer3_out[10460] <= layer2_out[7829];
     layer3_out[10461] <= ~layer2_out[8898];
     layer3_out[10462] <= ~(layer2_out[2666] & layer2_out[2667]);
     layer3_out[10463] <= layer2_out[1287];
     layer3_out[10464] <= ~layer2_out[6881];
     layer3_out[10465] <= layer2_out[11729] & ~layer2_out[11728];
     layer3_out[10466] <= layer2_out[3837];
     layer3_out[10467] <= layer2_out[7323];
     layer3_out[10468] <= ~(layer2_out[8453] | layer2_out[8454]);
     layer3_out[10469] <= ~layer2_out[1605];
     layer3_out[10470] <= layer2_out[3557];
     layer3_out[10471] <= layer2_out[4927];
     layer3_out[10472] <= layer2_out[9633] & ~layer2_out[9634];
     layer3_out[10473] <= ~layer2_out[8240];
     layer3_out[10474] <= layer2_out[6469];
     layer3_out[10475] <= layer2_out[1219];
     layer3_out[10476] <= layer2_out[7273];
     layer3_out[10477] <= layer2_out[10992] & ~layer2_out[10993];
     layer3_out[10478] <= ~(layer2_out[9777] & layer2_out[9778]);
     layer3_out[10479] <= layer2_out[117] & ~layer2_out[118];
     layer3_out[10480] <= ~layer2_out[7229] | layer2_out[7228];
     layer3_out[10481] <= ~(layer2_out[11549] | layer2_out[11550]);
     layer3_out[10482] <= ~layer2_out[6945];
     layer3_out[10483] <= ~layer2_out[412] | layer2_out[413];
     layer3_out[10484] <= layer2_out[8433] & ~layer2_out[8434];
     layer3_out[10485] <= layer2_out[4059];
     layer3_out[10486] <= layer2_out[8736] & ~layer2_out[8735];
     layer3_out[10487] <= layer2_out[1081] & ~layer2_out[1080];
     layer3_out[10488] <= layer2_out[483];
     layer3_out[10489] <= ~layer2_out[9191];
     layer3_out[10490] <= layer2_out[11548] & ~layer2_out[11549];
     layer3_out[10491] <= layer2_out[2369] & layer2_out[2370];
     layer3_out[10492] <= ~layer2_out[9657];
     layer3_out[10493] <= layer2_out[3599];
     layer3_out[10494] <= ~layer2_out[8946] | layer2_out[8945];
     layer3_out[10495] <= layer2_out[4458] & layer2_out[4459];
     layer3_out[10496] <= layer2_out[7932] & layer2_out[7933];
     layer3_out[10497] <= layer2_out[4918] & layer2_out[4919];
     layer3_out[10498] <= layer2_out[7572];
     layer3_out[10499] <= ~layer2_out[7064];
     layer3_out[10500] <= ~layer2_out[4440];
     layer3_out[10501] <= layer2_out[2150] & ~layer2_out[2149];
     layer3_out[10502] <= layer2_out[11782] & layer2_out[11783];
     layer3_out[10503] <= ~(layer2_out[8545] ^ layer2_out[8546]);
     layer3_out[10504] <= ~layer2_out[4388];
     layer3_out[10505] <= ~layer2_out[2236] | layer2_out[2235];
     layer3_out[10506] <= layer2_out[1039];
     layer3_out[10507] <= layer2_out[10799] & layer2_out[10800];
     layer3_out[10508] <= layer2_out[8949] & ~layer2_out[8950];
     layer3_out[10509] <= layer2_out[2535];
     layer3_out[10510] <= ~(layer2_out[194] | layer2_out[195]);
     layer3_out[10511] <= ~layer2_out[11028];
     layer3_out[10512] <= ~layer2_out[3852];
     layer3_out[10513] <= layer2_out[3887] & ~layer2_out[3888];
     layer3_out[10514] <= layer2_out[3527] ^ layer2_out[3528];
     layer3_out[10515] <= ~layer2_out[9454] | layer2_out[9453];
     layer3_out[10516] <= ~layer2_out[5013] | layer2_out[5014];
     layer3_out[10517] <= ~layer2_out[9280];
     layer3_out[10518] <= layer2_out[8872];
     layer3_out[10519] <= layer2_out[1378];
     layer3_out[10520] <= layer2_out[8954] & layer2_out[8955];
     layer3_out[10521] <= ~layer2_out[3158] | layer2_out[3157];
     layer3_out[10522] <= layer2_out[9120];
     layer3_out[10523] <= ~layer2_out[773];
     layer3_out[10524] <= ~layer2_out[4489];
     layer3_out[10525] <= ~(layer2_out[11745] | layer2_out[11746]);
     layer3_out[10526] <= layer2_out[8981];
     layer3_out[10527] <= layer2_out[7841];
     layer3_out[10528] <= layer2_out[7531];
     layer3_out[10529] <= layer2_out[3976];
     layer3_out[10530] <= layer2_out[5349] ^ layer2_out[5350];
     layer3_out[10531] <= layer2_out[11964];
     layer3_out[10532] <= ~(layer2_out[3516] ^ layer2_out[3517]);
     layer3_out[10533] <= ~(layer2_out[981] & layer2_out[982]);
     layer3_out[10534] <= layer2_out[1510];
     layer3_out[10535] <= ~(layer2_out[11647] | layer2_out[11648]);
     layer3_out[10536] <= layer2_out[5836] & ~layer2_out[5835];
     layer3_out[10537] <= layer2_out[2727] & ~layer2_out[2728];
     layer3_out[10538] <= layer2_out[435] ^ layer2_out[436];
     layer3_out[10539] <= ~(layer2_out[5428] ^ layer2_out[5429]);
     layer3_out[10540] <= ~layer2_out[2117];
     layer3_out[10541] <= ~(layer2_out[964] ^ layer2_out[965]);
     layer3_out[10542] <= ~layer2_out[11028];
     layer3_out[10543] <= ~layer2_out[2178] | layer2_out[2177];
     layer3_out[10544] <= layer2_out[6089] | layer2_out[6090];
     layer3_out[10545] <= ~(layer2_out[1416] ^ layer2_out[1417]);
     layer3_out[10546] <= ~(layer2_out[6407] ^ layer2_out[6408]);
     layer3_out[10547] <= layer2_out[3821] ^ layer2_out[3822];
     layer3_out[10548] <= layer2_out[4001] & layer2_out[4002];
     layer3_out[10549] <= layer2_out[9902] & ~layer2_out[9901];
     layer3_out[10550] <= layer2_out[1726] & ~layer2_out[1725];
     layer3_out[10551] <= ~layer2_out[3862];
     layer3_out[10552] <= layer2_out[9081] & ~layer2_out[9082];
     layer3_out[10553] <= ~(layer2_out[3636] | layer2_out[3637]);
     layer3_out[10554] <= layer2_out[6265] & ~layer2_out[6264];
     layer3_out[10555] <= ~(layer2_out[2423] | layer2_out[2424]);
     layer3_out[10556] <= ~(layer2_out[9217] ^ layer2_out[9218]);
     layer3_out[10557] <= ~layer2_out[2440] | layer2_out[2439];
     layer3_out[10558] <= ~layer2_out[7398];
     layer3_out[10559] <= layer2_out[9405];
     layer3_out[10560] <= layer2_out[9352] | layer2_out[9353];
     layer3_out[10561] <= layer2_out[6787];
     layer3_out[10562] <= layer2_out[8425];
     layer3_out[10563] <= ~layer2_out[7408];
     layer3_out[10564] <= layer2_out[4551] & ~layer2_out[4550];
     layer3_out[10565] <= layer2_out[9810] & ~layer2_out[9811];
     layer3_out[10566] <= ~layer2_out[5245];
     layer3_out[10567] <= layer2_out[4563] & ~layer2_out[4564];
     layer3_out[10568] <= layer2_out[5602];
     layer3_out[10569] <= layer2_out[9552];
     layer3_out[10570] <= ~layer2_out[3906];
     layer3_out[10571] <= ~layer2_out[5575];
     layer3_out[10572] <= layer2_out[1977] & layer2_out[1978];
     layer3_out[10573] <= layer2_out[2324];
     layer3_out[10574] <= ~layer2_out[15];
     layer3_out[10575] <= ~(layer2_out[9082] | layer2_out[9083]);
     layer3_out[10576] <= layer2_out[6590] & ~layer2_out[6589];
     layer3_out[10577] <= layer2_out[2960] & ~layer2_out[2961];
     layer3_out[10578] <= layer2_out[10524] & layer2_out[10525];
     layer3_out[10579] <= layer2_out[6335] ^ layer2_out[6336];
     layer3_out[10580] <= layer2_out[7515];
     layer3_out[10581] <= ~(layer2_out[5409] | layer2_out[5410]);
     layer3_out[10582] <= ~layer2_out[11850];
     layer3_out[10583] <= ~layer2_out[2870];
     layer3_out[10584] <= layer2_out[6006] & layer2_out[6007];
     layer3_out[10585] <= layer2_out[3205] & ~layer2_out[3206];
     layer3_out[10586] <= layer2_out[6631] ^ layer2_out[6632];
     layer3_out[10587] <= ~layer2_out[8288];
     layer3_out[10588] <= ~(layer2_out[1201] & layer2_out[1202]);
     layer3_out[10589] <= layer2_out[6439];
     layer3_out[10590] <= ~(layer2_out[2508] | layer2_out[2509]);
     layer3_out[10591] <= layer2_out[228];
     layer3_out[10592] <= layer2_out[8030] & ~layer2_out[8031];
     layer3_out[10593] <= ~(layer2_out[1107] | layer2_out[1108]);
     layer3_out[10594] <= layer2_out[10931];
     layer3_out[10595] <= layer2_out[4594] & ~layer2_out[4593];
     layer3_out[10596] <= ~layer2_out[2199];
     layer3_out[10597] <= layer2_out[11556] & ~layer2_out[11557];
     layer3_out[10598] <= layer2_out[6618];
     layer3_out[10599] <= layer2_out[4180] & layer2_out[4181];
     layer3_out[10600] <= layer2_out[11889];
     layer3_out[10601] <= ~layer2_out[1465];
     layer3_out[10602] <= layer2_out[11359];
     layer3_out[10603] <= layer2_out[4394];
     layer3_out[10604] <= ~layer2_out[2769];
     layer3_out[10605] <= layer2_out[8237] & layer2_out[8238];
     layer3_out[10606] <= layer2_out[8781];
     layer3_out[10607] <= ~layer2_out[342];
     layer3_out[10608] <= layer2_out[4802];
     layer3_out[10609] <= layer2_out[6373] | layer2_out[6374];
     layer3_out[10610] <= layer2_out[9984] ^ layer2_out[9985];
     layer3_out[10611] <= ~layer2_out[6579];
     layer3_out[10612] <= ~layer2_out[5082];
     layer3_out[10613] <= layer2_out[6928] & ~layer2_out[6929];
     layer3_out[10614] <= layer2_out[7281];
     layer3_out[10615] <= layer2_out[2046];
     layer3_out[10616] <= ~(layer2_out[923] | layer2_out[924]);
     layer3_out[10617] <= ~layer2_out[3518];
     layer3_out[10618] <= layer2_out[10753];
     layer3_out[10619] <= ~layer2_out[3161] | layer2_out[3162];
     layer3_out[10620] <= ~layer2_out[7102];
     layer3_out[10621] <= ~layer2_out[10996];
     layer3_out[10622] <= ~(layer2_out[7899] ^ layer2_out[7900]);
     layer3_out[10623] <= layer2_out[10441] & ~layer2_out[10442];
     layer3_out[10624] <= layer2_out[6630];
     layer3_out[10625] <= ~(layer2_out[6880] | layer2_out[6881]);
     layer3_out[10626] <= layer2_out[11536];
     layer3_out[10627] <= layer2_out[7987] ^ layer2_out[7988];
     layer3_out[10628] <= ~layer2_out[3110] | layer2_out[3111];
     layer3_out[10629] <= layer2_out[3089] ^ layer2_out[3090];
     layer3_out[10630] <= ~(layer2_out[3724] ^ layer2_out[3725]);
     layer3_out[10631] <= ~layer2_out[5264];
     layer3_out[10632] <= layer2_out[6597] & ~layer2_out[6598];
     layer3_out[10633] <= layer2_out[5067] ^ layer2_out[5068];
     layer3_out[10634] <= layer2_out[3179] & ~layer2_out[3178];
     layer3_out[10635] <= layer2_out[7913] & ~layer2_out[7912];
     layer3_out[10636] <= layer2_out[8605];
     layer3_out[10637] <= layer2_out[4921] & ~layer2_out[4920];
     layer3_out[10638] <= ~(layer2_out[8221] ^ layer2_out[8222]);
     layer3_out[10639] <= ~layer2_out[4052];
     layer3_out[10640] <= ~layer2_out[9570];
     layer3_out[10641] <= ~layer2_out[6370];
     layer3_out[10642] <= layer2_out[8661] & ~layer2_out[8662];
     layer3_out[10643] <= layer2_out[8566];
     layer3_out[10644] <= layer2_out[11621] ^ layer2_out[11622];
     layer3_out[10645] <= layer2_out[4951] & layer2_out[4952];
     layer3_out[10646] <= ~(layer2_out[3241] & layer2_out[3242]);
     layer3_out[10647] <= layer2_out[7209];
     layer3_out[10648] <= ~layer2_out[4467];
     layer3_out[10649] <= layer2_out[10322] ^ layer2_out[10323];
     layer3_out[10650] <= ~layer2_out[1152];
     layer3_out[10651] <= ~layer2_out[2060] | layer2_out[2061];
     layer3_out[10652] <= layer2_out[3488] | layer2_out[3489];
     layer3_out[10653] <= ~(layer2_out[8618] | layer2_out[8619]);
     layer3_out[10654] <= ~layer2_out[9928];
     layer3_out[10655] <= layer2_out[8835] & ~layer2_out[8836];
     layer3_out[10656] <= layer2_out[3557] & layer2_out[3558];
     layer3_out[10657] <= layer2_out[9182] & ~layer2_out[9181];
     layer3_out[10658] <= layer2_out[7457];
     layer3_out[10659] <= layer2_out[1547] ^ layer2_out[1548];
     layer3_out[10660] <= ~layer2_out[657];
     layer3_out[10661] <= layer2_out[1931];
     layer3_out[10662] <= ~layer2_out[10068];
     layer3_out[10663] <= layer2_out[3283] & ~layer2_out[3282];
     layer3_out[10664] <= layer2_out[1010] ^ layer2_out[1011];
     layer3_out[10665] <= layer2_out[2253] ^ layer2_out[2254];
     layer3_out[10666] <= ~(layer2_out[1616] | layer2_out[1617]);
     layer3_out[10667] <= ~(layer2_out[6384] ^ layer2_out[6385]);
     layer3_out[10668] <= ~layer2_out[7552] | layer2_out[7551];
     layer3_out[10669] <= ~layer2_out[8494];
     layer3_out[10670] <= ~(layer2_out[8446] | layer2_out[8447]);
     layer3_out[10671] <= ~layer2_out[8212];
     layer3_out[10672] <= ~(layer2_out[9017] ^ layer2_out[9018]);
     layer3_out[10673] <= ~layer2_out[11280] | layer2_out[11279];
     layer3_out[10674] <= ~(layer2_out[8268] ^ layer2_out[8269]);
     layer3_out[10675] <= layer2_out[10931];
     layer3_out[10676] <= ~layer2_out[4964];
     layer3_out[10677] <= layer2_out[9764];
     layer3_out[10678] <= ~layer2_out[10100] | layer2_out[10101];
     layer3_out[10679] <= layer2_out[7319];
     layer3_out[10680] <= ~layer2_out[2225] | layer2_out[2224];
     layer3_out[10681] <= ~(layer2_out[3280] | layer2_out[3281]);
     layer3_out[10682] <= ~layer2_out[3901];
     layer3_out[10683] <= ~(layer2_out[44] | layer2_out[45]);
     layer3_out[10684] <= ~(layer2_out[2452] | layer2_out[2453]);
     layer3_out[10685] <= ~(layer2_out[1907] | layer2_out[1908]);
     layer3_out[10686] <= ~layer2_out[2904] | layer2_out[2903];
     layer3_out[10687] <= ~layer2_out[9494];
     layer3_out[10688] <= ~layer2_out[5045] | layer2_out[5046];
     layer3_out[10689] <= ~(layer2_out[486] & layer2_out[487]);
     layer3_out[10690] <= layer2_out[8145];
     layer3_out[10691] <= ~(layer2_out[2521] | layer2_out[2522]);
     layer3_out[10692] <= layer2_out[5479] & layer2_out[5480];
     layer3_out[10693] <= layer2_out[1309] & ~layer2_out[1310];
     layer3_out[10694] <= layer2_out[3773] ^ layer2_out[3774];
     layer3_out[10695] <= layer2_out[2711];
     layer3_out[10696] <= ~layer2_out[5833];
     layer3_out[10697] <= layer2_out[5846] & ~layer2_out[5845];
     layer3_out[10698] <= layer2_out[88];
     layer3_out[10699] <= layer2_out[8401] | layer2_out[8402];
     layer3_out[10700] <= layer2_out[1763] & ~layer2_out[1764];
     layer3_out[10701] <= ~(layer2_out[2663] | layer2_out[2664]);
     layer3_out[10702] <= ~layer2_out[2147];
     layer3_out[10703] <= layer2_out[6521];
     layer3_out[10704] <= layer2_out[2137] & ~layer2_out[2136];
     layer3_out[10705] <= layer2_out[1140];
     layer3_out[10706] <= layer2_out[5567];
     layer3_out[10707] <= ~(layer2_out[10323] | layer2_out[10324]);
     layer3_out[10708] <= ~(layer2_out[5027] & layer2_out[5028]);
     layer3_out[10709] <= layer2_out[1142];
     layer3_out[10710] <= layer2_out[4084] & ~layer2_out[4085];
     layer3_out[10711] <= layer2_out[5251] & ~layer2_out[5250];
     layer3_out[10712] <= ~layer2_out[123];
     layer3_out[10713] <= ~layer2_out[9151] | layer2_out[9152];
     layer3_out[10714] <= layer2_out[2787];
     layer3_out[10715] <= ~layer2_out[9251];
     layer3_out[10716] <= layer2_out[5748];
     layer3_out[10717] <= ~layer2_out[9149];
     layer3_out[10718] <= layer2_out[3151];
     layer3_out[10719] <= layer2_out[1503];
     layer3_out[10720] <= ~layer2_out[10000];
     layer3_out[10721] <= ~layer2_out[4606];
     layer3_out[10722] <= layer2_out[11691] & layer2_out[11692];
     layer3_out[10723] <= layer2_out[9934];
     layer3_out[10724] <= ~(layer2_out[2214] | layer2_out[2215]);
     layer3_out[10725] <= ~layer2_out[7618] | layer2_out[7619];
     layer3_out[10726] <= layer2_out[8310] & layer2_out[8311];
     layer3_out[10727] <= ~layer2_out[3743] | layer2_out[3742];
     layer3_out[10728] <= layer2_out[6804] & ~layer2_out[6803];
     layer3_out[10729] <= ~layer2_out[11019];
     layer3_out[10730] <= layer2_out[7973];
     layer3_out[10731] <= ~(layer2_out[4879] | layer2_out[4880]);
     layer3_out[10732] <= ~layer2_out[2957];
     layer3_out[10733] <= ~(layer2_out[2624] | layer2_out[2625]);
     layer3_out[10734] <= layer2_out[8442];
     layer3_out[10735] <= layer2_out[11305];
     layer3_out[10736] <= ~(layer2_out[8581] | layer2_out[8582]);
     layer3_out[10737] <= layer2_out[4181] ^ layer2_out[4182];
     layer3_out[10738] <= layer2_out[7087] & ~layer2_out[7088];
     layer3_out[10739] <= ~layer2_out[770];
     layer3_out[10740] <= layer2_out[9629] & layer2_out[9630];
     layer3_out[10741] <= ~layer2_out[3984];
     layer3_out[10742] <= ~layer2_out[7483];
     layer3_out[10743] <= ~(layer2_out[3581] & layer2_out[3582]);
     layer3_out[10744] <= ~layer2_out[10946];
     layer3_out[10745] <= ~layer2_out[7753];
     layer3_out[10746] <= ~(layer2_out[4904] | layer2_out[4905]);
     layer3_out[10747] <= layer2_out[7632] & ~layer2_out[7631];
     layer3_out[10748] <= ~layer2_out[7081] | layer2_out[7080];
     layer3_out[10749] <= layer2_out[458] ^ layer2_out[459];
     layer3_out[10750] <= layer2_out[11774];
     layer3_out[10751] <= layer2_out[3855] & layer2_out[3856];
     layer3_out[10752] <= ~layer2_out[8489];
     layer3_out[10753] <= layer2_out[3588] & ~layer2_out[3587];
     layer3_out[10754] <= ~layer2_out[11553];
     layer3_out[10755] <= layer2_out[6772];
     layer3_out[10756] <= layer2_out[6259] & layer2_out[6260];
     layer3_out[10757] <= layer2_out[9013];
     layer3_out[10758] <= layer2_out[1783] & ~layer2_out[1782];
     layer3_out[10759] <= ~layer2_out[10289];
     layer3_out[10760] <= layer2_out[11010] & layer2_out[11011];
     layer3_out[10761] <= layer2_out[517] & ~layer2_out[516];
     layer3_out[10762] <= layer2_out[5181];
     layer3_out[10763] <= ~layer2_out[4883] | layer2_out[4882];
     layer3_out[10764] <= layer2_out[2813] ^ layer2_out[2814];
     layer3_out[10765] <= ~layer2_out[11341];
     layer3_out[10766] <= layer2_out[1391] ^ layer2_out[1392];
     layer3_out[10767] <= ~layer2_out[443];
     layer3_out[10768] <= layer2_out[11623];
     layer3_out[10769] <= layer2_out[7498];
     layer3_out[10770] <= layer2_out[3867];
     layer3_out[10771] <= layer2_out[11844] & ~layer2_out[11843];
     layer3_out[10772] <= ~layer2_out[4431];
     layer3_out[10773] <= layer2_out[5976] & ~layer2_out[5975];
     layer3_out[10774] <= ~layer2_out[7637];
     layer3_out[10775] <= ~layer2_out[3651];
     layer3_out[10776] <= layer2_out[53] & ~layer2_out[54];
     layer3_out[10777] <= layer2_out[2388] & layer2_out[2389];
     layer3_out[10778] <= layer2_out[6319] & ~layer2_out[6320];
     layer3_out[10779] <= ~layer2_out[4254];
     layer3_out[10780] <= layer2_out[6256] & ~layer2_out[6257];
     layer3_out[10781] <= ~layer2_out[2516];
     layer3_out[10782] <= ~(layer2_out[7045] ^ layer2_out[7046]);
     layer3_out[10783] <= ~(layer2_out[7401] | layer2_out[7402]);
     layer3_out[10784] <= ~(layer2_out[3505] | layer2_out[3506]);
     layer3_out[10785] <= layer2_out[1664];
     layer3_out[10786] <= ~layer2_out[9147];
     layer3_out[10787] <= ~(layer2_out[7315] | layer2_out[7316]);
     layer3_out[10788] <= layer2_out[4319];
     layer3_out[10789] <= layer2_out[3732] & ~layer2_out[3733];
     layer3_out[10790] <= ~(layer2_out[256] ^ layer2_out[257]);
     layer3_out[10791] <= ~layer2_out[5699];
     layer3_out[10792] <= layer2_out[7108];
     layer3_out[10793] <= layer2_out[4207];
     layer3_out[10794] <= layer2_out[993] & ~layer2_out[994];
     layer3_out[10795] <= ~(layer2_out[11974] | layer2_out[11975]);
     layer3_out[10796] <= layer2_out[9902] & ~layer2_out[9903];
     layer3_out[10797] <= ~(layer2_out[5107] ^ layer2_out[5108]);
     layer3_out[10798] <= layer2_out[4645] & layer2_out[4646];
     layer3_out[10799] <= layer2_out[5873] & layer2_out[5874];
     layer3_out[10800] <= ~layer2_out[10353] | layer2_out[10352];
     layer3_out[10801] <= ~(layer2_out[4546] ^ layer2_out[4547]);
     layer3_out[10802] <= ~layer2_out[594] | layer2_out[595];
     layer3_out[10803] <= layer2_out[6912] & layer2_out[6913];
     layer3_out[10804] <= ~(layer2_out[9427] | layer2_out[9428]);
     layer3_out[10805] <= layer2_out[2322];
     layer3_out[10806] <= layer2_out[3203] & ~layer2_out[3204];
     layer3_out[10807] <= ~(layer2_out[3480] ^ layer2_out[3481]);
     layer3_out[10808] <= ~layer2_out[388];
     layer3_out[10809] <= layer2_out[6597];
     layer3_out[10810] <= layer2_out[4263] | layer2_out[4264];
     layer3_out[10811] <= ~layer2_out[1123] | layer2_out[1124];
     layer3_out[10812] <= layer2_out[7538];
     layer3_out[10813] <= ~(layer2_out[6901] & layer2_out[6902]);
     layer3_out[10814] <= layer2_out[3695] & layer2_out[3696];
     layer3_out[10815] <= ~layer2_out[2464] | layer2_out[2465];
     layer3_out[10816] <= ~layer2_out[1431];
     layer3_out[10817] <= ~(layer2_out[10202] | layer2_out[10203]);
     layer3_out[10818] <= ~(layer2_out[4745] & layer2_out[4746]);
     layer3_out[10819] <= layer2_out[9926] ^ layer2_out[9927];
     layer3_out[10820] <= layer2_out[6774] ^ layer2_out[6775];
     layer3_out[10821] <= layer2_out[9282] & ~layer2_out[9283];
     layer3_out[10822] <= ~(layer2_out[3805] ^ layer2_out[3806]);
     layer3_out[10823] <= ~(layer2_out[9998] & layer2_out[9999]);
     layer3_out[10824] <= ~layer2_out[1612] | layer2_out[1611];
     layer3_out[10825] <= ~layer2_out[11809] | layer2_out[11810];
     layer3_out[10826] <= ~layer2_out[864];
     layer3_out[10827] <= layer2_out[8510];
     layer3_out[10828] <= ~layer2_out[10744];
     layer3_out[10829] <= layer2_out[9306] & ~layer2_out[9305];
     layer3_out[10830] <= ~layer2_out[1540] | layer2_out[1539];
     layer3_out[10831] <= layer2_out[9618];
     layer3_out[10832] <= layer2_out[6322] & layer2_out[6323];
     layer3_out[10833] <= layer2_out[10367];
     layer3_out[10834] <= layer2_out[6110];
     layer3_out[10835] <= ~(layer2_out[9487] | layer2_out[9488]);
     layer3_out[10836] <= ~layer2_out[10929];
     layer3_out[10837] <= layer2_out[7223] ^ layer2_out[7224];
     layer3_out[10838] <= layer2_out[4426];
     layer3_out[10839] <= layer2_out[7301];
     layer3_out[10840] <= ~layer2_out[6103];
     layer3_out[10841] <= layer2_out[2818] & layer2_out[2819];
     layer3_out[10842] <= ~layer2_out[7678];
     layer3_out[10843] <= ~(layer2_out[7885] | layer2_out[7886]);
     layer3_out[10844] <= ~layer2_out[1550];
     layer3_out[10845] <= layer2_out[699] ^ layer2_out[700];
     layer3_out[10846] <= ~(layer2_out[11919] ^ layer2_out[11920]);
     layer3_out[10847] <= ~layer2_out[10476];
     layer3_out[10848] <= layer2_out[11173];
     layer3_out[10849] <= layer2_out[9618];
     layer3_out[10850] <= ~(layer2_out[11529] & layer2_out[11530]);
     layer3_out[10851] <= ~layer2_out[3996] | layer2_out[3997];
     layer3_out[10852] <= ~(layer2_out[3754] ^ layer2_out[3755]);
     layer3_out[10853] <= ~(layer2_out[8810] | layer2_out[8811]);
     layer3_out[10854] <= ~layer2_out[4496];
     layer3_out[10855] <= layer2_out[4797];
     layer3_out[10856] <= layer2_out[5998] ^ layer2_out[5999];
     layer3_out[10857] <= ~layer2_out[11199];
     layer3_out[10858] <= layer2_out[1171];
     layer3_out[10859] <= ~layer2_out[2709];
     layer3_out[10860] <= layer2_out[8956];
     layer3_out[10861] <= layer2_out[1730];
     layer3_out[10862] <= layer2_out[3577] & ~layer2_out[3578];
     layer3_out[10863] <= ~layer2_out[5002];
     layer3_out[10864] <= layer2_out[3570] | layer2_out[3571];
     layer3_out[10865] <= ~layer2_out[11377];
     layer3_out[10866] <= layer2_out[6859];
     layer3_out[10867] <= layer2_out[10403] ^ layer2_out[10404];
     layer3_out[10868] <= layer2_out[2168];
     layer3_out[10869] <= ~layer2_out[1949] | layer2_out[1950];
     layer3_out[10870] <= layer2_out[6582] ^ layer2_out[6583];
     layer3_out[10871] <= layer2_out[11205] & ~layer2_out[11206];
     layer3_out[10872] <= layer2_out[5312] & ~layer2_out[5313];
     layer3_out[10873] <= layer2_out[10680];
     layer3_out[10874] <= layer2_out[3546];
     layer3_out[10875] <= layer2_out[6606];
     layer3_out[10876] <= layer2_out[3541];
     layer3_out[10877] <= layer2_out[9060] ^ layer2_out[9061];
     layer3_out[10878] <= ~layer2_out[156] | layer2_out[157];
     layer3_out[10879] <= ~(layer2_out[5731] & layer2_out[5732]);
     layer3_out[10880] <= layer2_out[2337];
     layer3_out[10881] <= layer2_out[10775] & layer2_out[10776];
     layer3_out[10882] <= layer2_out[11933];
     layer3_out[10883] <= layer2_out[9749];
     layer3_out[10884] <= layer2_out[5885];
     layer3_out[10885] <= layer2_out[8317] ^ layer2_out[8318];
     layer3_out[10886] <= layer2_out[4552] & layer2_out[4553];
     layer3_out[10887] <= layer2_out[7230];
     layer3_out[10888] <= ~(layer2_out[9670] & layer2_out[9671]);
     layer3_out[10889] <= ~(layer2_out[2951] | layer2_out[2952]);
     layer3_out[10890] <= ~layer2_out[952];
     layer3_out[10891] <= ~layer2_out[4402];
     layer3_out[10892] <= ~(layer2_out[6519] & layer2_out[6520]);
     layer3_out[10893] <= ~layer2_out[2153];
     layer3_out[10894] <= ~layer2_out[10010];
     layer3_out[10895] <= ~layer2_out[10796];
     layer3_out[10896] <= ~(layer2_out[5727] ^ layer2_out[5728]);
     layer3_out[10897] <= layer2_out[5817];
     layer3_out[10898] <= layer2_out[6951] & ~layer2_out[6950];
     layer3_out[10899] <= ~layer2_out[2357];
     layer3_out[10900] <= ~layer2_out[8576];
     layer3_out[10901] <= ~layer2_out[849];
     layer3_out[10902] <= ~layer2_out[479];
     layer3_out[10903] <= layer2_out[3735] ^ layer2_out[3736];
     layer3_out[10904] <= layer2_out[3741] | layer2_out[3742];
     layer3_out[10905] <= ~layer2_out[8882] | layer2_out[8881];
     layer3_out[10906] <= ~layer2_out[8928];
     layer3_out[10907] <= ~layer2_out[1903] | layer2_out[1902];
     layer3_out[10908] <= layer2_out[3602] ^ layer2_out[3603];
     layer3_out[10909] <= layer2_out[6280];
     layer3_out[10910] <= ~layer2_out[10902];
     layer3_out[10911] <= layer2_out[8922];
     layer3_out[10912] <= layer2_out[8131] | layer2_out[8132];
     layer3_out[10913] <= ~(layer2_out[1296] ^ layer2_out[1297]);
     layer3_out[10914] <= ~layer2_out[81] | layer2_out[82];
     layer3_out[10915] <= ~layer2_out[2810];
     layer3_out[10916] <= layer2_out[9625] ^ layer2_out[9626];
     layer3_out[10917] <= layer2_out[6499];
     layer3_out[10918] <= ~layer2_out[8710] | layer2_out[8709];
     layer3_out[10919] <= ~layer2_out[408] | layer2_out[409];
     layer3_out[10920] <= layer2_out[1666];
     layer3_out[10921] <= layer2_out[9443] & ~layer2_out[9444];
     layer3_out[10922] <= layer2_out[9417];
     layer3_out[10923] <= ~layer2_out[4975] | layer2_out[4976];
     layer3_out[10924] <= layer2_out[3260];
     layer3_out[10925] <= layer2_out[1679] ^ layer2_out[1680];
     layer3_out[10926] <= ~layer2_out[747];
     layer3_out[10927] <= layer2_out[3801];
     layer3_out[10928] <= layer2_out[8387] & layer2_out[8388];
     layer3_out[10929] <= ~layer2_out[2852];
     layer3_out[10930] <= layer2_out[4259] ^ layer2_out[4260];
     layer3_out[10931] <= layer2_out[11994] & layer2_out[11995];
     layer3_out[10932] <= layer2_out[1605] & ~layer2_out[1606];
     layer3_out[10933] <= layer2_out[10475];
     layer3_out[10934] <= layer2_out[5166];
     layer3_out[10935] <= ~layer2_out[11288] | layer2_out[11287];
     layer3_out[10936] <= ~layer2_out[6051] | layer2_out[6050];
     layer3_out[10937] <= ~layer2_out[3661] | layer2_out[3662];
     layer3_out[10938] <= ~(layer2_out[11170] ^ layer2_out[11171]);
     layer3_out[10939] <= ~(layer2_out[821] & layer2_out[822]);
     layer3_out[10940] <= layer2_out[11932];
     layer3_out[10941] <= layer2_out[4158];
     layer3_out[10942] <= layer2_out[10417];
     layer3_out[10943] <= ~(layer2_out[4291] & layer2_out[4292]);
     layer3_out[10944] <= ~(layer2_out[3383] & layer2_out[3384]);
     layer3_out[10945] <= ~(layer2_out[3090] ^ layer2_out[3091]);
     layer3_out[10946] <= ~layer2_out[6443];
     layer3_out[10947] <= layer2_out[8116];
     layer3_out[10948] <= ~layer2_out[6352];
     layer3_out[10949] <= layer2_out[8919] & ~layer2_out[8918];
     layer3_out[10950] <= layer2_out[1957];
     layer3_out[10951] <= ~layer2_out[7255] | layer2_out[7256];
     layer3_out[10952] <= ~(layer2_out[10327] ^ layer2_out[10328]);
     layer3_out[10953] <= ~layer2_out[6296];
     layer3_out[10954] <= ~(layer2_out[8873] & layer2_out[8874]);
     layer3_out[10955] <= ~layer2_out[4861];
     layer3_out[10956] <= layer2_out[4484] & ~layer2_out[4483];
     layer3_out[10957] <= ~layer2_out[6605] | layer2_out[6604];
     layer3_out[10958] <= ~layer2_out[2890] | layer2_out[2889];
     layer3_out[10959] <= layer2_out[1805];
     layer3_out[10960] <= ~layer2_out[7337];
     layer3_out[10961] <= layer2_out[4828] ^ layer2_out[4829];
     layer3_out[10962] <= ~(layer2_out[2458] ^ layer2_out[2459]);
     layer3_out[10963] <= layer2_out[8286];
     layer3_out[10964] <= layer2_out[2306];
     layer3_out[10965] <= layer2_out[2451];
     layer3_out[10966] <= ~layer2_out[2404];
     layer3_out[10967] <= ~(layer2_out[9056] ^ layer2_out[9057]);
     layer3_out[10968] <= layer2_out[4441] & layer2_out[4442];
     layer3_out[10969] <= layer2_out[1635] & ~layer2_out[1636];
     layer3_out[10970] <= ~layer2_out[3145];
     layer3_out[10971] <= ~(layer2_out[3761] | layer2_out[3762]);
     layer3_out[10972] <= ~layer2_out[8973];
     layer3_out[10973] <= ~(layer2_out[9937] & layer2_out[9938]);
     layer3_out[10974] <= layer2_out[7832];
     layer3_out[10975] <= layer2_out[2720];
     layer3_out[10976] <= ~layer2_out[2609];
     layer3_out[10977] <= ~(layer2_out[11872] ^ layer2_out[11873]);
     layer3_out[10978] <= ~(layer2_out[7561] & layer2_out[7562]);
     layer3_out[10979] <= layer2_out[8302];
     layer3_out[10980] <= layer2_out[10855];
     layer3_out[10981] <= layer2_out[941];
     layer3_out[10982] <= layer2_out[10563];
     layer3_out[10983] <= ~(layer2_out[5586] | layer2_out[5587]);
     layer3_out[10984] <= ~layer2_out[10166];
     layer3_out[10985] <= ~(layer2_out[8483] | layer2_out[8484]);
     layer3_out[10986] <= layer2_out[4527];
     layer3_out[10987] <= ~(layer2_out[1439] & layer2_out[1440]);
     layer3_out[10988] <= layer2_out[4350] & ~layer2_out[4349];
     layer3_out[10989] <= ~layer2_out[10311];
     layer3_out[10990] <= layer2_out[5987];
     layer3_out[10991] <= layer2_out[9365] | layer2_out[9366];
     layer3_out[10992] <= ~layer2_out[5267];
     layer3_out[10993] <= layer2_out[11829] | layer2_out[11830];
     layer3_out[10994] <= ~(layer2_out[8232] | layer2_out[8233]);
     layer3_out[10995] <= layer2_out[1345] ^ layer2_out[1346];
     layer3_out[10996] <= layer2_out[2998] | layer2_out[2999];
     layer3_out[10997] <= ~layer2_out[2461];
     layer3_out[10998] <= layer2_out[5258] & ~layer2_out[5257];
     layer3_out[10999] <= ~(layer2_out[7253] | layer2_out[7254]);
     layer3_out[11000] <= layer2_out[6430];
     layer3_out[11001] <= layer2_out[1157] & ~layer2_out[1156];
     layer3_out[11002] <= ~layer2_out[5116];
     layer3_out[11003] <= layer2_out[8432] & layer2_out[8433];
     layer3_out[11004] <= layer2_out[4726];
     layer3_out[11005] <= layer2_out[9188] & ~layer2_out[9187];
     layer3_out[11006] <= layer2_out[8931] & ~layer2_out[8930];
     layer3_out[11007] <= layer2_out[2272] ^ layer2_out[2273];
     layer3_out[11008] <= layer2_out[2939];
     layer3_out[11009] <= ~(layer2_out[3551] | layer2_out[3552]);
     layer3_out[11010] <= layer2_out[6357] & ~layer2_out[6356];
     layer3_out[11011] <= ~(layer2_out[10364] ^ layer2_out[10365]);
     layer3_out[11012] <= layer2_out[6019];
     layer3_out[11013] <= ~(layer2_out[1019] ^ layer2_out[1020]);
     layer3_out[11014] <= ~(layer2_out[8159] & layer2_out[8160]);
     layer3_out[11015] <= ~layer2_out[5353];
     layer3_out[11016] <= layer2_out[7167] | layer2_out[7168];
     layer3_out[11017] <= layer2_out[11759] & ~layer2_out[11760];
     layer3_out[11018] <= layer2_out[9195] & ~layer2_out[9194];
     layer3_out[11019] <= ~(layer2_out[4993] & layer2_out[4994]);
     layer3_out[11020] <= ~layer2_out[2263] | layer2_out[2264];
     layer3_out[11021] <= layer2_out[8626] ^ layer2_out[8627];
     layer3_out[11022] <= ~layer2_out[1461] | layer2_out[1462];
     layer3_out[11023] <= ~layer2_out[5869];
     layer3_out[11024] <= layer2_out[287];
     layer3_out[11025] <= ~layer2_out[5325] | layer2_out[5324];
     layer3_out[11026] <= ~layer2_out[9058];
     layer3_out[11027] <= layer2_out[2040];
     layer3_out[11028] <= ~layer2_out[417];
     layer3_out[11029] <= layer2_out[10832] & ~layer2_out[10831];
     layer3_out[11030] <= layer2_out[3764];
     layer3_out[11031] <= layer2_out[8828];
     layer3_out[11032] <= ~layer2_out[1];
     layer3_out[11033] <= layer2_out[11395] ^ layer2_out[11396];
     layer3_out[11034] <= layer2_out[11573] | layer2_out[11574];
     layer3_out[11035] <= layer2_out[3937] & ~layer2_out[3938];
     layer3_out[11036] <= layer2_out[4472];
     layer3_out[11037] <= layer2_out[1694] & ~layer2_out[1693];
     layer3_out[11038] <= layer2_out[9644];
     layer3_out[11039] <= layer2_out[7640] & ~layer2_out[7639];
     layer3_out[11040] <= ~layer2_out[1430] | layer2_out[1429];
     layer3_out[11041] <= layer2_out[8064] & ~layer2_out[8063];
     layer3_out[11042] <= layer2_out[11726] & ~layer2_out[11725];
     layer3_out[11043] <= ~(layer2_out[5907] ^ layer2_out[5908]);
     layer3_out[11044] <= ~layer2_out[8261];
     layer3_out[11045] <= ~layer2_out[7077];
     layer3_out[11046] <= ~layer2_out[2591];
     layer3_out[11047] <= layer2_out[1720];
     layer3_out[11048] <= layer2_out[4539] | layer2_out[4540];
     layer3_out[11049] <= ~(layer2_out[10719] ^ layer2_out[10720]);
     layer3_out[11050] <= layer2_out[2579];
     layer3_out[11051] <= layer2_out[5420] | layer2_out[5421];
     layer3_out[11052] <= ~(layer2_out[11477] ^ layer2_out[11478]);
     layer3_out[11053] <= ~layer2_out[6675] | layer2_out[6674];
     layer3_out[11054] <= ~(layer2_out[9738] | layer2_out[9739]);
     layer3_out[11055] <= layer2_out[10191];
     layer3_out[11056] <= ~layer2_out[3488];
     layer3_out[11057] <= layer2_out[575] | layer2_out[576];
     layer3_out[11058] <= layer2_out[9696] & ~layer2_out[9695];
     layer3_out[11059] <= ~(layer2_out[4934] & layer2_out[4935]);
     layer3_out[11060] <= layer2_out[8944] & ~layer2_out[8945];
     layer3_out[11061] <= ~(layer2_out[5461] | layer2_out[5462]);
     layer3_out[11062] <= layer2_out[2346];
     layer3_out[11063] <= ~(layer2_out[7814] & layer2_out[7815]);
     layer3_out[11064] <= ~layer2_out[295];
     layer3_out[11065] <= layer2_out[395];
     layer3_out[11066] <= layer2_out[10597] ^ layer2_out[10598];
     layer3_out[11067] <= layer2_out[915] ^ layer2_out[916];
     layer3_out[11068] <= ~layer2_out[1267] | layer2_out[1266];
     layer3_out[11069] <= ~layer2_out[2567];
     layer3_out[11070] <= layer2_out[7436] | layer2_out[7437];
     layer3_out[11071] <= ~layer2_out[5966] | layer2_out[5965];
     layer3_out[11072] <= ~layer2_out[6381];
     layer3_out[11073] <= layer2_out[145] & ~layer2_out[146];
     layer3_out[11074] <= layer2_out[3099] ^ layer2_out[3100];
     layer3_out[11075] <= layer2_out[3055];
     layer3_out[11076] <= ~(layer2_out[10197] ^ layer2_out[10198]);
     layer3_out[11077] <= ~layer2_out[1389];
     layer3_out[11078] <= layer2_out[9690] & ~layer2_out[9689];
     layer3_out[11079] <= layer2_out[9681] | layer2_out[9682];
     layer3_out[11080] <= ~layer2_out[9341];
     layer3_out[11081] <= layer2_out[6543];
     layer3_out[11082] <= ~layer2_out[3681];
     layer3_out[11083] <= ~layer2_out[9835] | layer2_out[9836];
     layer3_out[11084] <= ~layer2_out[4349] | layer2_out[4348];
     layer3_out[11085] <= ~layer2_out[5456];
     layer3_out[11086] <= ~layer2_out[6341] | layer2_out[6342];
     layer3_out[11087] <= layer2_out[11629] & ~layer2_out[11630];
     layer3_out[11088] <= ~(layer2_out[10731] & layer2_out[10732]);
     layer3_out[11089] <= ~layer2_out[5861];
     layer3_out[11090] <= layer2_out[11437];
     layer3_out[11091] <= ~(layer2_out[6968] ^ layer2_out[6969]);
     layer3_out[11092] <= ~layer2_out[6586] | layer2_out[6587];
     layer3_out[11093] <= ~layer2_out[3338];
     layer3_out[11094] <= ~layer2_out[10732];
     layer3_out[11095] <= layer2_out[5288];
     layer3_out[11096] <= layer2_out[8660] ^ layer2_out[8661];
     layer3_out[11097] <= layer2_out[1771] & layer2_out[1772];
     layer3_out[11098] <= ~layer2_out[10545];
     layer3_out[11099] <= layer2_out[11213];
     layer3_out[11100] <= ~(layer2_out[1951] & layer2_out[1952]);
     layer3_out[11101] <= ~layer2_out[8469];
     layer3_out[11102] <= layer2_out[11537] | layer2_out[11538];
     layer3_out[11103] <= layer2_out[712];
     layer3_out[11104] <= ~(layer2_out[10030] & layer2_out[10031]);
     layer3_out[11105] <= ~(layer2_out[5413] | layer2_out[5414]);
     layer3_out[11106] <= layer2_out[7746] ^ layer2_out[7747];
     layer3_out[11107] <= layer2_out[4970] | layer2_out[4971];
     layer3_out[11108] <= layer2_out[5852] & ~layer2_out[5853];
     layer3_out[11109] <= layer2_out[183];
     layer3_out[11110] <= ~layer2_out[11682];
     layer3_out[11111] <= layer2_out[9952];
     layer3_out[11112] <= layer2_out[6543] & ~layer2_out[6544];
     layer3_out[11113] <= ~(layer2_out[2487] & layer2_out[2488]);
     layer3_out[11114] <= ~(layer2_out[7153] ^ layer2_out[7154]);
     layer3_out[11115] <= layer2_out[9438] & ~layer2_out[9437];
     layer3_out[11116] <= layer2_out[4023] & layer2_out[4024];
     layer3_out[11117] <= layer2_out[1964];
     layer3_out[11118] <= layer2_out[11763];
     layer3_out[11119] <= ~(layer2_out[6564] ^ layer2_out[6565]);
     layer3_out[11120] <= layer2_out[1028];
     layer3_out[11121] <= layer2_out[2180];
     layer3_out[11122] <= layer2_out[198] & layer2_out[199];
     layer3_out[11123] <= layer2_out[2532] & layer2_out[2533];
     layer3_out[11124] <= ~layer2_out[5399];
     layer3_out[11125] <= layer2_out[9762] ^ layer2_out[9763];
     layer3_out[11126] <= ~layer2_out[633];
     layer3_out[11127] <= layer2_out[10819] | layer2_out[10820];
     layer3_out[11128] <= ~layer2_out[3137] | layer2_out[3136];
     layer3_out[11129] <= ~(layer2_out[7097] | layer2_out[7098]);
     layer3_out[11130] <= layer2_out[6841] & ~layer2_out[6840];
     layer3_out[11131] <= layer2_out[8151];
     layer3_out[11132] <= ~(layer2_out[9592] ^ layer2_out[9593]);
     layer3_out[11133] <= ~(layer2_out[3972] ^ layer2_out[3973]);
     layer3_out[11134] <= layer2_out[4509] | layer2_out[4510];
     layer3_out[11135] <= layer2_out[5296];
     layer3_out[11136] <= layer2_out[870] | layer2_out[871];
     layer3_out[11137] <= layer2_out[9936];
     layer3_out[11138] <= layer2_out[11121];
     layer3_out[11139] <= layer2_out[2362] | layer2_out[2363];
     layer3_out[11140] <= layer2_out[8178];
     layer3_out[11141] <= ~layer2_out[7805];
     layer3_out[11142] <= layer2_out[5392] ^ layer2_out[5393];
     layer3_out[11143] <= ~layer2_out[3646];
     layer3_out[11144] <= ~layer2_out[5792];
     layer3_out[11145] <= layer2_out[5535];
     layer3_out[11146] <= layer2_out[869] | layer2_out[870];
     layer3_out[11147] <= ~(layer2_out[828] ^ layer2_out[829]);
     layer3_out[11148] <= ~layer2_out[7869] | layer2_out[7870];
     layer3_out[11149] <= layer2_out[11729] ^ layer2_out[11730];
     layer3_out[11150] <= ~(layer2_out[513] & layer2_out[514]);
     layer3_out[11151] <= ~layer2_out[2315];
     layer3_out[11152] <= layer2_out[7688] & layer2_out[7689];
     layer3_out[11153] <= ~layer2_out[3578];
     layer3_out[11154] <= layer2_out[858];
     layer3_out[11155] <= layer2_out[10555] & ~layer2_out[10556];
     layer3_out[11156] <= layer2_out[7637] ^ layer2_out[7638];
     layer3_out[11157] <= layer2_out[4756] ^ layer2_out[4757];
     layer3_out[11158] <= layer2_out[11366] ^ layer2_out[11367];
     layer3_out[11159] <= layer2_out[1713] & ~layer2_out[1714];
     layer3_out[11160] <= ~(layer2_out[219] ^ layer2_out[220]);
     layer3_out[11161] <= ~layer2_out[7503];
     layer3_out[11162] <= ~layer2_out[5368];
     layer3_out[11163] <= ~layer2_out[10925];
     layer3_out[11164] <= layer2_out[11082] & ~layer2_out[11083];
     layer3_out[11165] <= layer2_out[1450] ^ layer2_out[1451];
     layer3_out[11166] <= ~layer2_out[4232];
     layer3_out[11167] <= ~(layer2_out[2821] ^ layer2_out[2822]);
     layer3_out[11168] <= ~layer2_out[6117];
     layer3_out[11169] <= ~layer2_out[3869] | layer2_out[3870];
     layer3_out[11170] <= layer2_out[9071];
     layer3_out[11171] <= ~layer2_out[5113];
     layer3_out[11172] <= ~layer2_out[5680] | layer2_out[5679];
     layer3_out[11173] <= layer2_out[1498] & ~layer2_out[1497];
     layer3_out[11174] <= ~(layer2_out[5116] ^ layer2_out[5117]);
     layer3_out[11175] <= layer2_out[11343];
     layer3_out[11176] <= ~(layer2_out[5039] ^ layer2_out[5040]);
     layer3_out[11177] <= layer2_out[11020] & ~layer2_out[11019];
     layer3_out[11178] <= ~(layer2_out[7078] ^ layer2_out[7079]);
     layer3_out[11179] <= layer2_out[7821] | layer2_out[7822];
     layer3_out[11180] <= ~(layer2_out[9329] & layer2_out[9330]);
     layer3_out[11181] <= layer2_out[1161];
     layer3_out[11182] <= ~layer2_out[881] | layer2_out[880];
     layer3_out[11183] <= layer2_out[5733];
     layer3_out[11184] <= layer2_out[8354] & ~layer2_out[8353];
     layer3_out[11185] <= layer2_out[2679];
     layer3_out[11186] <= layer2_out[4739];
     layer3_out[11187] <= layer2_out[6679];
     layer3_out[11188] <= ~layer2_out[2076];
     layer3_out[11189] <= layer2_out[840];
     layer3_out[11190] <= ~layer2_out[1941];
     layer3_out[11191] <= ~(layer2_out[3036] ^ layer2_out[3037]);
     layer3_out[11192] <= ~(layer2_out[8684] ^ layer2_out[8685]);
     layer3_out[11193] <= layer2_out[9246];
     layer3_out[11194] <= ~(layer2_out[3586] ^ layer2_out[3587]);
     layer3_out[11195] <= layer2_out[11461];
     layer3_out[11196] <= layer2_out[11381] & ~layer2_out[11382];
     layer3_out[11197] <= ~layer2_out[8007];
     layer3_out[11198] <= layer2_out[6001];
     layer3_out[11199] <= ~layer2_out[2911];
     layer3_out[11200] <= ~(layer2_out[7767] ^ layer2_out[7768]);
     layer3_out[11201] <= layer2_out[216] & layer2_out[217];
     layer3_out[11202] <= ~layer2_out[7471] | layer2_out[7470];
     layer3_out[11203] <= layer2_out[11989] ^ layer2_out[11990];
     layer3_out[11204] <= layer2_out[1399];
     layer3_out[11205] <= layer2_out[2730];
     layer3_out[11206] <= layer2_out[9469];
     layer3_out[11207] <= ~(layer2_out[7751] | layer2_out[7752]);
     layer3_out[11208] <= layer2_out[1750] | layer2_out[1751];
     layer3_out[11209] <= layer2_out[6228];
     layer3_out[11210] <= layer2_out[10444];
     layer3_out[11211] <= ~layer2_out[4213];
     layer3_out[11212] <= ~layer2_out[7797];
     layer3_out[11213] <= layer2_out[7487] ^ layer2_out[7488];
     layer3_out[11214] <= ~(layer2_out[6244] | layer2_out[6245]);
     layer3_out[11215] <= ~layer2_out[11451];
     layer3_out[11216] <= layer2_out[1666];
     layer3_out[11217] <= ~(layer2_out[5547] ^ layer2_out[5548]);
     layer3_out[11218] <= layer2_out[11181] & ~layer2_out[11182];
     layer3_out[11219] <= layer2_out[10595] | layer2_out[10596];
     layer3_out[11220] <= layer2_out[7237] & layer2_out[7238];
     layer3_out[11221] <= layer2_out[4940];
     layer3_out[11222] <= layer2_out[11757] & layer2_out[11758];
     layer3_out[11223] <= layer2_out[6465] | layer2_out[6466];
     layer3_out[11224] <= layer2_out[6946];
     layer3_out[11225] <= layer2_out[7386] & ~layer2_out[7387];
     layer3_out[11226] <= layer2_out[5068];
     layer3_out[11227] <= ~layer2_out[3081];
     layer3_out[11228] <= ~(layer2_out[6057] & layer2_out[6058]);
     layer3_out[11229] <= ~layer2_out[7074] | layer2_out[7075];
     layer3_out[11230] <= ~(layer2_out[3794] ^ layer2_out[3795]);
     layer3_out[11231] <= ~layer2_out[2574];
     layer3_out[11232] <= ~layer2_out[6172];
     layer3_out[11233] <= ~(layer2_out[1273] & layer2_out[1274]);
     layer3_out[11234] <= layer2_out[11613] ^ layer2_out[11614];
     layer3_out[11235] <= layer2_out[7039] & layer2_out[7040];
     layer3_out[11236] <= ~layer2_out[11644];
     layer3_out[11237] <= ~layer2_out[11273] | layer2_out[11272];
     layer3_out[11238] <= layer2_out[5615];
     layer3_out[11239] <= layer2_out[11312];
     layer3_out[11240] <= ~(layer2_out[5993] & layer2_out[5994]);
     layer3_out[11241] <= ~(layer2_out[9311] ^ layer2_out[9312]);
     layer3_out[11242] <= ~(layer2_out[6195] & layer2_out[6196]);
     layer3_out[11243] <= layer2_out[3524] | layer2_out[3525];
     layer3_out[11244] <= layer2_out[568] & layer2_out[569];
     layer3_out[11245] <= layer2_out[6604];
     layer3_out[11246] <= layer2_out[10373] & ~layer2_out[10372];
     layer3_out[11247] <= ~(layer2_out[10805] ^ layer2_out[10806]);
     layer3_out[11248] <= layer2_out[5147] & ~layer2_out[5146];
     layer3_out[11249] <= layer2_out[1222];
     layer3_out[11250] <= layer2_out[11988];
     layer3_out[11251] <= ~(layer2_out[8445] ^ layer2_out[8446]);
     layer3_out[11252] <= layer2_out[8978];
     layer3_out[11253] <= ~layer2_out[11730] | layer2_out[11731];
     layer3_out[11254] <= ~(layer2_out[6894] ^ layer2_out[6895]);
     layer3_out[11255] <= layer2_out[9745] & layer2_out[9746];
     layer3_out[11256] <= layer2_out[5124] & ~layer2_out[5125];
     layer3_out[11257] <= ~(layer2_out[5633] | layer2_out[5634]);
     layer3_out[11258] <= layer2_out[955] & ~layer2_out[956];
     layer3_out[11259] <= layer2_out[3532] ^ layer2_out[3533];
     layer3_out[11260] <= ~(layer2_out[6733] ^ layer2_out[6734]);
     layer3_out[11261] <= layer2_out[11423];
     layer3_out[11262] <= layer2_out[6954] ^ layer2_out[6955];
     layer3_out[11263] <= ~layer2_out[8248];
     layer3_out[11264] <= ~layer2_out[1476];
     layer3_out[11265] <= ~layer2_out[8696];
     layer3_out[11266] <= ~layer2_out[5669];
     layer3_out[11267] <= layer2_out[2183];
     layer3_out[11268] <= ~(layer2_out[9316] & layer2_out[9317]);
     layer3_out[11269] <= ~layer2_out[5656];
     layer3_out[11270] <= layer2_out[531];
     layer3_out[11271] <= ~(layer2_out[1904] ^ layer2_out[1905]);
     layer3_out[11272] <= ~layer2_out[10613];
     layer3_out[11273] <= layer2_out[7215] ^ layer2_out[7216];
     layer3_out[11274] <= ~layer2_out[9659];
     layer3_out[11275] <= layer2_out[2551];
     layer3_out[11276] <= ~layer2_out[3467] | layer2_out[3468];
     layer3_out[11277] <= ~(layer2_out[1244] | layer2_out[1245]);
     layer3_out[11278] <= ~(layer2_out[1610] | layer2_out[1611]);
     layer3_out[11279] <= layer2_out[4472] & ~layer2_out[4471];
     layer3_out[11280] <= layer2_out[8344] & layer2_out[8345];
     layer3_out[11281] <= ~layer2_out[22];
     layer3_out[11282] <= layer2_out[3197] | layer2_out[3198];
     layer3_out[11283] <= ~layer2_out[9878];
     layer3_out[11284] <= ~layer2_out[72];
     layer3_out[11285] <= layer2_out[11009];
     layer3_out[11286] <= layer2_out[3133];
     layer3_out[11287] <= ~(layer2_out[4572] | layer2_out[4573]);
     layer3_out[11288] <= layer2_out[6299];
     layer3_out[11289] <= ~layer2_out[3644];
     layer3_out[11290] <= layer2_out[7437] ^ layer2_out[7438];
     layer3_out[11291] <= layer2_out[10939];
     layer3_out[11292] <= ~layer2_out[8621];
     layer3_out[11293] <= ~layer2_out[1665] | layer2_out[1664];
     layer3_out[11294] <= layer2_out[8383] ^ layer2_out[8384];
     layer3_out[11295] <= layer2_out[684] ^ layer2_out[685];
     layer3_out[11296] <= ~(layer2_out[9254] ^ layer2_out[9255]);
     layer3_out[11297] <= layer2_out[324];
     layer3_out[11298] <= ~layer2_out[3094];
     layer3_out[11299] <= ~(layer2_out[3631] & layer2_out[3632]);
     layer3_out[11300] <= ~layer2_out[8278] | layer2_out[8277];
     layer3_out[11301] <= ~(layer2_out[7141] | layer2_out[7142]);
     layer3_out[11302] <= ~(layer2_out[3454] | layer2_out[3455]);
     layer3_out[11303] <= ~layer2_out[8201];
     layer3_out[11304] <= layer2_out[7863] | layer2_out[7864];
     layer3_out[11305] <= ~(layer2_out[10830] & layer2_out[10831]);
     layer3_out[11306] <= ~layer2_out[5351];
     layer3_out[11307] <= layer2_out[558] | layer2_out[559];
     layer3_out[11308] <= layer2_out[3236] ^ layer2_out[3237];
     layer3_out[11309] <= layer2_out[1099] & ~layer2_out[1100];
     layer3_out[11310] <= ~layer2_out[3725];
     layer3_out[11311] <= layer2_out[2735] & ~layer2_out[2734];
     layer3_out[11312] <= ~layer2_out[11922];
     layer3_out[11313] <= ~layer2_out[7425];
     layer3_out[11314] <= layer2_out[5917] & layer2_out[5918];
     layer3_out[11315] <= layer2_out[9649] & ~layer2_out[9648];
     layer3_out[11316] <= layer2_out[4299] & ~layer2_out[4300];
     layer3_out[11317] <= ~layer2_out[668] | layer2_out[669];
     layer3_out[11318] <= ~layer2_out[7485];
     layer3_out[11319] <= layer2_out[8920] & layer2_out[8921];
     layer3_out[11320] <= layer2_out[1293] ^ layer2_out[1294];
     layer3_out[11321] <= layer2_out[8194];
     layer3_out[11322] <= ~layer2_out[3193];
     layer3_out[11323] <= ~layer2_out[3311] | layer2_out[3310];
     layer3_out[11324] <= layer2_out[970];
     layer3_out[11325] <= ~(layer2_out[7477] | layer2_out[7478]);
     layer3_out[11326] <= layer2_out[5913] & ~layer2_out[5912];
     layer3_out[11327] <= ~(layer2_out[5069] & layer2_out[5070]);
     layer3_out[11328] <= layer2_out[9891];
     layer3_out[11329] <= ~layer2_out[2779];
     layer3_out[11330] <= layer2_out[9459] | layer2_out[9460];
     layer3_out[11331] <= ~layer2_out[2937];
     layer3_out[11332] <= ~(layer2_out[3175] ^ layer2_out[3176]);
     layer3_out[11333] <= ~(layer2_out[5379] ^ layer2_out[5380]);
     layer3_out[11334] <= ~layer2_out[4275] | layer2_out[4276];
     layer3_out[11335] <= ~layer2_out[9031];
     layer3_out[11336] <= layer2_out[7749] ^ layer2_out[7750];
     layer3_out[11337] <= layer2_out[7111];
     layer3_out[11338] <= ~(layer2_out[3616] | layer2_out[3617]);
     layer3_out[11339] <= layer2_out[80] & ~layer2_out[79];
     layer3_out[11340] <= ~(layer2_out[9677] | layer2_out[9678]);
     layer3_out[11341] <= ~(layer2_out[3975] ^ layer2_out[3976]);
     layer3_out[11342] <= layer2_out[909] & ~layer2_out[910];
     layer3_out[11343] <= ~layer2_out[9640];
     layer3_out[11344] <= layer2_out[8033] & ~layer2_out[8034];
     layer3_out[11345] <= ~(layer2_out[928] | layer2_out[929]);
     layer3_out[11346] <= ~layer2_out[8109];
     layer3_out[11347] <= ~layer2_out[8860];
     layer3_out[11348] <= ~layer2_out[8743] | layer2_out[8742];
     layer3_out[11349] <= ~layer2_out[6569];
     layer3_out[11350] <= layer2_out[5709] ^ layer2_out[5710];
     layer3_out[11351] <= layer2_out[629];
     layer3_out[11352] <= ~(layer2_out[10262] ^ layer2_out[10263]);
     layer3_out[11353] <= ~layer2_out[8124];
     layer3_out[11354] <= ~layer2_out[6684];
     layer3_out[11355] <= layer2_out[8975];
     layer3_out[11356] <= ~layer2_out[11427] | layer2_out[11428];
     layer3_out[11357] <= ~layer2_out[5092];
     layer3_out[11358] <= ~layer2_out[4701] | layer2_out[4700];
     layer3_out[11359] <= ~layer2_out[5433];
     layer3_out[11360] <= ~layer2_out[8349];
     layer3_out[11361] <= ~layer2_out[4209];
     layer3_out[11362] <= ~layer2_out[10071];
     layer3_out[11363] <= ~layer2_out[817] | layer2_out[818];
     layer3_out[11364] <= ~layer2_out[7600];
     layer3_out[11365] <= ~layer2_out[1568] | layer2_out[1569];
     layer3_out[11366] <= layer2_out[8541] & ~layer2_out[8542];
     layer3_out[11367] <= layer2_out[2898];
     layer3_out[11368] <= layer2_out[4324] & layer2_out[4325];
     layer3_out[11369] <= ~layer2_out[7306] | layer2_out[7305];
     layer3_out[11370] <= layer2_out[4626];
     layer3_out[11371] <= ~(layer2_out[11580] & layer2_out[11581]);
     layer3_out[11372] <= ~(layer2_out[8843] & layer2_out[8844]);
     layer3_out[11373] <= layer2_out[5205] | layer2_out[5206];
     layer3_out[11374] <= layer2_out[9127] & ~layer2_out[9126];
     layer3_out[11375] <= layer2_out[4984] ^ layer2_out[4985];
     layer3_out[11376] <= layer2_out[1373] ^ layer2_out[1374];
     layer3_out[11377] <= ~layer2_out[7681];
     layer3_out[11378] <= layer2_out[5571];
     layer3_out[11379] <= layer2_out[8828] & ~layer2_out[8829];
     layer3_out[11380] <= layer2_out[6440];
     layer3_out[11381] <= ~layer2_out[7555] | layer2_out[7556];
     layer3_out[11382] <= ~layer2_out[4953];
     layer3_out[11383] <= ~layer2_out[10359];
     layer3_out[11384] <= layer2_out[8534];
     layer3_out[11385] <= ~(layer2_out[7776] | layer2_out[7777]);
     layer3_out[11386] <= layer2_out[6307];
     layer3_out[11387] <= layer2_out[1283];
     layer3_out[11388] <= ~layer2_out[9299];
     layer3_out[11389] <= ~layer2_out[5919] | layer2_out[5920];
     layer3_out[11390] <= layer2_out[403];
     layer3_out[11391] <= layer2_out[197] & layer2_out[198];
     layer3_out[11392] <= layer2_out[3521];
     layer3_out[11393] <= ~(layer2_out[206] ^ layer2_out[207]);
     layer3_out[11394] <= ~layer2_out[1103];
     layer3_out[11395] <= ~layer2_out[10104];
     layer3_out[11396] <= ~layer2_out[3345] | layer2_out[3346];
     layer3_out[11397] <= ~(layer2_out[3785] & layer2_out[3786]);
     layer3_out[11398] <= layer2_out[10463] & ~layer2_out[10464];
     layer3_out[11399] <= layer2_out[542];
     layer3_out[11400] <= layer2_out[7684] & ~layer2_out[7685];
     layer3_out[11401] <= layer2_out[4264] ^ layer2_out[4265];
     layer3_out[11402] <= layer2_out[9123] ^ layer2_out[9124];
     layer3_out[11403] <= ~layer2_out[7109];
     layer3_out[11404] <= layer2_out[10351];
     layer3_out[11405] <= layer2_out[10499];
     layer3_out[11406] <= ~layer2_out[5762];
     layer3_out[11407] <= ~layer2_out[10256] | layer2_out[10257];
     layer3_out[11408] <= ~layer2_out[2142];
     layer3_out[11409] <= layer2_out[7612] | layer2_out[7613];
     layer3_out[11410] <= layer2_out[10073];
     layer3_out[11411] <= ~(layer2_out[10902] & layer2_out[10903]);
     layer3_out[11412] <= ~(layer2_out[7218] & layer2_out[7219]);
     layer3_out[11413] <= layer2_out[7730];
     layer3_out[11414] <= layer2_out[84] & ~layer2_out[83];
     layer3_out[11415] <= layer2_out[2016];
     layer3_out[11416] <= layer2_out[8465];
     layer3_out[11417] <= layer2_out[2253];
     layer3_out[11418] <= ~layer2_out[3852];
     layer3_out[11419] <= ~layer2_out[2087];
     layer3_out[11420] <= layer2_out[7104];
     layer3_out[11421] <= layer2_out[6160] | layer2_out[6161];
     layer3_out[11422] <= ~layer2_out[7063];
     layer3_out[11423] <= ~layer2_out[502] | layer2_out[503];
     layer3_out[11424] <= layer2_out[7908] ^ layer2_out[7909];
     layer3_out[11425] <= layer2_out[1971];
     layer3_out[11426] <= layer2_out[4892];
     layer3_out[11427] <= ~layer2_out[8962];
     layer3_out[11428] <= ~layer2_out[8822];
     layer3_out[11429] <= layer2_out[2036];
     layer3_out[11430] <= layer2_out[10114];
     layer3_out[11431] <= layer2_out[4944];
     layer3_out[11432] <= ~(layer2_out[8733] & layer2_out[8734]);
     layer3_out[11433] <= layer2_out[5274];
     layer3_out[11434] <= ~layer2_out[3932];
     layer3_out[11435] <= layer2_out[11104] | layer2_out[11105];
     layer3_out[11436] <= ~layer2_out[5344] | layer2_out[5345];
     layer3_out[11437] <= ~layer2_out[4932];
     layer3_out[11438] <= ~(layer2_out[6460] ^ layer2_out[6461]);
     layer3_out[11439] <= layer2_out[7185] ^ layer2_out[7186];
     layer3_out[11440] <= ~layer2_out[9734];
     layer3_out[11441] <= layer2_out[7587];
     layer3_out[11442] <= ~layer2_out[11967] | layer2_out[11968];
     layer3_out[11443] <= layer2_out[1537];
     layer3_out[11444] <= ~layer2_out[30];
     layer3_out[11445] <= ~(layer2_out[9173] & layer2_out[9174]);
     layer3_out[11446] <= layer2_out[6247];
     layer3_out[11447] <= ~(layer2_out[3214] ^ layer2_out[3215]);
     layer3_out[11448] <= layer2_out[10036] ^ layer2_out[10037];
     layer3_out[11449] <= layer2_out[2281] ^ layer2_out[2282];
     layer3_out[11450] <= layer2_out[8058];
     layer3_out[11451] <= layer2_out[8425];
     layer3_out[11452] <= layer2_out[9886];
     layer3_out[11453] <= ~(layer2_out[7811] ^ layer2_out[7812]);
     layer3_out[11454] <= ~layer2_out[5786] | layer2_out[5787];
     layer3_out[11455] <= layer2_out[608] & ~layer2_out[607];
     layer3_out[11456] <= layer2_out[10409] | layer2_out[10410];
     layer3_out[11457] <= layer2_out[9559];
     layer3_out[11458] <= layer2_out[4527];
     layer3_out[11459] <= layer2_out[9499] | layer2_out[9500];
     layer3_out[11460] <= layer2_out[5934];
     layer3_out[11461] <= ~layer2_out[8744];
     layer3_out[11462] <= ~(layer2_out[997] & layer2_out[998]);
     layer3_out[11463] <= ~layer2_out[3018] | layer2_out[3017];
     layer3_out[11464] <= ~layer2_out[2797];
     layer3_out[11465] <= ~(layer2_out[3886] & layer2_out[3887]);
     layer3_out[11466] <= ~(layer2_out[1138] | layer2_out[1139]);
     layer3_out[11467] <= ~layer2_out[10755];
     layer3_out[11468] <= layer2_out[11177] & layer2_out[11178];
     layer3_out[11469] <= layer2_out[8435] & layer2_out[8436];
     layer3_out[11470] <= layer2_out[9109] | layer2_out[9110];
     layer3_out[11471] <= layer2_out[1854] & layer2_out[1855];
     layer3_out[11472] <= layer2_out[5613] & ~layer2_out[5612];
     layer3_out[11473] <= layer2_out[1776];
     layer3_out[11474] <= ~layer2_out[3476] | layer2_out[3475];
     layer3_out[11475] <= layer2_out[11132] | layer2_out[11133];
     layer3_out[11476] <= layer2_out[3359] ^ layer2_out[3360];
     layer3_out[11477] <= ~layer2_out[5281] | layer2_out[5282];
     layer3_out[11478] <= layer2_out[4534] & ~layer2_out[4535];
     layer3_out[11479] <= layer2_out[5914] | layer2_out[5915];
     layer3_out[11480] <= layer2_out[6084];
     layer3_out[11481] <= layer2_out[2260] & layer2_out[2261];
     layer3_out[11482] <= ~layer2_out[7528] | layer2_out[7529];
     layer3_out[11483] <= ~layer2_out[3770];
     layer3_out[11484] <= ~(layer2_out[9846] ^ layer2_out[9847]);
     layer3_out[11485] <= layer2_out[3213] ^ layer2_out[3214];
     layer3_out[11486] <= layer2_out[10037] | layer2_out[10038];
     layer3_out[11487] <= layer2_out[3962] & layer2_out[3963];
     layer3_out[11488] <= layer2_out[482];
     layer3_out[11489] <= layer2_out[6290] | layer2_out[6291];
     layer3_out[11490] <= ~(layer2_out[2562] ^ layer2_out[2563]);
     layer3_out[11491] <= ~layer2_out[727] | layer2_out[728];
     layer3_out[11492] <= layer2_out[8892];
     layer3_out[11493] <= layer2_out[7438];
     layer3_out[11494] <= layer2_out[11161];
     layer3_out[11495] <= layer2_out[2244] ^ layer2_out[2245];
     layer3_out[11496] <= ~layer2_out[11851];
     layer3_out[11497] <= ~layer2_out[3394] | layer2_out[3393];
     layer3_out[11498] <= layer2_out[4131] & ~layer2_out[4132];
     layer3_out[11499] <= ~layer2_out[4415];
     layer3_out[11500] <= layer2_out[4079] & ~layer2_out[4078];
     layer3_out[11501] <= ~layer2_out[2885] | layer2_out[2886];
     layer3_out[11502] <= ~(layer2_out[7856] ^ layer2_out[7857]);
     layer3_out[11503] <= ~layer2_out[4179] | layer2_out[4178];
     layer3_out[11504] <= ~(layer2_out[661] ^ layer2_out[662]);
     layer3_out[11505] <= ~layer2_out[8473];
     layer3_out[11506] <= layer2_out[6736];
     layer3_out[11507] <= layer2_out[5677];
     layer3_out[11508] <= ~layer2_out[7579];
     layer3_out[11509] <= ~layer2_out[4524];
     layer3_out[11510] <= ~(layer2_out[5836] & layer2_out[5837]);
     layer3_out[11511] <= layer2_out[2164];
     layer3_out[11512] <= layer2_out[8987];
     layer3_out[11513] <= ~layer2_out[3871];
     layer3_out[11514] <= layer2_out[11123] | layer2_out[11124];
     layer3_out[11515] <= ~layer2_out[218] | layer2_out[219];
     layer3_out[11516] <= layer2_out[2392] ^ layer2_out[2393];
     layer3_out[11517] <= ~layer2_out[10869];
     layer3_out[11518] <= ~(layer2_out[7197] & layer2_out[7198]);
     layer3_out[11519] <= layer2_out[10115] & ~layer2_out[10116];
     layer3_out[11520] <= ~layer2_out[6087];
     layer3_out[11521] <= ~layer2_out[11654] | layer2_out[11655];
     layer3_out[11522] <= layer2_out[8012] | layer2_out[8013];
     layer3_out[11523] <= layer2_out[494] ^ layer2_out[495];
     layer3_out[11524] <= ~layer2_out[1256] | layer2_out[1255];
     layer3_out[11525] <= layer2_out[7686] & ~layer2_out[7685];
     layer3_out[11526] <= ~layer2_out[8770] | layer2_out[8771];
     layer3_out[11527] <= ~layer2_out[11062];
     layer3_out[11528] <= layer2_out[2071] & ~layer2_out[2070];
     layer3_out[11529] <= ~layer2_out[7672];
     layer3_out[11530] <= ~layer2_out[9526];
     layer3_out[11531] <= layer2_out[6307];
     layer3_out[11532] <= layer2_out[7100] & ~layer2_out[7101];
     layer3_out[11533] <= layer2_out[11998];
     layer3_out[11534] <= ~layer2_out[4601];
     layer3_out[11535] <= ~layer2_out[8853];
     layer3_out[11536] <= ~(layer2_out[9336] ^ layer2_out[9337]);
     layer3_out[11537] <= ~layer2_out[11062];
     layer3_out[11538] <= layer2_out[3139] ^ layer2_out[3140];
     layer3_out[11539] <= layer2_out[10505];
     layer3_out[11540] <= layer2_out[3112];
     layer3_out[11541] <= ~layer2_out[4687] | layer2_out[4688];
     layer3_out[11542] <= layer2_out[6540];
     layer3_out[11543] <= layer2_out[4377] & layer2_out[4378];
     layer3_out[11544] <= layer2_out[4797];
     layer3_out[11545] <= layer2_out[8359] & ~layer2_out[8358];
     layer3_out[11546] <= ~layer2_out[7503];
     layer3_out[11547] <= ~(layer2_out[155] | layer2_out[156]);
     layer3_out[11548] <= layer2_out[3131];
     layer3_out[11549] <= layer2_out[11308];
     layer3_out[11550] <= ~(layer2_out[6270] & layer2_out[6271]);
     layer3_out[11551] <= ~layer2_out[7712];
     layer3_out[11552] <= layer2_out[4586] & layer2_out[4587];
     layer3_out[11553] <= ~(layer2_out[11471] ^ layer2_out[11472]);
     layer3_out[11554] <= ~layer2_out[5729];
     layer3_out[11555] <= layer2_out[7139] & ~layer2_out[7140];
     layer3_out[11556] <= ~(layer2_out[509] ^ layer2_out[510]);
     layer3_out[11557] <= layer2_out[2322];
     layer3_out[11558] <= ~layer2_out[2304] | layer2_out[2305];
     layer3_out[11559] <= layer2_out[8804] & layer2_out[8805];
     layer3_out[11560] <= ~layer2_out[3608];
     layer3_out[11561] <= ~(layer2_out[11760] | layer2_out[11761]);
     layer3_out[11562] <= ~layer2_out[1760] | layer2_out[1759];
     layer3_out[11563] <= ~(layer2_out[5648] | layer2_out[5649]);
     layer3_out[11564] <= ~(layer2_out[4130] ^ layer2_out[4131]);
     layer3_out[11565] <= ~layer2_out[3076];
     layer3_out[11566] <= ~layer2_out[5174];
     layer3_out[11567] <= ~(layer2_out[7560] ^ layer2_out[7561]);
     layer3_out[11568] <= ~(layer2_out[2461] & layer2_out[2462]);
     layer3_out[11569] <= ~(layer2_out[273] ^ layer2_out[274]);
     layer3_out[11570] <= ~(layer2_out[11583] & layer2_out[11584]);
     layer3_out[11571] <= ~layer2_out[3299] | layer2_out[3300];
     layer3_out[11572] <= ~layer2_out[5297];
     layer3_out[11573] <= ~layer2_out[3174];
     layer3_out[11574] <= ~(layer2_out[11227] & layer2_out[11228]);
     layer3_out[11575] <= ~layer2_out[3210];
     layer3_out[11576] <= ~(layer2_out[5452] ^ layer2_out[5453]);
     layer3_out[11577] <= ~layer2_out[378];
     layer3_out[11578] <= ~layer2_out[4224];
     layer3_out[11579] <= layer2_out[6192] | layer2_out[6193];
     layer3_out[11580] <= ~(layer2_out[375] ^ layer2_out[376]);
     layer3_out[11581] <= ~layer2_out[8396];
     layer3_out[11582] <= 1'b1;
     layer3_out[11583] <= layer2_out[11716];
     layer3_out[11584] <= layer2_out[5595] & layer2_out[5596];
     layer3_out[11585] <= layer2_out[6382];
     layer3_out[11586] <= layer2_out[11329];
     layer3_out[11587] <= layer2_out[11224];
     layer3_out[11588] <= ~layer2_out[5906];
     layer3_out[11589] <= layer2_out[1588] | layer2_out[1589];
     layer3_out[11590] <= ~layer2_out[10886];
     layer3_out[11591] <= layer2_out[7696] ^ layer2_out[7697];
     layer3_out[11592] <= ~layer2_out[3135] | layer2_out[3136];
     layer3_out[11593] <= layer2_out[571] & ~layer2_out[572];
     layer3_out[11594] <= layer2_out[4013] | layer2_out[4014];
     layer3_out[11595] <= ~(layer2_out[114] & layer2_out[115]);
     layer3_out[11596] <= ~layer2_out[1856];
     layer3_out[11597] <= ~layer2_out[3702];
     layer3_out[11598] <= layer2_out[4626];
     layer3_out[11599] <= ~layer2_out[9719];
     layer3_out[11600] <= ~layer2_out[8621] | layer2_out[8622];
     layer3_out[11601] <= layer2_out[4273];
     layer3_out[11602] <= layer2_out[8263];
     layer3_out[11603] <= layer2_out[808] | layer2_out[809];
     layer3_out[11604] <= layer2_out[9051] & layer2_out[9052];
     layer3_out[11605] <= layer2_out[3462] | layer2_out[3463];
     layer3_out[11606] <= ~layer2_out[9359] | layer2_out[9358];
     layer3_out[11607] <= ~layer2_out[3616] | layer2_out[3615];
     layer3_out[11608] <= layer2_out[429];
     layer3_out[11609] <= layer2_out[8876];
     layer3_out[11610] <= ~layer2_out[2265];
     layer3_out[11611] <= ~layer2_out[3728];
     layer3_out[11612] <= layer2_out[10790];
     layer3_out[11613] <= layer2_out[6021] & layer2_out[6022];
     layer3_out[11614] <= ~layer2_out[11849] | layer2_out[11848];
     layer3_out[11615] <= layer2_out[5722] ^ layer2_out[5723];
     layer3_out[11616] <= ~layer2_out[5391] | layer2_out[5392];
     layer3_out[11617] <= ~layer2_out[3980] | layer2_out[3979];
     layer3_out[11618] <= layer2_out[8005];
     layer3_out[11619] <= ~layer2_out[10812];
     layer3_out[11620] <= ~layer2_out[2748] | layer2_out[2747];
     layer3_out[11621] <= layer2_out[10084];
     layer3_out[11622] <= layer2_out[5486];
     layer3_out[11623] <= ~(layer2_out[10228] & layer2_out[10229]);
     layer3_out[11624] <= ~layer2_out[6187];
     layer3_out[11625] <= ~layer2_out[6011];
     layer3_out[11626] <= ~(layer2_out[1124] ^ layer2_out[1125]);
     layer3_out[11627] <= ~layer2_out[2172];
     layer3_out[11628] <= ~layer2_out[2327];
     layer3_out[11629] <= ~layer2_out[788];
     layer3_out[11630] <= layer2_out[3128] ^ layer2_out[3129];
     layer3_out[11631] <= layer2_out[9114];
     layer3_out[11632] <= ~layer2_out[4204];
     layer3_out[11633] <= layer2_out[1731] & layer2_out[1732];
     layer3_out[11634] <= layer2_out[94] | layer2_out[95];
     layer3_out[11635] <= ~layer2_out[8235];
     layer3_out[11636] <= layer2_out[3356];
     layer3_out[11637] <= layer2_out[10975] & layer2_out[10976];
     layer3_out[11638] <= ~(layer2_out[10268] & layer2_out[10269]);
     layer3_out[11639] <= layer2_out[7989];
     layer3_out[11640] <= ~layer2_out[10649] | layer2_out[10648];
     layer3_out[11641] <= layer2_out[2785] & layer2_out[2786];
     layer3_out[11642] <= ~layer2_out[4496];
     layer3_out[11643] <= layer2_out[11456] | layer2_out[11457];
     layer3_out[11644] <= layer2_out[326] & layer2_out[327];
     layer3_out[11645] <= ~layer2_out[8173];
     layer3_out[11646] <= layer2_out[9822];
     layer3_out[11647] <= ~layer2_out[4549];
     layer3_out[11648] <= ~(layer2_out[8184] | layer2_out[8185]);
     layer3_out[11649] <= ~layer2_out[1899] | layer2_out[1898];
     layer3_out[11650] <= ~(layer2_out[11973] ^ layer2_out[11974]);
     layer3_out[11651] <= layer2_out[9419];
     layer3_out[11652] <= ~layer2_out[7493];
     layer3_out[11653] <= ~layer2_out[9908];
     layer3_out[11654] <= layer2_out[8916] & ~layer2_out[8915];
     layer3_out[11655] <= layer2_out[1651] & layer2_out[1652];
     layer3_out[11656] <= layer2_out[4030] & ~layer2_out[4029];
     layer3_out[11657] <= layer2_out[6410];
     layer3_out[11658] <= layer2_out[5935];
     layer3_out[11659] <= ~layer2_out[10897];
     layer3_out[11660] <= layer2_out[4509];
     layer3_out[11661] <= layer2_out[8838];
     layer3_out[11662] <= layer2_out[9597] ^ layer2_out[9598];
     layer3_out[11663] <= ~layer2_out[748];
     layer3_out[11664] <= ~layer2_out[7635] | layer2_out[7636];
     layer3_out[11665] <= ~layer2_out[4749] | layer2_out[4748];
     layer3_out[11666] <= layer2_out[10369];
     layer3_out[11667] <= ~layer2_out[187] | layer2_out[188];
     layer3_out[11668] <= layer2_out[3172] & ~layer2_out[3171];
     layer3_out[11669] <= ~layer2_out[8950];
     layer3_out[11670] <= ~layer2_out[1960] | layer2_out[1959];
     layer3_out[11671] <= ~layer2_out[11217];
     layer3_out[11672] <= layer2_out[5652] & layer2_out[5653];
     layer3_out[11673] <= layer2_out[7170];
     layer3_out[11674] <= layer2_out[2439];
     layer3_out[11675] <= layer2_out[7066];
     layer3_out[11676] <= layer2_out[9226];
     layer3_out[11677] <= layer2_out[10623] ^ layer2_out[10624];
     layer3_out[11678] <= layer2_out[5272] & ~layer2_out[5271];
     layer3_out[11679] <= ~(layer2_out[1861] & layer2_out[1862]);
     layer3_out[11680] <= ~(layer2_out[9412] | layer2_out[9413]);
     layer3_out[11681] <= ~layer2_out[5161];
     layer3_out[11682] <= layer2_out[9784] & layer2_out[9785];
     layer3_out[11683] <= ~(layer2_out[2478] ^ layer2_out[2479]);
     layer3_out[11684] <= layer2_out[2856];
     layer3_out[11685] <= ~layer2_out[3238] | layer2_out[3237];
     layer3_out[11686] <= layer2_out[4913] & ~layer2_out[4912];
     layer3_out[11687] <= layer2_out[11125] | layer2_out[11126];
     layer3_out[11688] <= layer2_out[8405];
     layer3_out[11689] <= ~layer2_out[6195];
     layer3_out[11690] <= ~layer2_out[7350];
     layer3_out[11691] <= ~(layer2_out[1563] & layer2_out[1564]);
     layer3_out[11692] <= ~layer2_out[1156];
     layer3_out[11693] <= ~layer2_out[7759];
     layer3_out[11694] <= ~layer2_out[2698];
     layer3_out[11695] <= ~layer2_out[5190] | layer2_out[5189];
     layer3_out[11696] <= layer2_out[6748];
     layer3_out[11697] <= layer2_out[6956];
     layer3_out[11698] <= layer2_out[3536];
     layer3_out[11699] <= ~layer2_out[6646];
     layer3_out[11700] <= ~layer2_out[10942];
     layer3_out[11701] <= ~layer2_out[4827] | layer2_out[4828];
     layer3_out[11702] <= ~layer2_out[3479] | layer2_out[3480];
     layer3_out[11703] <= layer2_out[10954] & layer2_out[10955];
     layer3_out[11704] <= layer2_out[10271] | layer2_out[10272];
     layer3_out[11705] <= ~(layer2_out[9136] ^ layer2_out[9137]);
     layer3_out[11706] <= layer2_out[4119] & ~layer2_out[4120];
     layer3_out[11707] <= layer2_out[2501] | layer2_out[2502];
     layer3_out[11708] <= ~layer2_out[5696];
     layer3_out[11709] <= ~layer2_out[6338];
     layer3_out[11710] <= ~(layer2_out[9286] & layer2_out[9287]);
     layer3_out[11711] <= ~(layer2_out[4010] & layer2_out[4011]);
     layer3_out[11712] <= ~(layer2_out[4775] | layer2_out[4776]);
     layer3_out[11713] <= ~(layer2_out[7697] & layer2_out[7698]);
     layer3_out[11714] <= ~layer2_out[5921] | layer2_out[5922];
     layer3_out[11715] <= layer2_out[287];
     layer3_out[11716] <= layer2_out[8334] ^ layer2_out[8335];
     layer3_out[11717] <= layer2_out[7902] & ~layer2_out[7901];
     layer3_out[11718] <= layer2_out[5661];
     layer3_out[11719] <= ~(layer2_out[9382] ^ layer2_out[9383]);
     layer3_out[11720] <= layer2_out[10169] & ~layer2_out[10168];
     layer3_out[11721] <= ~(layer2_out[707] & layer2_out[708]);
     layer3_out[11722] <= layer2_out[3163];
     layer3_out[11723] <= layer2_out[5247];
     layer3_out[11724] <= layer2_out[5437] ^ layer2_out[5438];
     layer3_out[11725] <= ~layer2_out[2564];
     layer3_out[11726] <= layer2_out[1053];
     layer3_out[11727] <= ~(layer2_out[8852] & layer2_out[8853]);
     layer3_out[11728] <= ~(layer2_out[6709] ^ layer2_out[6710]);
     layer3_out[11729] <= layer2_out[11322] & layer2_out[11323];
     layer3_out[11730] <= ~layer2_out[2462];
     layer3_out[11731] <= layer2_out[5752];
     layer3_out[11732] <= ~layer2_out[5841];
     layer3_out[11733] <= ~(layer2_out[10140] & layer2_out[10141]);
     layer3_out[11734] <= ~layer2_out[10599];
     layer3_out[11735] <= layer2_out[11038];
     layer3_out[11736] <= layer2_out[7073] ^ layer2_out[7074];
     layer3_out[11737] <= ~(layer2_out[9674] | layer2_out[9675]);
     layer3_out[11738] <= ~(layer2_out[11092] | layer2_out[11093]);
     layer3_out[11739] <= layer2_out[8046] | layer2_out[8047];
     layer3_out[11740] <= ~(layer2_out[7581] | layer2_out[7582]);
     layer3_out[11741] <= layer2_out[5407] ^ layer2_out[5408];
     layer3_out[11742] <= ~layer2_out[8620] | layer2_out[8619];
     layer3_out[11743] <= ~(layer2_out[1682] ^ layer2_out[1683]);
     layer3_out[11744] <= ~(layer2_out[1172] | layer2_out[1173]);
     layer3_out[11745] <= layer2_out[1396];
     layer3_out[11746] <= layer2_out[2451];
     layer3_out[11747] <= ~layer2_out[11364] | layer2_out[11363];
     layer3_out[11748] <= layer2_out[347];
     layer3_out[11749] <= ~(layer2_out[5519] & layer2_out[5520]);
     layer3_out[11750] <= ~layer2_out[5896] | layer2_out[5895];
     layer3_out[11751] <= layer2_out[6422] | layer2_out[6423];
     layer3_out[11752] <= layer2_out[4706] & ~layer2_out[4707];
     layer3_out[11753] <= layer2_out[6986];
     layer3_out[11754] <= layer2_out[8766];
     layer3_out[11755] <= layer2_out[7640];
     layer3_out[11756] <= layer2_out[5932] & layer2_out[5933];
     layer3_out[11757] <= ~layer2_out[2030];
     layer3_out[11758] <= ~layer2_out[6836];
     layer3_out[11759] <= layer2_out[8038] & layer2_out[8039];
     layer3_out[11760] <= layer2_out[6314] ^ layer2_out[6315];
     layer3_out[11761] <= ~layer2_out[372];
     layer3_out[11762] <= layer2_out[9315];
     layer3_out[11763] <= layer2_out[1772];
     layer3_out[11764] <= layer2_out[2018] | layer2_out[2019];
     layer3_out[11765] <= layer2_out[7947];
     layer3_out[11766] <= layer2_out[11039];
     layer3_out[11767] <= ~layer2_out[790];
     layer3_out[11768] <= ~layer2_out[3681];
     layer3_out[11769] <= layer2_out[10815];
     layer3_out[11770] <= layer2_out[3986] & layer2_out[3987];
     layer3_out[11771] <= layer2_out[2683];
     layer3_out[11772] <= ~layer2_out[3646];
     layer3_out[11773] <= ~layer2_out[7914] | layer2_out[7915];
     layer3_out[11774] <= ~layer2_out[8120];
     layer3_out[11775] <= ~layer2_out[2788];
     layer3_out[11776] <= ~(layer2_out[9826] & layer2_out[9827]);
     layer3_out[11777] <= ~layer2_out[8954] | layer2_out[8953];
     layer3_out[11778] <= ~(layer2_out[9290] ^ layer2_out[9291]);
     layer3_out[11779] <= layer2_out[8569];
     layer3_out[11780] <= ~layer2_out[10107] | layer2_out[10108];
     layer3_out[11781] <= layer2_out[11915];
     layer3_out[11782] <= layer2_out[10990];
     layer3_out[11783] <= ~layer2_out[11826];
     layer3_out[11784] <= layer2_out[7394] & ~layer2_out[7395];
     layer3_out[11785] <= ~(layer2_out[5857] & layer2_out[5858]);
     layer3_out[11786] <= layer2_out[3506] & ~layer2_out[3507];
     layer3_out[11787] <= layer2_out[9300] & ~layer2_out[9301];
     layer3_out[11788] <= layer2_out[1518] | layer2_out[1519];
     layer3_out[11789] <= ~(layer2_out[2382] ^ layer2_out[2383]);
     layer3_out[11790] <= layer2_out[5828];
     layer3_out[11791] <= layer2_out[6124] ^ layer2_out[6125];
     layer3_out[11792] <= layer2_out[8274] ^ layer2_out[8275];
     layer3_out[11793] <= ~(layer2_out[5565] ^ layer2_out[5566]);
     layer3_out[11794] <= ~(layer2_out[10269] & layer2_out[10270]);
     layer3_out[11795] <= ~layer2_out[11693] | layer2_out[11694];
     layer3_out[11796] <= ~layer2_out[6332] | layer2_out[6331];
     layer3_out[11797] <= layer2_out[6272] & ~layer2_out[6273];
     layer3_out[11798] <= ~layer2_out[9132] | layer2_out[9131];
     layer3_out[11799] <= layer2_out[3326];
     layer3_out[11800] <= ~layer2_out[10658] | layer2_out[10659];
     layer3_out[11801] <= layer2_out[4147];
     layer3_out[11802] <= ~layer2_out[39];
     layer3_out[11803] <= ~layer2_out[4974];
     layer3_out[11804] <= ~layer2_out[11476] | layer2_out[11475];
     layer3_out[11805] <= layer2_out[1906];
     layer3_out[11806] <= ~layer2_out[5827] | layer2_out[5828];
     layer3_out[11807] <= ~layer2_out[8506];
     layer3_out[11808] <= ~(layer2_out[3768] | layer2_out[3769]);
     layer3_out[11809] <= layer2_out[2684] & layer2_out[2685];
     layer3_out[11810] <= layer2_out[5818];
     layer3_out[11811] <= layer2_out[2974];
     layer3_out[11812] <= ~layer2_out[3959];
     layer3_out[11813] <= ~layer2_out[2876];
     layer3_out[11814] <= ~layer2_out[10172];
     layer3_out[11815] <= layer2_out[8354];
     layer3_out[11816] <= ~layer2_out[1254];
     layer3_out[11817] <= layer2_out[10065];
     layer3_out[11818] <= layer2_out[7971];
     layer3_out[11819] <= layer2_out[6401];
     layer3_out[11820] <= layer2_out[6798] & ~layer2_out[6797];
     layer3_out[11821] <= ~layer2_out[1352];
     layer3_out[11822] <= layer2_out[6748];
     layer3_out[11823] <= ~layer2_out[5703];
     layer3_out[11824] <= layer2_out[7596];
     layer3_out[11825] <= ~(layer2_out[9534] ^ layer2_out[9535]);
     layer3_out[11826] <= ~layer2_out[10300];
     layer3_out[11827] <= ~layer2_out[9576] | layer2_out[9575];
     layer3_out[11828] <= layer2_out[8290] & ~layer2_out[8289];
     layer3_out[11829] <= ~layer2_out[9925] | layer2_out[9924];
     layer3_out[11830] <= ~layer2_out[5962];
     layer3_out[11831] <= layer2_out[5597];
     layer3_out[11832] <= ~layer2_out[6201];
     layer3_out[11833] <= layer2_out[7173];
     layer3_out[11834] <= ~(layer2_out[5879] & layer2_out[5880]);
     layer3_out[11835] <= ~layer2_out[11262] | layer2_out[11263];
     layer3_out[11836] <= ~(layer2_out[1640] ^ layer2_out[1641]);
     layer3_out[11837] <= layer2_out[1378] & layer2_out[1379];
     layer3_out[11838] <= layer2_out[2310];
     layer3_out[11839] <= ~(layer2_out[390] | layer2_out[391]);
     layer3_out[11840] <= layer2_out[4737];
     layer3_out[11841] <= layer2_out[4879] & ~layer2_out[4878];
     layer3_out[11842] <= layer2_out[1660];
     layer3_out[11843] <= layer2_out[2997] | layer2_out[2998];
     layer3_out[11844] <= layer2_out[4073];
     layer3_out[11845] <= layer2_out[4241] & ~layer2_out[4242];
     layer3_out[11846] <= ~layer2_out[5074];
     layer3_out[11847] <= layer2_out[521];
     layer3_out[11848] <= ~(layer2_out[9520] & layer2_out[9521]);
     layer3_out[11849] <= layer2_out[909];
     layer3_out[11850] <= layer2_out[11854] & ~layer2_out[11855];
     layer3_out[11851] <= ~layer2_out[4717];
     layer3_out[11852] <= ~(layer2_out[5707] ^ layer2_out[5708]);
     layer3_out[11853] <= layer2_out[11767] & ~layer2_out[11766];
     layer3_out[11854] <= layer2_out[69] | layer2_out[70];
     layer3_out[11855] <= ~layer2_out[9450] | layer2_out[9451];
     layer3_out[11856] <= ~(layer2_out[7810] | layer2_out[7811]);
     layer3_out[11857] <= ~layer2_out[7805];
     layer3_out[11858] <= ~(layer2_out[5057] ^ layer2_out[5058]);
     layer3_out[11859] <= ~layer2_out[7861];
     layer3_out[11860] <= layer2_out[3055];
     layer3_out[11861] <= layer2_out[3698] & ~layer2_out[3699];
     layer3_out[11862] <= layer2_out[6859];
     layer3_out[11863] <= layer2_out[2268];
     layer3_out[11864] <= layer2_out[9652];
     layer3_out[11865] <= ~layer2_out[3596];
     layer3_out[11866] <= ~layer2_out[9384];
     layer3_out[11867] <= layer2_out[7623];
     layer3_out[11868] <= layer2_out[7441];
     layer3_out[11869] <= ~layer2_out[648] | layer2_out[647];
     layer3_out[11870] <= layer2_out[10907] ^ layer2_out[10908];
     layer3_out[11871] <= layer2_out[1589];
     layer3_out[11872] <= ~layer2_out[3923] | layer2_out[3924];
     layer3_out[11873] <= ~layer2_out[8642] | layer2_out[8643];
     layer3_out[11874] <= ~layer2_out[5074];
     layer3_out[11875] <= layer2_out[1634];
     layer3_out[11876] <= layer2_out[2651];
     layer3_out[11877] <= ~layer2_out[10634] | layer2_out[10633];
     layer3_out[11878] <= layer2_out[5992] & ~layer2_out[5993];
     layer3_out[11879] <= ~(layer2_out[3992] ^ layer2_out[3993]);
     layer3_out[11880] <= layer2_out[5170] ^ layer2_out[5171];
     layer3_out[11881] <= ~(layer2_out[5032] & layer2_out[5033]);
     layer3_out[11882] <= layer2_out[11767] & layer2_out[11768];
     layer3_out[11883] <= ~layer2_out[1508] | layer2_out[1507];
     layer3_out[11884] <= layer2_out[398] & ~layer2_out[397];
     layer3_out[11885] <= layer2_out[8344];
     layer3_out[11886] <= ~layer2_out[9464];
     layer3_out[11887] <= ~(layer2_out[9558] ^ layer2_out[9559]);
     layer3_out[11888] <= ~layer2_out[5371] | layer2_out[5372];
     layer3_out[11889] <= ~layer2_out[1425] | layer2_out[1424];
     layer3_out[11890] <= layer2_out[11555] & layer2_out[11556];
     layer3_out[11891] <= layer2_out[5127] ^ layer2_out[5128];
     layer3_out[11892] <= layer2_out[10453] ^ layer2_out[10454];
     layer3_out[11893] <= layer2_out[9595];
     layer3_out[11894] <= ~layer2_out[5419];
     layer3_out[11895] <= ~layer2_out[6744];
     layer3_out[11896] <= ~layer2_out[3728];
     layer3_out[11897] <= ~layer2_out[4581] | layer2_out[4582];
     layer3_out[11898] <= layer2_out[10305] ^ layer2_out[10306];
     layer3_out[11899] <= ~layer2_out[9031];
     layer3_out[11900] <= ~layer2_out[7887];
     layer3_out[11901] <= layer2_out[5219];
     layer3_out[11902] <= layer2_out[6649] & ~layer2_out[6650];
     layer3_out[11903] <= layer2_out[11643] & ~layer2_out[11644];
     layer3_out[11904] <= ~layer2_out[9284];
     layer3_out[11905] <= ~layer2_out[8925];
     layer3_out[11906] <= ~(layer2_out[8597] | layer2_out[8598]);
     layer3_out[11907] <= ~layer2_out[8092];
     layer3_out[11908] <= ~layer2_out[7771];
     layer3_out[11909] <= layer2_out[10239] & layer2_out[10240];
     layer3_out[11910] <= ~layer2_out[5849];
     layer3_out[11911] <= layer2_out[1283];
     layer3_out[11912] <= layer2_out[307];
     layer3_out[11913] <= layer2_out[7149];
     layer3_out[11914] <= ~layer2_out[7086];
     layer3_out[11915] <= ~layer2_out[9830] | layer2_out[9831];
     layer3_out[11916] <= layer2_out[5425] & layer2_out[5426];
     layer3_out[11917] <= ~(layer2_out[4331] ^ layer2_out[4332]);
     layer3_out[11918] <= layer2_out[5089] & ~layer2_out[5090];
     layer3_out[11919] <= ~layer2_out[10494];
     layer3_out[11920] <= ~layer2_out[2831] | layer2_out[2830];
     layer3_out[11921] <= layer2_out[5305];
     layer3_out[11922] <= ~layer2_out[2171];
     layer3_out[11923] <= ~layer2_out[5961];
     layer3_out[11924] <= ~layer2_out[1977];
     layer3_out[11925] <= ~layer2_out[6230];
     layer3_out[11926] <= ~(layer2_out[2626] | layer2_out[2627]);
     layer3_out[11927] <= ~(layer2_out[45] ^ layer2_out[46]);
     layer3_out[11928] <= ~(layer2_out[3344] ^ layer2_out[3345]);
     layer3_out[11929] <= layer2_out[7690];
     layer3_out[11930] <= ~layer2_out[10738] | layer2_out[10739];
     layer3_out[11931] <= ~layer2_out[8634];
     layer3_out[11932] <= layer2_out[3627];
     layer3_out[11933] <= layer2_out[11415];
     layer3_out[11934] <= layer2_out[6876];
     layer3_out[11935] <= layer2_out[517] & layer2_out[518];
     layer3_out[11936] <= layer2_out[7876];
     layer3_out[11937] <= layer2_out[9761] | layer2_out[9762];
     layer3_out[11938] <= layer2_out[3104] | layer2_out[3105];
     layer3_out[11939] <= layer2_out[3185];
     layer3_out[11940] <= layer2_out[6480] ^ layer2_out[6481];
     layer3_out[11941] <= layer2_out[11744];
     layer3_out[11942] <= ~layer2_out[5678] | layer2_out[5677];
     layer3_out[11943] <= ~layer2_out[3457] | layer2_out[3456];
     layer3_out[11944] <= ~layer2_out[6475];
     layer3_out[11945] <= layer2_out[6860] & ~layer2_out[6861];
     layer3_out[11946] <= layer2_out[338] & ~layer2_out[337];
     layer3_out[11947] <= ~layer2_out[10306];
     layer3_out[11948] <= layer2_out[8143];
     layer3_out[11949] <= ~layer2_out[1824] | layer2_out[1823];
     layer3_out[11950] <= ~(layer2_out[2156] & layer2_out[2157]);
     layer3_out[11951] <= ~(layer2_out[10770] & layer2_out[10771]);
     layer3_out[11952] <= ~layer2_out[7630];
     layer3_out[11953] <= ~layer2_out[9939] | layer2_out[9940];
     layer3_out[11954] <= ~(layer2_out[5390] & layer2_out[5391]);
     layer3_out[11955] <= layer2_out[11906] | layer2_out[11907];
     layer3_out[11956] <= ~(layer2_out[10522] & layer2_out[10523]);
     layer3_out[11957] <= layer2_out[190] ^ layer2_out[191];
     layer3_out[11958] <= layer2_out[1942] & ~layer2_out[1941];
     layer3_out[11959] <= layer2_out[1831] | layer2_out[1832];
     layer3_out[11960] <= layer2_out[4818];
     layer3_out[11961] <= layer2_out[10734] & layer2_out[10735];
     layer3_out[11962] <= ~(layer2_out[7898] | layer2_out[7899]);
     layer3_out[11963] <= ~layer2_out[4053] | layer2_out[4054];
     layer3_out[11964] <= ~layer2_out[11897];
     layer3_out[11965] <= ~(layer2_out[6923] ^ layer2_out[6924]);
     layer3_out[11966] <= layer2_out[8919];
     layer3_out[11967] <= layer2_out[8023] & layer2_out[8024];
     layer3_out[11968] <= ~layer2_out[113] | layer2_out[112];
     layer3_out[11969] <= ~layer2_out[7681];
     layer3_out[11970] <= layer2_out[6972] & layer2_out[6973];
     layer3_out[11971] <= ~layer2_out[10912];
     layer3_out[11972] <= layer2_out[6568] ^ layer2_out[6569];
     layer3_out[11973] <= layer2_out[7663] & ~layer2_out[7662];
     layer3_out[11974] <= layer2_out[7056];
     layer3_out[11975] <= ~(layer2_out[2022] ^ layer2_out[2023]);
     layer3_out[11976] <= ~layer2_out[435] | layer2_out[434];
     layer3_out[11977] <= ~layer2_out[1196];
     layer3_out[11978] <= ~layer2_out[1966];
     layer3_out[11979] <= ~layer2_out[5365] | layer2_out[5366];
     layer3_out[11980] <= ~layer2_out[8927] | layer2_out[8926];
     layer3_out[11981] <= layer2_out[7479];
     layer3_out[11982] <= layer2_out[4638];
     layer3_out[11983] <= layer2_out[2009] & layer2_out[2010];
     layer3_out[11984] <= ~(layer2_out[1714] | layer2_out[1715]);
     layer3_out[11985] <= layer2_out[3818];
     layer3_out[11986] <= ~layer2_out[5269];
     layer3_out[11987] <= layer2_out[2534] ^ layer2_out[2535];
     layer3_out[11988] <= ~(layer2_out[9263] & layer2_out[9264]);
     layer3_out[11989] <= ~layer2_out[10937];
     layer3_out[11990] <= layer2_out[11834];
     layer3_out[11991] <= layer2_out[10183];
     layer3_out[11992] <= ~(layer2_out[6818] & layer2_out[6819]);
     layer3_out[11993] <= layer2_out[9110];
     layer3_out[11994] <= ~layer2_out[3064];
     layer3_out[11995] <= layer2_out[8836] | layer2_out[8837];
     layer3_out[11996] <= ~(layer2_out[432] | layer2_out[433]);
     layer3_out[11997] <= ~layer2_out[4538];
     layer3_out[11998] <= ~(layer2_out[9359] & layer2_out[9360]);
     layer3_out[11999] <= layer2_out[7983] | layer2_out[7984];
      last_layer_output <= layer3_out;

      result[0] <= last_layer_output[0] + last_layer_output[1] + last_layer_output[2] + last_layer_output[3] + last_layer_output[4] + last_layer_output[5] + last_layer_output[6] + last_layer_output[7] + last_layer_output[8] + last_layer_output[9] + last_layer_output[10] + last_layer_output[11] + last_layer_output[12] + last_layer_output[13] + last_layer_output[14] + last_layer_output[15] + last_layer_output[16] + last_layer_output[17] + last_layer_output[18] + last_layer_output[19] + last_layer_output[20] + last_layer_output[21] + last_layer_output[22] + last_layer_output[23] + last_layer_output[24] + last_layer_output[25] + last_layer_output[26] + last_layer_output[27] + last_layer_output[28] + last_layer_output[29] + last_layer_output[30] + last_layer_output[31] + last_layer_output[32] + last_layer_output[33] + last_layer_output[34] + last_layer_output[35] + last_layer_output[36] + last_layer_output[37] + last_layer_output[38] + last_layer_output[39] + last_layer_output[40] + last_layer_output[41] + last_layer_output[42] + last_layer_output[43] + last_layer_output[44] + last_layer_output[45] + last_layer_output[46] + last_layer_output[47] + last_layer_output[48] + last_layer_output[49] + last_layer_output[50] + last_layer_output[51] + last_layer_output[52] + last_layer_output[53] + last_layer_output[54] + last_layer_output[55] + last_layer_output[56] + last_layer_output[57] + last_layer_output[58] + last_layer_output[59] + last_layer_output[60] + last_layer_output[61] + last_layer_output[62] + last_layer_output[63] + last_layer_output[64] + last_layer_output[65] + last_layer_output[66] + last_layer_output[67] + last_layer_output[68] + last_layer_output[69] + last_layer_output[70] + last_layer_output[71] + last_layer_output[72] + last_layer_output[73] + last_layer_output[74] + last_layer_output[75] + last_layer_output[76] + last_layer_output[77] + last_layer_output[78] + last_layer_output[79] + last_layer_output[80] + last_layer_output[81] + last_layer_output[82] + last_layer_output[83] + last_layer_output[84] + last_layer_output[85] + last_layer_output[86] + last_layer_output[87] + last_layer_output[88] + last_layer_output[89] + last_layer_output[90] + last_layer_output[91] + last_layer_output[92] + last_layer_output[93] + last_layer_output[94] + last_layer_output[95] + last_layer_output[96] + last_layer_output[97] + last_layer_output[98] + last_layer_output[99] + last_layer_output[100] + last_layer_output[101] + last_layer_output[102] + last_layer_output[103] + last_layer_output[104] + last_layer_output[105] + last_layer_output[106] + last_layer_output[107] + last_layer_output[108] + last_layer_output[109] + last_layer_output[110] + last_layer_output[111] + last_layer_output[112] + last_layer_output[113] + last_layer_output[114] + last_layer_output[115] + last_layer_output[116] + last_layer_output[117] + last_layer_output[118] + last_layer_output[119] + last_layer_output[120] + last_layer_output[121] + last_layer_output[122] + last_layer_output[123] + last_layer_output[124] + last_layer_output[125] + last_layer_output[126] + last_layer_output[127] + last_layer_output[128] + last_layer_output[129] + last_layer_output[130] + last_layer_output[131] + last_layer_output[132] + last_layer_output[133] + last_layer_output[134] + last_layer_output[135] + last_layer_output[136] + last_layer_output[137] + last_layer_output[138] + last_layer_output[139] + last_layer_output[140] + last_layer_output[141] + last_layer_output[142] + last_layer_output[143] + last_layer_output[144] + last_layer_output[145] + last_layer_output[146] + last_layer_output[147] + last_layer_output[148] + last_layer_output[149] + last_layer_output[150] + last_layer_output[151] + last_layer_output[152] + last_layer_output[153] + last_layer_output[154] + last_layer_output[155] + last_layer_output[156] + last_layer_output[157] + last_layer_output[158] + last_layer_output[159] + last_layer_output[160] + last_layer_output[161] + last_layer_output[162] + last_layer_output[163] + last_layer_output[164] + last_layer_output[165] + last_layer_output[166] + last_layer_output[167] + last_layer_output[168] + last_layer_output[169] + last_layer_output[170] + last_layer_output[171] + last_layer_output[172] + last_layer_output[173] + last_layer_output[174] + last_layer_output[175] + last_layer_output[176] + last_layer_output[177] + last_layer_output[178] + last_layer_output[179] + last_layer_output[180] + last_layer_output[181] + last_layer_output[182] + last_layer_output[183] + last_layer_output[184] + last_layer_output[185] + last_layer_output[186] + last_layer_output[187] + last_layer_output[188] + last_layer_output[189] + last_layer_output[190] + last_layer_output[191] + last_layer_output[192] + last_layer_output[193] + last_layer_output[194] + last_layer_output[195] + last_layer_output[196] + last_layer_output[197] + last_layer_output[198] + last_layer_output[199] + last_layer_output[200] + last_layer_output[201] + last_layer_output[202] + last_layer_output[203] + last_layer_output[204] + last_layer_output[205] + last_layer_output[206] + last_layer_output[207] + last_layer_output[208] + last_layer_output[209] + last_layer_output[210] + last_layer_output[211] + last_layer_output[212] + last_layer_output[213] + last_layer_output[214] + last_layer_output[215] + last_layer_output[216] + last_layer_output[217] + last_layer_output[218] + last_layer_output[219] + last_layer_output[220] + last_layer_output[221] + last_layer_output[222] + last_layer_output[223] + last_layer_output[224] + last_layer_output[225] + last_layer_output[226] + last_layer_output[227] + last_layer_output[228] + last_layer_output[229] + last_layer_output[230] + last_layer_output[231] + last_layer_output[232] + last_layer_output[233] + last_layer_output[234] + last_layer_output[235] + last_layer_output[236] + last_layer_output[237] + last_layer_output[238] + last_layer_output[239] + last_layer_output[240] + last_layer_output[241] + last_layer_output[242] + last_layer_output[243] + last_layer_output[244] + last_layer_output[245] + last_layer_output[246] + last_layer_output[247] + last_layer_output[248] + last_layer_output[249] + last_layer_output[250] + last_layer_output[251] + last_layer_output[252] + last_layer_output[253] + last_layer_output[254] + last_layer_output[255] + last_layer_output[256] + last_layer_output[257] + last_layer_output[258] + last_layer_output[259] + last_layer_output[260] + last_layer_output[261] + last_layer_output[262] + last_layer_output[263] + last_layer_output[264] + last_layer_output[265] + last_layer_output[266] + last_layer_output[267] + last_layer_output[268] + last_layer_output[269] + last_layer_output[270] + last_layer_output[271] + last_layer_output[272] + last_layer_output[273] + last_layer_output[274] + last_layer_output[275] + last_layer_output[276] + last_layer_output[277] + last_layer_output[278] + last_layer_output[279] + last_layer_output[280] + last_layer_output[281] + last_layer_output[282] + last_layer_output[283] + last_layer_output[284] + last_layer_output[285] + last_layer_output[286] + last_layer_output[287] + last_layer_output[288] + last_layer_output[289] + last_layer_output[290] + last_layer_output[291] + last_layer_output[292] + last_layer_output[293] + last_layer_output[294] + last_layer_output[295] + last_layer_output[296] + last_layer_output[297] + last_layer_output[298] + last_layer_output[299] + last_layer_output[300] + last_layer_output[301] + last_layer_output[302] + last_layer_output[303] + last_layer_output[304] + last_layer_output[305] + last_layer_output[306] + last_layer_output[307] + last_layer_output[308] + last_layer_output[309] + last_layer_output[310] + last_layer_output[311] + last_layer_output[312] + last_layer_output[313] + last_layer_output[314] + last_layer_output[315] + last_layer_output[316] + last_layer_output[317] + last_layer_output[318] + last_layer_output[319] + last_layer_output[320] + last_layer_output[321] + last_layer_output[322] + last_layer_output[323] + last_layer_output[324] + last_layer_output[325] + last_layer_output[326] + last_layer_output[327] + last_layer_output[328] + last_layer_output[329] + last_layer_output[330] + last_layer_output[331] + last_layer_output[332] + last_layer_output[333] + last_layer_output[334] + last_layer_output[335] + last_layer_output[336] + last_layer_output[337] + last_layer_output[338] + last_layer_output[339] + last_layer_output[340] + last_layer_output[341] + last_layer_output[342] + last_layer_output[343] + last_layer_output[344] + last_layer_output[345] + last_layer_output[346] + last_layer_output[347] + last_layer_output[348] + last_layer_output[349] + last_layer_output[350] + last_layer_output[351] + last_layer_output[352] + last_layer_output[353] + last_layer_output[354] + last_layer_output[355] + last_layer_output[356] + last_layer_output[357] + last_layer_output[358] + last_layer_output[359] + last_layer_output[360] + last_layer_output[361] + last_layer_output[362] + last_layer_output[363] + last_layer_output[364] + last_layer_output[365] + last_layer_output[366] + last_layer_output[367] + last_layer_output[368] + last_layer_output[369] + last_layer_output[370] + last_layer_output[371] + last_layer_output[372] + last_layer_output[373] + last_layer_output[374] + last_layer_output[375] + last_layer_output[376] + last_layer_output[377] + last_layer_output[378] + last_layer_output[379] + last_layer_output[380] + last_layer_output[381] + last_layer_output[382] + last_layer_output[383] + last_layer_output[384] + last_layer_output[385] + last_layer_output[386] + last_layer_output[387] + last_layer_output[388] + last_layer_output[389] + last_layer_output[390] + last_layer_output[391] + last_layer_output[392] + last_layer_output[393] + last_layer_output[394] + last_layer_output[395] + last_layer_output[396] + last_layer_output[397] + last_layer_output[398] + last_layer_output[399] + last_layer_output[400] + last_layer_output[401] + last_layer_output[402] + last_layer_output[403] + last_layer_output[404] + last_layer_output[405] + last_layer_output[406] + last_layer_output[407] + last_layer_output[408] + last_layer_output[409] + last_layer_output[410] + last_layer_output[411] + last_layer_output[412] + last_layer_output[413] + last_layer_output[414] + last_layer_output[415] + last_layer_output[416] + last_layer_output[417] + last_layer_output[418] + last_layer_output[419] + last_layer_output[420] + last_layer_output[421] + last_layer_output[422] + last_layer_output[423] + last_layer_output[424] + last_layer_output[425] + last_layer_output[426] + last_layer_output[427] + last_layer_output[428] + last_layer_output[429] + last_layer_output[430] + last_layer_output[431] + last_layer_output[432] + last_layer_output[433] + last_layer_output[434] + last_layer_output[435] + last_layer_output[436] + last_layer_output[437] + last_layer_output[438] + last_layer_output[439] + last_layer_output[440] + last_layer_output[441] + last_layer_output[442] + last_layer_output[443] + last_layer_output[444] + last_layer_output[445] + last_layer_output[446] + last_layer_output[447] + last_layer_output[448] + last_layer_output[449] + last_layer_output[450] + last_layer_output[451] + last_layer_output[452] + last_layer_output[453] + last_layer_output[454] + last_layer_output[455] + last_layer_output[456] + last_layer_output[457] + last_layer_output[458] + last_layer_output[459] + last_layer_output[460] + last_layer_output[461] + last_layer_output[462] + last_layer_output[463] + last_layer_output[464] + last_layer_output[465] + last_layer_output[466] + last_layer_output[467] + last_layer_output[468] + last_layer_output[469] + last_layer_output[470] + last_layer_output[471] + last_layer_output[472] + last_layer_output[473] + last_layer_output[474] + last_layer_output[475] + last_layer_output[476] + last_layer_output[477] + last_layer_output[478] + last_layer_output[479] + last_layer_output[480] + last_layer_output[481] + last_layer_output[482] + last_layer_output[483] + last_layer_output[484] + last_layer_output[485] + last_layer_output[486] + last_layer_output[487] + last_layer_output[488] + last_layer_output[489] + last_layer_output[490] + last_layer_output[491] + last_layer_output[492] + last_layer_output[493] + last_layer_output[494] + last_layer_output[495] + last_layer_output[496] + last_layer_output[497] + last_layer_output[498] + last_layer_output[499] + last_layer_output[500] + last_layer_output[501] + last_layer_output[502] + last_layer_output[503] + last_layer_output[504] + last_layer_output[505] + last_layer_output[506] + last_layer_output[507] + last_layer_output[508] + last_layer_output[509] + last_layer_output[510] + last_layer_output[511] + last_layer_output[512] + last_layer_output[513] + last_layer_output[514] + last_layer_output[515] + last_layer_output[516] + last_layer_output[517] + last_layer_output[518] + last_layer_output[519] + last_layer_output[520] + last_layer_output[521] + last_layer_output[522] + last_layer_output[523] + last_layer_output[524] + last_layer_output[525] + last_layer_output[526] + last_layer_output[527] + last_layer_output[528] + last_layer_output[529] + last_layer_output[530] + last_layer_output[531] + last_layer_output[532] + last_layer_output[533] + last_layer_output[534] + last_layer_output[535] + last_layer_output[536] + last_layer_output[537] + last_layer_output[538] + last_layer_output[539] + last_layer_output[540] + last_layer_output[541] + last_layer_output[542] + last_layer_output[543] + last_layer_output[544] + last_layer_output[545] + last_layer_output[546] + last_layer_output[547] + last_layer_output[548] + last_layer_output[549] + last_layer_output[550] + last_layer_output[551] + last_layer_output[552] + last_layer_output[553] + last_layer_output[554] + last_layer_output[555] + last_layer_output[556] + last_layer_output[557] + last_layer_output[558] + last_layer_output[559] + last_layer_output[560] + last_layer_output[561] + last_layer_output[562] + last_layer_output[563] + last_layer_output[564] + last_layer_output[565] + last_layer_output[566] + last_layer_output[567] + last_layer_output[568] + last_layer_output[569] + last_layer_output[570] + last_layer_output[571] + last_layer_output[572] + last_layer_output[573] + last_layer_output[574] + last_layer_output[575] + last_layer_output[576] + last_layer_output[577] + last_layer_output[578] + last_layer_output[579] + last_layer_output[580] + last_layer_output[581] + last_layer_output[582] + last_layer_output[583] + last_layer_output[584] + last_layer_output[585] + last_layer_output[586] + last_layer_output[587] + last_layer_output[588] + last_layer_output[589] + last_layer_output[590] + last_layer_output[591] + last_layer_output[592] + last_layer_output[593] + last_layer_output[594] + last_layer_output[595] + last_layer_output[596] + last_layer_output[597] + last_layer_output[598] + last_layer_output[599] + last_layer_output[600] + last_layer_output[601] + last_layer_output[602] + last_layer_output[603] + last_layer_output[604] + last_layer_output[605] + last_layer_output[606] + last_layer_output[607] + last_layer_output[608] + last_layer_output[609] + last_layer_output[610] + last_layer_output[611] + last_layer_output[612] + last_layer_output[613] + last_layer_output[614] + last_layer_output[615] + last_layer_output[616] + last_layer_output[617] + last_layer_output[618] + last_layer_output[619] + last_layer_output[620] + last_layer_output[621] + last_layer_output[622] + last_layer_output[623] + last_layer_output[624] + last_layer_output[625] + last_layer_output[626] + last_layer_output[627] + last_layer_output[628] + last_layer_output[629] + last_layer_output[630] + last_layer_output[631] + last_layer_output[632] + last_layer_output[633] + last_layer_output[634] + last_layer_output[635] + last_layer_output[636] + last_layer_output[637] + last_layer_output[638] + last_layer_output[639] + last_layer_output[640] + last_layer_output[641] + last_layer_output[642] + last_layer_output[643] + last_layer_output[644] + last_layer_output[645] + last_layer_output[646] + last_layer_output[647] + last_layer_output[648] + last_layer_output[649] + last_layer_output[650] + last_layer_output[651] + last_layer_output[652] + last_layer_output[653] + last_layer_output[654] + last_layer_output[655] + last_layer_output[656] + last_layer_output[657] + last_layer_output[658] + last_layer_output[659] + last_layer_output[660] + last_layer_output[661] + last_layer_output[662] + last_layer_output[663] + last_layer_output[664] + last_layer_output[665] + last_layer_output[666] + last_layer_output[667] + last_layer_output[668] + last_layer_output[669] + last_layer_output[670] + last_layer_output[671] + last_layer_output[672] + last_layer_output[673] + last_layer_output[674] + last_layer_output[675] + last_layer_output[676] + last_layer_output[677] + last_layer_output[678] + last_layer_output[679] + last_layer_output[680] + last_layer_output[681] + last_layer_output[682] + last_layer_output[683] + last_layer_output[684] + last_layer_output[685] + last_layer_output[686] + last_layer_output[687] + last_layer_output[688] + last_layer_output[689] + last_layer_output[690] + last_layer_output[691] + last_layer_output[692] + last_layer_output[693] + last_layer_output[694] + last_layer_output[695] + last_layer_output[696] + last_layer_output[697] + last_layer_output[698] + last_layer_output[699] + last_layer_output[700] + last_layer_output[701] + last_layer_output[702] + last_layer_output[703] + last_layer_output[704] + last_layer_output[705] + last_layer_output[706] + last_layer_output[707] + last_layer_output[708] + last_layer_output[709] + last_layer_output[710] + last_layer_output[711] + last_layer_output[712] + last_layer_output[713] + last_layer_output[714] + last_layer_output[715] + last_layer_output[716] + last_layer_output[717] + last_layer_output[718] + last_layer_output[719] + last_layer_output[720] + last_layer_output[721] + last_layer_output[722] + last_layer_output[723] + last_layer_output[724] + last_layer_output[725] + last_layer_output[726] + last_layer_output[727] + last_layer_output[728] + last_layer_output[729] + last_layer_output[730] + last_layer_output[731] + last_layer_output[732] + last_layer_output[733] + last_layer_output[734] + last_layer_output[735] + last_layer_output[736] + last_layer_output[737] + last_layer_output[738] + last_layer_output[739] + last_layer_output[740] + last_layer_output[741] + last_layer_output[742] + last_layer_output[743] + last_layer_output[744] + last_layer_output[745] + last_layer_output[746] + last_layer_output[747] + last_layer_output[748] + last_layer_output[749] + last_layer_output[750] + last_layer_output[751] + last_layer_output[752] + last_layer_output[753] + last_layer_output[754] + last_layer_output[755] + last_layer_output[756] + last_layer_output[757] + last_layer_output[758] + last_layer_output[759] + last_layer_output[760] + last_layer_output[761] + last_layer_output[762] + last_layer_output[763] + last_layer_output[764] + last_layer_output[765] + last_layer_output[766] + last_layer_output[767] + last_layer_output[768] + last_layer_output[769] + last_layer_output[770] + last_layer_output[771] + last_layer_output[772] + last_layer_output[773] + last_layer_output[774] + last_layer_output[775] + last_layer_output[776] + last_layer_output[777] + last_layer_output[778] + last_layer_output[779] + last_layer_output[780] + last_layer_output[781] + last_layer_output[782] + last_layer_output[783] + last_layer_output[784] + last_layer_output[785] + last_layer_output[786] + last_layer_output[787] + last_layer_output[788] + last_layer_output[789] + last_layer_output[790] + last_layer_output[791] + last_layer_output[792] + last_layer_output[793] + last_layer_output[794] + last_layer_output[795] + last_layer_output[796] + last_layer_output[797] + last_layer_output[798] + last_layer_output[799] + last_layer_output[800] + last_layer_output[801] + last_layer_output[802] + last_layer_output[803] + last_layer_output[804] + last_layer_output[805] + last_layer_output[806] + last_layer_output[807] + last_layer_output[808] + last_layer_output[809] + last_layer_output[810] + last_layer_output[811] + last_layer_output[812] + last_layer_output[813] + last_layer_output[814] + last_layer_output[815] + last_layer_output[816] + last_layer_output[817] + last_layer_output[818] + last_layer_output[819] + last_layer_output[820] + last_layer_output[821] + last_layer_output[822] + last_layer_output[823] + last_layer_output[824] + last_layer_output[825] + last_layer_output[826] + last_layer_output[827] + last_layer_output[828] + last_layer_output[829] + last_layer_output[830] + last_layer_output[831] + last_layer_output[832] + last_layer_output[833] + last_layer_output[834] + last_layer_output[835] + last_layer_output[836] + last_layer_output[837] + last_layer_output[838] + last_layer_output[839] + last_layer_output[840] + last_layer_output[841] + last_layer_output[842] + last_layer_output[843] + last_layer_output[844] + last_layer_output[845] + last_layer_output[846] + last_layer_output[847] + last_layer_output[848] + last_layer_output[849] + last_layer_output[850] + last_layer_output[851] + last_layer_output[852] + last_layer_output[853] + last_layer_output[854] + last_layer_output[855] + last_layer_output[856] + last_layer_output[857] + last_layer_output[858] + last_layer_output[859] + last_layer_output[860] + last_layer_output[861] + last_layer_output[862] + last_layer_output[863] + last_layer_output[864] + last_layer_output[865] + last_layer_output[866] + last_layer_output[867] + last_layer_output[868] + last_layer_output[869] + last_layer_output[870] + last_layer_output[871] + last_layer_output[872] + last_layer_output[873] + last_layer_output[874] + last_layer_output[875] + last_layer_output[876] + last_layer_output[877] + last_layer_output[878] + last_layer_output[879] + last_layer_output[880] + last_layer_output[881] + last_layer_output[882] + last_layer_output[883] + last_layer_output[884] + last_layer_output[885] + last_layer_output[886] + last_layer_output[887] + last_layer_output[888] + last_layer_output[889] + last_layer_output[890] + last_layer_output[891] + last_layer_output[892] + last_layer_output[893] + last_layer_output[894] + last_layer_output[895] + last_layer_output[896] + last_layer_output[897] + last_layer_output[898] + last_layer_output[899] + last_layer_output[900] + last_layer_output[901] + last_layer_output[902] + last_layer_output[903] + last_layer_output[904] + last_layer_output[905] + last_layer_output[906] + last_layer_output[907] + last_layer_output[908] + last_layer_output[909] + last_layer_output[910] + last_layer_output[911] + last_layer_output[912] + last_layer_output[913] + last_layer_output[914] + last_layer_output[915] + last_layer_output[916] + last_layer_output[917] + last_layer_output[918] + last_layer_output[919] + last_layer_output[920] + last_layer_output[921] + last_layer_output[922] + last_layer_output[923] + last_layer_output[924] + last_layer_output[925] + last_layer_output[926] + last_layer_output[927] + last_layer_output[928] + last_layer_output[929] + last_layer_output[930] + last_layer_output[931] + last_layer_output[932] + last_layer_output[933] + last_layer_output[934] + last_layer_output[935] + last_layer_output[936] + last_layer_output[937] + last_layer_output[938] + last_layer_output[939] + last_layer_output[940] + last_layer_output[941] + last_layer_output[942] + last_layer_output[943] + last_layer_output[944] + last_layer_output[945] + last_layer_output[946] + last_layer_output[947] + last_layer_output[948] + last_layer_output[949] + last_layer_output[950] + last_layer_output[951] + last_layer_output[952] + last_layer_output[953] + last_layer_output[954] + last_layer_output[955] + last_layer_output[956] + last_layer_output[957] + last_layer_output[958] + last_layer_output[959] + last_layer_output[960] + last_layer_output[961] + last_layer_output[962] + last_layer_output[963] + last_layer_output[964] + last_layer_output[965] + last_layer_output[966] + last_layer_output[967] + last_layer_output[968] + last_layer_output[969] + last_layer_output[970] + last_layer_output[971] + last_layer_output[972] + last_layer_output[973] + last_layer_output[974] + last_layer_output[975] + last_layer_output[976] + last_layer_output[977] + last_layer_output[978] + last_layer_output[979] + last_layer_output[980] + last_layer_output[981] + last_layer_output[982] + last_layer_output[983] + last_layer_output[984] + last_layer_output[985] + last_layer_output[986] + last_layer_output[987] + last_layer_output[988] + last_layer_output[989] + last_layer_output[990] + last_layer_output[991] + last_layer_output[992] + last_layer_output[993] + last_layer_output[994] + last_layer_output[995] + last_layer_output[996] + last_layer_output[997] + last_layer_output[998] + last_layer_output[999] + last_layer_output[1000] + last_layer_output[1001] + last_layer_output[1002] + last_layer_output[1003] + last_layer_output[1004] + last_layer_output[1005] + last_layer_output[1006] + last_layer_output[1007] + last_layer_output[1008] + last_layer_output[1009] + last_layer_output[1010] + last_layer_output[1011] + last_layer_output[1012] + last_layer_output[1013] + last_layer_output[1014] + last_layer_output[1015] + last_layer_output[1016] + last_layer_output[1017] + last_layer_output[1018] + last_layer_output[1019] + last_layer_output[1020] + last_layer_output[1021] + last_layer_output[1022] + last_layer_output[1023] + last_layer_output[1024] + last_layer_output[1025] + last_layer_output[1026] + last_layer_output[1027] + last_layer_output[1028] + last_layer_output[1029] + last_layer_output[1030] + last_layer_output[1031] + last_layer_output[1032] + last_layer_output[1033] + last_layer_output[1034] + last_layer_output[1035] + last_layer_output[1036] + last_layer_output[1037] + last_layer_output[1038] + last_layer_output[1039] + last_layer_output[1040] + last_layer_output[1041] + last_layer_output[1042] + last_layer_output[1043] + last_layer_output[1044] + last_layer_output[1045] + last_layer_output[1046] + last_layer_output[1047] + last_layer_output[1048] + last_layer_output[1049] + last_layer_output[1050] + last_layer_output[1051] + last_layer_output[1052] + last_layer_output[1053] + last_layer_output[1054] + last_layer_output[1055] + last_layer_output[1056] + last_layer_output[1057] + last_layer_output[1058] + last_layer_output[1059] + last_layer_output[1060] + last_layer_output[1061] + last_layer_output[1062] + last_layer_output[1063] + last_layer_output[1064] + last_layer_output[1065] + last_layer_output[1066] + last_layer_output[1067] + last_layer_output[1068] + last_layer_output[1069] + last_layer_output[1070] + last_layer_output[1071] + last_layer_output[1072] + last_layer_output[1073] + last_layer_output[1074] + last_layer_output[1075] + last_layer_output[1076] + last_layer_output[1077] + last_layer_output[1078] + last_layer_output[1079] + last_layer_output[1080] + last_layer_output[1081] + last_layer_output[1082] + last_layer_output[1083] + last_layer_output[1084] + last_layer_output[1085] + last_layer_output[1086] + last_layer_output[1087] + last_layer_output[1088] + last_layer_output[1089] + last_layer_output[1090] + last_layer_output[1091] + last_layer_output[1092] + last_layer_output[1093] + last_layer_output[1094] + last_layer_output[1095] + last_layer_output[1096] + last_layer_output[1097] + last_layer_output[1098] + last_layer_output[1099] + last_layer_output[1100] + last_layer_output[1101] + last_layer_output[1102] + last_layer_output[1103] + last_layer_output[1104] + last_layer_output[1105] + last_layer_output[1106] + last_layer_output[1107] + last_layer_output[1108] + last_layer_output[1109] + last_layer_output[1110] + last_layer_output[1111] + last_layer_output[1112] + last_layer_output[1113] + last_layer_output[1114] + last_layer_output[1115] + last_layer_output[1116] + last_layer_output[1117] + last_layer_output[1118] + last_layer_output[1119] + last_layer_output[1120] + last_layer_output[1121] + last_layer_output[1122] + last_layer_output[1123] + last_layer_output[1124] + last_layer_output[1125] + last_layer_output[1126] + last_layer_output[1127] + last_layer_output[1128] + last_layer_output[1129] + last_layer_output[1130] + last_layer_output[1131] + last_layer_output[1132] + last_layer_output[1133] + last_layer_output[1134] + last_layer_output[1135] + last_layer_output[1136] + last_layer_output[1137] + last_layer_output[1138] + last_layer_output[1139] + last_layer_output[1140] + last_layer_output[1141] + last_layer_output[1142] + last_layer_output[1143] + last_layer_output[1144] + last_layer_output[1145] + last_layer_output[1146] + last_layer_output[1147] + last_layer_output[1148] + last_layer_output[1149] + last_layer_output[1150] + last_layer_output[1151] + last_layer_output[1152] + last_layer_output[1153] + last_layer_output[1154] + last_layer_output[1155] + last_layer_output[1156] + last_layer_output[1157] + last_layer_output[1158] + last_layer_output[1159] + last_layer_output[1160] + last_layer_output[1161] + last_layer_output[1162] + last_layer_output[1163] + last_layer_output[1164] + last_layer_output[1165] + last_layer_output[1166] + last_layer_output[1167] + last_layer_output[1168] + last_layer_output[1169] + last_layer_output[1170] + last_layer_output[1171] + last_layer_output[1172] + last_layer_output[1173] + last_layer_output[1174] + last_layer_output[1175] + last_layer_output[1176] + last_layer_output[1177] + last_layer_output[1178] + last_layer_output[1179] + last_layer_output[1180] + last_layer_output[1181] + last_layer_output[1182] + last_layer_output[1183] + last_layer_output[1184] + last_layer_output[1185] + last_layer_output[1186] + last_layer_output[1187] + last_layer_output[1188] + last_layer_output[1189] + last_layer_output[1190] + last_layer_output[1191] + last_layer_output[1192] + last_layer_output[1193] + last_layer_output[1194] + last_layer_output[1195] + last_layer_output[1196] + last_layer_output[1197] + last_layer_output[1198] + last_layer_output[1199];
      result[1] <= last_layer_output[1200] + last_layer_output[1201] + last_layer_output[1202] + last_layer_output[1203] + last_layer_output[1204] + last_layer_output[1205] + last_layer_output[1206] + last_layer_output[1207] + last_layer_output[1208] + last_layer_output[1209] + last_layer_output[1210] + last_layer_output[1211] + last_layer_output[1212] + last_layer_output[1213] + last_layer_output[1214] + last_layer_output[1215] + last_layer_output[1216] + last_layer_output[1217] + last_layer_output[1218] + last_layer_output[1219] + last_layer_output[1220] + last_layer_output[1221] + last_layer_output[1222] + last_layer_output[1223] + last_layer_output[1224] + last_layer_output[1225] + last_layer_output[1226] + last_layer_output[1227] + last_layer_output[1228] + last_layer_output[1229] + last_layer_output[1230] + last_layer_output[1231] + last_layer_output[1232] + last_layer_output[1233] + last_layer_output[1234] + last_layer_output[1235] + last_layer_output[1236] + last_layer_output[1237] + last_layer_output[1238] + last_layer_output[1239] + last_layer_output[1240] + last_layer_output[1241] + last_layer_output[1242] + last_layer_output[1243] + last_layer_output[1244] + last_layer_output[1245] + last_layer_output[1246] + last_layer_output[1247] + last_layer_output[1248] + last_layer_output[1249] + last_layer_output[1250] + last_layer_output[1251] + last_layer_output[1252] + last_layer_output[1253] + last_layer_output[1254] + last_layer_output[1255] + last_layer_output[1256] + last_layer_output[1257] + last_layer_output[1258] + last_layer_output[1259] + last_layer_output[1260] + last_layer_output[1261] + last_layer_output[1262] + last_layer_output[1263] + last_layer_output[1264] + last_layer_output[1265] + last_layer_output[1266] + last_layer_output[1267] + last_layer_output[1268] + last_layer_output[1269] + last_layer_output[1270] + last_layer_output[1271] + last_layer_output[1272] + last_layer_output[1273] + last_layer_output[1274] + last_layer_output[1275] + last_layer_output[1276] + last_layer_output[1277] + last_layer_output[1278] + last_layer_output[1279] + last_layer_output[1280] + last_layer_output[1281] + last_layer_output[1282] + last_layer_output[1283] + last_layer_output[1284] + last_layer_output[1285] + last_layer_output[1286] + last_layer_output[1287] + last_layer_output[1288] + last_layer_output[1289] + last_layer_output[1290] + last_layer_output[1291] + last_layer_output[1292] + last_layer_output[1293] + last_layer_output[1294] + last_layer_output[1295] + last_layer_output[1296] + last_layer_output[1297] + last_layer_output[1298] + last_layer_output[1299] + last_layer_output[1300] + last_layer_output[1301] + last_layer_output[1302] + last_layer_output[1303] + last_layer_output[1304] + last_layer_output[1305] + last_layer_output[1306] + last_layer_output[1307] + last_layer_output[1308] + last_layer_output[1309] + last_layer_output[1310] + last_layer_output[1311] + last_layer_output[1312] + last_layer_output[1313] + last_layer_output[1314] + last_layer_output[1315] + last_layer_output[1316] + last_layer_output[1317] + last_layer_output[1318] + last_layer_output[1319] + last_layer_output[1320] + last_layer_output[1321] + last_layer_output[1322] + last_layer_output[1323] + last_layer_output[1324] + last_layer_output[1325] + last_layer_output[1326] + last_layer_output[1327] + last_layer_output[1328] + last_layer_output[1329] + last_layer_output[1330] + last_layer_output[1331] + last_layer_output[1332] + last_layer_output[1333] + last_layer_output[1334] + last_layer_output[1335] + last_layer_output[1336] + last_layer_output[1337] + last_layer_output[1338] + last_layer_output[1339] + last_layer_output[1340] + last_layer_output[1341] + last_layer_output[1342] + last_layer_output[1343] + last_layer_output[1344] + last_layer_output[1345] + last_layer_output[1346] + last_layer_output[1347] + last_layer_output[1348] + last_layer_output[1349] + last_layer_output[1350] + last_layer_output[1351] + last_layer_output[1352] + last_layer_output[1353] + last_layer_output[1354] + last_layer_output[1355] + last_layer_output[1356] + last_layer_output[1357] + last_layer_output[1358] + last_layer_output[1359] + last_layer_output[1360] + last_layer_output[1361] + last_layer_output[1362] + last_layer_output[1363] + last_layer_output[1364] + last_layer_output[1365] + last_layer_output[1366] + last_layer_output[1367] + last_layer_output[1368] + last_layer_output[1369] + last_layer_output[1370] + last_layer_output[1371] + last_layer_output[1372] + last_layer_output[1373] + last_layer_output[1374] + last_layer_output[1375] + last_layer_output[1376] + last_layer_output[1377] + last_layer_output[1378] + last_layer_output[1379] + last_layer_output[1380] + last_layer_output[1381] + last_layer_output[1382] + last_layer_output[1383] + last_layer_output[1384] + last_layer_output[1385] + last_layer_output[1386] + last_layer_output[1387] + last_layer_output[1388] + last_layer_output[1389] + last_layer_output[1390] + last_layer_output[1391] + last_layer_output[1392] + last_layer_output[1393] + last_layer_output[1394] + last_layer_output[1395] + last_layer_output[1396] + last_layer_output[1397] + last_layer_output[1398] + last_layer_output[1399] + last_layer_output[1400] + last_layer_output[1401] + last_layer_output[1402] + last_layer_output[1403] + last_layer_output[1404] + last_layer_output[1405] + last_layer_output[1406] + last_layer_output[1407] + last_layer_output[1408] + last_layer_output[1409] + last_layer_output[1410] + last_layer_output[1411] + last_layer_output[1412] + last_layer_output[1413] + last_layer_output[1414] + last_layer_output[1415] + last_layer_output[1416] + last_layer_output[1417] + last_layer_output[1418] + last_layer_output[1419] + last_layer_output[1420] + last_layer_output[1421] + last_layer_output[1422] + last_layer_output[1423] + last_layer_output[1424] + last_layer_output[1425] + last_layer_output[1426] + last_layer_output[1427] + last_layer_output[1428] + last_layer_output[1429] + last_layer_output[1430] + last_layer_output[1431] + last_layer_output[1432] + last_layer_output[1433] + last_layer_output[1434] + last_layer_output[1435] + last_layer_output[1436] + last_layer_output[1437] + last_layer_output[1438] + last_layer_output[1439] + last_layer_output[1440] + last_layer_output[1441] + last_layer_output[1442] + last_layer_output[1443] + last_layer_output[1444] + last_layer_output[1445] + last_layer_output[1446] + last_layer_output[1447] + last_layer_output[1448] + last_layer_output[1449] + last_layer_output[1450] + last_layer_output[1451] + last_layer_output[1452] + last_layer_output[1453] + last_layer_output[1454] + last_layer_output[1455] + last_layer_output[1456] + last_layer_output[1457] + last_layer_output[1458] + last_layer_output[1459] + last_layer_output[1460] + last_layer_output[1461] + last_layer_output[1462] + last_layer_output[1463] + last_layer_output[1464] + last_layer_output[1465] + last_layer_output[1466] + last_layer_output[1467] + last_layer_output[1468] + last_layer_output[1469] + last_layer_output[1470] + last_layer_output[1471] + last_layer_output[1472] + last_layer_output[1473] + last_layer_output[1474] + last_layer_output[1475] + last_layer_output[1476] + last_layer_output[1477] + last_layer_output[1478] + last_layer_output[1479] + last_layer_output[1480] + last_layer_output[1481] + last_layer_output[1482] + last_layer_output[1483] + last_layer_output[1484] + last_layer_output[1485] + last_layer_output[1486] + last_layer_output[1487] + last_layer_output[1488] + last_layer_output[1489] + last_layer_output[1490] + last_layer_output[1491] + last_layer_output[1492] + last_layer_output[1493] + last_layer_output[1494] + last_layer_output[1495] + last_layer_output[1496] + last_layer_output[1497] + last_layer_output[1498] + last_layer_output[1499] + last_layer_output[1500] + last_layer_output[1501] + last_layer_output[1502] + last_layer_output[1503] + last_layer_output[1504] + last_layer_output[1505] + last_layer_output[1506] + last_layer_output[1507] + last_layer_output[1508] + last_layer_output[1509] + last_layer_output[1510] + last_layer_output[1511] + last_layer_output[1512] + last_layer_output[1513] + last_layer_output[1514] + last_layer_output[1515] + last_layer_output[1516] + last_layer_output[1517] + last_layer_output[1518] + last_layer_output[1519] + last_layer_output[1520] + last_layer_output[1521] + last_layer_output[1522] + last_layer_output[1523] + last_layer_output[1524] + last_layer_output[1525] + last_layer_output[1526] + last_layer_output[1527] + last_layer_output[1528] + last_layer_output[1529] + last_layer_output[1530] + last_layer_output[1531] + last_layer_output[1532] + last_layer_output[1533] + last_layer_output[1534] + last_layer_output[1535] + last_layer_output[1536] + last_layer_output[1537] + last_layer_output[1538] + last_layer_output[1539] + last_layer_output[1540] + last_layer_output[1541] + last_layer_output[1542] + last_layer_output[1543] + last_layer_output[1544] + last_layer_output[1545] + last_layer_output[1546] + last_layer_output[1547] + last_layer_output[1548] + last_layer_output[1549] + last_layer_output[1550] + last_layer_output[1551] + last_layer_output[1552] + last_layer_output[1553] + last_layer_output[1554] + last_layer_output[1555] + last_layer_output[1556] + last_layer_output[1557] + last_layer_output[1558] + last_layer_output[1559] + last_layer_output[1560] + last_layer_output[1561] + last_layer_output[1562] + last_layer_output[1563] + last_layer_output[1564] + last_layer_output[1565] + last_layer_output[1566] + last_layer_output[1567] + last_layer_output[1568] + last_layer_output[1569] + last_layer_output[1570] + last_layer_output[1571] + last_layer_output[1572] + last_layer_output[1573] + last_layer_output[1574] + last_layer_output[1575] + last_layer_output[1576] + last_layer_output[1577] + last_layer_output[1578] + last_layer_output[1579] + last_layer_output[1580] + last_layer_output[1581] + last_layer_output[1582] + last_layer_output[1583] + last_layer_output[1584] + last_layer_output[1585] + last_layer_output[1586] + last_layer_output[1587] + last_layer_output[1588] + last_layer_output[1589] + last_layer_output[1590] + last_layer_output[1591] + last_layer_output[1592] + last_layer_output[1593] + last_layer_output[1594] + last_layer_output[1595] + last_layer_output[1596] + last_layer_output[1597] + last_layer_output[1598] + last_layer_output[1599] + last_layer_output[1600] + last_layer_output[1601] + last_layer_output[1602] + last_layer_output[1603] + last_layer_output[1604] + last_layer_output[1605] + last_layer_output[1606] + last_layer_output[1607] + last_layer_output[1608] + last_layer_output[1609] + last_layer_output[1610] + last_layer_output[1611] + last_layer_output[1612] + last_layer_output[1613] + last_layer_output[1614] + last_layer_output[1615] + last_layer_output[1616] + last_layer_output[1617] + last_layer_output[1618] + last_layer_output[1619] + last_layer_output[1620] + last_layer_output[1621] + last_layer_output[1622] + last_layer_output[1623] + last_layer_output[1624] + last_layer_output[1625] + last_layer_output[1626] + last_layer_output[1627] + last_layer_output[1628] + last_layer_output[1629] + last_layer_output[1630] + last_layer_output[1631] + last_layer_output[1632] + last_layer_output[1633] + last_layer_output[1634] + last_layer_output[1635] + last_layer_output[1636] + last_layer_output[1637] + last_layer_output[1638] + last_layer_output[1639] + last_layer_output[1640] + last_layer_output[1641] + last_layer_output[1642] + last_layer_output[1643] + last_layer_output[1644] + last_layer_output[1645] + last_layer_output[1646] + last_layer_output[1647] + last_layer_output[1648] + last_layer_output[1649] + last_layer_output[1650] + last_layer_output[1651] + last_layer_output[1652] + last_layer_output[1653] + last_layer_output[1654] + last_layer_output[1655] + last_layer_output[1656] + last_layer_output[1657] + last_layer_output[1658] + last_layer_output[1659] + last_layer_output[1660] + last_layer_output[1661] + last_layer_output[1662] + last_layer_output[1663] + last_layer_output[1664] + last_layer_output[1665] + last_layer_output[1666] + last_layer_output[1667] + last_layer_output[1668] + last_layer_output[1669] + last_layer_output[1670] + last_layer_output[1671] + last_layer_output[1672] + last_layer_output[1673] + last_layer_output[1674] + last_layer_output[1675] + last_layer_output[1676] + last_layer_output[1677] + last_layer_output[1678] + last_layer_output[1679] + last_layer_output[1680] + last_layer_output[1681] + last_layer_output[1682] + last_layer_output[1683] + last_layer_output[1684] + last_layer_output[1685] + last_layer_output[1686] + last_layer_output[1687] + last_layer_output[1688] + last_layer_output[1689] + last_layer_output[1690] + last_layer_output[1691] + last_layer_output[1692] + last_layer_output[1693] + last_layer_output[1694] + last_layer_output[1695] + last_layer_output[1696] + last_layer_output[1697] + last_layer_output[1698] + last_layer_output[1699] + last_layer_output[1700] + last_layer_output[1701] + last_layer_output[1702] + last_layer_output[1703] + last_layer_output[1704] + last_layer_output[1705] + last_layer_output[1706] + last_layer_output[1707] + last_layer_output[1708] + last_layer_output[1709] + last_layer_output[1710] + last_layer_output[1711] + last_layer_output[1712] + last_layer_output[1713] + last_layer_output[1714] + last_layer_output[1715] + last_layer_output[1716] + last_layer_output[1717] + last_layer_output[1718] + last_layer_output[1719] + last_layer_output[1720] + last_layer_output[1721] + last_layer_output[1722] + last_layer_output[1723] + last_layer_output[1724] + last_layer_output[1725] + last_layer_output[1726] + last_layer_output[1727] + last_layer_output[1728] + last_layer_output[1729] + last_layer_output[1730] + last_layer_output[1731] + last_layer_output[1732] + last_layer_output[1733] + last_layer_output[1734] + last_layer_output[1735] + last_layer_output[1736] + last_layer_output[1737] + last_layer_output[1738] + last_layer_output[1739] + last_layer_output[1740] + last_layer_output[1741] + last_layer_output[1742] + last_layer_output[1743] + last_layer_output[1744] + last_layer_output[1745] + last_layer_output[1746] + last_layer_output[1747] + last_layer_output[1748] + last_layer_output[1749] + last_layer_output[1750] + last_layer_output[1751] + last_layer_output[1752] + last_layer_output[1753] + last_layer_output[1754] + last_layer_output[1755] + last_layer_output[1756] + last_layer_output[1757] + last_layer_output[1758] + last_layer_output[1759] + last_layer_output[1760] + last_layer_output[1761] + last_layer_output[1762] + last_layer_output[1763] + last_layer_output[1764] + last_layer_output[1765] + last_layer_output[1766] + last_layer_output[1767] + last_layer_output[1768] + last_layer_output[1769] + last_layer_output[1770] + last_layer_output[1771] + last_layer_output[1772] + last_layer_output[1773] + last_layer_output[1774] + last_layer_output[1775] + last_layer_output[1776] + last_layer_output[1777] + last_layer_output[1778] + last_layer_output[1779] + last_layer_output[1780] + last_layer_output[1781] + last_layer_output[1782] + last_layer_output[1783] + last_layer_output[1784] + last_layer_output[1785] + last_layer_output[1786] + last_layer_output[1787] + last_layer_output[1788] + last_layer_output[1789] + last_layer_output[1790] + last_layer_output[1791] + last_layer_output[1792] + last_layer_output[1793] + last_layer_output[1794] + last_layer_output[1795] + last_layer_output[1796] + last_layer_output[1797] + last_layer_output[1798] + last_layer_output[1799] + last_layer_output[1800] + last_layer_output[1801] + last_layer_output[1802] + last_layer_output[1803] + last_layer_output[1804] + last_layer_output[1805] + last_layer_output[1806] + last_layer_output[1807] + last_layer_output[1808] + last_layer_output[1809] + last_layer_output[1810] + last_layer_output[1811] + last_layer_output[1812] + last_layer_output[1813] + last_layer_output[1814] + last_layer_output[1815] + last_layer_output[1816] + last_layer_output[1817] + last_layer_output[1818] + last_layer_output[1819] + last_layer_output[1820] + last_layer_output[1821] + last_layer_output[1822] + last_layer_output[1823] + last_layer_output[1824] + last_layer_output[1825] + last_layer_output[1826] + last_layer_output[1827] + last_layer_output[1828] + last_layer_output[1829] + last_layer_output[1830] + last_layer_output[1831] + last_layer_output[1832] + last_layer_output[1833] + last_layer_output[1834] + last_layer_output[1835] + last_layer_output[1836] + last_layer_output[1837] + last_layer_output[1838] + last_layer_output[1839] + last_layer_output[1840] + last_layer_output[1841] + last_layer_output[1842] + last_layer_output[1843] + last_layer_output[1844] + last_layer_output[1845] + last_layer_output[1846] + last_layer_output[1847] + last_layer_output[1848] + last_layer_output[1849] + last_layer_output[1850] + last_layer_output[1851] + last_layer_output[1852] + last_layer_output[1853] + last_layer_output[1854] + last_layer_output[1855] + last_layer_output[1856] + last_layer_output[1857] + last_layer_output[1858] + last_layer_output[1859] + last_layer_output[1860] + last_layer_output[1861] + last_layer_output[1862] + last_layer_output[1863] + last_layer_output[1864] + last_layer_output[1865] + last_layer_output[1866] + last_layer_output[1867] + last_layer_output[1868] + last_layer_output[1869] + last_layer_output[1870] + last_layer_output[1871] + last_layer_output[1872] + last_layer_output[1873] + last_layer_output[1874] + last_layer_output[1875] + last_layer_output[1876] + last_layer_output[1877] + last_layer_output[1878] + last_layer_output[1879] + last_layer_output[1880] + last_layer_output[1881] + last_layer_output[1882] + last_layer_output[1883] + last_layer_output[1884] + last_layer_output[1885] + last_layer_output[1886] + last_layer_output[1887] + last_layer_output[1888] + last_layer_output[1889] + last_layer_output[1890] + last_layer_output[1891] + last_layer_output[1892] + last_layer_output[1893] + last_layer_output[1894] + last_layer_output[1895] + last_layer_output[1896] + last_layer_output[1897] + last_layer_output[1898] + last_layer_output[1899] + last_layer_output[1900] + last_layer_output[1901] + last_layer_output[1902] + last_layer_output[1903] + last_layer_output[1904] + last_layer_output[1905] + last_layer_output[1906] + last_layer_output[1907] + last_layer_output[1908] + last_layer_output[1909] + last_layer_output[1910] + last_layer_output[1911] + last_layer_output[1912] + last_layer_output[1913] + last_layer_output[1914] + last_layer_output[1915] + last_layer_output[1916] + last_layer_output[1917] + last_layer_output[1918] + last_layer_output[1919] + last_layer_output[1920] + last_layer_output[1921] + last_layer_output[1922] + last_layer_output[1923] + last_layer_output[1924] + last_layer_output[1925] + last_layer_output[1926] + last_layer_output[1927] + last_layer_output[1928] + last_layer_output[1929] + last_layer_output[1930] + last_layer_output[1931] + last_layer_output[1932] + last_layer_output[1933] + last_layer_output[1934] + last_layer_output[1935] + last_layer_output[1936] + last_layer_output[1937] + last_layer_output[1938] + last_layer_output[1939] + last_layer_output[1940] + last_layer_output[1941] + last_layer_output[1942] + last_layer_output[1943] + last_layer_output[1944] + last_layer_output[1945] + last_layer_output[1946] + last_layer_output[1947] + last_layer_output[1948] + last_layer_output[1949] + last_layer_output[1950] + last_layer_output[1951] + last_layer_output[1952] + last_layer_output[1953] + last_layer_output[1954] + last_layer_output[1955] + last_layer_output[1956] + last_layer_output[1957] + last_layer_output[1958] + last_layer_output[1959] + last_layer_output[1960] + last_layer_output[1961] + last_layer_output[1962] + last_layer_output[1963] + last_layer_output[1964] + last_layer_output[1965] + last_layer_output[1966] + last_layer_output[1967] + last_layer_output[1968] + last_layer_output[1969] + last_layer_output[1970] + last_layer_output[1971] + last_layer_output[1972] + last_layer_output[1973] + last_layer_output[1974] + last_layer_output[1975] + last_layer_output[1976] + last_layer_output[1977] + last_layer_output[1978] + last_layer_output[1979] + last_layer_output[1980] + last_layer_output[1981] + last_layer_output[1982] + last_layer_output[1983] + last_layer_output[1984] + last_layer_output[1985] + last_layer_output[1986] + last_layer_output[1987] + last_layer_output[1988] + last_layer_output[1989] + last_layer_output[1990] + last_layer_output[1991] + last_layer_output[1992] + last_layer_output[1993] + last_layer_output[1994] + last_layer_output[1995] + last_layer_output[1996] + last_layer_output[1997] + last_layer_output[1998] + last_layer_output[1999] + last_layer_output[2000] + last_layer_output[2001] + last_layer_output[2002] + last_layer_output[2003] + last_layer_output[2004] + last_layer_output[2005] + last_layer_output[2006] + last_layer_output[2007] + last_layer_output[2008] + last_layer_output[2009] + last_layer_output[2010] + last_layer_output[2011] + last_layer_output[2012] + last_layer_output[2013] + last_layer_output[2014] + last_layer_output[2015] + last_layer_output[2016] + last_layer_output[2017] + last_layer_output[2018] + last_layer_output[2019] + last_layer_output[2020] + last_layer_output[2021] + last_layer_output[2022] + last_layer_output[2023] + last_layer_output[2024] + last_layer_output[2025] + last_layer_output[2026] + last_layer_output[2027] + last_layer_output[2028] + last_layer_output[2029] + last_layer_output[2030] + last_layer_output[2031] + last_layer_output[2032] + last_layer_output[2033] + last_layer_output[2034] + last_layer_output[2035] + last_layer_output[2036] + last_layer_output[2037] + last_layer_output[2038] + last_layer_output[2039] + last_layer_output[2040] + last_layer_output[2041] + last_layer_output[2042] + last_layer_output[2043] + last_layer_output[2044] + last_layer_output[2045] + last_layer_output[2046] + last_layer_output[2047] + last_layer_output[2048] + last_layer_output[2049] + last_layer_output[2050] + last_layer_output[2051] + last_layer_output[2052] + last_layer_output[2053] + last_layer_output[2054] + last_layer_output[2055] + last_layer_output[2056] + last_layer_output[2057] + last_layer_output[2058] + last_layer_output[2059] + last_layer_output[2060] + last_layer_output[2061] + last_layer_output[2062] + last_layer_output[2063] + last_layer_output[2064] + last_layer_output[2065] + last_layer_output[2066] + last_layer_output[2067] + last_layer_output[2068] + last_layer_output[2069] + last_layer_output[2070] + last_layer_output[2071] + last_layer_output[2072] + last_layer_output[2073] + last_layer_output[2074] + last_layer_output[2075] + last_layer_output[2076] + last_layer_output[2077] + last_layer_output[2078] + last_layer_output[2079] + last_layer_output[2080] + last_layer_output[2081] + last_layer_output[2082] + last_layer_output[2083] + last_layer_output[2084] + last_layer_output[2085] + last_layer_output[2086] + last_layer_output[2087] + last_layer_output[2088] + last_layer_output[2089] + last_layer_output[2090] + last_layer_output[2091] + last_layer_output[2092] + last_layer_output[2093] + last_layer_output[2094] + last_layer_output[2095] + last_layer_output[2096] + last_layer_output[2097] + last_layer_output[2098] + last_layer_output[2099] + last_layer_output[2100] + last_layer_output[2101] + last_layer_output[2102] + last_layer_output[2103] + last_layer_output[2104] + last_layer_output[2105] + last_layer_output[2106] + last_layer_output[2107] + last_layer_output[2108] + last_layer_output[2109] + last_layer_output[2110] + last_layer_output[2111] + last_layer_output[2112] + last_layer_output[2113] + last_layer_output[2114] + last_layer_output[2115] + last_layer_output[2116] + last_layer_output[2117] + last_layer_output[2118] + last_layer_output[2119] + last_layer_output[2120] + last_layer_output[2121] + last_layer_output[2122] + last_layer_output[2123] + last_layer_output[2124] + last_layer_output[2125] + last_layer_output[2126] + last_layer_output[2127] + last_layer_output[2128] + last_layer_output[2129] + last_layer_output[2130] + last_layer_output[2131] + last_layer_output[2132] + last_layer_output[2133] + last_layer_output[2134] + last_layer_output[2135] + last_layer_output[2136] + last_layer_output[2137] + last_layer_output[2138] + last_layer_output[2139] + last_layer_output[2140] + last_layer_output[2141] + last_layer_output[2142] + last_layer_output[2143] + last_layer_output[2144] + last_layer_output[2145] + last_layer_output[2146] + last_layer_output[2147] + last_layer_output[2148] + last_layer_output[2149] + last_layer_output[2150] + last_layer_output[2151] + last_layer_output[2152] + last_layer_output[2153] + last_layer_output[2154] + last_layer_output[2155] + last_layer_output[2156] + last_layer_output[2157] + last_layer_output[2158] + last_layer_output[2159] + last_layer_output[2160] + last_layer_output[2161] + last_layer_output[2162] + last_layer_output[2163] + last_layer_output[2164] + last_layer_output[2165] + last_layer_output[2166] + last_layer_output[2167] + last_layer_output[2168] + last_layer_output[2169] + last_layer_output[2170] + last_layer_output[2171] + last_layer_output[2172] + last_layer_output[2173] + last_layer_output[2174] + last_layer_output[2175] + last_layer_output[2176] + last_layer_output[2177] + last_layer_output[2178] + last_layer_output[2179] + last_layer_output[2180] + last_layer_output[2181] + last_layer_output[2182] + last_layer_output[2183] + last_layer_output[2184] + last_layer_output[2185] + last_layer_output[2186] + last_layer_output[2187] + last_layer_output[2188] + last_layer_output[2189] + last_layer_output[2190] + last_layer_output[2191] + last_layer_output[2192] + last_layer_output[2193] + last_layer_output[2194] + last_layer_output[2195] + last_layer_output[2196] + last_layer_output[2197] + last_layer_output[2198] + last_layer_output[2199] + last_layer_output[2200] + last_layer_output[2201] + last_layer_output[2202] + last_layer_output[2203] + last_layer_output[2204] + last_layer_output[2205] + last_layer_output[2206] + last_layer_output[2207] + last_layer_output[2208] + last_layer_output[2209] + last_layer_output[2210] + last_layer_output[2211] + last_layer_output[2212] + last_layer_output[2213] + last_layer_output[2214] + last_layer_output[2215] + last_layer_output[2216] + last_layer_output[2217] + last_layer_output[2218] + last_layer_output[2219] + last_layer_output[2220] + last_layer_output[2221] + last_layer_output[2222] + last_layer_output[2223] + last_layer_output[2224] + last_layer_output[2225] + last_layer_output[2226] + last_layer_output[2227] + last_layer_output[2228] + last_layer_output[2229] + last_layer_output[2230] + last_layer_output[2231] + last_layer_output[2232] + last_layer_output[2233] + last_layer_output[2234] + last_layer_output[2235] + last_layer_output[2236] + last_layer_output[2237] + last_layer_output[2238] + last_layer_output[2239] + last_layer_output[2240] + last_layer_output[2241] + last_layer_output[2242] + last_layer_output[2243] + last_layer_output[2244] + last_layer_output[2245] + last_layer_output[2246] + last_layer_output[2247] + last_layer_output[2248] + last_layer_output[2249] + last_layer_output[2250] + last_layer_output[2251] + last_layer_output[2252] + last_layer_output[2253] + last_layer_output[2254] + last_layer_output[2255] + last_layer_output[2256] + last_layer_output[2257] + last_layer_output[2258] + last_layer_output[2259] + last_layer_output[2260] + last_layer_output[2261] + last_layer_output[2262] + last_layer_output[2263] + last_layer_output[2264] + last_layer_output[2265] + last_layer_output[2266] + last_layer_output[2267] + last_layer_output[2268] + last_layer_output[2269] + last_layer_output[2270] + last_layer_output[2271] + last_layer_output[2272] + last_layer_output[2273] + last_layer_output[2274] + last_layer_output[2275] + last_layer_output[2276] + last_layer_output[2277] + last_layer_output[2278] + last_layer_output[2279] + last_layer_output[2280] + last_layer_output[2281] + last_layer_output[2282] + last_layer_output[2283] + last_layer_output[2284] + last_layer_output[2285] + last_layer_output[2286] + last_layer_output[2287] + last_layer_output[2288] + last_layer_output[2289] + last_layer_output[2290] + last_layer_output[2291] + last_layer_output[2292] + last_layer_output[2293] + last_layer_output[2294] + last_layer_output[2295] + last_layer_output[2296] + last_layer_output[2297] + last_layer_output[2298] + last_layer_output[2299] + last_layer_output[2300] + last_layer_output[2301] + last_layer_output[2302] + last_layer_output[2303] + last_layer_output[2304] + last_layer_output[2305] + last_layer_output[2306] + last_layer_output[2307] + last_layer_output[2308] + last_layer_output[2309] + last_layer_output[2310] + last_layer_output[2311] + last_layer_output[2312] + last_layer_output[2313] + last_layer_output[2314] + last_layer_output[2315] + last_layer_output[2316] + last_layer_output[2317] + last_layer_output[2318] + last_layer_output[2319] + last_layer_output[2320] + last_layer_output[2321] + last_layer_output[2322] + last_layer_output[2323] + last_layer_output[2324] + last_layer_output[2325] + last_layer_output[2326] + last_layer_output[2327] + last_layer_output[2328] + last_layer_output[2329] + last_layer_output[2330] + last_layer_output[2331] + last_layer_output[2332] + last_layer_output[2333] + last_layer_output[2334] + last_layer_output[2335] + last_layer_output[2336] + last_layer_output[2337] + last_layer_output[2338] + last_layer_output[2339] + last_layer_output[2340] + last_layer_output[2341] + last_layer_output[2342] + last_layer_output[2343] + last_layer_output[2344] + last_layer_output[2345] + last_layer_output[2346] + last_layer_output[2347] + last_layer_output[2348] + last_layer_output[2349] + last_layer_output[2350] + last_layer_output[2351] + last_layer_output[2352] + last_layer_output[2353] + last_layer_output[2354] + last_layer_output[2355] + last_layer_output[2356] + last_layer_output[2357] + last_layer_output[2358] + last_layer_output[2359] + last_layer_output[2360] + last_layer_output[2361] + last_layer_output[2362] + last_layer_output[2363] + last_layer_output[2364] + last_layer_output[2365] + last_layer_output[2366] + last_layer_output[2367] + last_layer_output[2368] + last_layer_output[2369] + last_layer_output[2370] + last_layer_output[2371] + last_layer_output[2372] + last_layer_output[2373] + last_layer_output[2374] + last_layer_output[2375] + last_layer_output[2376] + last_layer_output[2377] + last_layer_output[2378] + last_layer_output[2379] + last_layer_output[2380] + last_layer_output[2381] + last_layer_output[2382] + last_layer_output[2383] + last_layer_output[2384] + last_layer_output[2385] + last_layer_output[2386] + last_layer_output[2387] + last_layer_output[2388] + last_layer_output[2389] + last_layer_output[2390] + last_layer_output[2391] + last_layer_output[2392] + last_layer_output[2393] + last_layer_output[2394] + last_layer_output[2395] + last_layer_output[2396] + last_layer_output[2397] + last_layer_output[2398] + last_layer_output[2399];
      result[2] <= last_layer_output[2400] + last_layer_output[2401] + last_layer_output[2402] + last_layer_output[2403] + last_layer_output[2404] + last_layer_output[2405] + last_layer_output[2406] + last_layer_output[2407] + last_layer_output[2408] + last_layer_output[2409] + last_layer_output[2410] + last_layer_output[2411] + last_layer_output[2412] + last_layer_output[2413] + last_layer_output[2414] + last_layer_output[2415] + last_layer_output[2416] + last_layer_output[2417] + last_layer_output[2418] + last_layer_output[2419] + last_layer_output[2420] + last_layer_output[2421] + last_layer_output[2422] + last_layer_output[2423] + last_layer_output[2424] + last_layer_output[2425] + last_layer_output[2426] + last_layer_output[2427] + last_layer_output[2428] + last_layer_output[2429] + last_layer_output[2430] + last_layer_output[2431] + last_layer_output[2432] + last_layer_output[2433] + last_layer_output[2434] + last_layer_output[2435] + last_layer_output[2436] + last_layer_output[2437] + last_layer_output[2438] + last_layer_output[2439] + last_layer_output[2440] + last_layer_output[2441] + last_layer_output[2442] + last_layer_output[2443] + last_layer_output[2444] + last_layer_output[2445] + last_layer_output[2446] + last_layer_output[2447] + last_layer_output[2448] + last_layer_output[2449] + last_layer_output[2450] + last_layer_output[2451] + last_layer_output[2452] + last_layer_output[2453] + last_layer_output[2454] + last_layer_output[2455] + last_layer_output[2456] + last_layer_output[2457] + last_layer_output[2458] + last_layer_output[2459] + last_layer_output[2460] + last_layer_output[2461] + last_layer_output[2462] + last_layer_output[2463] + last_layer_output[2464] + last_layer_output[2465] + last_layer_output[2466] + last_layer_output[2467] + last_layer_output[2468] + last_layer_output[2469] + last_layer_output[2470] + last_layer_output[2471] + last_layer_output[2472] + last_layer_output[2473] + last_layer_output[2474] + last_layer_output[2475] + last_layer_output[2476] + last_layer_output[2477] + last_layer_output[2478] + last_layer_output[2479] + last_layer_output[2480] + last_layer_output[2481] + last_layer_output[2482] + last_layer_output[2483] + last_layer_output[2484] + last_layer_output[2485] + last_layer_output[2486] + last_layer_output[2487] + last_layer_output[2488] + last_layer_output[2489] + last_layer_output[2490] + last_layer_output[2491] + last_layer_output[2492] + last_layer_output[2493] + last_layer_output[2494] + last_layer_output[2495] + last_layer_output[2496] + last_layer_output[2497] + last_layer_output[2498] + last_layer_output[2499] + last_layer_output[2500] + last_layer_output[2501] + last_layer_output[2502] + last_layer_output[2503] + last_layer_output[2504] + last_layer_output[2505] + last_layer_output[2506] + last_layer_output[2507] + last_layer_output[2508] + last_layer_output[2509] + last_layer_output[2510] + last_layer_output[2511] + last_layer_output[2512] + last_layer_output[2513] + last_layer_output[2514] + last_layer_output[2515] + last_layer_output[2516] + last_layer_output[2517] + last_layer_output[2518] + last_layer_output[2519] + last_layer_output[2520] + last_layer_output[2521] + last_layer_output[2522] + last_layer_output[2523] + last_layer_output[2524] + last_layer_output[2525] + last_layer_output[2526] + last_layer_output[2527] + last_layer_output[2528] + last_layer_output[2529] + last_layer_output[2530] + last_layer_output[2531] + last_layer_output[2532] + last_layer_output[2533] + last_layer_output[2534] + last_layer_output[2535] + last_layer_output[2536] + last_layer_output[2537] + last_layer_output[2538] + last_layer_output[2539] + last_layer_output[2540] + last_layer_output[2541] + last_layer_output[2542] + last_layer_output[2543] + last_layer_output[2544] + last_layer_output[2545] + last_layer_output[2546] + last_layer_output[2547] + last_layer_output[2548] + last_layer_output[2549] + last_layer_output[2550] + last_layer_output[2551] + last_layer_output[2552] + last_layer_output[2553] + last_layer_output[2554] + last_layer_output[2555] + last_layer_output[2556] + last_layer_output[2557] + last_layer_output[2558] + last_layer_output[2559] + last_layer_output[2560] + last_layer_output[2561] + last_layer_output[2562] + last_layer_output[2563] + last_layer_output[2564] + last_layer_output[2565] + last_layer_output[2566] + last_layer_output[2567] + last_layer_output[2568] + last_layer_output[2569] + last_layer_output[2570] + last_layer_output[2571] + last_layer_output[2572] + last_layer_output[2573] + last_layer_output[2574] + last_layer_output[2575] + last_layer_output[2576] + last_layer_output[2577] + last_layer_output[2578] + last_layer_output[2579] + last_layer_output[2580] + last_layer_output[2581] + last_layer_output[2582] + last_layer_output[2583] + last_layer_output[2584] + last_layer_output[2585] + last_layer_output[2586] + last_layer_output[2587] + last_layer_output[2588] + last_layer_output[2589] + last_layer_output[2590] + last_layer_output[2591] + last_layer_output[2592] + last_layer_output[2593] + last_layer_output[2594] + last_layer_output[2595] + last_layer_output[2596] + last_layer_output[2597] + last_layer_output[2598] + last_layer_output[2599] + last_layer_output[2600] + last_layer_output[2601] + last_layer_output[2602] + last_layer_output[2603] + last_layer_output[2604] + last_layer_output[2605] + last_layer_output[2606] + last_layer_output[2607] + last_layer_output[2608] + last_layer_output[2609] + last_layer_output[2610] + last_layer_output[2611] + last_layer_output[2612] + last_layer_output[2613] + last_layer_output[2614] + last_layer_output[2615] + last_layer_output[2616] + last_layer_output[2617] + last_layer_output[2618] + last_layer_output[2619] + last_layer_output[2620] + last_layer_output[2621] + last_layer_output[2622] + last_layer_output[2623] + last_layer_output[2624] + last_layer_output[2625] + last_layer_output[2626] + last_layer_output[2627] + last_layer_output[2628] + last_layer_output[2629] + last_layer_output[2630] + last_layer_output[2631] + last_layer_output[2632] + last_layer_output[2633] + last_layer_output[2634] + last_layer_output[2635] + last_layer_output[2636] + last_layer_output[2637] + last_layer_output[2638] + last_layer_output[2639] + last_layer_output[2640] + last_layer_output[2641] + last_layer_output[2642] + last_layer_output[2643] + last_layer_output[2644] + last_layer_output[2645] + last_layer_output[2646] + last_layer_output[2647] + last_layer_output[2648] + last_layer_output[2649] + last_layer_output[2650] + last_layer_output[2651] + last_layer_output[2652] + last_layer_output[2653] + last_layer_output[2654] + last_layer_output[2655] + last_layer_output[2656] + last_layer_output[2657] + last_layer_output[2658] + last_layer_output[2659] + last_layer_output[2660] + last_layer_output[2661] + last_layer_output[2662] + last_layer_output[2663] + last_layer_output[2664] + last_layer_output[2665] + last_layer_output[2666] + last_layer_output[2667] + last_layer_output[2668] + last_layer_output[2669] + last_layer_output[2670] + last_layer_output[2671] + last_layer_output[2672] + last_layer_output[2673] + last_layer_output[2674] + last_layer_output[2675] + last_layer_output[2676] + last_layer_output[2677] + last_layer_output[2678] + last_layer_output[2679] + last_layer_output[2680] + last_layer_output[2681] + last_layer_output[2682] + last_layer_output[2683] + last_layer_output[2684] + last_layer_output[2685] + last_layer_output[2686] + last_layer_output[2687] + last_layer_output[2688] + last_layer_output[2689] + last_layer_output[2690] + last_layer_output[2691] + last_layer_output[2692] + last_layer_output[2693] + last_layer_output[2694] + last_layer_output[2695] + last_layer_output[2696] + last_layer_output[2697] + last_layer_output[2698] + last_layer_output[2699] + last_layer_output[2700] + last_layer_output[2701] + last_layer_output[2702] + last_layer_output[2703] + last_layer_output[2704] + last_layer_output[2705] + last_layer_output[2706] + last_layer_output[2707] + last_layer_output[2708] + last_layer_output[2709] + last_layer_output[2710] + last_layer_output[2711] + last_layer_output[2712] + last_layer_output[2713] + last_layer_output[2714] + last_layer_output[2715] + last_layer_output[2716] + last_layer_output[2717] + last_layer_output[2718] + last_layer_output[2719] + last_layer_output[2720] + last_layer_output[2721] + last_layer_output[2722] + last_layer_output[2723] + last_layer_output[2724] + last_layer_output[2725] + last_layer_output[2726] + last_layer_output[2727] + last_layer_output[2728] + last_layer_output[2729] + last_layer_output[2730] + last_layer_output[2731] + last_layer_output[2732] + last_layer_output[2733] + last_layer_output[2734] + last_layer_output[2735] + last_layer_output[2736] + last_layer_output[2737] + last_layer_output[2738] + last_layer_output[2739] + last_layer_output[2740] + last_layer_output[2741] + last_layer_output[2742] + last_layer_output[2743] + last_layer_output[2744] + last_layer_output[2745] + last_layer_output[2746] + last_layer_output[2747] + last_layer_output[2748] + last_layer_output[2749] + last_layer_output[2750] + last_layer_output[2751] + last_layer_output[2752] + last_layer_output[2753] + last_layer_output[2754] + last_layer_output[2755] + last_layer_output[2756] + last_layer_output[2757] + last_layer_output[2758] + last_layer_output[2759] + last_layer_output[2760] + last_layer_output[2761] + last_layer_output[2762] + last_layer_output[2763] + last_layer_output[2764] + last_layer_output[2765] + last_layer_output[2766] + last_layer_output[2767] + last_layer_output[2768] + last_layer_output[2769] + last_layer_output[2770] + last_layer_output[2771] + last_layer_output[2772] + last_layer_output[2773] + last_layer_output[2774] + last_layer_output[2775] + last_layer_output[2776] + last_layer_output[2777] + last_layer_output[2778] + last_layer_output[2779] + last_layer_output[2780] + last_layer_output[2781] + last_layer_output[2782] + last_layer_output[2783] + last_layer_output[2784] + last_layer_output[2785] + last_layer_output[2786] + last_layer_output[2787] + last_layer_output[2788] + last_layer_output[2789] + last_layer_output[2790] + last_layer_output[2791] + last_layer_output[2792] + last_layer_output[2793] + last_layer_output[2794] + last_layer_output[2795] + last_layer_output[2796] + last_layer_output[2797] + last_layer_output[2798] + last_layer_output[2799] + last_layer_output[2800] + last_layer_output[2801] + last_layer_output[2802] + last_layer_output[2803] + last_layer_output[2804] + last_layer_output[2805] + last_layer_output[2806] + last_layer_output[2807] + last_layer_output[2808] + last_layer_output[2809] + last_layer_output[2810] + last_layer_output[2811] + last_layer_output[2812] + last_layer_output[2813] + last_layer_output[2814] + last_layer_output[2815] + last_layer_output[2816] + last_layer_output[2817] + last_layer_output[2818] + last_layer_output[2819] + last_layer_output[2820] + last_layer_output[2821] + last_layer_output[2822] + last_layer_output[2823] + last_layer_output[2824] + last_layer_output[2825] + last_layer_output[2826] + last_layer_output[2827] + last_layer_output[2828] + last_layer_output[2829] + last_layer_output[2830] + last_layer_output[2831] + last_layer_output[2832] + last_layer_output[2833] + last_layer_output[2834] + last_layer_output[2835] + last_layer_output[2836] + last_layer_output[2837] + last_layer_output[2838] + last_layer_output[2839] + last_layer_output[2840] + last_layer_output[2841] + last_layer_output[2842] + last_layer_output[2843] + last_layer_output[2844] + last_layer_output[2845] + last_layer_output[2846] + last_layer_output[2847] + last_layer_output[2848] + last_layer_output[2849] + last_layer_output[2850] + last_layer_output[2851] + last_layer_output[2852] + last_layer_output[2853] + last_layer_output[2854] + last_layer_output[2855] + last_layer_output[2856] + last_layer_output[2857] + last_layer_output[2858] + last_layer_output[2859] + last_layer_output[2860] + last_layer_output[2861] + last_layer_output[2862] + last_layer_output[2863] + last_layer_output[2864] + last_layer_output[2865] + last_layer_output[2866] + last_layer_output[2867] + last_layer_output[2868] + last_layer_output[2869] + last_layer_output[2870] + last_layer_output[2871] + last_layer_output[2872] + last_layer_output[2873] + last_layer_output[2874] + last_layer_output[2875] + last_layer_output[2876] + last_layer_output[2877] + last_layer_output[2878] + last_layer_output[2879] + last_layer_output[2880] + last_layer_output[2881] + last_layer_output[2882] + last_layer_output[2883] + last_layer_output[2884] + last_layer_output[2885] + last_layer_output[2886] + last_layer_output[2887] + last_layer_output[2888] + last_layer_output[2889] + last_layer_output[2890] + last_layer_output[2891] + last_layer_output[2892] + last_layer_output[2893] + last_layer_output[2894] + last_layer_output[2895] + last_layer_output[2896] + last_layer_output[2897] + last_layer_output[2898] + last_layer_output[2899] + last_layer_output[2900] + last_layer_output[2901] + last_layer_output[2902] + last_layer_output[2903] + last_layer_output[2904] + last_layer_output[2905] + last_layer_output[2906] + last_layer_output[2907] + last_layer_output[2908] + last_layer_output[2909] + last_layer_output[2910] + last_layer_output[2911] + last_layer_output[2912] + last_layer_output[2913] + last_layer_output[2914] + last_layer_output[2915] + last_layer_output[2916] + last_layer_output[2917] + last_layer_output[2918] + last_layer_output[2919] + last_layer_output[2920] + last_layer_output[2921] + last_layer_output[2922] + last_layer_output[2923] + last_layer_output[2924] + last_layer_output[2925] + last_layer_output[2926] + last_layer_output[2927] + last_layer_output[2928] + last_layer_output[2929] + last_layer_output[2930] + last_layer_output[2931] + last_layer_output[2932] + last_layer_output[2933] + last_layer_output[2934] + last_layer_output[2935] + last_layer_output[2936] + last_layer_output[2937] + last_layer_output[2938] + last_layer_output[2939] + last_layer_output[2940] + last_layer_output[2941] + last_layer_output[2942] + last_layer_output[2943] + last_layer_output[2944] + last_layer_output[2945] + last_layer_output[2946] + last_layer_output[2947] + last_layer_output[2948] + last_layer_output[2949] + last_layer_output[2950] + last_layer_output[2951] + last_layer_output[2952] + last_layer_output[2953] + last_layer_output[2954] + last_layer_output[2955] + last_layer_output[2956] + last_layer_output[2957] + last_layer_output[2958] + last_layer_output[2959] + last_layer_output[2960] + last_layer_output[2961] + last_layer_output[2962] + last_layer_output[2963] + last_layer_output[2964] + last_layer_output[2965] + last_layer_output[2966] + last_layer_output[2967] + last_layer_output[2968] + last_layer_output[2969] + last_layer_output[2970] + last_layer_output[2971] + last_layer_output[2972] + last_layer_output[2973] + last_layer_output[2974] + last_layer_output[2975] + last_layer_output[2976] + last_layer_output[2977] + last_layer_output[2978] + last_layer_output[2979] + last_layer_output[2980] + last_layer_output[2981] + last_layer_output[2982] + last_layer_output[2983] + last_layer_output[2984] + last_layer_output[2985] + last_layer_output[2986] + last_layer_output[2987] + last_layer_output[2988] + last_layer_output[2989] + last_layer_output[2990] + last_layer_output[2991] + last_layer_output[2992] + last_layer_output[2993] + last_layer_output[2994] + last_layer_output[2995] + last_layer_output[2996] + last_layer_output[2997] + last_layer_output[2998] + last_layer_output[2999] + last_layer_output[3000] + last_layer_output[3001] + last_layer_output[3002] + last_layer_output[3003] + last_layer_output[3004] + last_layer_output[3005] + last_layer_output[3006] + last_layer_output[3007] + last_layer_output[3008] + last_layer_output[3009] + last_layer_output[3010] + last_layer_output[3011] + last_layer_output[3012] + last_layer_output[3013] + last_layer_output[3014] + last_layer_output[3015] + last_layer_output[3016] + last_layer_output[3017] + last_layer_output[3018] + last_layer_output[3019] + last_layer_output[3020] + last_layer_output[3021] + last_layer_output[3022] + last_layer_output[3023] + last_layer_output[3024] + last_layer_output[3025] + last_layer_output[3026] + last_layer_output[3027] + last_layer_output[3028] + last_layer_output[3029] + last_layer_output[3030] + last_layer_output[3031] + last_layer_output[3032] + last_layer_output[3033] + last_layer_output[3034] + last_layer_output[3035] + last_layer_output[3036] + last_layer_output[3037] + last_layer_output[3038] + last_layer_output[3039] + last_layer_output[3040] + last_layer_output[3041] + last_layer_output[3042] + last_layer_output[3043] + last_layer_output[3044] + last_layer_output[3045] + last_layer_output[3046] + last_layer_output[3047] + last_layer_output[3048] + last_layer_output[3049] + last_layer_output[3050] + last_layer_output[3051] + last_layer_output[3052] + last_layer_output[3053] + last_layer_output[3054] + last_layer_output[3055] + last_layer_output[3056] + last_layer_output[3057] + last_layer_output[3058] + last_layer_output[3059] + last_layer_output[3060] + last_layer_output[3061] + last_layer_output[3062] + last_layer_output[3063] + last_layer_output[3064] + last_layer_output[3065] + last_layer_output[3066] + last_layer_output[3067] + last_layer_output[3068] + last_layer_output[3069] + last_layer_output[3070] + last_layer_output[3071] + last_layer_output[3072] + last_layer_output[3073] + last_layer_output[3074] + last_layer_output[3075] + last_layer_output[3076] + last_layer_output[3077] + last_layer_output[3078] + last_layer_output[3079] + last_layer_output[3080] + last_layer_output[3081] + last_layer_output[3082] + last_layer_output[3083] + last_layer_output[3084] + last_layer_output[3085] + last_layer_output[3086] + last_layer_output[3087] + last_layer_output[3088] + last_layer_output[3089] + last_layer_output[3090] + last_layer_output[3091] + last_layer_output[3092] + last_layer_output[3093] + last_layer_output[3094] + last_layer_output[3095] + last_layer_output[3096] + last_layer_output[3097] + last_layer_output[3098] + last_layer_output[3099] + last_layer_output[3100] + last_layer_output[3101] + last_layer_output[3102] + last_layer_output[3103] + last_layer_output[3104] + last_layer_output[3105] + last_layer_output[3106] + last_layer_output[3107] + last_layer_output[3108] + last_layer_output[3109] + last_layer_output[3110] + last_layer_output[3111] + last_layer_output[3112] + last_layer_output[3113] + last_layer_output[3114] + last_layer_output[3115] + last_layer_output[3116] + last_layer_output[3117] + last_layer_output[3118] + last_layer_output[3119] + last_layer_output[3120] + last_layer_output[3121] + last_layer_output[3122] + last_layer_output[3123] + last_layer_output[3124] + last_layer_output[3125] + last_layer_output[3126] + last_layer_output[3127] + last_layer_output[3128] + last_layer_output[3129] + last_layer_output[3130] + last_layer_output[3131] + last_layer_output[3132] + last_layer_output[3133] + last_layer_output[3134] + last_layer_output[3135] + last_layer_output[3136] + last_layer_output[3137] + last_layer_output[3138] + last_layer_output[3139] + last_layer_output[3140] + last_layer_output[3141] + last_layer_output[3142] + last_layer_output[3143] + last_layer_output[3144] + last_layer_output[3145] + last_layer_output[3146] + last_layer_output[3147] + last_layer_output[3148] + last_layer_output[3149] + last_layer_output[3150] + last_layer_output[3151] + last_layer_output[3152] + last_layer_output[3153] + last_layer_output[3154] + last_layer_output[3155] + last_layer_output[3156] + last_layer_output[3157] + last_layer_output[3158] + last_layer_output[3159] + last_layer_output[3160] + last_layer_output[3161] + last_layer_output[3162] + last_layer_output[3163] + last_layer_output[3164] + last_layer_output[3165] + last_layer_output[3166] + last_layer_output[3167] + last_layer_output[3168] + last_layer_output[3169] + last_layer_output[3170] + last_layer_output[3171] + last_layer_output[3172] + last_layer_output[3173] + last_layer_output[3174] + last_layer_output[3175] + last_layer_output[3176] + last_layer_output[3177] + last_layer_output[3178] + last_layer_output[3179] + last_layer_output[3180] + last_layer_output[3181] + last_layer_output[3182] + last_layer_output[3183] + last_layer_output[3184] + last_layer_output[3185] + last_layer_output[3186] + last_layer_output[3187] + last_layer_output[3188] + last_layer_output[3189] + last_layer_output[3190] + last_layer_output[3191] + last_layer_output[3192] + last_layer_output[3193] + last_layer_output[3194] + last_layer_output[3195] + last_layer_output[3196] + last_layer_output[3197] + last_layer_output[3198] + last_layer_output[3199] + last_layer_output[3200] + last_layer_output[3201] + last_layer_output[3202] + last_layer_output[3203] + last_layer_output[3204] + last_layer_output[3205] + last_layer_output[3206] + last_layer_output[3207] + last_layer_output[3208] + last_layer_output[3209] + last_layer_output[3210] + last_layer_output[3211] + last_layer_output[3212] + last_layer_output[3213] + last_layer_output[3214] + last_layer_output[3215] + last_layer_output[3216] + last_layer_output[3217] + last_layer_output[3218] + last_layer_output[3219] + last_layer_output[3220] + last_layer_output[3221] + last_layer_output[3222] + last_layer_output[3223] + last_layer_output[3224] + last_layer_output[3225] + last_layer_output[3226] + last_layer_output[3227] + last_layer_output[3228] + last_layer_output[3229] + last_layer_output[3230] + last_layer_output[3231] + last_layer_output[3232] + last_layer_output[3233] + last_layer_output[3234] + last_layer_output[3235] + last_layer_output[3236] + last_layer_output[3237] + last_layer_output[3238] + last_layer_output[3239] + last_layer_output[3240] + last_layer_output[3241] + last_layer_output[3242] + last_layer_output[3243] + last_layer_output[3244] + last_layer_output[3245] + last_layer_output[3246] + last_layer_output[3247] + last_layer_output[3248] + last_layer_output[3249] + last_layer_output[3250] + last_layer_output[3251] + last_layer_output[3252] + last_layer_output[3253] + last_layer_output[3254] + last_layer_output[3255] + last_layer_output[3256] + last_layer_output[3257] + last_layer_output[3258] + last_layer_output[3259] + last_layer_output[3260] + last_layer_output[3261] + last_layer_output[3262] + last_layer_output[3263] + last_layer_output[3264] + last_layer_output[3265] + last_layer_output[3266] + last_layer_output[3267] + last_layer_output[3268] + last_layer_output[3269] + last_layer_output[3270] + last_layer_output[3271] + last_layer_output[3272] + last_layer_output[3273] + last_layer_output[3274] + last_layer_output[3275] + last_layer_output[3276] + last_layer_output[3277] + last_layer_output[3278] + last_layer_output[3279] + last_layer_output[3280] + last_layer_output[3281] + last_layer_output[3282] + last_layer_output[3283] + last_layer_output[3284] + last_layer_output[3285] + last_layer_output[3286] + last_layer_output[3287] + last_layer_output[3288] + last_layer_output[3289] + last_layer_output[3290] + last_layer_output[3291] + last_layer_output[3292] + last_layer_output[3293] + last_layer_output[3294] + last_layer_output[3295] + last_layer_output[3296] + last_layer_output[3297] + last_layer_output[3298] + last_layer_output[3299] + last_layer_output[3300] + last_layer_output[3301] + last_layer_output[3302] + last_layer_output[3303] + last_layer_output[3304] + last_layer_output[3305] + last_layer_output[3306] + last_layer_output[3307] + last_layer_output[3308] + last_layer_output[3309] + last_layer_output[3310] + last_layer_output[3311] + last_layer_output[3312] + last_layer_output[3313] + last_layer_output[3314] + last_layer_output[3315] + last_layer_output[3316] + last_layer_output[3317] + last_layer_output[3318] + last_layer_output[3319] + last_layer_output[3320] + last_layer_output[3321] + last_layer_output[3322] + last_layer_output[3323] + last_layer_output[3324] + last_layer_output[3325] + last_layer_output[3326] + last_layer_output[3327] + last_layer_output[3328] + last_layer_output[3329] + last_layer_output[3330] + last_layer_output[3331] + last_layer_output[3332] + last_layer_output[3333] + last_layer_output[3334] + last_layer_output[3335] + last_layer_output[3336] + last_layer_output[3337] + last_layer_output[3338] + last_layer_output[3339] + last_layer_output[3340] + last_layer_output[3341] + last_layer_output[3342] + last_layer_output[3343] + last_layer_output[3344] + last_layer_output[3345] + last_layer_output[3346] + last_layer_output[3347] + last_layer_output[3348] + last_layer_output[3349] + last_layer_output[3350] + last_layer_output[3351] + last_layer_output[3352] + last_layer_output[3353] + last_layer_output[3354] + last_layer_output[3355] + last_layer_output[3356] + last_layer_output[3357] + last_layer_output[3358] + last_layer_output[3359] + last_layer_output[3360] + last_layer_output[3361] + last_layer_output[3362] + last_layer_output[3363] + last_layer_output[3364] + last_layer_output[3365] + last_layer_output[3366] + last_layer_output[3367] + last_layer_output[3368] + last_layer_output[3369] + last_layer_output[3370] + last_layer_output[3371] + last_layer_output[3372] + last_layer_output[3373] + last_layer_output[3374] + last_layer_output[3375] + last_layer_output[3376] + last_layer_output[3377] + last_layer_output[3378] + last_layer_output[3379] + last_layer_output[3380] + last_layer_output[3381] + last_layer_output[3382] + last_layer_output[3383] + last_layer_output[3384] + last_layer_output[3385] + last_layer_output[3386] + last_layer_output[3387] + last_layer_output[3388] + last_layer_output[3389] + last_layer_output[3390] + last_layer_output[3391] + last_layer_output[3392] + last_layer_output[3393] + last_layer_output[3394] + last_layer_output[3395] + last_layer_output[3396] + last_layer_output[3397] + last_layer_output[3398] + last_layer_output[3399] + last_layer_output[3400] + last_layer_output[3401] + last_layer_output[3402] + last_layer_output[3403] + last_layer_output[3404] + last_layer_output[3405] + last_layer_output[3406] + last_layer_output[3407] + last_layer_output[3408] + last_layer_output[3409] + last_layer_output[3410] + last_layer_output[3411] + last_layer_output[3412] + last_layer_output[3413] + last_layer_output[3414] + last_layer_output[3415] + last_layer_output[3416] + last_layer_output[3417] + last_layer_output[3418] + last_layer_output[3419] + last_layer_output[3420] + last_layer_output[3421] + last_layer_output[3422] + last_layer_output[3423] + last_layer_output[3424] + last_layer_output[3425] + last_layer_output[3426] + last_layer_output[3427] + last_layer_output[3428] + last_layer_output[3429] + last_layer_output[3430] + last_layer_output[3431] + last_layer_output[3432] + last_layer_output[3433] + last_layer_output[3434] + last_layer_output[3435] + last_layer_output[3436] + last_layer_output[3437] + last_layer_output[3438] + last_layer_output[3439] + last_layer_output[3440] + last_layer_output[3441] + last_layer_output[3442] + last_layer_output[3443] + last_layer_output[3444] + last_layer_output[3445] + last_layer_output[3446] + last_layer_output[3447] + last_layer_output[3448] + last_layer_output[3449] + last_layer_output[3450] + last_layer_output[3451] + last_layer_output[3452] + last_layer_output[3453] + last_layer_output[3454] + last_layer_output[3455] + last_layer_output[3456] + last_layer_output[3457] + last_layer_output[3458] + last_layer_output[3459] + last_layer_output[3460] + last_layer_output[3461] + last_layer_output[3462] + last_layer_output[3463] + last_layer_output[3464] + last_layer_output[3465] + last_layer_output[3466] + last_layer_output[3467] + last_layer_output[3468] + last_layer_output[3469] + last_layer_output[3470] + last_layer_output[3471] + last_layer_output[3472] + last_layer_output[3473] + last_layer_output[3474] + last_layer_output[3475] + last_layer_output[3476] + last_layer_output[3477] + last_layer_output[3478] + last_layer_output[3479] + last_layer_output[3480] + last_layer_output[3481] + last_layer_output[3482] + last_layer_output[3483] + last_layer_output[3484] + last_layer_output[3485] + last_layer_output[3486] + last_layer_output[3487] + last_layer_output[3488] + last_layer_output[3489] + last_layer_output[3490] + last_layer_output[3491] + last_layer_output[3492] + last_layer_output[3493] + last_layer_output[3494] + last_layer_output[3495] + last_layer_output[3496] + last_layer_output[3497] + last_layer_output[3498] + last_layer_output[3499] + last_layer_output[3500] + last_layer_output[3501] + last_layer_output[3502] + last_layer_output[3503] + last_layer_output[3504] + last_layer_output[3505] + last_layer_output[3506] + last_layer_output[3507] + last_layer_output[3508] + last_layer_output[3509] + last_layer_output[3510] + last_layer_output[3511] + last_layer_output[3512] + last_layer_output[3513] + last_layer_output[3514] + last_layer_output[3515] + last_layer_output[3516] + last_layer_output[3517] + last_layer_output[3518] + last_layer_output[3519] + last_layer_output[3520] + last_layer_output[3521] + last_layer_output[3522] + last_layer_output[3523] + last_layer_output[3524] + last_layer_output[3525] + last_layer_output[3526] + last_layer_output[3527] + last_layer_output[3528] + last_layer_output[3529] + last_layer_output[3530] + last_layer_output[3531] + last_layer_output[3532] + last_layer_output[3533] + last_layer_output[3534] + last_layer_output[3535] + last_layer_output[3536] + last_layer_output[3537] + last_layer_output[3538] + last_layer_output[3539] + last_layer_output[3540] + last_layer_output[3541] + last_layer_output[3542] + last_layer_output[3543] + last_layer_output[3544] + last_layer_output[3545] + last_layer_output[3546] + last_layer_output[3547] + last_layer_output[3548] + last_layer_output[3549] + last_layer_output[3550] + last_layer_output[3551] + last_layer_output[3552] + last_layer_output[3553] + last_layer_output[3554] + last_layer_output[3555] + last_layer_output[3556] + last_layer_output[3557] + last_layer_output[3558] + last_layer_output[3559] + last_layer_output[3560] + last_layer_output[3561] + last_layer_output[3562] + last_layer_output[3563] + last_layer_output[3564] + last_layer_output[3565] + last_layer_output[3566] + last_layer_output[3567] + last_layer_output[3568] + last_layer_output[3569] + last_layer_output[3570] + last_layer_output[3571] + last_layer_output[3572] + last_layer_output[3573] + last_layer_output[3574] + last_layer_output[3575] + last_layer_output[3576] + last_layer_output[3577] + last_layer_output[3578] + last_layer_output[3579] + last_layer_output[3580] + last_layer_output[3581] + last_layer_output[3582] + last_layer_output[3583] + last_layer_output[3584] + last_layer_output[3585] + last_layer_output[3586] + last_layer_output[3587] + last_layer_output[3588] + last_layer_output[3589] + last_layer_output[3590] + last_layer_output[3591] + last_layer_output[3592] + last_layer_output[3593] + last_layer_output[3594] + last_layer_output[3595] + last_layer_output[3596] + last_layer_output[3597] + last_layer_output[3598] + last_layer_output[3599];
      result[3] <= last_layer_output[3600] + last_layer_output[3601] + last_layer_output[3602] + last_layer_output[3603] + last_layer_output[3604] + last_layer_output[3605] + last_layer_output[3606] + last_layer_output[3607] + last_layer_output[3608] + last_layer_output[3609] + last_layer_output[3610] + last_layer_output[3611] + last_layer_output[3612] + last_layer_output[3613] + last_layer_output[3614] + last_layer_output[3615] + last_layer_output[3616] + last_layer_output[3617] + last_layer_output[3618] + last_layer_output[3619] + last_layer_output[3620] + last_layer_output[3621] + last_layer_output[3622] + last_layer_output[3623] + last_layer_output[3624] + last_layer_output[3625] + last_layer_output[3626] + last_layer_output[3627] + last_layer_output[3628] + last_layer_output[3629] + last_layer_output[3630] + last_layer_output[3631] + last_layer_output[3632] + last_layer_output[3633] + last_layer_output[3634] + last_layer_output[3635] + last_layer_output[3636] + last_layer_output[3637] + last_layer_output[3638] + last_layer_output[3639] + last_layer_output[3640] + last_layer_output[3641] + last_layer_output[3642] + last_layer_output[3643] + last_layer_output[3644] + last_layer_output[3645] + last_layer_output[3646] + last_layer_output[3647] + last_layer_output[3648] + last_layer_output[3649] + last_layer_output[3650] + last_layer_output[3651] + last_layer_output[3652] + last_layer_output[3653] + last_layer_output[3654] + last_layer_output[3655] + last_layer_output[3656] + last_layer_output[3657] + last_layer_output[3658] + last_layer_output[3659] + last_layer_output[3660] + last_layer_output[3661] + last_layer_output[3662] + last_layer_output[3663] + last_layer_output[3664] + last_layer_output[3665] + last_layer_output[3666] + last_layer_output[3667] + last_layer_output[3668] + last_layer_output[3669] + last_layer_output[3670] + last_layer_output[3671] + last_layer_output[3672] + last_layer_output[3673] + last_layer_output[3674] + last_layer_output[3675] + last_layer_output[3676] + last_layer_output[3677] + last_layer_output[3678] + last_layer_output[3679] + last_layer_output[3680] + last_layer_output[3681] + last_layer_output[3682] + last_layer_output[3683] + last_layer_output[3684] + last_layer_output[3685] + last_layer_output[3686] + last_layer_output[3687] + last_layer_output[3688] + last_layer_output[3689] + last_layer_output[3690] + last_layer_output[3691] + last_layer_output[3692] + last_layer_output[3693] + last_layer_output[3694] + last_layer_output[3695] + last_layer_output[3696] + last_layer_output[3697] + last_layer_output[3698] + last_layer_output[3699] + last_layer_output[3700] + last_layer_output[3701] + last_layer_output[3702] + last_layer_output[3703] + last_layer_output[3704] + last_layer_output[3705] + last_layer_output[3706] + last_layer_output[3707] + last_layer_output[3708] + last_layer_output[3709] + last_layer_output[3710] + last_layer_output[3711] + last_layer_output[3712] + last_layer_output[3713] + last_layer_output[3714] + last_layer_output[3715] + last_layer_output[3716] + last_layer_output[3717] + last_layer_output[3718] + last_layer_output[3719] + last_layer_output[3720] + last_layer_output[3721] + last_layer_output[3722] + last_layer_output[3723] + last_layer_output[3724] + last_layer_output[3725] + last_layer_output[3726] + last_layer_output[3727] + last_layer_output[3728] + last_layer_output[3729] + last_layer_output[3730] + last_layer_output[3731] + last_layer_output[3732] + last_layer_output[3733] + last_layer_output[3734] + last_layer_output[3735] + last_layer_output[3736] + last_layer_output[3737] + last_layer_output[3738] + last_layer_output[3739] + last_layer_output[3740] + last_layer_output[3741] + last_layer_output[3742] + last_layer_output[3743] + last_layer_output[3744] + last_layer_output[3745] + last_layer_output[3746] + last_layer_output[3747] + last_layer_output[3748] + last_layer_output[3749] + last_layer_output[3750] + last_layer_output[3751] + last_layer_output[3752] + last_layer_output[3753] + last_layer_output[3754] + last_layer_output[3755] + last_layer_output[3756] + last_layer_output[3757] + last_layer_output[3758] + last_layer_output[3759] + last_layer_output[3760] + last_layer_output[3761] + last_layer_output[3762] + last_layer_output[3763] + last_layer_output[3764] + last_layer_output[3765] + last_layer_output[3766] + last_layer_output[3767] + last_layer_output[3768] + last_layer_output[3769] + last_layer_output[3770] + last_layer_output[3771] + last_layer_output[3772] + last_layer_output[3773] + last_layer_output[3774] + last_layer_output[3775] + last_layer_output[3776] + last_layer_output[3777] + last_layer_output[3778] + last_layer_output[3779] + last_layer_output[3780] + last_layer_output[3781] + last_layer_output[3782] + last_layer_output[3783] + last_layer_output[3784] + last_layer_output[3785] + last_layer_output[3786] + last_layer_output[3787] + last_layer_output[3788] + last_layer_output[3789] + last_layer_output[3790] + last_layer_output[3791] + last_layer_output[3792] + last_layer_output[3793] + last_layer_output[3794] + last_layer_output[3795] + last_layer_output[3796] + last_layer_output[3797] + last_layer_output[3798] + last_layer_output[3799] + last_layer_output[3800] + last_layer_output[3801] + last_layer_output[3802] + last_layer_output[3803] + last_layer_output[3804] + last_layer_output[3805] + last_layer_output[3806] + last_layer_output[3807] + last_layer_output[3808] + last_layer_output[3809] + last_layer_output[3810] + last_layer_output[3811] + last_layer_output[3812] + last_layer_output[3813] + last_layer_output[3814] + last_layer_output[3815] + last_layer_output[3816] + last_layer_output[3817] + last_layer_output[3818] + last_layer_output[3819] + last_layer_output[3820] + last_layer_output[3821] + last_layer_output[3822] + last_layer_output[3823] + last_layer_output[3824] + last_layer_output[3825] + last_layer_output[3826] + last_layer_output[3827] + last_layer_output[3828] + last_layer_output[3829] + last_layer_output[3830] + last_layer_output[3831] + last_layer_output[3832] + last_layer_output[3833] + last_layer_output[3834] + last_layer_output[3835] + last_layer_output[3836] + last_layer_output[3837] + last_layer_output[3838] + last_layer_output[3839] + last_layer_output[3840] + last_layer_output[3841] + last_layer_output[3842] + last_layer_output[3843] + last_layer_output[3844] + last_layer_output[3845] + last_layer_output[3846] + last_layer_output[3847] + last_layer_output[3848] + last_layer_output[3849] + last_layer_output[3850] + last_layer_output[3851] + last_layer_output[3852] + last_layer_output[3853] + last_layer_output[3854] + last_layer_output[3855] + last_layer_output[3856] + last_layer_output[3857] + last_layer_output[3858] + last_layer_output[3859] + last_layer_output[3860] + last_layer_output[3861] + last_layer_output[3862] + last_layer_output[3863] + last_layer_output[3864] + last_layer_output[3865] + last_layer_output[3866] + last_layer_output[3867] + last_layer_output[3868] + last_layer_output[3869] + last_layer_output[3870] + last_layer_output[3871] + last_layer_output[3872] + last_layer_output[3873] + last_layer_output[3874] + last_layer_output[3875] + last_layer_output[3876] + last_layer_output[3877] + last_layer_output[3878] + last_layer_output[3879] + last_layer_output[3880] + last_layer_output[3881] + last_layer_output[3882] + last_layer_output[3883] + last_layer_output[3884] + last_layer_output[3885] + last_layer_output[3886] + last_layer_output[3887] + last_layer_output[3888] + last_layer_output[3889] + last_layer_output[3890] + last_layer_output[3891] + last_layer_output[3892] + last_layer_output[3893] + last_layer_output[3894] + last_layer_output[3895] + last_layer_output[3896] + last_layer_output[3897] + last_layer_output[3898] + last_layer_output[3899] + last_layer_output[3900] + last_layer_output[3901] + last_layer_output[3902] + last_layer_output[3903] + last_layer_output[3904] + last_layer_output[3905] + last_layer_output[3906] + last_layer_output[3907] + last_layer_output[3908] + last_layer_output[3909] + last_layer_output[3910] + last_layer_output[3911] + last_layer_output[3912] + last_layer_output[3913] + last_layer_output[3914] + last_layer_output[3915] + last_layer_output[3916] + last_layer_output[3917] + last_layer_output[3918] + last_layer_output[3919] + last_layer_output[3920] + last_layer_output[3921] + last_layer_output[3922] + last_layer_output[3923] + last_layer_output[3924] + last_layer_output[3925] + last_layer_output[3926] + last_layer_output[3927] + last_layer_output[3928] + last_layer_output[3929] + last_layer_output[3930] + last_layer_output[3931] + last_layer_output[3932] + last_layer_output[3933] + last_layer_output[3934] + last_layer_output[3935] + last_layer_output[3936] + last_layer_output[3937] + last_layer_output[3938] + last_layer_output[3939] + last_layer_output[3940] + last_layer_output[3941] + last_layer_output[3942] + last_layer_output[3943] + last_layer_output[3944] + last_layer_output[3945] + last_layer_output[3946] + last_layer_output[3947] + last_layer_output[3948] + last_layer_output[3949] + last_layer_output[3950] + last_layer_output[3951] + last_layer_output[3952] + last_layer_output[3953] + last_layer_output[3954] + last_layer_output[3955] + last_layer_output[3956] + last_layer_output[3957] + last_layer_output[3958] + last_layer_output[3959] + last_layer_output[3960] + last_layer_output[3961] + last_layer_output[3962] + last_layer_output[3963] + last_layer_output[3964] + last_layer_output[3965] + last_layer_output[3966] + last_layer_output[3967] + last_layer_output[3968] + last_layer_output[3969] + last_layer_output[3970] + last_layer_output[3971] + last_layer_output[3972] + last_layer_output[3973] + last_layer_output[3974] + last_layer_output[3975] + last_layer_output[3976] + last_layer_output[3977] + last_layer_output[3978] + last_layer_output[3979] + last_layer_output[3980] + last_layer_output[3981] + last_layer_output[3982] + last_layer_output[3983] + last_layer_output[3984] + last_layer_output[3985] + last_layer_output[3986] + last_layer_output[3987] + last_layer_output[3988] + last_layer_output[3989] + last_layer_output[3990] + last_layer_output[3991] + last_layer_output[3992] + last_layer_output[3993] + last_layer_output[3994] + last_layer_output[3995] + last_layer_output[3996] + last_layer_output[3997] + last_layer_output[3998] + last_layer_output[3999] + last_layer_output[4000] + last_layer_output[4001] + last_layer_output[4002] + last_layer_output[4003] + last_layer_output[4004] + last_layer_output[4005] + last_layer_output[4006] + last_layer_output[4007] + last_layer_output[4008] + last_layer_output[4009] + last_layer_output[4010] + last_layer_output[4011] + last_layer_output[4012] + last_layer_output[4013] + last_layer_output[4014] + last_layer_output[4015] + last_layer_output[4016] + last_layer_output[4017] + last_layer_output[4018] + last_layer_output[4019] + last_layer_output[4020] + last_layer_output[4021] + last_layer_output[4022] + last_layer_output[4023] + last_layer_output[4024] + last_layer_output[4025] + last_layer_output[4026] + last_layer_output[4027] + last_layer_output[4028] + last_layer_output[4029] + last_layer_output[4030] + last_layer_output[4031] + last_layer_output[4032] + last_layer_output[4033] + last_layer_output[4034] + last_layer_output[4035] + last_layer_output[4036] + last_layer_output[4037] + last_layer_output[4038] + last_layer_output[4039] + last_layer_output[4040] + last_layer_output[4041] + last_layer_output[4042] + last_layer_output[4043] + last_layer_output[4044] + last_layer_output[4045] + last_layer_output[4046] + last_layer_output[4047] + last_layer_output[4048] + last_layer_output[4049] + last_layer_output[4050] + last_layer_output[4051] + last_layer_output[4052] + last_layer_output[4053] + last_layer_output[4054] + last_layer_output[4055] + last_layer_output[4056] + last_layer_output[4057] + last_layer_output[4058] + last_layer_output[4059] + last_layer_output[4060] + last_layer_output[4061] + last_layer_output[4062] + last_layer_output[4063] + last_layer_output[4064] + last_layer_output[4065] + last_layer_output[4066] + last_layer_output[4067] + last_layer_output[4068] + last_layer_output[4069] + last_layer_output[4070] + last_layer_output[4071] + last_layer_output[4072] + last_layer_output[4073] + last_layer_output[4074] + last_layer_output[4075] + last_layer_output[4076] + last_layer_output[4077] + last_layer_output[4078] + last_layer_output[4079] + last_layer_output[4080] + last_layer_output[4081] + last_layer_output[4082] + last_layer_output[4083] + last_layer_output[4084] + last_layer_output[4085] + last_layer_output[4086] + last_layer_output[4087] + last_layer_output[4088] + last_layer_output[4089] + last_layer_output[4090] + last_layer_output[4091] + last_layer_output[4092] + last_layer_output[4093] + last_layer_output[4094] + last_layer_output[4095] + last_layer_output[4096] + last_layer_output[4097] + last_layer_output[4098] + last_layer_output[4099] + last_layer_output[4100] + last_layer_output[4101] + last_layer_output[4102] + last_layer_output[4103] + last_layer_output[4104] + last_layer_output[4105] + last_layer_output[4106] + last_layer_output[4107] + last_layer_output[4108] + last_layer_output[4109] + last_layer_output[4110] + last_layer_output[4111] + last_layer_output[4112] + last_layer_output[4113] + last_layer_output[4114] + last_layer_output[4115] + last_layer_output[4116] + last_layer_output[4117] + last_layer_output[4118] + last_layer_output[4119] + last_layer_output[4120] + last_layer_output[4121] + last_layer_output[4122] + last_layer_output[4123] + last_layer_output[4124] + last_layer_output[4125] + last_layer_output[4126] + last_layer_output[4127] + last_layer_output[4128] + last_layer_output[4129] + last_layer_output[4130] + last_layer_output[4131] + last_layer_output[4132] + last_layer_output[4133] + last_layer_output[4134] + last_layer_output[4135] + last_layer_output[4136] + last_layer_output[4137] + last_layer_output[4138] + last_layer_output[4139] + last_layer_output[4140] + last_layer_output[4141] + last_layer_output[4142] + last_layer_output[4143] + last_layer_output[4144] + last_layer_output[4145] + last_layer_output[4146] + last_layer_output[4147] + last_layer_output[4148] + last_layer_output[4149] + last_layer_output[4150] + last_layer_output[4151] + last_layer_output[4152] + last_layer_output[4153] + last_layer_output[4154] + last_layer_output[4155] + last_layer_output[4156] + last_layer_output[4157] + last_layer_output[4158] + last_layer_output[4159] + last_layer_output[4160] + last_layer_output[4161] + last_layer_output[4162] + last_layer_output[4163] + last_layer_output[4164] + last_layer_output[4165] + last_layer_output[4166] + last_layer_output[4167] + last_layer_output[4168] + last_layer_output[4169] + last_layer_output[4170] + last_layer_output[4171] + last_layer_output[4172] + last_layer_output[4173] + last_layer_output[4174] + last_layer_output[4175] + last_layer_output[4176] + last_layer_output[4177] + last_layer_output[4178] + last_layer_output[4179] + last_layer_output[4180] + last_layer_output[4181] + last_layer_output[4182] + last_layer_output[4183] + last_layer_output[4184] + last_layer_output[4185] + last_layer_output[4186] + last_layer_output[4187] + last_layer_output[4188] + last_layer_output[4189] + last_layer_output[4190] + last_layer_output[4191] + last_layer_output[4192] + last_layer_output[4193] + last_layer_output[4194] + last_layer_output[4195] + last_layer_output[4196] + last_layer_output[4197] + last_layer_output[4198] + last_layer_output[4199] + last_layer_output[4200] + last_layer_output[4201] + last_layer_output[4202] + last_layer_output[4203] + last_layer_output[4204] + last_layer_output[4205] + last_layer_output[4206] + last_layer_output[4207] + last_layer_output[4208] + last_layer_output[4209] + last_layer_output[4210] + last_layer_output[4211] + last_layer_output[4212] + last_layer_output[4213] + last_layer_output[4214] + last_layer_output[4215] + last_layer_output[4216] + last_layer_output[4217] + last_layer_output[4218] + last_layer_output[4219] + last_layer_output[4220] + last_layer_output[4221] + last_layer_output[4222] + last_layer_output[4223] + last_layer_output[4224] + last_layer_output[4225] + last_layer_output[4226] + last_layer_output[4227] + last_layer_output[4228] + last_layer_output[4229] + last_layer_output[4230] + last_layer_output[4231] + last_layer_output[4232] + last_layer_output[4233] + last_layer_output[4234] + last_layer_output[4235] + last_layer_output[4236] + last_layer_output[4237] + last_layer_output[4238] + last_layer_output[4239] + last_layer_output[4240] + last_layer_output[4241] + last_layer_output[4242] + last_layer_output[4243] + last_layer_output[4244] + last_layer_output[4245] + last_layer_output[4246] + last_layer_output[4247] + last_layer_output[4248] + last_layer_output[4249] + last_layer_output[4250] + last_layer_output[4251] + last_layer_output[4252] + last_layer_output[4253] + last_layer_output[4254] + last_layer_output[4255] + last_layer_output[4256] + last_layer_output[4257] + last_layer_output[4258] + last_layer_output[4259] + last_layer_output[4260] + last_layer_output[4261] + last_layer_output[4262] + last_layer_output[4263] + last_layer_output[4264] + last_layer_output[4265] + last_layer_output[4266] + last_layer_output[4267] + last_layer_output[4268] + last_layer_output[4269] + last_layer_output[4270] + last_layer_output[4271] + last_layer_output[4272] + last_layer_output[4273] + last_layer_output[4274] + last_layer_output[4275] + last_layer_output[4276] + last_layer_output[4277] + last_layer_output[4278] + last_layer_output[4279] + last_layer_output[4280] + last_layer_output[4281] + last_layer_output[4282] + last_layer_output[4283] + last_layer_output[4284] + last_layer_output[4285] + last_layer_output[4286] + last_layer_output[4287] + last_layer_output[4288] + last_layer_output[4289] + last_layer_output[4290] + last_layer_output[4291] + last_layer_output[4292] + last_layer_output[4293] + last_layer_output[4294] + last_layer_output[4295] + last_layer_output[4296] + last_layer_output[4297] + last_layer_output[4298] + last_layer_output[4299] + last_layer_output[4300] + last_layer_output[4301] + last_layer_output[4302] + last_layer_output[4303] + last_layer_output[4304] + last_layer_output[4305] + last_layer_output[4306] + last_layer_output[4307] + last_layer_output[4308] + last_layer_output[4309] + last_layer_output[4310] + last_layer_output[4311] + last_layer_output[4312] + last_layer_output[4313] + last_layer_output[4314] + last_layer_output[4315] + last_layer_output[4316] + last_layer_output[4317] + last_layer_output[4318] + last_layer_output[4319] + last_layer_output[4320] + last_layer_output[4321] + last_layer_output[4322] + last_layer_output[4323] + last_layer_output[4324] + last_layer_output[4325] + last_layer_output[4326] + last_layer_output[4327] + last_layer_output[4328] + last_layer_output[4329] + last_layer_output[4330] + last_layer_output[4331] + last_layer_output[4332] + last_layer_output[4333] + last_layer_output[4334] + last_layer_output[4335] + last_layer_output[4336] + last_layer_output[4337] + last_layer_output[4338] + last_layer_output[4339] + last_layer_output[4340] + last_layer_output[4341] + last_layer_output[4342] + last_layer_output[4343] + last_layer_output[4344] + last_layer_output[4345] + last_layer_output[4346] + last_layer_output[4347] + last_layer_output[4348] + last_layer_output[4349] + last_layer_output[4350] + last_layer_output[4351] + last_layer_output[4352] + last_layer_output[4353] + last_layer_output[4354] + last_layer_output[4355] + last_layer_output[4356] + last_layer_output[4357] + last_layer_output[4358] + last_layer_output[4359] + last_layer_output[4360] + last_layer_output[4361] + last_layer_output[4362] + last_layer_output[4363] + last_layer_output[4364] + last_layer_output[4365] + last_layer_output[4366] + last_layer_output[4367] + last_layer_output[4368] + last_layer_output[4369] + last_layer_output[4370] + last_layer_output[4371] + last_layer_output[4372] + last_layer_output[4373] + last_layer_output[4374] + last_layer_output[4375] + last_layer_output[4376] + last_layer_output[4377] + last_layer_output[4378] + last_layer_output[4379] + last_layer_output[4380] + last_layer_output[4381] + last_layer_output[4382] + last_layer_output[4383] + last_layer_output[4384] + last_layer_output[4385] + last_layer_output[4386] + last_layer_output[4387] + last_layer_output[4388] + last_layer_output[4389] + last_layer_output[4390] + last_layer_output[4391] + last_layer_output[4392] + last_layer_output[4393] + last_layer_output[4394] + last_layer_output[4395] + last_layer_output[4396] + last_layer_output[4397] + last_layer_output[4398] + last_layer_output[4399] + last_layer_output[4400] + last_layer_output[4401] + last_layer_output[4402] + last_layer_output[4403] + last_layer_output[4404] + last_layer_output[4405] + last_layer_output[4406] + last_layer_output[4407] + last_layer_output[4408] + last_layer_output[4409] + last_layer_output[4410] + last_layer_output[4411] + last_layer_output[4412] + last_layer_output[4413] + last_layer_output[4414] + last_layer_output[4415] + last_layer_output[4416] + last_layer_output[4417] + last_layer_output[4418] + last_layer_output[4419] + last_layer_output[4420] + last_layer_output[4421] + last_layer_output[4422] + last_layer_output[4423] + last_layer_output[4424] + last_layer_output[4425] + last_layer_output[4426] + last_layer_output[4427] + last_layer_output[4428] + last_layer_output[4429] + last_layer_output[4430] + last_layer_output[4431] + last_layer_output[4432] + last_layer_output[4433] + last_layer_output[4434] + last_layer_output[4435] + last_layer_output[4436] + last_layer_output[4437] + last_layer_output[4438] + last_layer_output[4439] + last_layer_output[4440] + last_layer_output[4441] + last_layer_output[4442] + last_layer_output[4443] + last_layer_output[4444] + last_layer_output[4445] + last_layer_output[4446] + last_layer_output[4447] + last_layer_output[4448] + last_layer_output[4449] + last_layer_output[4450] + last_layer_output[4451] + last_layer_output[4452] + last_layer_output[4453] + last_layer_output[4454] + last_layer_output[4455] + last_layer_output[4456] + last_layer_output[4457] + last_layer_output[4458] + last_layer_output[4459] + last_layer_output[4460] + last_layer_output[4461] + last_layer_output[4462] + last_layer_output[4463] + last_layer_output[4464] + last_layer_output[4465] + last_layer_output[4466] + last_layer_output[4467] + last_layer_output[4468] + last_layer_output[4469] + last_layer_output[4470] + last_layer_output[4471] + last_layer_output[4472] + last_layer_output[4473] + last_layer_output[4474] + last_layer_output[4475] + last_layer_output[4476] + last_layer_output[4477] + last_layer_output[4478] + last_layer_output[4479] + last_layer_output[4480] + last_layer_output[4481] + last_layer_output[4482] + last_layer_output[4483] + last_layer_output[4484] + last_layer_output[4485] + last_layer_output[4486] + last_layer_output[4487] + last_layer_output[4488] + last_layer_output[4489] + last_layer_output[4490] + last_layer_output[4491] + last_layer_output[4492] + last_layer_output[4493] + last_layer_output[4494] + last_layer_output[4495] + last_layer_output[4496] + last_layer_output[4497] + last_layer_output[4498] + last_layer_output[4499] + last_layer_output[4500] + last_layer_output[4501] + last_layer_output[4502] + last_layer_output[4503] + last_layer_output[4504] + last_layer_output[4505] + last_layer_output[4506] + last_layer_output[4507] + last_layer_output[4508] + last_layer_output[4509] + last_layer_output[4510] + last_layer_output[4511] + last_layer_output[4512] + last_layer_output[4513] + last_layer_output[4514] + last_layer_output[4515] + last_layer_output[4516] + last_layer_output[4517] + last_layer_output[4518] + last_layer_output[4519] + last_layer_output[4520] + last_layer_output[4521] + last_layer_output[4522] + last_layer_output[4523] + last_layer_output[4524] + last_layer_output[4525] + last_layer_output[4526] + last_layer_output[4527] + last_layer_output[4528] + last_layer_output[4529] + last_layer_output[4530] + last_layer_output[4531] + last_layer_output[4532] + last_layer_output[4533] + last_layer_output[4534] + last_layer_output[4535] + last_layer_output[4536] + last_layer_output[4537] + last_layer_output[4538] + last_layer_output[4539] + last_layer_output[4540] + last_layer_output[4541] + last_layer_output[4542] + last_layer_output[4543] + last_layer_output[4544] + last_layer_output[4545] + last_layer_output[4546] + last_layer_output[4547] + last_layer_output[4548] + last_layer_output[4549] + last_layer_output[4550] + last_layer_output[4551] + last_layer_output[4552] + last_layer_output[4553] + last_layer_output[4554] + last_layer_output[4555] + last_layer_output[4556] + last_layer_output[4557] + last_layer_output[4558] + last_layer_output[4559] + last_layer_output[4560] + last_layer_output[4561] + last_layer_output[4562] + last_layer_output[4563] + last_layer_output[4564] + last_layer_output[4565] + last_layer_output[4566] + last_layer_output[4567] + last_layer_output[4568] + last_layer_output[4569] + last_layer_output[4570] + last_layer_output[4571] + last_layer_output[4572] + last_layer_output[4573] + last_layer_output[4574] + last_layer_output[4575] + last_layer_output[4576] + last_layer_output[4577] + last_layer_output[4578] + last_layer_output[4579] + last_layer_output[4580] + last_layer_output[4581] + last_layer_output[4582] + last_layer_output[4583] + last_layer_output[4584] + last_layer_output[4585] + last_layer_output[4586] + last_layer_output[4587] + last_layer_output[4588] + last_layer_output[4589] + last_layer_output[4590] + last_layer_output[4591] + last_layer_output[4592] + last_layer_output[4593] + last_layer_output[4594] + last_layer_output[4595] + last_layer_output[4596] + last_layer_output[4597] + last_layer_output[4598] + last_layer_output[4599] + last_layer_output[4600] + last_layer_output[4601] + last_layer_output[4602] + last_layer_output[4603] + last_layer_output[4604] + last_layer_output[4605] + last_layer_output[4606] + last_layer_output[4607] + last_layer_output[4608] + last_layer_output[4609] + last_layer_output[4610] + last_layer_output[4611] + last_layer_output[4612] + last_layer_output[4613] + last_layer_output[4614] + last_layer_output[4615] + last_layer_output[4616] + last_layer_output[4617] + last_layer_output[4618] + last_layer_output[4619] + last_layer_output[4620] + last_layer_output[4621] + last_layer_output[4622] + last_layer_output[4623] + last_layer_output[4624] + last_layer_output[4625] + last_layer_output[4626] + last_layer_output[4627] + last_layer_output[4628] + last_layer_output[4629] + last_layer_output[4630] + last_layer_output[4631] + last_layer_output[4632] + last_layer_output[4633] + last_layer_output[4634] + last_layer_output[4635] + last_layer_output[4636] + last_layer_output[4637] + last_layer_output[4638] + last_layer_output[4639] + last_layer_output[4640] + last_layer_output[4641] + last_layer_output[4642] + last_layer_output[4643] + last_layer_output[4644] + last_layer_output[4645] + last_layer_output[4646] + last_layer_output[4647] + last_layer_output[4648] + last_layer_output[4649] + last_layer_output[4650] + last_layer_output[4651] + last_layer_output[4652] + last_layer_output[4653] + last_layer_output[4654] + last_layer_output[4655] + last_layer_output[4656] + last_layer_output[4657] + last_layer_output[4658] + last_layer_output[4659] + last_layer_output[4660] + last_layer_output[4661] + last_layer_output[4662] + last_layer_output[4663] + last_layer_output[4664] + last_layer_output[4665] + last_layer_output[4666] + last_layer_output[4667] + last_layer_output[4668] + last_layer_output[4669] + last_layer_output[4670] + last_layer_output[4671] + last_layer_output[4672] + last_layer_output[4673] + last_layer_output[4674] + last_layer_output[4675] + last_layer_output[4676] + last_layer_output[4677] + last_layer_output[4678] + last_layer_output[4679] + last_layer_output[4680] + last_layer_output[4681] + last_layer_output[4682] + last_layer_output[4683] + last_layer_output[4684] + last_layer_output[4685] + last_layer_output[4686] + last_layer_output[4687] + last_layer_output[4688] + last_layer_output[4689] + last_layer_output[4690] + last_layer_output[4691] + last_layer_output[4692] + last_layer_output[4693] + last_layer_output[4694] + last_layer_output[4695] + last_layer_output[4696] + last_layer_output[4697] + last_layer_output[4698] + last_layer_output[4699] + last_layer_output[4700] + last_layer_output[4701] + last_layer_output[4702] + last_layer_output[4703] + last_layer_output[4704] + last_layer_output[4705] + last_layer_output[4706] + last_layer_output[4707] + last_layer_output[4708] + last_layer_output[4709] + last_layer_output[4710] + last_layer_output[4711] + last_layer_output[4712] + last_layer_output[4713] + last_layer_output[4714] + last_layer_output[4715] + last_layer_output[4716] + last_layer_output[4717] + last_layer_output[4718] + last_layer_output[4719] + last_layer_output[4720] + last_layer_output[4721] + last_layer_output[4722] + last_layer_output[4723] + last_layer_output[4724] + last_layer_output[4725] + last_layer_output[4726] + last_layer_output[4727] + last_layer_output[4728] + last_layer_output[4729] + last_layer_output[4730] + last_layer_output[4731] + last_layer_output[4732] + last_layer_output[4733] + last_layer_output[4734] + last_layer_output[4735] + last_layer_output[4736] + last_layer_output[4737] + last_layer_output[4738] + last_layer_output[4739] + last_layer_output[4740] + last_layer_output[4741] + last_layer_output[4742] + last_layer_output[4743] + last_layer_output[4744] + last_layer_output[4745] + last_layer_output[4746] + last_layer_output[4747] + last_layer_output[4748] + last_layer_output[4749] + last_layer_output[4750] + last_layer_output[4751] + last_layer_output[4752] + last_layer_output[4753] + last_layer_output[4754] + last_layer_output[4755] + last_layer_output[4756] + last_layer_output[4757] + last_layer_output[4758] + last_layer_output[4759] + last_layer_output[4760] + last_layer_output[4761] + last_layer_output[4762] + last_layer_output[4763] + last_layer_output[4764] + last_layer_output[4765] + last_layer_output[4766] + last_layer_output[4767] + last_layer_output[4768] + last_layer_output[4769] + last_layer_output[4770] + last_layer_output[4771] + last_layer_output[4772] + last_layer_output[4773] + last_layer_output[4774] + last_layer_output[4775] + last_layer_output[4776] + last_layer_output[4777] + last_layer_output[4778] + last_layer_output[4779] + last_layer_output[4780] + last_layer_output[4781] + last_layer_output[4782] + last_layer_output[4783] + last_layer_output[4784] + last_layer_output[4785] + last_layer_output[4786] + last_layer_output[4787] + last_layer_output[4788] + last_layer_output[4789] + last_layer_output[4790] + last_layer_output[4791] + last_layer_output[4792] + last_layer_output[4793] + last_layer_output[4794] + last_layer_output[4795] + last_layer_output[4796] + last_layer_output[4797] + last_layer_output[4798] + last_layer_output[4799];
      result[4] <= last_layer_output[4800] + last_layer_output[4801] + last_layer_output[4802] + last_layer_output[4803] + last_layer_output[4804] + last_layer_output[4805] + last_layer_output[4806] + last_layer_output[4807] + last_layer_output[4808] + last_layer_output[4809] + last_layer_output[4810] + last_layer_output[4811] + last_layer_output[4812] + last_layer_output[4813] + last_layer_output[4814] + last_layer_output[4815] + last_layer_output[4816] + last_layer_output[4817] + last_layer_output[4818] + last_layer_output[4819] + last_layer_output[4820] + last_layer_output[4821] + last_layer_output[4822] + last_layer_output[4823] + last_layer_output[4824] + last_layer_output[4825] + last_layer_output[4826] + last_layer_output[4827] + last_layer_output[4828] + last_layer_output[4829] + last_layer_output[4830] + last_layer_output[4831] + last_layer_output[4832] + last_layer_output[4833] + last_layer_output[4834] + last_layer_output[4835] + last_layer_output[4836] + last_layer_output[4837] + last_layer_output[4838] + last_layer_output[4839] + last_layer_output[4840] + last_layer_output[4841] + last_layer_output[4842] + last_layer_output[4843] + last_layer_output[4844] + last_layer_output[4845] + last_layer_output[4846] + last_layer_output[4847] + last_layer_output[4848] + last_layer_output[4849] + last_layer_output[4850] + last_layer_output[4851] + last_layer_output[4852] + last_layer_output[4853] + last_layer_output[4854] + last_layer_output[4855] + last_layer_output[4856] + last_layer_output[4857] + last_layer_output[4858] + last_layer_output[4859] + last_layer_output[4860] + last_layer_output[4861] + last_layer_output[4862] + last_layer_output[4863] + last_layer_output[4864] + last_layer_output[4865] + last_layer_output[4866] + last_layer_output[4867] + last_layer_output[4868] + last_layer_output[4869] + last_layer_output[4870] + last_layer_output[4871] + last_layer_output[4872] + last_layer_output[4873] + last_layer_output[4874] + last_layer_output[4875] + last_layer_output[4876] + last_layer_output[4877] + last_layer_output[4878] + last_layer_output[4879] + last_layer_output[4880] + last_layer_output[4881] + last_layer_output[4882] + last_layer_output[4883] + last_layer_output[4884] + last_layer_output[4885] + last_layer_output[4886] + last_layer_output[4887] + last_layer_output[4888] + last_layer_output[4889] + last_layer_output[4890] + last_layer_output[4891] + last_layer_output[4892] + last_layer_output[4893] + last_layer_output[4894] + last_layer_output[4895] + last_layer_output[4896] + last_layer_output[4897] + last_layer_output[4898] + last_layer_output[4899] + last_layer_output[4900] + last_layer_output[4901] + last_layer_output[4902] + last_layer_output[4903] + last_layer_output[4904] + last_layer_output[4905] + last_layer_output[4906] + last_layer_output[4907] + last_layer_output[4908] + last_layer_output[4909] + last_layer_output[4910] + last_layer_output[4911] + last_layer_output[4912] + last_layer_output[4913] + last_layer_output[4914] + last_layer_output[4915] + last_layer_output[4916] + last_layer_output[4917] + last_layer_output[4918] + last_layer_output[4919] + last_layer_output[4920] + last_layer_output[4921] + last_layer_output[4922] + last_layer_output[4923] + last_layer_output[4924] + last_layer_output[4925] + last_layer_output[4926] + last_layer_output[4927] + last_layer_output[4928] + last_layer_output[4929] + last_layer_output[4930] + last_layer_output[4931] + last_layer_output[4932] + last_layer_output[4933] + last_layer_output[4934] + last_layer_output[4935] + last_layer_output[4936] + last_layer_output[4937] + last_layer_output[4938] + last_layer_output[4939] + last_layer_output[4940] + last_layer_output[4941] + last_layer_output[4942] + last_layer_output[4943] + last_layer_output[4944] + last_layer_output[4945] + last_layer_output[4946] + last_layer_output[4947] + last_layer_output[4948] + last_layer_output[4949] + last_layer_output[4950] + last_layer_output[4951] + last_layer_output[4952] + last_layer_output[4953] + last_layer_output[4954] + last_layer_output[4955] + last_layer_output[4956] + last_layer_output[4957] + last_layer_output[4958] + last_layer_output[4959] + last_layer_output[4960] + last_layer_output[4961] + last_layer_output[4962] + last_layer_output[4963] + last_layer_output[4964] + last_layer_output[4965] + last_layer_output[4966] + last_layer_output[4967] + last_layer_output[4968] + last_layer_output[4969] + last_layer_output[4970] + last_layer_output[4971] + last_layer_output[4972] + last_layer_output[4973] + last_layer_output[4974] + last_layer_output[4975] + last_layer_output[4976] + last_layer_output[4977] + last_layer_output[4978] + last_layer_output[4979] + last_layer_output[4980] + last_layer_output[4981] + last_layer_output[4982] + last_layer_output[4983] + last_layer_output[4984] + last_layer_output[4985] + last_layer_output[4986] + last_layer_output[4987] + last_layer_output[4988] + last_layer_output[4989] + last_layer_output[4990] + last_layer_output[4991] + last_layer_output[4992] + last_layer_output[4993] + last_layer_output[4994] + last_layer_output[4995] + last_layer_output[4996] + last_layer_output[4997] + last_layer_output[4998] + last_layer_output[4999] + last_layer_output[5000] + last_layer_output[5001] + last_layer_output[5002] + last_layer_output[5003] + last_layer_output[5004] + last_layer_output[5005] + last_layer_output[5006] + last_layer_output[5007] + last_layer_output[5008] + last_layer_output[5009] + last_layer_output[5010] + last_layer_output[5011] + last_layer_output[5012] + last_layer_output[5013] + last_layer_output[5014] + last_layer_output[5015] + last_layer_output[5016] + last_layer_output[5017] + last_layer_output[5018] + last_layer_output[5019] + last_layer_output[5020] + last_layer_output[5021] + last_layer_output[5022] + last_layer_output[5023] + last_layer_output[5024] + last_layer_output[5025] + last_layer_output[5026] + last_layer_output[5027] + last_layer_output[5028] + last_layer_output[5029] + last_layer_output[5030] + last_layer_output[5031] + last_layer_output[5032] + last_layer_output[5033] + last_layer_output[5034] + last_layer_output[5035] + last_layer_output[5036] + last_layer_output[5037] + last_layer_output[5038] + last_layer_output[5039] + last_layer_output[5040] + last_layer_output[5041] + last_layer_output[5042] + last_layer_output[5043] + last_layer_output[5044] + last_layer_output[5045] + last_layer_output[5046] + last_layer_output[5047] + last_layer_output[5048] + last_layer_output[5049] + last_layer_output[5050] + last_layer_output[5051] + last_layer_output[5052] + last_layer_output[5053] + last_layer_output[5054] + last_layer_output[5055] + last_layer_output[5056] + last_layer_output[5057] + last_layer_output[5058] + last_layer_output[5059] + last_layer_output[5060] + last_layer_output[5061] + last_layer_output[5062] + last_layer_output[5063] + last_layer_output[5064] + last_layer_output[5065] + last_layer_output[5066] + last_layer_output[5067] + last_layer_output[5068] + last_layer_output[5069] + last_layer_output[5070] + last_layer_output[5071] + last_layer_output[5072] + last_layer_output[5073] + last_layer_output[5074] + last_layer_output[5075] + last_layer_output[5076] + last_layer_output[5077] + last_layer_output[5078] + last_layer_output[5079] + last_layer_output[5080] + last_layer_output[5081] + last_layer_output[5082] + last_layer_output[5083] + last_layer_output[5084] + last_layer_output[5085] + last_layer_output[5086] + last_layer_output[5087] + last_layer_output[5088] + last_layer_output[5089] + last_layer_output[5090] + last_layer_output[5091] + last_layer_output[5092] + last_layer_output[5093] + last_layer_output[5094] + last_layer_output[5095] + last_layer_output[5096] + last_layer_output[5097] + last_layer_output[5098] + last_layer_output[5099] + last_layer_output[5100] + last_layer_output[5101] + last_layer_output[5102] + last_layer_output[5103] + last_layer_output[5104] + last_layer_output[5105] + last_layer_output[5106] + last_layer_output[5107] + last_layer_output[5108] + last_layer_output[5109] + last_layer_output[5110] + last_layer_output[5111] + last_layer_output[5112] + last_layer_output[5113] + last_layer_output[5114] + last_layer_output[5115] + last_layer_output[5116] + last_layer_output[5117] + last_layer_output[5118] + last_layer_output[5119] + last_layer_output[5120] + last_layer_output[5121] + last_layer_output[5122] + last_layer_output[5123] + last_layer_output[5124] + last_layer_output[5125] + last_layer_output[5126] + last_layer_output[5127] + last_layer_output[5128] + last_layer_output[5129] + last_layer_output[5130] + last_layer_output[5131] + last_layer_output[5132] + last_layer_output[5133] + last_layer_output[5134] + last_layer_output[5135] + last_layer_output[5136] + last_layer_output[5137] + last_layer_output[5138] + last_layer_output[5139] + last_layer_output[5140] + last_layer_output[5141] + last_layer_output[5142] + last_layer_output[5143] + last_layer_output[5144] + last_layer_output[5145] + last_layer_output[5146] + last_layer_output[5147] + last_layer_output[5148] + last_layer_output[5149] + last_layer_output[5150] + last_layer_output[5151] + last_layer_output[5152] + last_layer_output[5153] + last_layer_output[5154] + last_layer_output[5155] + last_layer_output[5156] + last_layer_output[5157] + last_layer_output[5158] + last_layer_output[5159] + last_layer_output[5160] + last_layer_output[5161] + last_layer_output[5162] + last_layer_output[5163] + last_layer_output[5164] + last_layer_output[5165] + last_layer_output[5166] + last_layer_output[5167] + last_layer_output[5168] + last_layer_output[5169] + last_layer_output[5170] + last_layer_output[5171] + last_layer_output[5172] + last_layer_output[5173] + last_layer_output[5174] + last_layer_output[5175] + last_layer_output[5176] + last_layer_output[5177] + last_layer_output[5178] + last_layer_output[5179] + last_layer_output[5180] + last_layer_output[5181] + last_layer_output[5182] + last_layer_output[5183] + last_layer_output[5184] + last_layer_output[5185] + last_layer_output[5186] + last_layer_output[5187] + last_layer_output[5188] + last_layer_output[5189] + last_layer_output[5190] + last_layer_output[5191] + last_layer_output[5192] + last_layer_output[5193] + last_layer_output[5194] + last_layer_output[5195] + last_layer_output[5196] + last_layer_output[5197] + last_layer_output[5198] + last_layer_output[5199] + last_layer_output[5200] + last_layer_output[5201] + last_layer_output[5202] + last_layer_output[5203] + last_layer_output[5204] + last_layer_output[5205] + last_layer_output[5206] + last_layer_output[5207] + last_layer_output[5208] + last_layer_output[5209] + last_layer_output[5210] + last_layer_output[5211] + last_layer_output[5212] + last_layer_output[5213] + last_layer_output[5214] + last_layer_output[5215] + last_layer_output[5216] + last_layer_output[5217] + last_layer_output[5218] + last_layer_output[5219] + last_layer_output[5220] + last_layer_output[5221] + last_layer_output[5222] + last_layer_output[5223] + last_layer_output[5224] + last_layer_output[5225] + last_layer_output[5226] + last_layer_output[5227] + last_layer_output[5228] + last_layer_output[5229] + last_layer_output[5230] + last_layer_output[5231] + last_layer_output[5232] + last_layer_output[5233] + last_layer_output[5234] + last_layer_output[5235] + last_layer_output[5236] + last_layer_output[5237] + last_layer_output[5238] + last_layer_output[5239] + last_layer_output[5240] + last_layer_output[5241] + last_layer_output[5242] + last_layer_output[5243] + last_layer_output[5244] + last_layer_output[5245] + last_layer_output[5246] + last_layer_output[5247] + last_layer_output[5248] + last_layer_output[5249] + last_layer_output[5250] + last_layer_output[5251] + last_layer_output[5252] + last_layer_output[5253] + last_layer_output[5254] + last_layer_output[5255] + last_layer_output[5256] + last_layer_output[5257] + last_layer_output[5258] + last_layer_output[5259] + last_layer_output[5260] + last_layer_output[5261] + last_layer_output[5262] + last_layer_output[5263] + last_layer_output[5264] + last_layer_output[5265] + last_layer_output[5266] + last_layer_output[5267] + last_layer_output[5268] + last_layer_output[5269] + last_layer_output[5270] + last_layer_output[5271] + last_layer_output[5272] + last_layer_output[5273] + last_layer_output[5274] + last_layer_output[5275] + last_layer_output[5276] + last_layer_output[5277] + last_layer_output[5278] + last_layer_output[5279] + last_layer_output[5280] + last_layer_output[5281] + last_layer_output[5282] + last_layer_output[5283] + last_layer_output[5284] + last_layer_output[5285] + last_layer_output[5286] + last_layer_output[5287] + last_layer_output[5288] + last_layer_output[5289] + last_layer_output[5290] + last_layer_output[5291] + last_layer_output[5292] + last_layer_output[5293] + last_layer_output[5294] + last_layer_output[5295] + last_layer_output[5296] + last_layer_output[5297] + last_layer_output[5298] + last_layer_output[5299] + last_layer_output[5300] + last_layer_output[5301] + last_layer_output[5302] + last_layer_output[5303] + last_layer_output[5304] + last_layer_output[5305] + last_layer_output[5306] + last_layer_output[5307] + last_layer_output[5308] + last_layer_output[5309] + last_layer_output[5310] + last_layer_output[5311] + last_layer_output[5312] + last_layer_output[5313] + last_layer_output[5314] + last_layer_output[5315] + last_layer_output[5316] + last_layer_output[5317] + last_layer_output[5318] + last_layer_output[5319] + last_layer_output[5320] + last_layer_output[5321] + last_layer_output[5322] + last_layer_output[5323] + last_layer_output[5324] + last_layer_output[5325] + last_layer_output[5326] + last_layer_output[5327] + last_layer_output[5328] + last_layer_output[5329] + last_layer_output[5330] + last_layer_output[5331] + last_layer_output[5332] + last_layer_output[5333] + last_layer_output[5334] + last_layer_output[5335] + last_layer_output[5336] + last_layer_output[5337] + last_layer_output[5338] + last_layer_output[5339] + last_layer_output[5340] + last_layer_output[5341] + last_layer_output[5342] + last_layer_output[5343] + last_layer_output[5344] + last_layer_output[5345] + last_layer_output[5346] + last_layer_output[5347] + last_layer_output[5348] + last_layer_output[5349] + last_layer_output[5350] + last_layer_output[5351] + last_layer_output[5352] + last_layer_output[5353] + last_layer_output[5354] + last_layer_output[5355] + last_layer_output[5356] + last_layer_output[5357] + last_layer_output[5358] + last_layer_output[5359] + last_layer_output[5360] + last_layer_output[5361] + last_layer_output[5362] + last_layer_output[5363] + last_layer_output[5364] + last_layer_output[5365] + last_layer_output[5366] + last_layer_output[5367] + last_layer_output[5368] + last_layer_output[5369] + last_layer_output[5370] + last_layer_output[5371] + last_layer_output[5372] + last_layer_output[5373] + last_layer_output[5374] + last_layer_output[5375] + last_layer_output[5376] + last_layer_output[5377] + last_layer_output[5378] + last_layer_output[5379] + last_layer_output[5380] + last_layer_output[5381] + last_layer_output[5382] + last_layer_output[5383] + last_layer_output[5384] + last_layer_output[5385] + last_layer_output[5386] + last_layer_output[5387] + last_layer_output[5388] + last_layer_output[5389] + last_layer_output[5390] + last_layer_output[5391] + last_layer_output[5392] + last_layer_output[5393] + last_layer_output[5394] + last_layer_output[5395] + last_layer_output[5396] + last_layer_output[5397] + last_layer_output[5398] + last_layer_output[5399] + last_layer_output[5400] + last_layer_output[5401] + last_layer_output[5402] + last_layer_output[5403] + last_layer_output[5404] + last_layer_output[5405] + last_layer_output[5406] + last_layer_output[5407] + last_layer_output[5408] + last_layer_output[5409] + last_layer_output[5410] + last_layer_output[5411] + last_layer_output[5412] + last_layer_output[5413] + last_layer_output[5414] + last_layer_output[5415] + last_layer_output[5416] + last_layer_output[5417] + last_layer_output[5418] + last_layer_output[5419] + last_layer_output[5420] + last_layer_output[5421] + last_layer_output[5422] + last_layer_output[5423] + last_layer_output[5424] + last_layer_output[5425] + last_layer_output[5426] + last_layer_output[5427] + last_layer_output[5428] + last_layer_output[5429] + last_layer_output[5430] + last_layer_output[5431] + last_layer_output[5432] + last_layer_output[5433] + last_layer_output[5434] + last_layer_output[5435] + last_layer_output[5436] + last_layer_output[5437] + last_layer_output[5438] + last_layer_output[5439] + last_layer_output[5440] + last_layer_output[5441] + last_layer_output[5442] + last_layer_output[5443] + last_layer_output[5444] + last_layer_output[5445] + last_layer_output[5446] + last_layer_output[5447] + last_layer_output[5448] + last_layer_output[5449] + last_layer_output[5450] + last_layer_output[5451] + last_layer_output[5452] + last_layer_output[5453] + last_layer_output[5454] + last_layer_output[5455] + last_layer_output[5456] + last_layer_output[5457] + last_layer_output[5458] + last_layer_output[5459] + last_layer_output[5460] + last_layer_output[5461] + last_layer_output[5462] + last_layer_output[5463] + last_layer_output[5464] + last_layer_output[5465] + last_layer_output[5466] + last_layer_output[5467] + last_layer_output[5468] + last_layer_output[5469] + last_layer_output[5470] + last_layer_output[5471] + last_layer_output[5472] + last_layer_output[5473] + last_layer_output[5474] + last_layer_output[5475] + last_layer_output[5476] + last_layer_output[5477] + last_layer_output[5478] + last_layer_output[5479] + last_layer_output[5480] + last_layer_output[5481] + last_layer_output[5482] + last_layer_output[5483] + last_layer_output[5484] + last_layer_output[5485] + last_layer_output[5486] + last_layer_output[5487] + last_layer_output[5488] + last_layer_output[5489] + last_layer_output[5490] + last_layer_output[5491] + last_layer_output[5492] + last_layer_output[5493] + last_layer_output[5494] + last_layer_output[5495] + last_layer_output[5496] + last_layer_output[5497] + last_layer_output[5498] + last_layer_output[5499] + last_layer_output[5500] + last_layer_output[5501] + last_layer_output[5502] + last_layer_output[5503] + last_layer_output[5504] + last_layer_output[5505] + last_layer_output[5506] + last_layer_output[5507] + last_layer_output[5508] + last_layer_output[5509] + last_layer_output[5510] + last_layer_output[5511] + last_layer_output[5512] + last_layer_output[5513] + last_layer_output[5514] + last_layer_output[5515] + last_layer_output[5516] + last_layer_output[5517] + last_layer_output[5518] + last_layer_output[5519] + last_layer_output[5520] + last_layer_output[5521] + last_layer_output[5522] + last_layer_output[5523] + last_layer_output[5524] + last_layer_output[5525] + last_layer_output[5526] + last_layer_output[5527] + last_layer_output[5528] + last_layer_output[5529] + last_layer_output[5530] + last_layer_output[5531] + last_layer_output[5532] + last_layer_output[5533] + last_layer_output[5534] + last_layer_output[5535] + last_layer_output[5536] + last_layer_output[5537] + last_layer_output[5538] + last_layer_output[5539] + last_layer_output[5540] + last_layer_output[5541] + last_layer_output[5542] + last_layer_output[5543] + last_layer_output[5544] + last_layer_output[5545] + last_layer_output[5546] + last_layer_output[5547] + last_layer_output[5548] + last_layer_output[5549] + last_layer_output[5550] + last_layer_output[5551] + last_layer_output[5552] + last_layer_output[5553] + last_layer_output[5554] + last_layer_output[5555] + last_layer_output[5556] + last_layer_output[5557] + last_layer_output[5558] + last_layer_output[5559] + last_layer_output[5560] + last_layer_output[5561] + last_layer_output[5562] + last_layer_output[5563] + last_layer_output[5564] + last_layer_output[5565] + last_layer_output[5566] + last_layer_output[5567] + last_layer_output[5568] + last_layer_output[5569] + last_layer_output[5570] + last_layer_output[5571] + last_layer_output[5572] + last_layer_output[5573] + last_layer_output[5574] + last_layer_output[5575] + last_layer_output[5576] + last_layer_output[5577] + last_layer_output[5578] + last_layer_output[5579] + last_layer_output[5580] + last_layer_output[5581] + last_layer_output[5582] + last_layer_output[5583] + last_layer_output[5584] + last_layer_output[5585] + last_layer_output[5586] + last_layer_output[5587] + last_layer_output[5588] + last_layer_output[5589] + last_layer_output[5590] + last_layer_output[5591] + last_layer_output[5592] + last_layer_output[5593] + last_layer_output[5594] + last_layer_output[5595] + last_layer_output[5596] + last_layer_output[5597] + last_layer_output[5598] + last_layer_output[5599] + last_layer_output[5600] + last_layer_output[5601] + last_layer_output[5602] + last_layer_output[5603] + last_layer_output[5604] + last_layer_output[5605] + last_layer_output[5606] + last_layer_output[5607] + last_layer_output[5608] + last_layer_output[5609] + last_layer_output[5610] + last_layer_output[5611] + last_layer_output[5612] + last_layer_output[5613] + last_layer_output[5614] + last_layer_output[5615] + last_layer_output[5616] + last_layer_output[5617] + last_layer_output[5618] + last_layer_output[5619] + last_layer_output[5620] + last_layer_output[5621] + last_layer_output[5622] + last_layer_output[5623] + last_layer_output[5624] + last_layer_output[5625] + last_layer_output[5626] + last_layer_output[5627] + last_layer_output[5628] + last_layer_output[5629] + last_layer_output[5630] + last_layer_output[5631] + last_layer_output[5632] + last_layer_output[5633] + last_layer_output[5634] + last_layer_output[5635] + last_layer_output[5636] + last_layer_output[5637] + last_layer_output[5638] + last_layer_output[5639] + last_layer_output[5640] + last_layer_output[5641] + last_layer_output[5642] + last_layer_output[5643] + last_layer_output[5644] + last_layer_output[5645] + last_layer_output[5646] + last_layer_output[5647] + last_layer_output[5648] + last_layer_output[5649] + last_layer_output[5650] + last_layer_output[5651] + last_layer_output[5652] + last_layer_output[5653] + last_layer_output[5654] + last_layer_output[5655] + last_layer_output[5656] + last_layer_output[5657] + last_layer_output[5658] + last_layer_output[5659] + last_layer_output[5660] + last_layer_output[5661] + last_layer_output[5662] + last_layer_output[5663] + last_layer_output[5664] + last_layer_output[5665] + last_layer_output[5666] + last_layer_output[5667] + last_layer_output[5668] + last_layer_output[5669] + last_layer_output[5670] + last_layer_output[5671] + last_layer_output[5672] + last_layer_output[5673] + last_layer_output[5674] + last_layer_output[5675] + last_layer_output[5676] + last_layer_output[5677] + last_layer_output[5678] + last_layer_output[5679] + last_layer_output[5680] + last_layer_output[5681] + last_layer_output[5682] + last_layer_output[5683] + last_layer_output[5684] + last_layer_output[5685] + last_layer_output[5686] + last_layer_output[5687] + last_layer_output[5688] + last_layer_output[5689] + last_layer_output[5690] + last_layer_output[5691] + last_layer_output[5692] + last_layer_output[5693] + last_layer_output[5694] + last_layer_output[5695] + last_layer_output[5696] + last_layer_output[5697] + last_layer_output[5698] + last_layer_output[5699] + last_layer_output[5700] + last_layer_output[5701] + last_layer_output[5702] + last_layer_output[5703] + last_layer_output[5704] + last_layer_output[5705] + last_layer_output[5706] + last_layer_output[5707] + last_layer_output[5708] + last_layer_output[5709] + last_layer_output[5710] + last_layer_output[5711] + last_layer_output[5712] + last_layer_output[5713] + last_layer_output[5714] + last_layer_output[5715] + last_layer_output[5716] + last_layer_output[5717] + last_layer_output[5718] + last_layer_output[5719] + last_layer_output[5720] + last_layer_output[5721] + last_layer_output[5722] + last_layer_output[5723] + last_layer_output[5724] + last_layer_output[5725] + last_layer_output[5726] + last_layer_output[5727] + last_layer_output[5728] + last_layer_output[5729] + last_layer_output[5730] + last_layer_output[5731] + last_layer_output[5732] + last_layer_output[5733] + last_layer_output[5734] + last_layer_output[5735] + last_layer_output[5736] + last_layer_output[5737] + last_layer_output[5738] + last_layer_output[5739] + last_layer_output[5740] + last_layer_output[5741] + last_layer_output[5742] + last_layer_output[5743] + last_layer_output[5744] + last_layer_output[5745] + last_layer_output[5746] + last_layer_output[5747] + last_layer_output[5748] + last_layer_output[5749] + last_layer_output[5750] + last_layer_output[5751] + last_layer_output[5752] + last_layer_output[5753] + last_layer_output[5754] + last_layer_output[5755] + last_layer_output[5756] + last_layer_output[5757] + last_layer_output[5758] + last_layer_output[5759] + last_layer_output[5760] + last_layer_output[5761] + last_layer_output[5762] + last_layer_output[5763] + last_layer_output[5764] + last_layer_output[5765] + last_layer_output[5766] + last_layer_output[5767] + last_layer_output[5768] + last_layer_output[5769] + last_layer_output[5770] + last_layer_output[5771] + last_layer_output[5772] + last_layer_output[5773] + last_layer_output[5774] + last_layer_output[5775] + last_layer_output[5776] + last_layer_output[5777] + last_layer_output[5778] + last_layer_output[5779] + last_layer_output[5780] + last_layer_output[5781] + last_layer_output[5782] + last_layer_output[5783] + last_layer_output[5784] + last_layer_output[5785] + last_layer_output[5786] + last_layer_output[5787] + last_layer_output[5788] + last_layer_output[5789] + last_layer_output[5790] + last_layer_output[5791] + last_layer_output[5792] + last_layer_output[5793] + last_layer_output[5794] + last_layer_output[5795] + last_layer_output[5796] + last_layer_output[5797] + last_layer_output[5798] + last_layer_output[5799] + last_layer_output[5800] + last_layer_output[5801] + last_layer_output[5802] + last_layer_output[5803] + last_layer_output[5804] + last_layer_output[5805] + last_layer_output[5806] + last_layer_output[5807] + last_layer_output[5808] + last_layer_output[5809] + last_layer_output[5810] + last_layer_output[5811] + last_layer_output[5812] + last_layer_output[5813] + last_layer_output[5814] + last_layer_output[5815] + last_layer_output[5816] + last_layer_output[5817] + last_layer_output[5818] + last_layer_output[5819] + last_layer_output[5820] + last_layer_output[5821] + last_layer_output[5822] + last_layer_output[5823] + last_layer_output[5824] + last_layer_output[5825] + last_layer_output[5826] + last_layer_output[5827] + last_layer_output[5828] + last_layer_output[5829] + last_layer_output[5830] + last_layer_output[5831] + last_layer_output[5832] + last_layer_output[5833] + last_layer_output[5834] + last_layer_output[5835] + last_layer_output[5836] + last_layer_output[5837] + last_layer_output[5838] + last_layer_output[5839] + last_layer_output[5840] + last_layer_output[5841] + last_layer_output[5842] + last_layer_output[5843] + last_layer_output[5844] + last_layer_output[5845] + last_layer_output[5846] + last_layer_output[5847] + last_layer_output[5848] + last_layer_output[5849] + last_layer_output[5850] + last_layer_output[5851] + last_layer_output[5852] + last_layer_output[5853] + last_layer_output[5854] + last_layer_output[5855] + last_layer_output[5856] + last_layer_output[5857] + last_layer_output[5858] + last_layer_output[5859] + last_layer_output[5860] + last_layer_output[5861] + last_layer_output[5862] + last_layer_output[5863] + last_layer_output[5864] + last_layer_output[5865] + last_layer_output[5866] + last_layer_output[5867] + last_layer_output[5868] + last_layer_output[5869] + last_layer_output[5870] + last_layer_output[5871] + last_layer_output[5872] + last_layer_output[5873] + last_layer_output[5874] + last_layer_output[5875] + last_layer_output[5876] + last_layer_output[5877] + last_layer_output[5878] + last_layer_output[5879] + last_layer_output[5880] + last_layer_output[5881] + last_layer_output[5882] + last_layer_output[5883] + last_layer_output[5884] + last_layer_output[5885] + last_layer_output[5886] + last_layer_output[5887] + last_layer_output[5888] + last_layer_output[5889] + last_layer_output[5890] + last_layer_output[5891] + last_layer_output[5892] + last_layer_output[5893] + last_layer_output[5894] + last_layer_output[5895] + last_layer_output[5896] + last_layer_output[5897] + last_layer_output[5898] + last_layer_output[5899] + last_layer_output[5900] + last_layer_output[5901] + last_layer_output[5902] + last_layer_output[5903] + last_layer_output[5904] + last_layer_output[5905] + last_layer_output[5906] + last_layer_output[5907] + last_layer_output[5908] + last_layer_output[5909] + last_layer_output[5910] + last_layer_output[5911] + last_layer_output[5912] + last_layer_output[5913] + last_layer_output[5914] + last_layer_output[5915] + last_layer_output[5916] + last_layer_output[5917] + last_layer_output[5918] + last_layer_output[5919] + last_layer_output[5920] + last_layer_output[5921] + last_layer_output[5922] + last_layer_output[5923] + last_layer_output[5924] + last_layer_output[5925] + last_layer_output[5926] + last_layer_output[5927] + last_layer_output[5928] + last_layer_output[5929] + last_layer_output[5930] + last_layer_output[5931] + last_layer_output[5932] + last_layer_output[5933] + last_layer_output[5934] + last_layer_output[5935] + last_layer_output[5936] + last_layer_output[5937] + last_layer_output[5938] + last_layer_output[5939] + last_layer_output[5940] + last_layer_output[5941] + last_layer_output[5942] + last_layer_output[5943] + last_layer_output[5944] + last_layer_output[5945] + last_layer_output[5946] + last_layer_output[5947] + last_layer_output[5948] + last_layer_output[5949] + last_layer_output[5950] + last_layer_output[5951] + last_layer_output[5952] + last_layer_output[5953] + last_layer_output[5954] + last_layer_output[5955] + last_layer_output[5956] + last_layer_output[5957] + last_layer_output[5958] + last_layer_output[5959] + last_layer_output[5960] + last_layer_output[5961] + last_layer_output[5962] + last_layer_output[5963] + last_layer_output[5964] + last_layer_output[5965] + last_layer_output[5966] + last_layer_output[5967] + last_layer_output[5968] + last_layer_output[5969] + last_layer_output[5970] + last_layer_output[5971] + last_layer_output[5972] + last_layer_output[5973] + last_layer_output[5974] + last_layer_output[5975] + last_layer_output[5976] + last_layer_output[5977] + last_layer_output[5978] + last_layer_output[5979] + last_layer_output[5980] + last_layer_output[5981] + last_layer_output[5982] + last_layer_output[5983] + last_layer_output[5984] + last_layer_output[5985] + last_layer_output[5986] + last_layer_output[5987] + last_layer_output[5988] + last_layer_output[5989] + last_layer_output[5990] + last_layer_output[5991] + last_layer_output[5992] + last_layer_output[5993] + last_layer_output[5994] + last_layer_output[5995] + last_layer_output[5996] + last_layer_output[5997] + last_layer_output[5998] + last_layer_output[5999];
      result[5] <= last_layer_output[6000] + last_layer_output[6001] + last_layer_output[6002] + last_layer_output[6003] + last_layer_output[6004] + last_layer_output[6005] + last_layer_output[6006] + last_layer_output[6007] + last_layer_output[6008] + last_layer_output[6009] + last_layer_output[6010] + last_layer_output[6011] + last_layer_output[6012] + last_layer_output[6013] + last_layer_output[6014] + last_layer_output[6015] + last_layer_output[6016] + last_layer_output[6017] + last_layer_output[6018] + last_layer_output[6019] + last_layer_output[6020] + last_layer_output[6021] + last_layer_output[6022] + last_layer_output[6023] + last_layer_output[6024] + last_layer_output[6025] + last_layer_output[6026] + last_layer_output[6027] + last_layer_output[6028] + last_layer_output[6029] + last_layer_output[6030] + last_layer_output[6031] + last_layer_output[6032] + last_layer_output[6033] + last_layer_output[6034] + last_layer_output[6035] + last_layer_output[6036] + last_layer_output[6037] + last_layer_output[6038] + last_layer_output[6039] + last_layer_output[6040] + last_layer_output[6041] + last_layer_output[6042] + last_layer_output[6043] + last_layer_output[6044] + last_layer_output[6045] + last_layer_output[6046] + last_layer_output[6047] + last_layer_output[6048] + last_layer_output[6049] + last_layer_output[6050] + last_layer_output[6051] + last_layer_output[6052] + last_layer_output[6053] + last_layer_output[6054] + last_layer_output[6055] + last_layer_output[6056] + last_layer_output[6057] + last_layer_output[6058] + last_layer_output[6059] + last_layer_output[6060] + last_layer_output[6061] + last_layer_output[6062] + last_layer_output[6063] + last_layer_output[6064] + last_layer_output[6065] + last_layer_output[6066] + last_layer_output[6067] + last_layer_output[6068] + last_layer_output[6069] + last_layer_output[6070] + last_layer_output[6071] + last_layer_output[6072] + last_layer_output[6073] + last_layer_output[6074] + last_layer_output[6075] + last_layer_output[6076] + last_layer_output[6077] + last_layer_output[6078] + last_layer_output[6079] + last_layer_output[6080] + last_layer_output[6081] + last_layer_output[6082] + last_layer_output[6083] + last_layer_output[6084] + last_layer_output[6085] + last_layer_output[6086] + last_layer_output[6087] + last_layer_output[6088] + last_layer_output[6089] + last_layer_output[6090] + last_layer_output[6091] + last_layer_output[6092] + last_layer_output[6093] + last_layer_output[6094] + last_layer_output[6095] + last_layer_output[6096] + last_layer_output[6097] + last_layer_output[6098] + last_layer_output[6099] + last_layer_output[6100] + last_layer_output[6101] + last_layer_output[6102] + last_layer_output[6103] + last_layer_output[6104] + last_layer_output[6105] + last_layer_output[6106] + last_layer_output[6107] + last_layer_output[6108] + last_layer_output[6109] + last_layer_output[6110] + last_layer_output[6111] + last_layer_output[6112] + last_layer_output[6113] + last_layer_output[6114] + last_layer_output[6115] + last_layer_output[6116] + last_layer_output[6117] + last_layer_output[6118] + last_layer_output[6119] + last_layer_output[6120] + last_layer_output[6121] + last_layer_output[6122] + last_layer_output[6123] + last_layer_output[6124] + last_layer_output[6125] + last_layer_output[6126] + last_layer_output[6127] + last_layer_output[6128] + last_layer_output[6129] + last_layer_output[6130] + last_layer_output[6131] + last_layer_output[6132] + last_layer_output[6133] + last_layer_output[6134] + last_layer_output[6135] + last_layer_output[6136] + last_layer_output[6137] + last_layer_output[6138] + last_layer_output[6139] + last_layer_output[6140] + last_layer_output[6141] + last_layer_output[6142] + last_layer_output[6143] + last_layer_output[6144] + last_layer_output[6145] + last_layer_output[6146] + last_layer_output[6147] + last_layer_output[6148] + last_layer_output[6149] + last_layer_output[6150] + last_layer_output[6151] + last_layer_output[6152] + last_layer_output[6153] + last_layer_output[6154] + last_layer_output[6155] + last_layer_output[6156] + last_layer_output[6157] + last_layer_output[6158] + last_layer_output[6159] + last_layer_output[6160] + last_layer_output[6161] + last_layer_output[6162] + last_layer_output[6163] + last_layer_output[6164] + last_layer_output[6165] + last_layer_output[6166] + last_layer_output[6167] + last_layer_output[6168] + last_layer_output[6169] + last_layer_output[6170] + last_layer_output[6171] + last_layer_output[6172] + last_layer_output[6173] + last_layer_output[6174] + last_layer_output[6175] + last_layer_output[6176] + last_layer_output[6177] + last_layer_output[6178] + last_layer_output[6179] + last_layer_output[6180] + last_layer_output[6181] + last_layer_output[6182] + last_layer_output[6183] + last_layer_output[6184] + last_layer_output[6185] + last_layer_output[6186] + last_layer_output[6187] + last_layer_output[6188] + last_layer_output[6189] + last_layer_output[6190] + last_layer_output[6191] + last_layer_output[6192] + last_layer_output[6193] + last_layer_output[6194] + last_layer_output[6195] + last_layer_output[6196] + last_layer_output[6197] + last_layer_output[6198] + last_layer_output[6199] + last_layer_output[6200] + last_layer_output[6201] + last_layer_output[6202] + last_layer_output[6203] + last_layer_output[6204] + last_layer_output[6205] + last_layer_output[6206] + last_layer_output[6207] + last_layer_output[6208] + last_layer_output[6209] + last_layer_output[6210] + last_layer_output[6211] + last_layer_output[6212] + last_layer_output[6213] + last_layer_output[6214] + last_layer_output[6215] + last_layer_output[6216] + last_layer_output[6217] + last_layer_output[6218] + last_layer_output[6219] + last_layer_output[6220] + last_layer_output[6221] + last_layer_output[6222] + last_layer_output[6223] + last_layer_output[6224] + last_layer_output[6225] + last_layer_output[6226] + last_layer_output[6227] + last_layer_output[6228] + last_layer_output[6229] + last_layer_output[6230] + last_layer_output[6231] + last_layer_output[6232] + last_layer_output[6233] + last_layer_output[6234] + last_layer_output[6235] + last_layer_output[6236] + last_layer_output[6237] + last_layer_output[6238] + last_layer_output[6239] + last_layer_output[6240] + last_layer_output[6241] + last_layer_output[6242] + last_layer_output[6243] + last_layer_output[6244] + last_layer_output[6245] + last_layer_output[6246] + last_layer_output[6247] + last_layer_output[6248] + last_layer_output[6249] + last_layer_output[6250] + last_layer_output[6251] + last_layer_output[6252] + last_layer_output[6253] + last_layer_output[6254] + last_layer_output[6255] + last_layer_output[6256] + last_layer_output[6257] + last_layer_output[6258] + last_layer_output[6259] + last_layer_output[6260] + last_layer_output[6261] + last_layer_output[6262] + last_layer_output[6263] + last_layer_output[6264] + last_layer_output[6265] + last_layer_output[6266] + last_layer_output[6267] + last_layer_output[6268] + last_layer_output[6269] + last_layer_output[6270] + last_layer_output[6271] + last_layer_output[6272] + last_layer_output[6273] + last_layer_output[6274] + last_layer_output[6275] + last_layer_output[6276] + last_layer_output[6277] + last_layer_output[6278] + last_layer_output[6279] + last_layer_output[6280] + last_layer_output[6281] + last_layer_output[6282] + last_layer_output[6283] + last_layer_output[6284] + last_layer_output[6285] + last_layer_output[6286] + last_layer_output[6287] + last_layer_output[6288] + last_layer_output[6289] + last_layer_output[6290] + last_layer_output[6291] + last_layer_output[6292] + last_layer_output[6293] + last_layer_output[6294] + last_layer_output[6295] + last_layer_output[6296] + last_layer_output[6297] + last_layer_output[6298] + last_layer_output[6299] + last_layer_output[6300] + last_layer_output[6301] + last_layer_output[6302] + last_layer_output[6303] + last_layer_output[6304] + last_layer_output[6305] + last_layer_output[6306] + last_layer_output[6307] + last_layer_output[6308] + last_layer_output[6309] + last_layer_output[6310] + last_layer_output[6311] + last_layer_output[6312] + last_layer_output[6313] + last_layer_output[6314] + last_layer_output[6315] + last_layer_output[6316] + last_layer_output[6317] + last_layer_output[6318] + last_layer_output[6319] + last_layer_output[6320] + last_layer_output[6321] + last_layer_output[6322] + last_layer_output[6323] + last_layer_output[6324] + last_layer_output[6325] + last_layer_output[6326] + last_layer_output[6327] + last_layer_output[6328] + last_layer_output[6329] + last_layer_output[6330] + last_layer_output[6331] + last_layer_output[6332] + last_layer_output[6333] + last_layer_output[6334] + last_layer_output[6335] + last_layer_output[6336] + last_layer_output[6337] + last_layer_output[6338] + last_layer_output[6339] + last_layer_output[6340] + last_layer_output[6341] + last_layer_output[6342] + last_layer_output[6343] + last_layer_output[6344] + last_layer_output[6345] + last_layer_output[6346] + last_layer_output[6347] + last_layer_output[6348] + last_layer_output[6349] + last_layer_output[6350] + last_layer_output[6351] + last_layer_output[6352] + last_layer_output[6353] + last_layer_output[6354] + last_layer_output[6355] + last_layer_output[6356] + last_layer_output[6357] + last_layer_output[6358] + last_layer_output[6359] + last_layer_output[6360] + last_layer_output[6361] + last_layer_output[6362] + last_layer_output[6363] + last_layer_output[6364] + last_layer_output[6365] + last_layer_output[6366] + last_layer_output[6367] + last_layer_output[6368] + last_layer_output[6369] + last_layer_output[6370] + last_layer_output[6371] + last_layer_output[6372] + last_layer_output[6373] + last_layer_output[6374] + last_layer_output[6375] + last_layer_output[6376] + last_layer_output[6377] + last_layer_output[6378] + last_layer_output[6379] + last_layer_output[6380] + last_layer_output[6381] + last_layer_output[6382] + last_layer_output[6383] + last_layer_output[6384] + last_layer_output[6385] + last_layer_output[6386] + last_layer_output[6387] + last_layer_output[6388] + last_layer_output[6389] + last_layer_output[6390] + last_layer_output[6391] + last_layer_output[6392] + last_layer_output[6393] + last_layer_output[6394] + last_layer_output[6395] + last_layer_output[6396] + last_layer_output[6397] + last_layer_output[6398] + last_layer_output[6399] + last_layer_output[6400] + last_layer_output[6401] + last_layer_output[6402] + last_layer_output[6403] + last_layer_output[6404] + last_layer_output[6405] + last_layer_output[6406] + last_layer_output[6407] + last_layer_output[6408] + last_layer_output[6409] + last_layer_output[6410] + last_layer_output[6411] + last_layer_output[6412] + last_layer_output[6413] + last_layer_output[6414] + last_layer_output[6415] + last_layer_output[6416] + last_layer_output[6417] + last_layer_output[6418] + last_layer_output[6419] + last_layer_output[6420] + last_layer_output[6421] + last_layer_output[6422] + last_layer_output[6423] + last_layer_output[6424] + last_layer_output[6425] + last_layer_output[6426] + last_layer_output[6427] + last_layer_output[6428] + last_layer_output[6429] + last_layer_output[6430] + last_layer_output[6431] + last_layer_output[6432] + last_layer_output[6433] + last_layer_output[6434] + last_layer_output[6435] + last_layer_output[6436] + last_layer_output[6437] + last_layer_output[6438] + last_layer_output[6439] + last_layer_output[6440] + last_layer_output[6441] + last_layer_output[6442] + last_layer_output[6443] + last_layer_output[6444] + last_layer_output[6445] + last_layer_output[6446] + last_layer_output[6447] + last_layer_output[6448] + last_layer_output[6449] + last_layer_output[6450] + last_layer_output[6451] + last_layer_output[6452] + last_layer_output[6453] + last_layer_output[6454] + last_layer_output[6455] + last_layer_output[6456] + last_layer_output[6457] + last_layer_output[6458] + last_layer_output[6459] + last_layer_output[6460] + last_layer_output[6461] + last_layer_output[6462] + last_layer_output[6463] + last_layer_output[6464] + last_layer_output[6465] + last_layer_output[6466] + last_layer_output[6467] + last_layer_output[6468] + last_layer_output[6469] + last_layer_output[6470] + last_layer_output[6471] + last_layer_output[6472] + last_layer_output[6473] + last_layer_output[6474] + last_layer_output[6475] + last_layer_output[6476] + last_layer_output[6477] + last_layer_output[6478] + last_layer_output[6479] + last_layer_output[6480] + last_layer_output[6481] + last_layer_output[6482] + last_layer_output[6483] + last_layer_output[6484] + last_layer_output[6485] + last_layer_output[6486] + last_layer_output[6487] + last_layer_output[6488] + last_layer_output[6489] + last_layer_output[6490] + last_layer_output[6491] + last_layer_output[6492] + last_layer_output[6493] + last_layer_output[6494] + last_layer_output[6495] + last_layer_output[6496] + last_layer_output[6497] + last_layer_output[6498] + last_layer_output[6499] + last_layer_output[6500] + last_layer_output[6501] + last_layer_output[6502] + last_layer_output[6503] + last_layer_output[6504] + last_layer_output[6505] + last_layer_output[6506] + last_layer_output[6507] + last_layer_output[6508] + last_layer_output[6509] + last_layer_output[6510] + last_layer_output[6511] + last_layer_output[6512] + last_layer_output[6513] + last_layer_output[6514] + last_layer_output[6515] + last_layer_output[6516] + last_layer_output[6517] + last_layer_output[6518] + last_layer_output[6519] + last_layer_output[6520] + last_layer_output[6521] + last_layer_output[6522] + last_layer_output[6523] + last_layer_output[6524] + last_layer_output[6525] + last_layer_output[6526] + last_layer_output[6527] + last_layer_output[6528] + last_layer_output[6529] + last_layer_output[6530] + last_layer_output[6531] + last_layer_output[6532] + last_layer_output[6533] + last_layer_output[6534] + last_layer_output[6535] + last_layer_output[6536] + last_layer_output[6537] + last_layer_output[6538] + last_layer_output[6539] + last_layer_output[6540] + last_layer_output[6541] + last_layer_output[6542] + last_layer_output[6543] + last_layer_output[6544] + last_layer_output[6545] + last_layer_output[6546] + last_layer_output[6547] + last_layer_output[6548] + last_layer_output[6549] + last_layer_output[6550] + last_layer_output[6551] + last_layer_output[6552] + last_layer_output[6553] + last_layer_output[6554] + last_layer_output[6555] + last_layer_output[6556] + last_layer_output[6557] + last_layer_output[6558] + last_layer_output[6559] + last_layer_output[6560] + last_layer_output[6561] + last_layer_output[6562] + last_layer_output[6563] + last_layer_output[6564] + last_layer_output[6565] + last_layer_output[6566] + last_layer_output[6567] + last_layer_output[6568] + last_layer_output[6569] + last_layer_output[6570] + last_layer_output[6571] + last_layer_output[6572] + last_layer_output[6573] + last_layer_output[6574] + last_layer_output[6575] + last_layer_output[6576] + last_layer_output[6577] + last_layer_output[6578] + last_layer_output[6579] + last_layer_output[6580] + last_layer_output[6581] + last_layer_output[6582] + last_layer_output[6583] + last_layer_output[6584] + last_layer_output[6585] + last_layer_output[6586] + last_layer_output[6587] + last_layer_output[6588] + last_layer_output[6589] + last_layer_output[6590] + last_layer_output[6591] + last_layer_output[6592] + last_layer_output[6593] + last_layer_output[6594] + last_layer_output[6595] + last_layer_output[6596] + last_layer_output[6597] + last_layer_output[6598] + last_layer_output[6599] + last_layer_output[6600] + last_layer_output[6601] + last_layer_output[6602] + last_layer_output[6603] + last_layer_output[6604] + last_layer_output[6605] + last_layer_output[6606] + last_layer_output[6607] + last_layer_output[6608] + last_layer_output[6609] + last_layer_output[6610] + last_layer_output[6611] + last_layer_output[6612] + last_layer_output[6613] + last_layer_output[6614] + last_layer_output[6615] + last_layer_output[6616] + last_layer_output[6617] + last_layer_output[6618] + last_layer_output[6619] + last_layer_output[6620] + last_layer_output[6621] + last_layer_output[6622] + last_layer_output[6623] + last_layer_output[6624] + last_layer_output[6625] + last_layer_output[6626] + last_layer_output[6627] + last_layer_output[6628] + last_layer_output[6629] + last_layer_output[6630] + last_layer_output[6631] + last_layer_output[6632] + last_layer_output[6633] + last_layer_output[6634] + last_layer_output[6635] + last_layer_output[6636] + last_layer_output[6637] + last_layer_output[6638] + last_layer_output[6639] + last_layer_output[6640] + last_layer_output[6641] + last_layer_output[6642] + last_layer_output[6643] + last_layer_output[6644] + last_layer_output[6645] + last_layer_output[6646] + last_layer_output[6647] + last_layer_output[6648] + last_layer_output[6649] + last_layer_output[6650] + last_layer_output[6651] + last_layer_output[6652] + last_layer_output[6653] + last_layer_output[6654] + last_layer_output[6655] + last_layer_output[6656] + last_layer_output[6657] + last_layer_output[6658] + last_layer_output[6659] + last_layer_output[6660] + last_layer_output[6661] + last_layer_output[6662] + last_layer_output[6663] + last_layer_output[6664] + last_layer_output[6665] + last_layer_output[6666] + last_layer_output[6667] + last_layer_output[6668] + last_layer_output[6669] + last_layer_output[6670] + last_layer_output[6671] + last_layer_output[6672] + last_layer_output[6673] + last_layer_output[6674] + last_layer_output[6675] + last_layer_output[6676] + last_layer_output[6677] + last_layer_output[6678] + last_layer_output[6679] + last_layer_output[6680] + last_layer_output[6681] + last_layer_output[6682] + last_layer_output[6683] + last_layer_output[6684] + last_layer_output[6685] + last_layer_output[6686] + last_layer_output[6687] + last_layer_output[6688] + last_layer_output[6689] + last_layer_output[6690] + last_layer_output[6691] + last_layer_output[6692] + last_layer_output[6693] + last_layer_output[6694] + last_layer_output[6695] + last_layer_output[6696] + last_layer_output[6697] + last_layer_output[6698] + last_layer_output[6699] + last_layer_output[6700] + last_layer_output[6701] + last_layer_output[6702] + last_layer_output[6703] + last_layer_output[6704] + last_layer_output[6705] + last_layer_output[6706] + last_layer_output[6707] + last_layer_output[6708] + last_layer_output[6709] + last_layer_output[6710] + last_layer_output[6711] + last_layer_output[6712] + last_layer_output[6713] + last_layer_output[6714] + last_layer_output[6715] + last_layer_output[6716] + last_layer_output[6717] + last_layer_output[6718] + last_layer_output[6719] + last_layer_output[6720] + last_layer_output[6721] + last_layer_output[6722] + last_layer_output[6723] + last_layer_output[6724] + last_layer_output[6725] + last_layer_output[6726] + last_layer_output[6727] + last_layer_output[6728] + last_layer_output[6729] + last_layer_output[6730] + last_layer_output[6731] + last_layer_output[6732] + last_layer_output[6733] + last_layer_output[6734] + last_layer_output[6735] + last_layer_output[6736] + last_layer_output[6737] + last_layer_output[6738] + last_layer_output[6739] + last_layer_output[6740] + last_layer_output[6741] + last_layer_output[6742] + last_layer_output[6743] + last_layer_output[6744] + last_layer_output[6745] + last_layer_output[6746] + last_layer_output[6747] + last_layer_output[6748] + last_layer_output[6749] + last_layer_output[6750] + last_layer_output[6751] + last_layer_output[6752] + last_layer_output[6753] + last_layer_output[6754] + last_layer_output[6755] + last_layer_output[6756] + last_layer_output[6757] + last_layer_output[6758] + last_layer_output[6759] + last_layer_output[6760] + last_layer_output[6761] + last_layer_output[6762] + last_layer_output[6763] + last_layer_output[6764] + last_layer_output[6765] + last_layer_output[6766] + last_layer_output[6767] + last_layer_output[6768] + last_layer_output[6769] + last_layer_output[6770] + last_layer_output[6771] + last_layer_output[6772] + last_layer_output[6773] + last_layer_output[6774] + last_layer_output[6775] + last_layer_output[6776] + last_layer_output[6777] + last_layer_output[6778] + last_layer_output[6779] + last_layer_output[6780] + last_layer_output[6781] + last_layer_output[6782] + last_layer_output[6783] + last_layer_output[6784] + last_layer_output[6785] + last_layer_output[6786] + last_layer_output[6787] + last_layer_output[6788] + last_layer_output[6789] + last_layer_output[6790] + last_layer_output[6791] + last_layer_output[6792] + last_layer_output[6793] + last_layer_output[6794] + last_layer_output[6795] + last_layer_output[6796] + last_layer_output[6797] + last_layer_output[6798] + last_layer_output[6799] + last_layer_output[6800] + last_layer_output[6801] + last_layer_output[6802] + last_layer_output[6803] + last_layer_output[6804] + last_layer_output[6805] + last_layer_output[6806] + last_layer_output[6807] + last_layer_output[6808] + last_layer_output[6809] + last_layer_output[6810] + last_layer_output[6811] + last_layer_output[6812] + last_layer_output[6813] + last_layer_output[6814] + last_layer_output[6815] + last_layer_output[6816] + last_layer_output[6817] + last_layer_output[6818] + last_layer_output[6819] + last_layer_output[6820] + last_layer_output[6821] + last_layer_output[6822] + last_layer_output[6823] + last_layer_output[6824] + last_layer_output[6825] + last_layer_output[6826] + last_layer_output[6827] + last_layer_output[6828] + last_layer_output[6829] + last_layer_output[6830] + last_layer_output[6831] + last_layer_output[6832] + last_layer_output[6833] + last_layer_output[6834] + last_layer_output[6835] + last_layer_output[6836] + last_layer_output[6837] + last_layer_output[6838] + last_layer_output[6839] + last_layer_output[6840] + last_layer_output[6841] + last_layer_output[6842] + last_layer_output[6843] + last_layer_output[6844] + last_layer_output[6845] + last_layer_output[6846] + last_layer_output[6847] + last_layer_output[6848] + last_layer_output[6849] + last_layer_output[6850] + last_layer_output[6851] + last_layer_output[6852] + last_layer_output[6853] + last_layer_output[6854] + last_layer_output[6855] + last_layer_output[6856] + last_layer_output[6857] + last_layer_output[6858] + last_layer_output[6859] + last_layer_output[6860] + last_layer_output[6861] + last_layer_output[6862] + last_layer_output[6863] + last_layer_output[6864] + last_layer_output[6865] + last_layer_output[6866] + last_layer_output[6867] + last_layer_output[6868] + last_layer_output[6869] + last_layer_output[6870] + last_layer_output[6871] + last_layer_output[6872] + last_layer_output[6873] + last_layer_output[6874] + last_layer_output[6875] + last_layer_output[6876] + last_layer_output[6877] + last_layer_output[6878] + last_layer_output[6879] + last_layer_output[6880] + last_layer_output[6881] + last_layer_output[6882] + last_layer_output[6883] + last_layer_output[6884] + last_layer_output[6885] + last_layer_output[6886] + last_layer_output[6887] + last_layer_output[6888] + last_layer_output[6889] + last_layer_output[6890] + last_layer_output[6891] + last_layer_output[6892] + last_layer_output[6893] + last_layer_output[6894] + last_layer_output[6895] + last_layer_output[6896] + last_layer_output[6897] + last_layer_output[6898] + last_layer_output[6899] + last_layer_output[6900] + last_layer_output[6901] + last_layer_output[6902] + last_layer_output[6903] + last_layer_output[6904] + last_layer_output[6905] + last_layer_output[6906] + last_layer_output[6907] + last_layer_output[6908] + last_layer_output[6909] + last_layer_output[6910] + last_layer_output[6911] + last_layer_output[6912] + last_layer_output[6913] + last_layer_output[6914] + last_layer_output[6915] + last_layer_output[6916] + last_layer_output[6917] + last_layer_output[6918] + last_layer_output[6919] + last_layer_output[6920] + last_layer_output[6921] + last_layer_output[6922] + last_layer_output[6923] + last_layer_output[6924] + last_layer_output[6925] + last_layer_output[6926] + last_layer_output[6927] + last_layer_output[6928] + last_layer_output[6929] + last_layer_output[6930] + last_layer_output[6931] + last_layer_output[6932] + last_layer_output[6933] + last_layer_output[6934] + last_layer_output[6935] + last_layer_output[6936] + last_layer_output[6937] + last_layer_output[6938] + last_layer_output[6939] + last_layer_output[6940] + last_layer_output[6941] + last_layer_output[6942] + last_layer_output[6943] + last_layer_output[6944] + last_layer_output[6945] + last_layer_output[6946] + last_layer_output[6947] + last_layer_output[6948] + last_layer_output[6949] + last_layer_output[6950] + last_layer_output[6951] + last_layer_output[6952] + last_layer_output[6953] + last_layer_output[6954] + last_layer_output[6955] + last_layer_output[6956] + last_layer_output[6957] + last_layer_output[6958] + last_layer_output[6959] + last_layer_output[6960] + last_layer_output[6961] + last_layer_output[6962] + last_layer_output[6963] + last_layer_output[6964] + last_layer_output[6965] + last_layer_output[6966] + last_layer_output[6967] + last_layer_output[6968] + last_layer_output[6969] + last_layer_output[6970] + last_layer_output[6971] + last_layer_output[6972] + last_layer_output[6973] + last_layer_output[6974] + last_layer_output[6975] + last_layer_output[6976] + last_layer_output[6977] + last_layer_output[6978] + last_layer_output[6979] + last_layer_output[6980] + last_layer_output[6981] + last_layer_output[6982] + last_layer_output[6983] + last_layer_output[6984] + last_layer_output[6985] + last_layer_output[6986] + last_layer_output[6987] + last_layer_output[6988] + last_layer_output[6989] + last_layer_output[6990] + last_layer_output[6991] + last_layer_output[6992] + last_layer_output[6993] + last_layer_output[6994] + last_layer_output[6995] + last_layer_output[6996] + last_layer_output[6997] + last_layer_output[6998] + last_layer_output[6999] + last_layer_output[7000] + last_layer_output[7001] + last_layer_output[7002] + last_layer_output[7003] + last_layer_output[7004] + last_layer_output[7005] + last_layer_output[7006] + last_layer_output[7007] + last_layer_output[7008] + last_layer_output[7009] + last_layer_output[7010] + last_layer_output[7011] + last_layer_output[7012] + last_layer_output[7013] + last_layer_output[7014] + last_layer_output[7015] + last_layer_output[7016] + last_layer_output[7017] + last_layer_output[7018] + last_layer_output[7019] + last_layer_output[7020] + last_layer_output[7021] + last_layer_output[7022] + last_layer_output[7023] + last_layer_output[7024] + last_layer_output[7025] + last_layer_output[7026] + last_layer_output[7027] + last_layer_output[7028] + last_layer_output[7029] + last_layer_output[7030] + last_layer_output[7031] + last_layer_output[7032] + last_layer_output[7033] + last_layer_output[7034] + last_layer_output[7035] + last_layer_output[7036] + last_layer_output[7037] + last_layer_output[7038] + last_layer_output[7039] + last_layer_output[7040] + last_layer_output[7041] + last_layer_output[7042] + last_layer_output[7043] + last_layer_output[7044] + last_layer_output[7045] + last_layer_output[7046] + last_layer_output[7047] + last_layer_output[7048] + last_layer_output[7049] + last_layer_output[7050] + last_layer_output[7051] + last_layer_output[7052] + last_layer_output[7053] + last_layer_output[7054] + last_layer_output[7055] + last_layer_output[7056] + last_layer_output[7057] + last_layer_output[7058] + last_layer_output[7059] + last_layer_output[7060] + last_layer_output[7061] + last_layer_output[7062] + last_layer_output[7063] + last_layer_output[7064] + last_layer_output[7065] + last_layer_output[7066] + last_layer_output[7067] + last_layer_output[7068] + last_layer_output[7069] + last_layer_output[7070] + last_layer_output[7071] + last_layer_output[7072] + last_layer_output[7073] + last_layer_output[7074] + last_layer_output[7075] + last_layer_output[7076] + last_layer_output[7077] + last_layer_output[7078] + last_layer_output[7079] + last_layer_output[7080] + last_layer_output[7081] + last_layer_output[7082] + last_layer_output[7083] + last_layer_output[7084] + last_layer_output[7085] + last_layer_output[7086] + last_layer_output[7087] + last_layer_output[7088] + last_layer_output[7089] + last_layer_output[7090] + last_layer_output[7091] + last_layer_output[7092] + last_layer_output[7093] + last_layer_output[7094] + last_layer_output[7095] + last_layer_output[7096] + last_layer_output[7097] + last_layer_output[7098] + last_layer_output[7099] + last_layer_output[7100] + last_layer_output[7101] + last_layer_output[7102] + last_layer_output[7103] + last_layer_output[7104] + last_layer_output[7105] + last_layer_output[7106] + last_layer_output[7107] + last_layer_output[7108] + last_layer_output[7109] + last_layer_output[7110] + last_layer_output[7111] + last_layer_output[7112] + last_layer_output[7113] + last_layer_output[7114] + last_layer_output[7115] + last_layer_output[7116] + last_layer_output[7117] + last_layer_output[7118] + last_layer_output[7119] + last_layer_output[7120] + last_layer_output[7121] + last_layer_output[7122] + last_layer_output[7123] + last_layer_output[7124] + last_layer_output[7125] + last_layer_output[7126] + last_layer_output[7127] + last_layer_output[7128] + last_layer_output[7129] + last_layer_output[7130] + last_layer_output[7131] + last_layer_output[7132] + last_layer_output[7133] + last_layer_output[7134] + last_layer_output[7135] + last_layer_output[7136] + last_layer_output[7137] + last_layer_output[7138] + last_layer_output[7139] + last_layer_output[7140] + last_layer_output[7141] + last_layer_output[7142] + last_layer_output[7143] + last_layer_output[7144] + last_layer_output[7145] + last_layer_output[7146] + last_layer_output[7147] + last_layer_output[7148] + last_layer_output[7149] + last_layer_output[7150] + last_layer_output[7151] + last_layer_output[7152] + last_layer_output[7153] + last_layer_output[7154] + last_layer_output[7155] + last_layer_output[7156] + last_layer_output[7157] + last_layer_output[7158] + last_layer_output[7159] + last_layer_output[7160] + last_layer_output[7161] + last_layer_output[7162] + last_layer_output[7163] + last_layer_output[7164] + last_layer_output[7165] + last_layer_output[7166] + last_layer_output[7167] + last_layer_output[7168] + last_layer_output[7169] + last_layer_output[7170] + last_layer_output[7171] + last_layer_output[7172] + last_layer_output[7173] + last_layer_output[7174] + last_layer_output[7175] + last_layer_output[7176] + last_layer_output[7177] + last_layer_output[7178] + last_layer_output[7179] + last_layer_output[7180] + last_layer_output[7181] + last_layer_output[7182] + last_layer_output[7183] + last_layer_output[7184] + last_layer_output[7185] + last_layer_output[7186] + last_layer_output[7187] + last_layer_output[7188] + last_layer_output[7189] + last_layer_output[7190] + last_layer_output[7191] + last_layer_output[7192] + last_layer_output[7193] + last_layer_output[7194] + last_layer_output[7195] + last_layer_output[7196] + last_layer_output[7197] + last_layer_output[7198] + last_layer_output[7199];
      result[6] <= last_layer_output[7200] + last_layer_output[7201] + last_layer_output[7202] + last_layer_output[7203] + last_layer_output[7204] + last_layer_output[7205] + last_layer_output[7206] + last_layer_output[7207] + last_layer_output[7208] + last_layer_output[7209] + last_layer_output[7210] + last_layer_output[7211] + last_layer_output[7212] + last_layer_output[7213] + last_layer_output[7214] + last_layer_output[7215] + last_layer_output[7216] + last_layer_output[7217] + last_layer_output[7218] + last_layer_output[7219] + last_layer_output[7220] + last_layer_output[7221] + last_layer_output[7222] + last_layer_output[7223] + last_layer_output[7224] + last_layer_output[7225] + last_layer_output[7226] + last_layer_output[7227] + last_layer_output[7228] + last_layer_output[7229] + last_layer_output[7230] + last_layer_output[7231] + last_layer_output[7232] + last_layer_output[7233] + last_layer_output[7234] + last_layer_output[7235] + last_layer_output[7236] + last_layer_output[7237] + last_layer_output[7238] + last_layer_output[7239] + last_layer_output[7240] + last_layer_output[7241] + last_layer_output[7242] + last_layer_output[7243] + last_layer_output[7244] + last_layer_output[7245] + last_layer_output[7246] + last_layer_output[7247] + last_layer_output[7248] + last_layer_output[7249] + last_layer_output[7250] + last_layer_output[7251] + last_layer_output[7252] + last_layer_output[7253] + last_layer_output[7254] + last_layer_output[7255] + last_layer_output[7256] + last_layer_output[7257] + last_layer_output[7258] + last_layer_output[7259] + last_layer_output[7260] + last_layer_output[7261] + last_layer_output[7262] + last_layer_output[7263] + last_layer_output[7264] + last_layer_output[7265] + last_layer_output[7266] + last_layer_output[7267] + last_layer_output[7268] + last_layer_output[7269] + last_layer_output[7270] + last_layer_output[7271] + last_layer_output[7272] + last_layer_output[7273] + last_layer_output[7274] + last_layer_output[7275] + last_layer_output[7276] + last_layer_output[7277] + last_layer_output[7278] + last_layer_output[7279] + last_layer_output[7280] + last_layer_output[7281] + last_layer_output[7282] + last_layer_output[7283] + last_layer_output[7284] + last_layer_output[7285] + last_layer_output[7286] + last_layer_output[7287] + last_layer_output[7288] + last_layer_output[7289] + last_layer_output[7290] + last_layer_output[7291] + last_layer_output[7292] + last_layer_output[7293] + last_layer_output[7294] + last_layer_output[7295] + last_layer_output[7296] + last_layer_output[7297] + last_layer_output[7298] + last_layer_output[7299] + last_layer_output[7300] + last_layer_output[7301] + last_layer_output[7302] + last_layer_output[7303] + last_layer_output[7304] + last_layer_output[7305] + last_layer_output[7306] + last_layer_output[7307] + last_layer_output[7308] + last_layer_output[7309] + last_layer_output[7310] + last_layer_output[7311] + last_layer_output[7312] + last_layer_output[7313] + last_layer_output[7314] + last_layer_output[7315] + last_layer_output[7316] + last_layer_output[7317] + last_layer_output[7318] + last_layer_output[7319] + last_layer_output[7320] + last_layer_output[7321] + last_layer_output[7322] + last_layer_output[7323] + last_layer_output[7324] + last_layer_output[7325] + last_layer_output[7326] + last_layer_output[7327] + last_layer_output[7328] + last_layer_output[7329] + last_layer_output[7330] + last_layer_output[7331] + last_layer_output[7332] + last_layer_output[7333] + last_layer_output[7334] + last_layer_output[7335] + last_layer_output[7336] + last_layer_output[7337] + last_layer_output[7338] + last_layer_output[7339] + last_layer_output[7340] + last_layer_output[7341] + last_layer_output[7342] + last_layer_output[7343] + last_layer_output[7344] + last_layer_output[7345] + last_layer_output[7346] + last_layer_output[7347] + last_layer_output[7348] + last_layer_output[7349] + last_layer_output[7350] + last_layer_output[7351] + last_layer_output[7352] + last_layer_output[7353] + last_layer_output[7354] + last_layer_output[7355] + last_layer_output[7356] + last_layer_output[7357] + last_layer_output[7358] + last_layer_output[7359] + last_layer_output[7360] + last_layer_output[7361] + last_layer_output[7362] + last_layer_output[7363] + last_layer_output[7364] + last_layer_output[7365] + last_layer_output[7366] + last_layer_output[7367] + last_layer_output[7368] + last_layer_output[7369] + last_layer_output[7370] + last_layer_output[7371] + last_layer_output[7372] + last_layer_output[7373] + last_layer_output[7374] + last_layer_output[7375] + last_layer_output[7376] + last_layer_output[7377] + last_layer_output[7378] + last_layer_output[7379] + last_layer_output[7380] + last_layer_output[7381] + last_layer_output[7382] + last_layer_output[7383] + last_layer_output[7384] + last_layer_output[7385] + last_layer_output[7386] + last_layer_output[7387] + last_layer_output[7388] + last_layer_output[7389] + last_layer_output[7390] + last_layer_output[7391] + last_layer_output[7392] + last_layer_output[7393] + last_layer_output[7394] + last_layer_output[7395] + last_layer_output[7396] + last_layer_output[7397] + last_layer_output[7398] + last_layer_output[7399] + last_layer_output[7400] + last_layer_output[7401] + last_layer_output[7402] + last_layer_output[7403] + last_layer_output[7404] + last_layer_output[7405] + last_layer_output[7406] + last_layer_output[7407] + last_layer_output[7408] + last_layer_output[7409] + last_layer_output[7410] + last_layer_output[7411] + last_layer_output[7412] + last_layer_output[7413] + last_layer_output[7414] + last_layer_output[7415] + last_layer_output[7416] + last_layer_output[7417] + last_layer_output[7418] + last_layer_output[7419] + last_layer_output[7420] + last_layer_output[7421] + last_layer_output[7422] + last_layer_output[7423] + last_layer_output[7424] + last_layer_output[7425] + last_layer_output[7426] + last_layer_output[7427] + last_layer_output[7428] + last_layer_output[7429] + last_layer_output[7430] + last_layer_output[7431] + last_layer_output[7432] + last_layer_output[7433] + last_layer_output[7434] + last_layer_output[7435] + last_layer_output[7436] + last_layer_output[7437] + last_layer_output[7438] + last_layer_output[7439] + last_layer_output[7440] + last_layer_output[7441] + last_layer_output[7442] + last_layer_output[7443] + last_layer_output[7444] + last_layer_output[7445] + last_layer_output[7446] + last_layer_output[7447] + last_layer_output[7448] + last_layer_output[7449] + last_layer_output[7450] + last_layer_output[7451] + last_layer_output[7452] + last_layer_output[7453] + last_layer_output[7454] + last_layer_output[7455] + last_layer_output[7456] + last_layer_output[7457] + last_layer_output[7458] + last_layer_output[7459] + last_layer_output[7460] + last_layer_output[7461] + last_layer_output[7462] + last_layer_output[7463] + last_layer_output[7464] + last_layer_output[7465] + last_layer_output[7466] + last_layer_output[7467] + last_layer_output[7468] + last_layer_output[7469] + last_layer_output[7470] + last_layer_output[7471] + last_layer_output[7472] + last_layer_output[7473] + last_layer_output[7474] + last_layer_output[7475] + last_layer_output[7476] + last_layer_output[7477] + last_layer_output[7478] + last_layer_output[7479] + last_layer_output[7480] + last_layer_output[7481] + last_layer_output[7482] + last_layer_output[7483] + last_layer_output[7484] + last_layer_output[7485] + last_layer_output[7486] + last_layer_output[7487] + last_layer_output[7488] + last_layer_output[7489] + last_layer_output[7490] + last_layer_output[7491] + last_layer_output[7492] + last_layer_output[7493] + last_layer_output[7494] + last_layer_output[7495] + last_layer_output[7496] + last_layer_output[7497] + last_layer_output[7498] + last_layer_output[7499] + last_layer_output[7500] + last_layer_output[7501] + last_layer_output[7502] + last_layer_output[7503] + last_layer_output[7504] + last_layer_output[7505] + last_layer_output[7506] + last_layer_output[7507] + last_layer_output[7508] + last_layer_output[7509] + last_layer_output[7510] + last_layer_output[7511] + last_layer_output[7512] + last_layer_output[7513] + last_layer_output[7514] + last_layer_output[7515] + last_layer_output[7516] + last_layer_output[7517] + last_layer_output[7518] + last_layer_output[7519] + last_layer_output[7520] + last_layer_output[7521] + last_layer_output[7522] + last_layer_output[7523] + last_layer_output[7524] + last_layer_output[7525] + last_layer_output[7526] + last_layer_output[7527] + last_layer_output[7528] + last_layer_output[7529] + last_layer_output[7530] + last_layer_output[7531] + last_layer_output[7532] + last_layer_output[7533] + last_layer_output[7534] + last_layer_output[7535] + last_layer_output[7536] + last_layer_output[7537] + last_layer_output[7538] + last_layer_output[7539] + last_layer_output[7540] + last_layer_output[7541] + last_layer_output[7542] + last_layer_output[7543] + last_layer_output[7544] + last_layer_output[7545] + last_layer_output[7546] + last_layer_output[7547] + last_layer_output[7548] + last_layer_output[7549] + last_layer_output[7550] + last_layer_output[7551] + last_layer_output[7552] + last_layer_output[7553] + last_layer_output[7554] + last_layer_output[7555] + last_layer_output[7556] + last_layer_output[7557] + last_layer_output[7558] + last_layer_output[7559] + last_layer_output[7560] + last_layer_output[7561] + last_layer_output[7562] + last_layer_output[7563] + last_layer_output[7564] + last_layer_output[7565] + last_layer_output[7566] + last_layer_output[7567] + last_layer_output[7568] + last_layer_output[7569] + last_layer_output[7570] + last_layer_output[7571] + last_layer_output[7572] + last_layer_output[7573] + last_layer_output[7574] + last_layer_output[7575] + last_layer_output[7576] + last_layer_output[7577] + last_layer_output[7578] + last_layer_output[7579] + last_layer_output[7580] + last_layer_output[7581] + last_layer_output[7582] + last_layer_output[7583] + last_layer_output[7584] + last_layer_output[7585] + last_layer_output[7586] + last_layer_output[7587] + last_layer_output[7588] + last_layer_output[7589] + last_layer_output[7590] + last_layer_output[7591] + last_layer_output[7592] + last_layer_output[7593] + last_layer_output[7594] + last_layer_output[7595] + last_layer_output[7596] + last_layer_output[7597] + last_layer_output[7598] + last_layer_output[7599] + last_layer_output[7600] + last_layer_output[7601] + last_layer_output[7602] + last_layer_output[7603] + last_layer_output[7604] + last_layer_output[7605] + last_layer_output[7606] + last_layer_output[7607] + last_layer_output[7608] + last_layer_output[7609] + last_layer_output[7610] + last_layer_output[7611] + last_layer_output[7612] + last_layer_output[7613] + last_layer_output[7614] + last_layer_output[7615] + last_layer_output[7616] + last_layer_output[7617] + last_layer_output[7618] + last_layer_output[7619] + last_layer_output[7620] + last_layer_output[7621] + last_layer_output[7622] + last_layer_output[7623] + last_layer_output[7624] + last_layer_output[7625] + last_layer_output[7626] + last_layer_output[7627] + last_layer_output[7628] + last_layer_output[7629] + last_layer_output[7630] + last_layer_output[7631] + last_layer_output[7632] + last_layer_output[7633] + last_layer_output[7634] + last_layer_output[7635] + last_layer_output[7636] + last_layer_output[7637] + last_layer_output[7638] + last_layer_output[7639] + last_layer_output[7640] + last_layer_output[7641] + last_layer_output[7642] + last_layer_output[7643] + last_layer_output[7644] + last_layer_output[7645] + last_layer_output[7646] + last_layer_output[7647] + last_layer_output[7648] + last_layer_output[7649] + last_layer_output[7650] + last_layer_output[7651] + last_layer_output[7652] + last_layer_output[7653] + last_layer_output[7654] + last_layer_output[7655] + last_layer_output[7656] + last_layer_output[7657] + last_layer_output[7658] + last_layer_output[7659] + last_layer_output[7660] + last_layer_output[7661] + last_layer_output[7662] + last_layer_output[7663] + last_layer_output[7664] + last_layer_output[7665] + last_layer_output[7666] + last_layer_output[7667] + last_layer_output[7668] + last_layer_output[7669] + last_layer_output[7670] + last_layer_output[7671] + last_layer_output[7672] + last_layer_output[7673] + last_layer_output[7674] + last_layer_output[7675] + last_layer_output[7676] + last_layer_output[7677] + last_layer_output[7678] + last_layer_output[7679] + last_layer_output[7680] + last_layer_output[7681] + last_layer_output[7682] + last_layer_output[7683] + last_layer_output[7684] + last_layer_output[7685] + last_layer_output[7686] + last_layer_output[7687] + last_layer_output[7688] + last_layer_output[7689] + last_layer_output[7690] + last_layer_output[7691] + last_layer_output[7692] + last_layer_output[7693] + last_layer_output[7694] + last_layer_output[7695] + last_layer_output[7696] + last_layer_output[7697] + last_layer_output[7698] + last_layer_output[7699] + last_layer_output[7700] + last_layer_output[7701] + last_layer_output[7702] + last_layer_output[7703] + last_layer_output[7704] + last_layer_output[7705] + last_layer_output[7706] + last_layer_output[7707] + last_layer_output[7708] + last_layer_output[7709] + last_layer_output[7710] + last_layer_output[7711] + last_layer_output[7712] + last_layer_output[7713] + last_layer_output[7714] + last_layer_output[7715] + last_layer_output[7716] + last_layer_output[7717] + last_layer_output[7718] + last_layer_output[7719] + last_layer_output[7720] + last_layer_output[7721] + last_layer_output[7722] + last_layer_output[7723] + last_layer_output[7724] + last_layer_output[7725] + last_layer_output[7726] + last_layer_output[7727] + last_layer_output[7728] + last_layer_output[7729] + last_layer_output[7730] + last_layer_output[7731] + last_layer_output[7732] + last_layer_output[7733] + last_layer_output[7734] + last_layer_output[7735] + last_layer_output[7736] + last_layer_output[7737] + last_layer_output[7738] + last_layer_output[7739] + last_layer_output[7740] + last_layer_output[7741] + last_layer_output[7742] + last_layer_output[7743] + last_layer_output[7744] + last_layer_output[7745] + last_layer_output[7746] + last_layer_output[7747] + last_layer_output[7748] + last_layer_output[7749] + last_layer_output[7750] + last_layer_output[7751] + last_layer_output[7752] + last_layer_output[7753] + last_layer_output[7754] + last_layer_output[7755] + last_layer_output[7756] + last_layer_output[7757] + last_layer_output[7758] + last_layer_output[7759] + last_layer_output[7760] + last_layer_output[7761] + last_layer_output[7762] + last_layer_output[7763] + last_layer_output[7764] + last_layer_output[7765] + last_layer_output[7766] + last_layer_output[7767] + last_layer_output[7768] + last_layer_output[7769] + last_layer_output[7770] + last_layer_output[7771] + last_layer_output[7772] + last_layer_output[7773] + last_layer_output[7774] + last_layer_output[7775] + last_layer_output[7776] + last_layer_output[7777] + last_layer_output[7778] + last_layer_output[7779] + last_layer_output[7780] + last_layer_output[7781] + last_layer_output[7782] + last_layer_output[7783] + last_layer_output[7784] + last_layer_output[7785] + last_layer_output[7786] + last_layer_output[7787] + last_layer_output[7788] + last_layer_output[7789] + last_layer_output[7790] + last_layer_output[7791] + last_layer_output[7792] + last_layer_output[7793] + last_layer_output[7794] + last_layer_output[7795] + last_layer_output[7796] + last_layer_output[7797] + last_layer_output[7798] + last_layer_output[7799] + last_layer_output[7800] + last_layer_output[7801] + last_layer_output[7802] + last_layer_output[7803] + last_layer_output[7804] + last_layer_output[7805] + last_layer_output[7806] + last_layer_output[7807] + last_layer_output[7808] + last_layer_output[7809] + last_layer_output[7810] + last_layer_output[7811] + last_layer_output[7812] + last_layer_output[7813] + last_layer_output[7814] + last_layer_output[7815] + last_layer_output[7816] + last_layer_output[7817] + last_layer_output[7818] + last_layer_output[7819] + last_layer_output[7820] + last_layer_output[7821] + last_layer_output[7822] + last_layer_output[7823] + last_layer_output[7824] + last_layer_output[7825] + last_layer_output[7826] + last_layer_output[7827] + last_layer_output[7828] + last_layer_output[7829] + last_layer_output[7830] + last_layer_output[7831] + last_layer_output[7832] + last_layer_output[7833] + last_layer_output[7834] + last_layer_output[7835] + last_layer_output[7836] + last_layer_output[7837] + last_layer_output[7838] + last_layer_output[7839] + last_layer_output[7840] + last_layer_output[7841] + last_layer_output[7842] + last_layer_output[7843] + last_layer_output[7844] + last_layer_output[7845] + last_layer_output[7846] + last_layer_output[7847] + last_layer_output[7848] + last_layer_output[7849] + last_layer_output[7850] + last_layer_output[7851] + last_layer_output[7852] + last_layer_output[7853] + last_layer_output[7854] + last_layer_output[7855] + last_layer_output[7856] + last_layer_output[7857] + last_layer_output[7858] + last_layer_output[7859] + last_layer_output[7860] + last_layer_output[7861] + last_layer_output[7862] + last_layer_output[7863] + last_layer_output[7864] + last_layer_output[7865] + last_layer_output[7866] + last_layer_output[7867] + last_layer_output[7868] + last_layer_output[7869] + last_layer_output[7870] + last_layer_output[7871] + last_layer_output[7872] + last_layer_output[7873] + last_layer_output[7874] + last_layer_output[7875] + last_layer_output[7876] + last_layer_output[7877] + last_layer_output[7878] + last_layer_output[7879] + last_layer_output[7880] + last_layer_output[7881] + last_layer_output[7882] + last_layer_output[7883] + last_layer_output[7884] + last_layer_output[7885] + last_layer_output[7886] + last_layer_output[7887] + last_layer_output[7888] + last_layer_output[7889] + last_layer_output[7890] + last_layer_output[7891] + last_layer_output[7892] + last_layer_output[7893] + last_layer_output[7894] + last_layer_output[7895] + last_layer_output[7896] + last_layer_output[7897] + last_layer_output[7898] + last_layer_output[7899] + last_layer_output[7900] + last_layer_output[7901] + last_layer_output[7902] + last_layer_output[7903] + last_layer_output[7904] + last_layer_output[7905] + last_layer_output[7906] + last_layer_output[7907] + last_layer_output[7908] + last_layer_output[7909] + last_layer_output[7910] + last_layer_output[7911] + last_layer_output[7912] + last_layer_output[7913] + last_layer_output[7914] + last_layer_output[7915] + last_layer_output[7916] + last_layer_output[7917] + last_layer_output[7918] + last_layer_output[7919] + last_layer_output[7920] + last_layer_output[7921] + last_layer_output[7922] + last_layer_output[7923] + last_layer_output[7924] + last_layer_output[7925] + last_layer_output[7926] + last_layer_output[7927] + last_layer_output[7928] + last_layer_output[7929] + last_layer_output[7930] + last_layer_output[7931] + last_layer_output[7932] + last_layer_output[7933] + last_layer_output[7934] + last_layer_output[7935] + last_layer_output[7936] + last_layer_output[7937] + last_layer_output[7938] + last_layer_output[7939] + last_layer_output[7940] + last_layer_output[7941] + last_layer_output[7942] + last_layer_output[7943] + last_layer_output[7944] + last_layer_output[7945] + last_layer_output[7946] + last_layer_output[7947] + last_layer_output[7948] + last_layer_output[7949] + last_layer_output[7950] + last_layer_output[7951] + last_layer_output[7952] + last_layer_output[7953] + last_layer_output[7954] + last_layer_output[7955] + last_layer_output[7956] + last_layer_output[7957] + last_layer_output[7958] + last_layer_output[7959] + last_layer_output[7960] + last_layer_output[7961] + last_layer_output[7962] + last_layer_output[7963] + last_layer_output[7964] + last_layer_output[7965] + last_layer_output[7966] + last_layer_output[7967] + last_layer_output[7968] + last_layer_output[7969] + last_layer_output[7970] + last_layer_output[7971] + last_layer_output[7972] + last_layer_output[7973] + last_layer_output[7974] + last_layer_output[7975] + last_layer_output[7976] + last_layer_output[7977] + last_layer_output[7978] + last_layer_output[7979] + last_layer_output[7980] + last_layer_output[7981] + last_layer_output[7982] + last_layer_output[7983] + last_layer_output[7984] + last_layer_output[7985] + last_layer_output[7986] + last_layer_output[7987] + last_layer_output[7988] + last_layer_output[7989] + last_layer_output[7990] + last_layer_output[7991] + last_layer_output[7992] + last_layer_output[7993] + last_layer_output[7994] + last_layer_output[7995] + last_layer_output[7996] + last_layer_output[7997] + last_layer_output[7998] + last_layer_output[7999] + last_layer_output[8000] + last_layer_output[8001] + last_layer_output[8002] + last_layer_output[8003] + last_layer_output[8004] + last_layer_output[8005] + last_layer_output[8006] + last_layer_output[8007] + last_layer_output[8008] + last_layer_output[8009] + last_layer_output[8010] + last_layer_output[8011] + last_layer_output[8012] + last_layer_output[8013] + last_layer_output[8014] + last_layer_output[8015] + last_layer_output[8016] + last_layer_output[8017] + last_layer_output[8018] + last_layer_output[8019] + last_layer_output[8020] + last_layer_output[8021] + last_layer_output[8022] + last_layer_output[8023] + last_layer_output[8024] + last_layer_output[8025] + last_layer_output[8026] + last_layer_output[8027] + last_layer_output[8028] + last_layer_output[8029] + last_layer_output[8030] + last_layer_output[8031] + last_layer_output[8032] + last_layer_output[8033] + last_layer_output[8034] + last_layer_output[8035] + last_layer_output[8036] + last_layer_output[8037] + last_layer_output[8038] + last_layer_output[8039] + last_layer_output[8040] + last_layer_output[8041] + last_layer_output[8042] + last_layer_output[8043] + last_layer_output[8044] + last_layer_output[8045] + last_layer_output[8046] + last_layer_output[8047] + last_layer_output[8048] + last_layer_output[8049] + last_layer_output[8050] + last_layer_output[8051] + last_layer_output[8052] + last_layer_output[8053] + last_layer_output[8054] + last_layer_output[8055] + last_layer_output[8056] + last_layer_output[8057] + last_layer_output[8058] + last_layer_output[8059] + last_layer_output[8060] + last_layer_output[8061] + last_layer_output[8062] + last_layer_output[8063] + last_layer_output[8064] + last_layer_output[8065] + last_layer_output[8066] + last_layer_output[8067] + last_layer_output[8068] + last_layer_output[8069] + last_layer_output[8070] + last_layer_output[8071] + last_layer_output[8072] + last_layer_output[8073] + last_layer_output[8074] + last_layer_output[8075] + last_layer_output[8076] + last_layer_output[8077] + last_layer_output[8078] + last_layer_output[8079] + last_layer_output[8080] + last_layer_output[8081] + last_layer_output[8082] + last_layer_output[8083] + last_layer_output[8084] + last_layer_output[8085] + last_layer_output[8086] + last_layer_output[8087] + last_layer_output[8088] + last_layer_output[8089] + last_layer_output[8090] + last_layer_output[8091] + last_layer_output[8092] + last_layer_output[8093] + last_layer_output[8094] + last_layer_output[8095] + last_layer_output[8096] + last_layer_output[8097] + last_layer_output[8098] + last_layer_output[8099] + last_layer_output[8100] + last_layer_output[8101] + last_layer_output[8102] + last_layer_output[8103] + last_layer_output[8104] + last_layer_output[8105] + last_layer_output[8106] + last_layer_output[8107] + last_layer_output[8108] + last_layer_output[8109] + last_layer_output[8110] + last_layer_output[8111] + last_layer_output[8112] + last_layer_output[8113] + last_layer_output[8114] + last_layer_output[8115] + last_layer_output[8116] + last_layer_output[8117] + last_layer_output[8118] + last_layer_output[8119] + last_layer_output[8120] + last_layer_output[8121] + last_layer_output[8122] + last_layer_output[8123] + last_layer_output[8124] + last_layer_output[8125] + last_layer_output[8126] + last_layer_output[8127] + last_layer_output[8128] + last_layer_output[8129] + last_layer_output[8130] + last_layer_output[8131] + last_layer_output[8132] + last_layer_output[8133] + last_layer_output[8134] + last_layer_output[8135] + last_layer_output[8136] + last_layer_output[8137] + last_layer_output[8138] + last_layer_output[8139] + last_layer_output[8140] + last_layer_output[8141] + last_layer_output[8142] + last_layer_output[8143] + last_layer_output[8144] + last_layer_output[8145] + last_layer_output[8146] + last_layer_output[8147] + last_layer_output[8148] + last_layer_output[8149] + last_layer_output[8150] + last_layer_output[8151] + last_layer_output[8152] + last_layer_output[8153] + last_layer_output[8154] + last_layer_output[8155] + last_layer_output[8156] + last_layer_output[8157] + last_layer_output[8158] + last_layer_output[8159] + last_layer_output[8160] + last_layer_output[8161] + last_layer_output[8162] + last_layer_output[8163] + last_layer_output[8164] + last_layer_output[8165] + last_layer_output[8166] + last_layer_output[8167] + last_layer_output[8168] + last_layer_output[8169] + last_layer_output[8170] + last_layer_output[8171] + last_layer_output[8172] + last_layer_output[8173] + last_layer_output[8174] + last_layer_output[8175] + last_layer_output[8176] + last_layer_output[8177] + last_layer_output[8178] + last_layer_output[8179] + last_layer_output[8180] + last_layer_output[8181] + last_layer_output[8182] + last_layer_output[8183] + last_layer_output[8184] + last_layer_output[8185] + last_layer_output[8186] + last_layer_output[8187] + last_layer_output[8188] + last_layer_output[8189] + last_layer_output[8190] + last_layer_output[8191] + last_layer_output[8192] + last_layer_output[8193] + last_layer_output[8194] + last_layer_output[8195] + last_layer_output[8196] + last_layer_output[8197] + last_layer_output[8198] + last_layer_output[8199] + last_layer_output[8200] + last_layer_output[8201] + last_layer_output[8202] + last_layer_output[8203] + last_layer_output[8204] + last_layer_output[8205] + last_layer_output[8206] + last_layer_output[8207] + last_layer_output[8208] + last_layer_output[8209] + last_layer_output[8210] + last_layer_output[8211] + last_layer_output[8212] + last_layer_output[8213] + last_layer_output[8214] + last_layer_output[8215] + last_layer_output[8216] + last_layer_output[8217] + last_layer_output[8218] + last_layer_output[8219] + last_layer_output[8220] + last_layer_output[8221] + last_layer_output[8222] + last_layer_output[8223] + last_layer_output[8224] + last_layer_output[8225] + last_layer_output[8226] + last_layer_output[8227] + last_layer_output[8228] + last_layer_output[8229] + last_layer_output[8230] + last_layer_output[8231] + last_layer_output[8232] + last_layer_output[8233] + last_layer_output[8234] + last_layer_output[8235] + last_layer_output[8236] + last_layer_output[8237] + last_layer_output[8238] + last_layer_output[8239] + last_layer_output[8240] + last_layer_output[8241] + last_layer_output[8242] + last_layer_output[8243] + last_layer_output[8244] + last_layer_output[8245] + last_layer_output[8246] + last_layer_output[8247] + last_layer_output[8248] + last_layer_output[8249] + last_layer_output[8250] + last_layer_output[8251] + last_layer_output[8252] + last_layer_output[8253] + last_layer_output[8254] + last_layer_output[8255] + last_layer_output[8256] + last_layer_output[8257] + last_layer_output[8258] + last_layer_output[8259] + last_layer_output[8260] + last_layer_output[8261] + last_layer_output[8262] + last_layer_output[8263] + last_layer_output[8264] + last_layer_output[8265] + last_layer_output[8266] + last_layer_output[8267] + last_layer_output[8268] + last_layer_output[8269] + last_layer_output[8270] + last_layer_output[8271] + last_layer_output[8272] + last_layer_output[8273] + last_layer_output[8274] + last_layer_output[8275] + last_layer_output[8276] + last_layer_output[8277] + last_layer_output[8278] + last_layer_output[8279] + last_layer_output[8280] + last_layer_output[8281] + last_layer_output[8282] + last_layer_output[8283] + last_layer_output[8284] + last_layer_output[8285] + last_layer_output[8286] + last_layer_output[8287] + last_layer_output[8288] + last_layer_output[8289] + last_layer_output[8290] + last_layer_output[8291] + last_layer_output[8292] + last_layer_output[8293] + last_layer_output[8294] + last_layer_output[8295] + last_layer_output[8296] + last_layer_output[8297] + last_layer_output[8298] + last_layer_output[8299] + last_layer_output[8300] + last_layer_output[8301] + last_layer_output[8302] + last_layer_output[8303] + last_layer_output[8304] + last_layer_output[8305] + last_layer_output[8306] + last_layer_output[8307] + last_layer_output[8308] + last_layer_output[8309] + last_layer_output[8310] + last_layer_output[8311] + last_layer_output[8312] + last_layer_output[8313] + last_layer_output[8314] + last_layer_output[8315] + last_layer_output[8316] + last_layer_output[8317] + last_layer_output[8318] + last_layer_output[8319] + last_layer_output[8320] + last_layer_output[8321] + last_layer_output[8322] + last_layer_output[8323] + last_layer_output[8324] + last_layer_output[8325] + last_layer_output[8326] + last_layer_output[8327] + last_layer_output[8328] + last_layer_output[8329] + last_layer_output[8330] + last_layer_output[8331] + last_layer_output[8332] + last_layer_output[8333] + last_layer_output[8334] + last_layer_output[8335] + last_layer_output[8336] + last_layer_output[8337] + last_layer_output[8338] + last_layer_output[8339] + last_layer_output[8340] + last_layer_output[8341] + last_layer_output[8342] + last_layer_output[8343] + last_layer_output[8344] + last_layer_output[8345] + last_layer_output[8346] + last_layer_output[8347] + last_layer_output[8348] + last_layer_output[8349] + last_layer_output[8350] + last_layer_output[8351] + last_layer_output[8352] + last_layer_output[8353] + last_layer_output[8354] + last_layer_output[8355] + last_layer_output[8356] + last_layer_output[8357] + last_layer_output[8358] + last_layer_output[8359] + last_layer_output[8360] + last_layer_output[8361] + last_layer_output[8362] + last_layer_output[8363] + last_layer_output[8364] + last_layer_output[8365] + last_layer_output[8366] + last_layer_output[8367] + last_layer_output[8368] + last_layer_output[8369] + last_layer_output[8370] + last_layer_output[8371] + last_layer_output[8372] + last_layer_output[8373] + last_layer_output[8374] + last_layer_output[8375] + last_layer_output[8376] + last_layer_output[8377] + last_layer_output[8378] + last_layer_output[8379] + last_layer_output[8380] + last_layer_output[8381] + last_layer_output[8382] + last_layer_output[8383] + last_layer_output[8384] + last_layer_output[8385] + last_layer_output[8386] + last_layer_output[8387] + last_layer_output[8388] + last_layer_output[8389] + last_layer_output[8390] + last_layer_output[8391] + last_layer_output[8392] + last_layer_output[8393] + last_layer_output[8394] + last_layer_output[8395] + last_layer_output[8396] + last_layer_output[8397] + last_layer_output[8398] + last_layer_output[8399];
      result[7] <= last_layer_output[8400] + last_layer_output[8401] + last_layer_output[8402] + last_layer_output[8403] + last_layer_output[8404] + last_layer_output[8405] + last_layer_output[8406] + last_layer_output[8407] + last_layer_output[8408] + last_layer_output[8409] + last_layer_output[8410] + last_layer_output[8411] + last_layer_output[8412] + last_layer_output[8413] + last_layer_output[8414] + last_layer_output[8415] + last_layer_output[8416] + last_layer_output[8417] + last_layer_output[8418] + last_layer_output[8419] + last_layer_output[8420] + last_layer_output[8421] + last_layer_output[8422] + last_layer_output[8423] + last_layer_output[8424] + last_layer_output[8425] + last_layer_output[8426] + last_layer_output[8427] + last_layer_output[8428] + last_layer_output[8429] + last_layer_output[8430] + last_layer_output[8431] + last_layer_output[8432] + last_layer_output[8433] + last_layer_output[8434] + last_layer_output[8435] + last_layer_output[8436] + last_layer_output[8437] + last_layer_output[8438] + last_layer_output[8439] + last_layer_output[8440] + last_layer_output[8441] + last_layer_output[8442] + last_layer_output[8443] + last_layer_output[8444] + last_layer_output[8445] + last_layer_output[8446] + last_layer_output[8447] + last_layer_output[8448] + last_layer_output[8449] + last_layer_output[8450] + last_layer_output[8451] + last_layer_output[8452] + last_layer_output[8453] + last_layer_output[8454] + last_layer_output[8455] + last_layer_output[8456] + last_layer_output[8457] + last_layer_output[8458] + last_layer_output[8459] + last_layer_output[8460] + last_layer_output[8461] + last_layer_output[8462] + last_layer_output[8463] + last_layer_output[8464] + last_layer_output[8465] + last_layer_output[8466] + last_layer_output[8467] + last_layer_output[8468] + last_layer_output[8469] + last_layer_output[8470] + last_layer_output[8471] + last_layer_output[8472] + last_layer_output[8473] + last_layer_output[8474] + last_layer_output[8475] + last_layer_output[8476] + last_layer_output[8477] + last_layer_output[8478] + last_layer_output[8479] + last_layer_output[8480] + last_layer_output[8481] + last_layer_output[8482] + last_layer_output[8483] + last_layer_output[8484] + last_layer_output[8485] + last_layer_output[8486] + last_layer_output[8487] + last_layer_output[8488] + last_layer_output[8489] + last_layer_output[8490] + last_layer_output[8491] + last_layer_output[8492] + last_layer_output[8493] + last_layer_output[8494] + last_layer_output[8495] + last_layer_output[8496] + last_layer_output[8497] + last_layer_output[8498] + last_layer_output[8499] + last_layer_output[8500] + last_layer_output[8501] + last_layer_output[8502] + last_layer_output[8503] + last_layer_output[8504] + last_layer_output[8505] + last_layer_output[8506] + last_layer_output[8507] + last_layer_output[8508] + last_layer_output[8509] + last_layer_output[8510] + last_layer_output[8511] + last_layer_output[8512] + last_layer_output[8513] + last_layer_output[8514] + last_layer_output[8515] + last_layer_output[8516] + last_layer_output[8517] + last_layer_output[8518] + last_layer_output[8519] + last_layer_output[8520] + last_layer_output[8521] + last_layer_output[8522] + last_layer_output[8523] + last_layer_output[8524] + last_layer_output[8525] + last_layer_output[8526] + last_layer_output[8527] + last_layer_output[8528] + last_layer_output[8529] + last_layer_output[8530] + last_layer_output[8531] + last_layer_output[8532] + last_layer_output[8533] + last_layer_output[8534] + last_layer_output[8535] + last_layer_output[8536] + last_layer_output[8537] + last_layer_output[8538] + last_layer_output[8539] + last_layer_output[8540] + last_layer_output[8541] + last_layer_output[8542] + last_layer_output[8543] + last_layer_output[8544] + last_layer_output[8545] + last_layer_output[8546] + last_layer_output[8547] + last_layer_output[8548] + last_layer_output[8549] + last_layer_output[8550] + last_layer_output[8551] + last_layer_output[8552] + last_layer_output[8553] + last_layer_output[8554] + last_layer_output[8555] + last_layer_output[8556] + last_layer_output[8557] + last_layer_output[8558] + last_layer_output[8559] + last_layer_output[8560] + last_layer_output[8561] + last_layer_output[8562] + last_layer_output[8563] + last_layer_output[8564] + last_layer_output[8565] + last_layer_output[8566] + last_layer_output[8567] + last_layer_output[8568] + last_layer_output[8569] + last_layer_output[8570] + last_layer_output[8571] + last_layer_output[8572] + last_layer_output[8573] + last_layer_output[8574] + last_layer_output[8575] + last_layer_output[8576] + last_layer_output[8577] + last_layer_output[8578] + last_layer_output[8579] + last_layer_output[8580] + last_layer_output[8581] + last_layer_output[8582] + last_layer_output[8583] + last_layer_output[8584] + last_layer_output[8585] + last_layer_output[8586] + last_layer_output[8587] + last_layer_output[8588] + last_layer_output[8589] + last_layer_output[8590] + last_layer_output[8591] + last_layer_output[8592] + last_layer_output[8593] + last_layer_output[8594] + last_layer_output[8595] + last_layer_output[8596] + last_layer_output[8597] + last_layer_output[8598] + last_layer_output[8599] + last_layer_output[8600] + last_layer_output[8601] + last_layer_output[8602] + last_layer_output[8603] + last_layer_output[8604] + last_layer_output[8605] + last_layer_output[8606] + last_layer_output[8607] + last_layer_output[8608] + last_layer_output[8609] + last_layer_output[8610] + last_layer_output[8611] + last_layer_output[8612] + last_layer_output[8613] + last_layer_output[8614] + last_layer_output[8615] + last_layer_output[8616] + last_layer_output[8617] + last_layer_output[8618] + last_layer_output[8619] + last_layer_output[8620] + last_layer_output[8621] + last_layer_output[8622] + last_layer_output[8623] + last_layer_output[8624] + last_layer_output[8625] + last_layer_output[8626] + last_layer_output[8627] + last_layer_output[8628] + last_layer_output[8629] + last_layer_output[8630] + last_layer_output[8631] + last_layer_output[8632] + last_layer_output[8633] + last_layer_output[8634] + last_layer_output[8635] + last_layer_output[8636] + last_layer_output[8637] + last_layer_output[8638] + last_layer_output[8639] + last_layer_output[8640] + last_layer_output[8641] + last_layer_output[8642] + last_layer_output[8643] + last_layer_output[8644] + last_layer_output[8645] + last_layer_output[8646] + last_layer_output[8647] + last_layer_output[8648] + last_layer_output[8649] + last_layer_output[8650] + last_layer_output[8651] + last_layer_output[8652] + last_layer_output[8653] + last_layer_output[8654] + last_layer_output[8655] + last_layer_output[8656] + last_layer_output[8657] + last_layer_output[8658] + last_layer_output[8659] + last_layer_output[8660] + last_layer_output[8661] + last_layer_output[8662] + last_layer_output[8663] + last_layer_output[8664] + last_layer_output[8665] + last_layer_output[8666] + last_layer_output[8667] + last_layer_output[8668] + last_layer_output[8669] + last_layer_output[8670] + last_layer_output[8671] + last_layer_output[8672] + last_layer_output[8673] + last_layer_output[8674] + last_layer_output[8675] + last_layer_output[8676] + last_layer_output[8677] + last_layer_output[8678] + last_layer_output[8679] + last_layer_output[8680] + last_layer_output[8681] + last_layer_output[8682] + last_layer_output[8683] + last_layer_output[8684] + last_layer_output[8685] + last_layer_output[8686] + last_layer_output[8687] + last_layer_output[8688] + last_layer_output[8689] + last_layer_output[8690] + last_layer_output[8691] + last_layer_output[8692] + last_layer_output[8693] + last_layer_output[8694] + last_layer_output[8695] + last_layer_output[8696] + last_layer_output[8697] + last_layer_output[8698] + last_layer_output[8699] + last_layer_output[8700] + last_layer_output[8701] + last_layer_output[8702] + last_layer_output[8703] + last_layer_output[8704] + last_layer_output[8705] + last_layer_output[8706] + last_layer_output[8707] + last_layer_output[8708] + last_layer_output[8709] + last_layer_output[8710] + last_layer_output[8711] + last_layer_output[8712] + last_layer_output[8713] + last_layer_output[8714] + last_layer_output[8715] + last_layer_output[8716] + last_layer_output[8717] + last_layer_output[8718] + last_layer_output[8719] + last_layer_output[8720] + last_layer_output[8721] + last_layer_output[8722] + last_layer_output[8723] + last_layer_output[8724] + last_layer_output[8725] + last_layer_output[8726] + last_layer_output[8727] + last_layer_output[8728] + last_layer_output[8729] + last_layer_output[8730] + last_layer_output[8731] + last_layer_output[8732] + last_layer_output[8733] + last_layer_output[8734] + last_layer_output[8735] + last_layer_output[8736] + last_layer_output[8737] + last_layer_output[8738] + last_layer_output[8739] + last_layer_output[8740] + last_layer_output[8741] + last_layer_output[8742] + last_layer_output[8743] + last_layer_output[8744] + last_layer_output[8745] + last_layer_output[8746] + last_layer_output[8747] + last_layer_output[8748] + last_layer_output[8749] + last_layer_output[8750] + last_layer_output[8751] + last_layer_output[8752] + last_layer_output[8753] + last_layer_output[8754] + last_layer_output[8755] + last_layer_output[8756] + last_layer_output[8757] + last_layer_output[8758] + last_layer_output[8759] + last_layer_output[8760] + last_layer_output[8761] + last_layer_output[8762] + last_layer_output[8763] + last_layer_output[8764] + last_layer_output[8765] + last_layer_output[8766] + last_layer_output[8767] + last_layer_output[8768] + last_layer_output[8769] + last_layer_output[8770] + last_layer_output[8771] + last_layer_output[8772] + last_layer_output[8773] + last_layer_output[8774] + last_layer_output[8775] + last_layer_output[8776] + last_layer_output[8777] + last_layer_output[8778] + last_layer_output[8779] + last_layer_output[8780] + last_layer_output[8781] + last_layer_output[8782] + last_layer_output[8783] + last_layer_output[8784] + last_layer_output[8785] + last_layer_output[8786] + last_layer_output[8787] + last_layer_output[8788] + last_layer_output[8789] + last_layer_output[8790] + last_layer_output[8791] + last_layer_output[8792] + last_layer_output[8793] + last_layer_output[8794] + last_layer_output[8795] + last_layer_output[8796] + last_layer_output[8797] + last_layer_output[8798] + last_layer_output[8799] + last_layer_output[8800] + last_layer_output[8801] + last_layer_output[8802] + last_layer_output[8803] + last_layer_output[8804] + last_layer_output[8805] + last_layer_output[8806] + last_layer_output[8807] + last_layer_output[8808] + last_layer_output[8809] + last_layer_output[8810] + last_layer_output[8811] + last_layer_output[8812] + last_layer_output[8813] + last_layer_output[8814] + last_layer_output[8815] + last_layer_output[8816] + last_layer_output[8817] + last_layer_output[8818] + last_layer_output[8819] + last_layer_output[8820] + last_layer_output[8821] + last_layer_output[8822] + last_layer_output[8823] + last_layer_output[8824] + last_layer_output[8825] + last_layer_output[8826] + last_layer_output[8827] + last_layer_output[8828] + last_layer_output[8829] + last_layer_output[8830] + last_layer_output[8831] + last_layer_output[8832] + last_layer_output[8833] + last_layer_output[8834] + last_layer_output[8835] + last_layer_output[8836] + last_layer_output[8837] + last_layer_output[8838] + last_layer_output[8839] + last_layer_output[8840] + last_layer_output[8841] + last_layer_output[8842] + last_layer_output[8843] + last_layer_output[8844] + last_layer_output[8845] + last_layer_output[8846] + last_layer_output[8847] + last_layer_output[8848] + last_layer_output[8849] + last_layer_output[8850] + last_layer_output[8851] + last_layer_output[8852] + last_layer_output[8853] + last_layer_output[8854] + last_layer_output[8855] + last_layer_output[8856] + last_layer_output[8857] + last_layer_output[8858] + last_layer_output[8859] + last_layer_output[8860] + last_layer_output[8861] + last_layer_output[8862] + last_layer_output[8863] + last_layer_output[8864] + last_layer_output[8865] + last_layer_output[8866] + last_layer_output[8867] + last_layer_output[8868] + last_layer_output[8869] + last_layer_output[8870] + last_layer_output[8871] + last_layer_output[8872] + last_layer_output[8873] + last_layer_output[8874] + last_layer_output[8875] + last_layer_output[8876] + last_layer_output[8877] + last_layer_output[8878] + last_layer_output[8879] + last_layer_output[8880] + last_layer_output[8881] + last_layer_output[8882] + last_layer_output[8883] + last_layer_output[8884] + last_layer_output[8885] + last_layer_output[8886] + last_layer_output[8887] + last_layer_output[8888] + last_layer_output[8889] + last_layer_output[8890] + last_layer_output[8891] + last_layer_output[8892] + last_layer_output[8893] + last_layer_output[8894] + last_layer_output[8895] + last_layer_output[8896] + last_layer_output[8897] + last_layer_output[8898] + last_layer_output[8899] + last_layer_output[8900] + last_layer_output[8901] + last_layer_output[8902] + last_layer_output[8903] + last_layer_output[8904] + last_layer_output[8905] + last_layer_output[8906] + last_layer_output[8907] + last_layer_output[8908] + last_layer_output[8909] + last_layer_output[8910] + last_layer_output[8911] + last_layer_output[8912] + last_layer_output[8913] + last_layer_output[8914] + last_layer_output[8915] + last_layer_output[8916] + last_layer_output[8917] + last_layer_output[8918] + last_layer_output[8919] + last_layer_output[8920] + last_layer_output[8921] + last_layer_output[8922] + last_layer_output[8923] + last_layer_output[8924] + last_layer_output[8925] + last_layer_output[8926] + last_layer_output[8927] + last_layer_output[8928] + last_layer_output[8929] + last_layer_output[8930] + last_layer_output[8931] + last_layer_output[8932] + last_layer_output[8933] + last_layer_output[8934] + last_layer_output[8935] + last_layer_output[8936] + last_layer_output[8937] + last_layer_output[8938] + last_layer_output[8939] + last_layer_output[8940] + last_layer_output[8941] + last_layer_output[8942] + last_layer_output[8943] + last_layer_output[8944] + last_layer_output[8945] + last_layer_output[8946] + last_layer_output[8947] + last_layer_output[8948] + last_layer_output[8949] + last_layer_output[8950] + last_layer_output[8951] + last_layer_output[8952] + last_layer_output[8953] + last_layer_output[8954] + last_layer_output[8955] + last_layer_output[8956] + last_layer_output[8957] + last_layer_output[8958] + last_layer_output[8959] + last_layer_output[8960] + last_layer_output[8961] + last_layer_output[8962] + last_layer_output[8963] + last_layer_output[8964] + last_layer_output[8965] + last_layer_output[8966] + last_layer_output[8967] + last_layer_output[8968] + last_layer_output[8969] + last_layer_output[8970] + last_layer_output[8971] + last_layer_output[8972] + last_layer_output[8973] + last_layer_output[8974] + last_layer_output[8975] + last_layer_output[8976] + last_layer_output[8977] + last_layer_output[8978] + last_layer_output[8979] + last_layer_output[8980] + last_layer_output[8981] + last_layer_output[8982] + last_layer_output[8983] + last_layer_output[8984] + last_layer_output[8985] + last_layer_output[8986] + last_layer_output[8987] + last_layer_output[8988] + last_layer_output[8989] + last_layer_output[8990] + last_layer_output[8991] + last_layer_output[8992] + last_layer_output[8993] + last_layer_output[8994] + last_layer_output[8995] + last_layer_output[8996] + last_layer_output[8997] + last_layer_output[8998] + last_layer_output[8999] + last_layer_output[9000] + last_layer_output[9001] + last_layer_output[9002] + last_layer_output[9003] + last_layer_output[9004] + last_layer_output[9005] + last_layer_output[9006] + last_layer_output[9007] + last_layer_output[9008] + last_layer_output[9009] + last_layer_output[9010] + last_layer_output[9011] + last_layer_output[9012] + last_layer_output[9013] + last_layer_output[9014] + last_layer_output[9015] + last_layer_output[9016] + last_layer_output[9017] + last_layer_output[9018] + last_layer_output[9019] + last_layer_output[9020] + last_layer_output[9021] + last_layer_output[9022] + last_layer_output[9023] + last_layer_output[9024] + last_layer_output[9025] + last_layer_output[9026] + last_layer_output[9027] + last_layer_output[9028] + last_layer_output[9029] + last_layer_output[9030] + last_layer_output[9031] + last_layer_output[9032] + last_layer_output[9033] + last_layer_output[9034] + last_layer_output[9035] + last_layer_output[9036] + last_layer_output[9037] + last_layer_output[9038] + last_layer_output[9039] + last_layer_output[9040] + last_layer_output[9041] + last_layer_output[9042] + last_layer_output[9043] + last_layer_output[9044] + last_layer_output[9045] + last_layer_output[9046] + last_layer_output[9047] + last_layer_output[9048] + last_layer_output[9049] + last_layer_output[9050] + last_layer_output[9051] + last_layer_output[9052] + last_layer_output[9053] + last_layer_output[9054] + last_layer_output[9055] + last_layer_output[9056] + last_layer_output[9057] + last_layer_output[9058] + last_layer_output[9059] + last_layer_output[9060] + last_layer_output[9061] + last_layer_output[9062] + last_layer_output[9063] + last_layer_output[9064] + last_layer_output[9065] + last_layer_output[9066] + last_layer_output[9067] + last_layer_output[9068] + last_layer_output[9069] + last_layer_output[9070] + last_layer_output[9071] + last_layer_output[9072] + last_layer_output[9073] + last_layer_output[9074] + last_layer_output[9075] + last_layer_output[9076] + last_layer_output[9077] + last_layer_output[9078] + last_layer_output[9079] + last_layer_output[9080] + last_layer_output[9081] + last_layer_output[9082] + last_layer_output[9083] + last_layer_output[9084] + last_layer_output[9085] + last_layer_output[9086] + last_layer_output[9087] + last_layer_output[9088] + last_layer_output[9089] + last_layer_output[9090] + last_layer_output[9091] + last_layer_output[9092] + last_layer_output[9093] + last_layer_output[9094] + last_layer_output[9095] + last_layer_output[9096] + last_layer_output[9097] + last_layer_output[9098] + last_layer_output[9099] + last_layer_output[9100] + last_layer_output[9101] + last_layer_output[9102] + last_layer_output[9103] + last_layer_output[9104] + last_layer_output[9105] + last_layer_output[9106] + last_layer_output[9107] + last_layer_output[9108] + last_layer_output[9109] + last_layer_output[9110] + last_layer_output[9111] + last_layer_output[9112] + last_layer_output[9113] + last_layer_output[9114] + last_layer_output[9115] + last_layer_output[9116] + last_layer_output[9117] + last_layer_output[9118] + last_layer_output[9119] + last_layer_output[9120] + last_layer_output[9121] + last_layer_output[9122] + last_layer_output[9123] + last_layer_output[9124] + last_layer_output[9125] + last_layer_output[9126] + last_layer_output[9127] + last_layer_output[9128] + last_layer_output[9129] + last_layer_output[9130] + last_layer_output[9131] + last_layer_output[9132] + last_layer_output[9133] + last_layer_output[9134] + last_layer_output[9135] + last_layer_output[9136] + last_layer_output[9137] + last_layer_output[9138] + last_layer_output[9139] + last_layer_output[9140] + last_layer_output[9141] + last_layer_output[9142] + last_layer_output[9143] + last_layer_output[9144] + last_layer_output[9145] + last_layer_output[9146] + last_layer_output[9147] + last_layer_output[9148] + last_layer_output[9149] + last_layer_output[9150] + last_layer_output[9151] + last_layer_output[9152] + last_layer_output[9153] + last_layer_output[9154] + last_layer_output[9155] + last_layer_output[9156] + last_layer_output[9157] + last_layer_output[9158] + last_layer_output[9159] + last_layer_output[9160] + last_layer_output[9161] + last_layer_output[9162] + last_layer_output[9163] + last_layer_output[9164] + last_layer_output[9165] + last_layer_output[9166] + last_layer_output[9167] + last_layer_output[9168] + last_layer_output[9169] + last_layer_output[9170] + last_layer_output[9171] + last_layer_output[9172] + last_layer_output[9173] + last_layer_output[9174] + last_layer_output[9175] + last_layer_output[9176] + last_layer_output[9177] + last_layer_output[9178] + last_layer_output[9179] + last_layer_output[9180] + last_layer_output[9181] + last_layer_output[9182] + last_layer_output[9183] + last_layer_output[9184] + last_layer_output[9185] + last_layer_output[9186] + last_layer_output[9187] + last_layer_output[9188] + last_layer_output[9189] + last_layer_output[9190] + last_layer_output[9191] + last_layer_output[9192] + last_layer_output[9193] + last_layer_output[9194] + last_layer_output[9195] + last_layer_output[9196] + last_layer_output[9197] + last_layer_output[9198] + last_layer_output[9199] + last_layer_output[9200] + last_layer_output[9201] + last_layer_output[9202] + last_layer_output[9203] + last_layer_output[9204] + last_layer_output[9205] + last_layer_output[9206] + last_layer_output[9207] + last_layer_output[9208] + last_layer_output[9209] + last_layer_output[9210] + last_layer_output[9211] + last_layer_output[9212] + last_layer_output[9213] + last_layer_output[9214] + last_layer_output[9215] + last_layer_output[9216] + last_layer_output[9217] + last_layer_output[9218] + last_layer_output[9219] + last_layer_output[9220] + last_layer_output[9221] + last_layer_output[9222] + last_layer_output[9223] + last_layer_output[9224] + last_layer_output[9225] + last_layer_output[9226] + last_layer_output[9227] + last_layer_output[9228] + last_layer_output[9229] + last_layer_output[9230] + last_layer_output[9231] + last_layer_output[9232] + last_layer_output[9233] + last_layer_output[9234] + last_layer_output[9235] + last_layer_output[9236] + last_layer_output[9237] + last_layer_output[9238] + last_layer_output[9239] + last_layer_output[9240] + last_layer_output[9241] + last_layer_output[9242] + last_layer_output[9243] + last_layer_output[9244] + last_layer_output[9245] + last_layer_output[9246] + last_layer_output[9247] + last_layer_output[9248] + last_layer_output[9249] + last_layer_output[9250] + last_layer_output[9251] + last_layer_output[9252] + last_layer_output[9253] + last_layer_output[9254] + last_layer_output[9255] + last_layer_output[9256] + last_layer_output[9257] + last_layer_output[9258] + last_layer_output[9259] + last_layer_output[9260] + last_layer_output[9261] + last_layer_output[9262] + last_layer_output[9263] + last_layer_output[9264] + last_layer_output[9265] + last_layer_output[9266] + last_layer_output[9267] + last_layer_output[9268] + last_layer_output[9269] + last_layer_output[9270] + last_layer_output[9271] + last_layer_output[9272] + last_layer_output[9273] + last_layer_output[9274] + last_layer_output[9275] + last_layer_output[9276] + last_layer_output[9277] + last_layer_output[9278] + last_layer_output[9279] + last_layer_output[9280] + last_layer_output[9281] + last_layer_output[9282] + last_layer_output[9283] + last_layer_output[9284] + last_layer_output[9285] + last_layer_output[9286] + last_layer_output[9287] + last_layer_output[9288] + last_layer_output[9289] + last_layer_output[9290] + last_layer_output[9291] + last_layer_output[9292] + last_layer_output[9293] + last_layer_output[9294] + last_layer_output[9295] + last_layer_output[9296] + last_layer_output[9297] + last_layer_output[9298] + last_layer_output[9299] + last_layer_output[9300] + last_layer_output[9301] + last_layer_output[9302] + last_layer_output[9303] + last_layer_output[9304] + last_layer_output[9305] + last_layer_output[9306] + last_layer_output[9307] + last_layer_output[9308] + last_layer_output[9309] + last_layer_output[9310] + last_layer_output[9311] + last_layer_output[9312] + last_layer_output[9313] + last_layer_output[9314] + last_layer_output[9315] + last_layer_output[9316] + last_layer_output[9317] + last_layer_output[9318] + last_layer_output[9319] + last_layer_output[9320] + last_layer_output[9321] + last_layer_output[9322] + last_layer_output[9323] + last_layer_output[9324] + last_layer_output[9325] + last_layer_output[9326] + last_layer_output[9327] + last_layer_output[9328] + last_layer_output[9329] + last_layer_output[9330] + last_layer_output[9331] + last_layer_output[9332] + last_layer_output[9333] + last_layer_output[9334] + last_layer_output[9335] + last_layer_output[9336] + last_layer_output[9337] + last_layer_output[9338] + last_layer_output[9339] + last_layer_output[9340] + last_layer_output[9341] + last_layer_output[9342] + last_layer_output[9343] + last_layer_output[9344] + last_layer_output[9345] + last_layer_output[9346] + last_layer_output[9347] + last_layer_output[9348] + last_layer_output[9349] + last_layer_output[9350] + last_layer_output[9351] + last_layer_output[9352] + last_layer_output[9353] + last_layer_output[9354] + last_layer_output[9355] + last_layer_output[9356] + last_layer_output[9357] + last_layer_output[9358] + last_layer_output[9359] + last_layer_output[9360] + last_layer_output[9361] + last_layer_output[9362] + last_layer_output[9363] + last_layer_output[9364] + last_layer_output[9365] + last_layer_output[9366] + last_layer_output[9367] + last_layer_output[9368] + last_layer_output[9369] + last_layer_output[9370] + last_layer_output[9371] + last_layer_output[9372] + last_layer_output[9373] + last_layer_output[9374] + last_layer_output[9375] + last_layer_output[9376] + last_layer_output[9377] + last_layer_output[9378] + last_layer_output[9379] + last_layer_output[9380] + last_layer_output[9381] + last_layer_output[9382] + last_layer_output[9383] + last_layer_output[9384] + last_layer_output[9385] + last_layer_output[9386] + last_layer_output[9387] + last_layer_output[9388] + last_layer_output[9389] + last_layer_output[9390] + last_layer_output[9391] + last_layer_output[9392] + last_layer_output[9393] + last_layer_output[9394] + last_layer_output[9395] + last_layer_output[9396] + last_layer_output[9397] + last_layer_output[9398] + last_layer_output[9399] + last_layer_output[9400] + last_layer_output[9401] + last_layer_output[9402] + last_layer_output[9403] + last_layer_output[9404] + last_layer_output[9405] + last_layer_output[9406] + last_layer_output[9407] + last_layer_output[9408] + last_layer_output[9409] + last_layer_output[9410] + last_layer_output[9411] + last_layer_output[9412] + last_layer_output[9413] + last_layer_output[9414] + last_layer_output[9415] + last_layer_output[9416] + last_layer_output[9417] + last_layer_output[9418] + last_layer_output[9419] + last_layer_output[9420] + last_layer_output[9421] + last_layer_output[9422] + last_layer_output[9423] + last_layer_output[9424] + last_layer_output[9425] + last_layer_output[9426] + last_layer_output[9427] + last_layer_output[9428] + last_layer_output[9429] + last_layer_output[9430] + last_layer_output[9431] + last_layer_output[9432] + last_layer_output[9433] + last_layer_output[9434] + last_layer_output[9435] + last_layer_output[9436] + last_layer_output[9437] + last_layer_output[9438] + last_layer_output[9439] + last_layer_output[9440] + last_layer_output[9441] + last_layer_output[9442] + last_layer_output[9443] + last_layer_output[9444] + last_layer_output[9445] + last_layer_output[9446] + last_layer_output[9447] + last_layer_output[9448] + last_layer_output[9449] + last_layer_output[9450] + last_layer_output[9451] + last_layer_output[9452] + last_layer_output[9453] + last_layer_output[9454] + last_layer_output[9455] + last_layer_output[9456] + last_layer_output[9457] + last_layer_output[9458] + last_layer_output[9459] + last_layer_output[9460] + last_layer_output[9461] + last_layer_output[9462] + last_layer_output[9463] + last_layer_output[9464] + last_layer_output[9465] + last_layer_output[9466] + last_layer_output[9467] + last_layer_output[9468] + last_layer_output[9469] + last_layer_output[9470] + last_layer_output[9471] + last_layer_output[9472] + last_layer_output[9473] + last_layer_output[9474] + last_layer_output[9475] + last_layer_output[9476] + last_layer_output[9477] + last_layer_output[9478] + last_layer_output[9479] + last_layer_output[9480] + last_layer_output[9481] + last_layer_output[9482] + last_layer_output[9483] + last_layer_output[9484] + last_layer_output[9485] + last_layer_output[9486] + last_layer_output[9487] + last_layer_output[9488] + last_layer_output[9489] + last_layer_output[9490] + last_layer_output[9491] + last_layer_output[9492] + last_layer_output[9493] + last_layer_output[9494] + last_layer_output[9495] + last_layer_output[9496] + last_layer_output[9497] + last_layer_output[9498] + last_layer_output[9499] + last_layer_output[9500] + last_layer_output[9501] + last_layer_output[9502] + last_layer_output[9503] + last_layer_output[9504] + last_layer_output[9505] + last_layer_output[9506] + last_layer_output[9507] + last_layer_output[9508] + last_layer_output[9509] + last_layer_output[9510] + last_layer_output[9511] + last_layer_output[9512] + last_layer_output[9513] + last_layer_output[9514] + last_layer_output[9515] + last_layer_output[9516] + last_layer_output[9517] + last_layer_output[9518] + last_layer_output[9519] + last_layer_output[9520] + last_layer_output[9521] + last_layer_output[9522] + last_layer_output[9523] + last_layer_output[9524] + last_layer_output[9525] + last_layer_output[9526] + last_layer_output[9527] + last_layer_output[9528] + last_layer_output[9529] + last_layer_output[9530] + last_layer_output[9531] + last_layer_output[9532] + last_layer_output[9533] + last_layer_output[9534] + last_layer_output[9535] + last_layer_output[9536] + last_layer_output[9537] + last_layer_output[9538] + last_layer_output[9539] + last_layer_output[9540] + last_layer_output[9541] + last_layer_output[9542] + last_layer_output[9543] + last_layer_output[9544] + last_layer_output[9545] + last_layer_output[9546] + last_layer_output[9547] + last_layer_output[9548] + last_layer_output[9549] + last_layer_output[9550] + last_layer_output[9551] + last_layer_output[9552] + last_layer_output[9553] + last_layer_output[9554] + last_layer_output[9555] + last_layer_output[9556] + last_layer_output[9557] + last_layer_output[9558] + last_layer_output[9559] + last_layer_output[9560] + last_layer_output[9561] + last_layer_output[9562] + last_layer_output[9563] + last_layer_output[9564] + last_layer_output[9565] + last_layer_output[9566] + last_layer_output[9567] + last_layer_output[9568] + last_layer_output[9569] + last_layer_output[9570] + last_layer_output[9571] + last_layer_output[9572] + last_layer_output[9573] + last_layer_output[9574] + last_layer_output[9575] + last_layer_output[9576] + last_layer_output[9577] + last_layer_output[9578] + last_layer_output[9579] + last_layer_output[9580] + last_layer_output[9581] + last_layer_output[9582] + last_layer_output[9583] + last_layer_output[9584] + last_layer_output[9585] + last_layer_output[9586] + last_layer_output[9587] + last_layer_output[9588] + last_layer_output[9589] + last_layer_output[9590] + last_layer_output[9591] + last_layer_output[9592] + last_layer_output[9593] + last_layer_output[9594] + last_layer_output[9595] + last_layer_output[9596] + last_layer_output[9597] + last_layer_output[9598] + last_layer_output[9599];
      result[8] <= last_layer_output[9600] + last_layer_output[9601] + last_layer_output[9602] + last_layer_output[9603] + last_layer_output[9604] + last_layer_output[9605] + last_layer_output[9606] + last_layer_output[9607] + last_layer_output[9608] + last_layer_output[9609] + last_layer_output[9610] + last_layer_output[9611] + last_layer_output[9612] + last_layer_output[9613] + last_layer_output[9614] + last_layer_output[9615] + last_layer_output[9616] + last_layer_output[9617] + last_layer_output[9618] + last_layer_output[9619] + last_layer_output[9620] + last_layer_output[9621] + last_layer_output[9622] + last_layer_output[9623] + last_layer_output[9624] + last_layer_output[9625] + last_layer_output[9626] + last_layer_output[9627] + last_layer_output[9628] + last_layer_output[9629] + last_layer_output[9630] + last_layer_output[9631] + last_layer_output[9632] + last_layer_output[9633] + last_layer_output[9634] + last_layer_output[9635] + last_layer_output[9636] + last_layer_output[9637] + last_layer_output[9638] + last_layer_output[9639] + last_layer_output[9640] + last_layer_output[9641] + last_layer_output[9642] + last_layer_output[9643] + last_layer_output[9644] + last_layer_output[9645] + last_layer_output[9646] + last_layer_output[9647] + last_layer_output[9648] + last_layer_output[9649] + last_layer_output[9650] + last_layer_output[9651] + last_layer_output[9652] + last_layer_output[9653] + last_layer_output[9654] + last_layer_output[9655] + last_layer_output[9656] + last_layer_output[9657] + last_layer_output[9658] + last_layer_output[9659] + last_layer_output[9660] + last_layer_output[9661] + last_layer_output[9662] + last_layer_output[9663] + last_layer_output[9664] + last_layer_output[9665] + last_layer_output[9666] + last_layer_output[9667] + last_layer_output[9668] + last_layer_output[9669] + last_layer_output[9670] + last_layer_output[9671] + last_layer_output[9672] + last_layer_output[9673] + last_layer_output[9674] + last_layer_output[9675] + last_layer_output[9676] + last_layer_output[9677] + last_layer_output[9678] + last_layer_output[9679] + last_layer_output[9680] + last_layer_output[9681] + last_layer_output[9682] + last_layer_output[9683] + last_layer_output[9684] + last_layer_output[9685] + last_layer_output[9686] + last_layer_output[9687] + last_layer_output[9688] + last_layer_output[9689] + last_layer_output[9690] + last_layer_output[9691] + last_layer_output[9692] + last_layer_output[9693] + last_layer_output[9694] + last_layer_output[9695] + last_layer_output[9696] + last_layer_output[9697] + last_layer_output[9698] + last_layer_output[9699] + last_layer_output[9700] + last_layer_output[9701] + last_layer_output[9702] + last_layer_output[9703] + last_layer_output[9704] + last_layer_output[9705] + last_layer_output[9706] + last_layer_output[9707] + last_layer_output[9708] + last_layer_output[9709] + last_layer_output[9710] + last_layer_output[9711] + last_layer_output[9712] + last_layer_output[9713] + last_layer_output[9714] + last_layer_output[9715] + last_layer_output[9716] + last_layer_output[9717] + last_layer_output[9718] + last_layer_output[9719] + last_layer_output[9720] + last_layer_output[9721] + last_layer_output[9722] + last_layer_output[9723] + last_layer_output[9724] + last_layer_output[9725] + last_layer_output[9726] + last_layer_output[9727] + last_layer_output[9728] + last_layer_output[9729] + last_layer_output[9730] + last_layer_output[9731] + last_layer_output[9732] + last_layer_output[9733] + last_layer_output[9734] + last_layer_output[9735] + last_layer_output[9736] + last_layer_output[9737] + last_layer_output[9738] + last_layer_output[9739] + last_layer_output[9740] + last_layer_output[9741] + last_layer_output[9742] + last_layer_output[9743] + last_layer_output[9744] + last_layer_output[9745] + last_layer_output[9746] + last_layer_output[9747] + last_layer_output[9748] + last_layer_output[9749] + last_layer_output[9750] + last_layer_output[9751] + last_layer_output[9752] + last_layer_output[9753] + last_layer_output[9754] + last_layer_output[9755] + last_layer_output[9756] + last_layer_output[9757] + last_layer_output[9758] + last_layer_output[9759] + last_layer_output[9760] + last_layer_output[9761] + last_layer_output[9762] + last_layer_output[9763] + last_layer_output[9764] + last_layer_output[9765] + last_layer_output[9766] + last_layer_output[9767] + last_layer_output[9768] + last_layer_output[9769] + last_layer_output[9770] + last_layer_output[9771] + last_layer_output[9772] + last_layer_output[9773] + last_layer_output[9774] + last_layer_output[9775] + last_layer_output[9776] + last_layer_output[9777] + last_layer_output[9778] + last_layer_output[9779] + last_layer_output[9780] + last_layer_output[9781] + last_layer_output[9782] + last_layer_output[9783] + last_layer_output[9784] + last_layer_output[9785] + last_layer_output[9786] + last_layer_output[9787] + last_layer_output[9788] + last_layer_output[9789] + last_layer_output[9790] + last_layer_output[9791] + last_layer_output[9792] + last_layer_output[9793] + last_layer_output[9794] + last_layer_output[9795] + last_layer_output[9796] + last_layer_output[9797] + last_layer_output[9798] + last_layer_output[9799] + last_layer_output[9800] + last_layer_output[9801] + last_layer_output[9802] + last_layer_output[9803] + last_layer_output[9804] + last_layer_output[9805] + last_layer_output[9806] + last_layer_output[9807] + last_layer_output[9808] + last_layer_output[9809] + last_layer_output[9810] + last_layer_output[9811] + last_layer_output[9812] + last_layer_output[9813] + last_layer_output[9814] + last_layer_output[9815] + last_layer_output[9816] + last_layer_output[9817] + last_layer_output[9818] + last_layer_output[9819] + last_layer_output[9820] + last_layer_output[9821] + last_layer_output[9822] + last_layer_output[9823] + last_layer_output[9824] + last_layer_output[9825] + last_layer_output[9826] + last_layer_output[9827] + last_layer_output[9828] + last_layer_output[9829] + last_layer_output[9830] + last_layer_output[9831] + last_layer_output[9832] + last_layer_output[9833] + last_layer_output[9834] + last_layer_output[9835] + last_layer_output[9836] + last_layer_output[9837] + last_layer_output[9838] + last_layer_output[9839] + last_layer_output[9840] + last_layer_output[9841] + last_layer_output[9842] + last_layer_output[9843] + last_layer_output[9844] + last_layer_output[9845] + last_layer_output[9846] + last_layer_output[9847] + last_layer_output[9848] + last_layer_output[9849] + last_layer_output[9850] + last_layer_output[9851] + last_layer_output[9852] + last_layer_output[9853] + last_layer_output[9854] + last_layer_output[9855] + last_layer_output[9856] + last_layer_output[9857] + last_layer_output[9858] + last_layer_output[9859] + last_layer_output[9860] + last_layer_output[9861] + last_layer_output[9862] + last_layer_output[9863] + last_layer_output[9864] + last_layer_output[9865] + last_layer_output[9866] + last_layer_output[9867] + last_layer_output[9868] + last_layer_output[9869] + last_layer_output[9870] + last_layer_output[9871] + last_layer_output[9872] + last_layer_output[9873] + last_layer_output[9874] + last_layer_output[9875] + last_layer_output[9876] + last_layer_output[9877] + last_layer_output[9878] + last_layer_output[9879] + last_layer_output[9880] + last_layer_output[9881] + last_layer_output[9882] + last_layer_output[9883] + last_layer_output[9884] + last_layer_output[9885] + last_layer_output[9886] + last_layer_output[9887] + last_layer_output[9888] + last_layer_output[9889] + last_layer_output[9890] + last_layer_output[9891] + last_layer_output[9892] + last_layer_output[9893] + last_layer_output[9894] + last_layer_output[9895] + last_layer_output[9896] + last_layer_output[9897] + last_layer_output[9898] + last_layer_output[9899] + last_layer_output[9900] + last_layer_output[9901] + last_layer_output[9902] + last_layer_output[9903] + last_layer_output[9904] + last_layer_output[9905] + last_layer_output[9906] + last_layer_output[9907] + last_layer_output[9908] + last_layer_output[9909] + last_layer_output[9910] + last_layer_output[9911] + last_layer_output[9912] + last_layer_output[9913] + last_layer_output[9914] + last_layer_output[9915] + last_layer_output[9916] + last_layer_output[9917] + last_layer_output[9918] + last_layer_output[9919] + last_layer_output[9920] + last_layer_output[9921] + last_layer_output[9922] + last_layer_output[9923] + last_layer_output[9924] + last_layer_output[9925] + last_layer_output[9926] + last_layer_output[9927] + last_layer_output[9928] + last_layer_output[9929] + last_layer_output[9930] + last_layer_output[9931] + last_layer_output[9932] + last_layer_output[9933] + last_layer_output[9934] + last_layer_output[9935] + last_layer_output[9936] + last_layer_output[9937] + last_layer_output[9938] + last_layer_output[9939] + last_layer_output[9940] + last_layer_output[9941] + last_layer_output[9942] + last_layer_output[9943] + last_layer_output[9944] + last_layer_output[9945] + last_layer_output[9946] + last_layer_output[9947] + last_layer_output[9948] + last_layer_output[9949] + last_layer_output[9950] + last_layer_output[9951] + last_layer_output[9952] + last_layer_output[9953] + last_layer_output[9954] + last_layer_output[9955] + last_layer_output[9956] + last_layer_output[9957] + last_layer_output[9958] + last_layer_output[9959] + last_layer_output[9960] + last_layer_output[9961] + last_layer_output[9962] + last_layer_output[9963] + last_layer_output[9964] + last_layer_output[9965] + last_layer_output[9966] + last_layer_output[9967] + last_layer_output[9968] + last_layer_output[9969] + last_layer_output[9970] + last_layer_output[9971] + last_layer_output[9972] + last_layer_output[9973] + last_layer_output[9974] + last_layer_output[9975] + last_layer_output[9976] + last_layer_output[9977] + last_layer_output[9978] + last_layer_output[9979] + last_layer_output[9980] + last_layer_output[9981] + last_layer_output[9982] + last_layer_output[9983] + last_layer_output[9984] + last_layer_output[9985] + last_layer_output[9986] + last_layer_output[9987] + last_layer_output[9988] + last_layer_output[9989] + last_layer_output[9990] + last_layer_output[9991] + last_layer_output[9992] + last_layer_output[9993] + last_layer_output[9994] + last_layer_output[9995] + last_layer_output[9996] + last_layer_output[9997] + last_layer_output[9998] + last_layer_output[9999] + last_layer_output[10000] + last_layer_output[10001] + last_layer_output[10002] + last_layer_output[10003] + last_layer_output[10004] + last_layer_output[10005] + last_layer_output[10006] + last_layer_output[10007] + last_layer_output[10008] + last_layer_output[10009] + last_layer_output[10010] + last_layer_output[10011] + last_layer_output[10012] + last_layer_output[10013] + last_layer_output[10014] + last_layer_output[10015] + last_layer_output[10016] + last_layer_output[10017] + last_layer_output[10018] + last_layer_output[10019] + last_layer_output[10020] + last_layer_output[10021] + last_layer_output[10022] + last_layer_output[10023] + last_layer_output[10024] + last_layer_output[10025] + last_layer_output[10026] + last_layer_output[10027] + last_layer_output[10028] + last_layer_output[10029] + last_layer_output[10030] + last_layer_output[10031] + last_layer_output[10032] + last_layer_output[10033] + last_layer_output[10034] + last_layer_output[10035] + last_layer_output[10036] + last_layer_output[10037] + last_layer_output[10038] + last_layer_output[10039] + last_layer_output[10040] + last_layer_output[10041] + last_layer_output[10042] + last_layer_output[10043] + last_layer_output[10044] + last_layer_output[10045] + last_layer_output[10046] + last_layer_output[10047] + last_layer_output[10048] + last_layer_output[10049] + last_layer_output[10050] + last_layer_output[10051] + last_layer_output[10052] + last_layer_output[10053] + last_layer_output[10054] + last_layer_output[10055] + last_layer_output[10056] + last_layer_output[10057] + last_layer_output[10058] + last_layer_output[10059] + last_layer_output[10060] + last_layer_output[10061] + last_layer_output[10062] + last_layer_output[10063] + last_layer_output[10064] + last_layer_output[10065] + last_layer_output[10066] + last_layer_output[10067] + last_layer_output[10068] + last_layer_output[10069] + last_layer_output[10070] + last_layer_output[10071] + last_layer_output[10072] + last_layer_output[10073] + last_layer_output[10074] + last_layer_output[10075] + last_layer_output[10076] + last_layer_output[10077] + last_layer_output[10078] + last_layer_output[10079] + last_layer_output[10080] + last_layer_output[10081] + last_layer_output[10082] + last_layer_output[10083] + last_layer_output[10084] + last_layer_output[10085] + last_layer_output[10086] + last_layer_output[10087] + last_layer_output[10088] + last_layer_output[10089] + last_layer_output[10090] + last_layer_output[10091] + last_layer_output[10092] + last_layer_output[10093] + last_layer_output[10094] + last_layer_output[10095] + last_layer_output[10096] + last_layer_output[10097] + last_layer_output[10098] + last_layer_output[10099] + last_layer_output[10100] + last_layer_output[10101] + last_layer_output[10102] + last_layer_output[10103] + last_layer_output[10104] + last_layer_output[10105] + last_layer_output[10106] + last_layer_output[10107] + last_layer_output[10108] + last_layer_output[10109] + last_layer_output[10110] + last_layer_output[10111] + last_layer_output[10112] + last_layer_output[10113] + last_layer_output[10114] + last_layer_output[10115] + last_layer_output[10116] + last_layer_output[10117] + last_layer_output[10118] + last_layer_output[10119] + last_layer_output[10120] + last_layer_output[10121] + last_layer_output[10122] + last_layer_output[10123] + last_layer_output[10124] + last_layer_output[10125] + last_layer_output[10126] + last_layer_output[10127] + last_layer_output[10128] + last_layer_output[10129] + last_layer_output[10130] + last_layer_output[10131] + last_layer_output[10132] + last_layer_output[10133] + last_layer_output[10134] + last_layer_output[10135] + last_layer_output[10136] + last_layer_output[10137] + last_layer_output[10138] + last_layer_output[10139] + last_layer_output[10140] + last_layer_output[10141] + last_layer_output[10142] + last_layer_output[10143] + last_layer_output[10144] + last_layer_output[10145] + last_layer_output[10146] + last_layer_output[10147] + last_layer_output[10148] + last_layer_output[10149] + last_layer_output[10150] + last_layer_output[10151] + last_layer_output[10152] + last_layer_output[10153] + last_layer_output[10154] + last_layer_output[10155] + last_layer_output[10156] + last_layer_output[10157] + last_layer_output[10158] + last_layer_output[10159] + last_layer_output[10160] + last_layer_output[10161] + last_layer_output[10162] + last_layer_output[10163] + last_layer_output[10164] + last_layer_output[10165] + last_layer_output[10166] + last_layer_output[10167] + last_layer_output[10168] + last_layer_output[10169] + last_layer_output[10170] + last_layer_output[10171] + last_layer_output[10172] + last_layer_output[10173] + last_layer_output[10174] + last_layer_output[10175] + last_layer_output[10176] + last_layer_output[10177] + last_layer_output[10178] + last_layer_output[10179] + last_layer_output[10180] + last_layer_output[10181] + last_layer_output[10182] + last_layer_output[10183] + last_layer_output[10184] + last_layer_output[10185] + last_layer_output[10186] + last_layer_output[10187] + last_layer_output[10188] + last_layer_output[10189] + last_layer_output[10190] + last_layer_output[10191] + last_layer_output[10192] + last_layer_output[10193] + last_layer_output[10194] + last_layer_output[10195] + last_layer_output[10196] + last_layer_output[10197] + last_layer_output[10198] + last_layer_output[10199] + last_layer_output[10200] + last_layer_output[10201] + last_layer_output[10202] + last_layer_output[10203] + last_layer_output[10204] + last_layer_output[10205] + last_layer_output[10206] + last_layer_output[10207] + last_layer_output[10208] + last_layer_output[10209] + last_layer_output[10210] + last_layer_output[10211] + last_layer_output[10212] + last_layer_output[10213] + last_layer_output[10214] + last_layer_output[10215] + last_layer_output[10216] + last_layer_output[10217] + last_layer_output[10218] + last_layer_output[10219] + last_layer_output[10220] + last_layer_output[10221] + last_layer_output[10222] + last_layer_output[10223] + last_layer_output[10224] + last_layer_output[10225] + last_layer_output[10226] + last_layer_output[10227] + last_layer_output[10228] + last_layer_output[10229] + last_layer_output[10230] + last_layer_output[10231] + last_layer_output[10232] + last_layer_output[10233] + last_layer_output[10234] + last_layer_output[10235] + last_layer_output[10236] + last_layer_output[10237] + last_layer_output[10238] + last_layer_output[10239] + last_layer_output[10240] + last_layer_output[10241] + last_layer_output[10242] + last_layer_output[10243] + last_layer_output[10244] + last_layer_output[10245] + last_layer_output[10246] + last_layer_output[10247] + last_layer_output[10248] + last_layer_output[10249] + last_layer_output[10250] + last_layer_output[10251] + last_layer_output[10252] + last_layer_output[10253] + last_layer_output[10254] + last_layer_output[10255] + last_layer_output[10256] + last_layer_output[10257] + last_layer_output[10258] + last_layer_output[10259] + last_layer_output[10260] + last_layer_output[10261] + last_layer_output[10262] + last_layer_output[10263] + last_layer_output[10264] + last_layer_output[10265] + last_layer_output[10266] + last_layer_output[10267] + last_layer_output[10268] + last_layer_output[10269] + last_layer_output[10270] + last_layer_output[10271] + last_layer_output[10272] + last_layer_output[10273] + last_layer_output[10274] + last_layer_output[10275] + last_layer_output[10276] + last_layer_output[10277] + last_layer_output[10278] + last_layer_output[10279] + last_layer_output[10280] + last_layer_output[10281] + last_layer_output[10282] + last_layer_output[10283] + last_layer_output[10284] + last_layer_output[10285] + last_layer_output[10286] + last_layer_output[10287] + last_layer_output[10288] + last_layer_output[10289] + last_layer_output[10290] + last_layer_output[10291] + last_layer_output[10292] + last_layer_output[10293] + last_layer_output[10294] + last_layer_output[10295] + last_layer_output[10296] + last_layer_output[10297] + last_layer_output[10298] + last_layer_output[10299] + last_layer_output[10300] + last_layer_output[10301] + last_layer_output[10302] + last_layer_output[10303] + last_layer_output[10304] + last_layer_output[10305] + last_layer_output[10306] + last_layer_output[10307] + last_layer_output[10308] + last_layer_output[10309] + last_layer_output[10310] + last_layer_output[10311] + last_layer_output[10312] + last_layer_output[10313] + last_layer_output[10314] + last_layer_output[10315] + last_layer_output[10316] + last_layer_output[10317] + last_layer_output[10318] + last_layer_output[10319] + last_layer_output[10320] + last_layer_output[10321] + last_layer_output[10322] + last_layer_output[10323] + last_layer_output[10324] + last_layer_output[10325] + last_layer_output[10326] + last_layer_output[10327] + last_layer_output[10328] + last_layer_output[10329] + last_layer_output[10330] + last_layer_output[10331] + last_layer_output[10332] + last_layer_output[10333] + last_layer_output[10334] + last_layer_output[10335] + last_layer_output[10336] + last_layer_output[10337] + last_layer_output[10338] + last_layer_output[10339] + last_layer_output[10340] + last_layer_output[10341] + last_layer_output[10342] + last_layer_output[10343] + last_layer_output[10344] + last_layer_output[10345] + last_layer_output[10346] + last_layer_output[10347] + last_layer_output[10348] + last_layer_output[10349] + last_layer_output[10350] + last_layer_output[10351] + last_layer_output[10352] + last_layer_output[10353] + last_layer_output[10354] + last_layer_output[10355] + last_layer_output[10356] + last_layer_output[10357] + last_layer_output[10358] + last_layer_output[10359] + last_layer_output[10360] + last_layer_output[10361] + last_layer_output[10362] + last_layer_output[10363] + last_layer_output[10364] + last_layer_output[10365] + last_layer_output[10366] + last_layer_output[10367] + last_layer_output[10368] + last_layer_output[10369] + last_layer_output[10370] + last_layer_output[10371] + last_layer_output[10372] + last_layer_output[10373] + last_layer_output[10374] + last_layer_output[10375] + last_layer_output[10376] + last_layer_output[10377] + last_layer_output[10378] + last_layer_output[10379] + last_layer_output[10380] + last_layer_output[10381] + last_layer_output[10382] + last_layer_output[10383] + last_layer_output[10384] + last_layer_output[10385] + last_layer_output[10386] + last_layer_output[10387] + last_layer_output[10388] + last_layer_output[10389] + last_layer_output[10390] + last_layer_output[10391] + last_layer_output[10392] + last_layer_output[10393] + last_layer_output[10394] + last_layer_output[10395] + last_layer_output[10396] + last_layer_output[10397] + last_layer_output[10398] + last_layer_output[10399] + last_layer_output[10400] + last_layer_output[10401] + last_layer_output[10402] + last_layer_output[10403] + last_layer_output[10404] + last_layer_output[10405] + last_layer_output[10406] + last_layer_output[10407] + last_layer_output[10408] + last_layer_output[10409] + last_layer_output[10410] + last_layer_output[10411] + last_layer_output[10412] + last_layer_output[10413] + last_layer_output[10414] + last_layer_output[10415] + last_layer_output[10416] + last_layer_output[10417] + last_layer_output[10418] + last_layer_output[10419] + last_layer_output[10420] + last_layer_output[10421] + last_layer_output[10422] + last_layer_output[10423] + last_layer_output[10424] + last_layer_output[10425] + last_layer_output[10426] + last_layer_output[10427] + last_layer_output[10428] + last_layer_output[10429] + last_layer_output[10430] + last_layer_output[10431] + last_layer_output[10432] + last_layer_output[10433] + last_layer_output[10434] + last_layer_output[10435] + last_layer_output[10436] + last_layer_output[10437] + last_layer_output[10438] + last_layer_output[10439] + last_layer_output[10440] + last_layer_output[10441] + last_layer_output[10442] + last_layer_output[10443] + last_layer_output[10444] + last_layer_output[10445] + last_layer_output[10446] + last_layer_output[10447] + last_layer_output[10448] + last_layer_output[10449] + last_layer_output[10450] + last_layer_output[10451] + last_layer_output[10452] + last_layer_output[10453] + last_layer_output[10454] + last_layer_output[10455] + last_layer_output[10456] + last_layer_output[10457] + last_layer_output[10458] + last_layer_output[10459] + last_layer_output[10460] + last_layer_output[10461] + last_layer_output[10462] + last_layer_output[10463] + last_layer_output[10464] + last_layer_output[10465] + last_layer_output[10466] + last_layer_output[10467] + last_layer_output[10468] + last_layer_output[10469] + last_layer_output[10470] + last_layer_output[10471] + last_layer_output[10472] + last_layer_output[10473] + last_layer_output[10474] + last_layer_output[10475] + last_layer_output[10476] + last_layer_output[10477] + last_layer_output[10478] + last_layer_output[10479] + last_layer_output[10480] + last_layer_output[10481] + last_layer_output[10482] + last_layer_output[10483] + last_layer_output[10484] + last_layer_output[10485] + last_layer_output[10486] + last_layer_output[10487] + last_layer_output[10488] + last_layer_output[10489] + last_layer_output[10490] + last_layer_output[10491] + last_layer_output[10492] + last_layer_output[10493] + last_layer_output[10494] + last_layer_output[10495] + last_layer_output[10496] + last_layer_output[10497] + last_layer_output[10498] + last_layer_output[10499] + last_layer_output[10500] + last_layer_output[10501] + last_layer_output[10502] + last_layer_output[10503] + last_layer_output[10504] + last_layer_output[10505] + last_layer_output[10506] + last_layer_output[10507] + last_layer_output[10508] + last_layer_output[10509] + last_layer_output[10510] + last_layer_output[10511] + last_layer_output[10512] + last_layer_output[10513] + last_layer_output[10514] + last_layer_output[10515] + last_layer_output[10516] + last_layer_output[10517] + last_layer_output[10518] + last_layer_output[10519] + last_layer_output[10520] + last_layer_output[10521] + last_layer_output[10522] + last_layer_output[10523] + last_layer_output[10524] + last_layer_output[10525] + last_layer_output[10526] + last_layer_output[10527] + last_layer_output[10528] + last_layer_output[10529] + last_layer_output[10530] + last_layer_output[10531] + last_layer_output[10532] + last_layer_output[10533] + last_layer_output[10534] + last_layer_output[10535] + last_layer_output[10536] + last_layer_output[10537] + last_layer_output[10538] + last_layer_output[10539] + last_layer_output[10540] + last_layer_output[10541] + last_layer_output[10542] + last_layer_output[10543] + last_layer_output[10544] + last_layer_output[10545] + last_layer_output[10546] + last_layer_output[10547] + last_layer_output[10548] + last_layer_output[10549] + last_layer_output[10550] + last_layer_output[10551] + last_layer_output[10552] + last_layer_output[10553] + last_layer_output[10554] + last_layer_output[10555] + last_layer_output[10556] + last_layer_output[10557] + last_layer_output[10558] + last_layer_output[10559] + last_layer_output[10560] + last_layer_output[10561] + last_layer_output[10562] + last_layer_output[10563] + last_layer_output[10564] + last_layer_output[10565] + last_layer_output[10566] + last_layer_output[10567] + last_layer_output[10568] + last_layer_output[10569] + last_layer_output[10570] + last_layer_output[10571] + last_layer_output[10572] + last_layer_output[10573] + last_layer_output[10574] + last_layer_output[10575] + last_layer_output[10576] + last_layer_output[10577] + last_layer_output[10578] + last_layer_output[10579] + last_layer_output[10580] + last_layer_output[10581] + last_layer_output[10582] + last_layer_output[10583] + last_layer_output[10584] + last_layer_output[10585] + last_layer_output[10586] + last_layer_output[10587] + last_layer_output[10588] + last_layer_output[10589] + last_layer_output[10590] + last_layer_output[10591] + last_layer_output[10592] + last_layer_output[10593] + last_layer_output[10594] + last_layer_output[10595] + last_layer_output[10596] + last_layer_output[10597] + last_layer_output[10598] + last_layer_output[10599] + last_layer_output[10600] + last_layer_output[10601] + last_layer_output[10602] + last_layer_output[10603] + last_layer_output[10604] + last_layer_output[10605] + last_layer_output[10606] + last_layer_output[10607] + last_layer_output[10608] + last_layer_output[10609] + last_layer_output[10610] + last_layer_output[10611] + last_layer_output[10612] + last_layer_output[10613] + last_layer_output[10614] + last_layer_output[10615] + last_layer_output[10616] + last_layer_output[10617] + last_layer_output[10618] + last_layer_output[10619] + last_layer_output[10620] + last_layer_output[10621] + last_layer_output[10622] + last_layer_output[10623] + last_layer_output[10624] + last_layer_output[10625] + last_layer_output[10626] + last_layer_output[10627] + last_layer_output[10628] + last_layer_output[10629] + last_layer_output[10630] + last_layer_output[10631] + last_layer_output[10632] + last_layer_output[10633] + last_layer_output[10634] + last_layer_output[10635] + last_layer_output[10636] + last_layer_output[10637] + last_layer_output[10638] + last_layer_output[10639] + last_layer_output[10640] + last_layer_output[10641] + last_layer_output[10642] + last_layer_output[10643] + last_layer_output[10644] + last_layer_output[10645] + last_layer_output[10646] + last_layer_output[10647] + last_layer_output[10648] + last_layer_output[10649] + last_layer_output[10650] + last_layer_output[10651] + last_layer_output[10652] + last_layer_output[10653] + last_layer_output[10654] + last_layer_output[10655] + last_layer_output[10656] + last_layer_output[10657] + last_layer_output[10658] + last_layer_output[10659] + last_layer_output[10660] + last_layer_output[10661] + last_layer_output[10662] + last_layer_output[10663] + last_layer_output[10664] + last_layer_output[10665] + last_layer_output[10666] + last_layer_output[10667] + last_layer_output[10668] + last_layer_output[10669] + last_layer_output[10670] + last_layer_output[10671] + last_layer_output[10672] + last_layer_output[10673] + last_layer_output[10674] + last_layer_output[10675] + last_layer_output[10676] + last_layer_output[10677] + last_layer_output[10678] + last_layer_output[10679] + last_layer_output[10680] + last_layer_output[10681] + last_layer_output[10682] + last_layer_output[10683] + last_layer_output[10684] + last_layer_output[10685] + last_layer_output[10686] + last_layer_output[10687] + last_layer_output[10688] + last_layer_output[10689] + last_layer_output[10690] + last_layer_output[10691] + last_layer_output[10692] + last_layer_output[10693] + last_layer_output[10694] + last_layer_output[10695] + last_layer_output[10696] + last_layer_output[10697] + last_layer_output[10698] + last_layer_output[10699] + last_layer_output[10700] + last_layer_output[10701] + last_layer_output[10702] + last_layer_output[10703] + last_layer_output[10704] + last_layer_output[10705] + last_layer_output[10706] + last_layer_output[10707] + last_layer_output[10708] + last_layer_output[10709] + last_layer_output[10710] + last_layer_output[10711] + last_layer_output[10712] + last_layer_output[10713] + last_layer_output[10714] + last_layer_output[10715] + last_layer_output[10716] + last_layer_output[10717] + last_layer_output[10718] + last_layer_output[10719] + last_layer_output[10720] + last_layer_output[10721] + last_layer_output[10722] + last_layer_output[10723] + last_layer_output[10724] + last_layer_output[10725] + last_layer_output[10726] + last_layer_output[10727] + last_layer_output[10728] + last_layer_output[10729] + last_layer_output[10730] + last_layer_output[10731] + last_layer_output[10732] + last_layer_output[10733] + last_layer_output[10734] + last_layer_output[10735] + last_layer_output[10736] + last_layer_output[10737] + last_layer_output[10738] + last_layer_output[10739] + last_layer_output[10740] + last_layer_output[10741] + last_layer_output[10742] + last_layer_output[10743] + last_layer_output[10744] + last_layer_output[10745] + last_layer_output[10746] + last_layer_output[10747] + last_layer_output[10748] + last_layer_output[10749] + last_layer_output[10750] + last_layer_output[10751] + last_layer_output[10752] + last_layer_output[10753] + last_layer_output[10754] + last_layer_output[10755] + last_layer_output[10756] + last_layer_output[10757] + last_layer_output[10758] + last_layer_output[10759] + last_layer_output[10760] + last_layer_output[10761] + last_layer_output[10762] + last_layer_output[10763] + last_layer_output[10764] + last_layer_output[10765] + last_layer_output[10766] + last_layer_output[10767] + last_layer_output[10768] + last_layer_output[10769] + last_layer_output[10770] + last_layer_output[10771] + last_layer_output[10772] + last_layer_output[10773] + last_layer_output[10774] + last_layer_output[10775] + last_layer_output[10776] + last_layer_output[10777] + last_layer_output[10778] + last_layer_output[10779] + last_layer_output[10780] + last_layer_output[10781] + last_layer_output[10782] + last_layer_output[10783] + last_layer_output[10784] + last_layer_output[10785] + last_layer_output[10786] + last_layer_output[10787] + last_layer_output[10788] + last_layer_output[10789] + last_layer_output[10790] + last_layer_output[10791] + last_layer_output[10792] + last_layer_output[10793] + last_layer_output[10794] + last_layer_output[10795] + last_layer_output[10796] + last_layer_output[10797] + last_layer_output[10798] + last_layer_output[10799];
      result[9] <= last_layer_output[10800] + last_layer_output[10801] + last_layer_output[10802] + last_layer_output[10803] + last_layer_output[10804] + last_layer_output[10805] + last_layer_output[10806] + last_layer_output[10807] + last_layer_output[10808] + last_layer_output[10809] + last_layer_output[10810] + last_layer_output[10811] + last_layer_output[10812] + last_layer_output[10813] + last_layer_output[10814] + last_layer_output[10815] + last_layer_output[10816] + last_layer_output[10817] + last_layer_output[10818] + last_layer_output[10819] + last_layer_output[10820] + last_layer_output[10821] + last_layer_output[10822] + last_layer_output[10823] + last_layer_output[10824] + last_layer_output[10825] + last_layer_output[10826] + last_layer_output[10827] + last_layer_output[10828] + last_layer_output[10829] + last_layer_output[10830] + last_layer_output[10831] + last_layer_output[10832] + last_layer_output[10833] + last_layer_output[10834] + last_layer_output[10835] + last_layer_output[10836] + last_layer_output[10837] + last_layer_output[10838] + last_layer_output[10839] + last_layer_output[10840] + last_layer_output[10841] + last_layer_output[10842] + last_layer_output[10843] + last_layer_output[10844] + last_layer_output[10845] + last_layer_output[10846] + last_layer_output[10847] + last_layer_output[10848] + last_layer_output[10849] + last_layer_output[10850] + last_layer_output[10851] + last_layer_output[10852] + last_layer_output[10853] + last_layer_output[10854] + last_layer_output[10855] + last_layer_output[10856] + last_layer_output[10857] + last_layer_output[10858] + last_layer_output[10859] + last_layer_output[10860] + last_layer_output[10861] + last_layer_output[10862] + last_layer_output[10863] + last_layer_output[10864] + last_layer_output[10865] + last_layer_output[10866] + last_layer_output[10867] + last_layer_output[10868] + last_layer_output[10869] + last_layer_output[10870] + last_layer_output[10871] + last_layer_output[10872] + last_layer_output[10873] + last_layer_output[10874] + last_layer_output[10875] + last_layer_output[10876] + last_layer_output[10877] + last_layer_output[10878] + last_layer_output[10879] + last_layer_output[10880] + last_layer_output[10881] + last_layer_output[10882] + last_layer_output[10883] + last_layer_output[10884] + last_layer_output[10885] + last_layer_output[10886] + last_layer_output[10887] + last_layer_output[10888] + last_layer_output[10889] + last_layer_output[10890] + last_layer_output[10891] + last_layer_output[10892] + last_layer_output[10893] + last_layer_output[10894] + last_layer_output[10895] + last_layer_output[10896] + last_layer_output[10897] + last_layer_output[10898] + last_layer_output[10899] + last_layer_output[10900] + last_layer_output[10901] + last_layer_output[10902] + last_layer_output[10903] + last_layer_output[10904] + last_layer_output[10905] + last_layer_output[10906] + last_layer_output[10907] + last_layer_output[10908] + last_layer_output[10909] + last_layer_output[10910] + last_layer_output[10911] + last_layer_output[10912] + last_layer_output[10913] + last_layer_output[10914] + last_layer_output[10915] + last_layer_output[10916] + last_layer_output[10917] + last_layer_output[10918] + last_layer_output[10919] + last_layer_output[10920] + last_layer_output[10921] + last_layer_output[10922] + last_layer_output[10923] + last_layer_output[10924] + last_layer_output[10925] + last_layer_output[10926] + last_layer_output[10927] + last_layer_output[10928] + last_layer_output[10929] + last_layer_output[10930] + last_layer_output[10931] + last_layer_output[10932] + last_layer_output[10933] + last_layer_output[10934] + last_layer_output[10935] + last_layer_output[10936] + last_layer_output[10937] + last_layer_output[10938] + last_layer_output[10939] + last_layer_output[10940] + last_layer_output[10941] + last_layer_output[10942] + last_layer_output[10943] + last_layer_output[10944] + last_layer_output[10945] + last_layer_output[10946] + last_layer_output[10947] + last_layer_output[10948] + last_layer_output[10949] + last_layer_output[10950] + last_layer_output[10951] + last_layer_output[10952] + last_layer_output[10953] + last_layer_output[10954] + last_layer_output[10955] + last_layer_output[10956] + last_layer_output[10957] + last_layer_output[10958] + last_layer_output[10959] + last_layer_output[10960] + last_layer_output[10961] + last_layer_output[10962] + last_layer_output[10963] + last_layer_output[10964] + last_layer_output[10965] + last_layer_output[10966] + last_layer_output[10967] + last_layer_output[10968] + last_layer_output[10969] + last_layer_output[10970] + last_layer_output[10971] + last_layer_output[10972] + last_layer_output[10973] + last_layer_output[10974] + last_layer_output[10975] + last_layer_output[10976] + last_layer_output[10977] + last_layer_output[10978] + last_layer_output[10979] + last_layer_output[10980] + last_layer_output[10981] + last_layer_output[10982] + last_layer_output[10983] + last_layer_output[10984] + last_layer_output[10985] + last_layer_output[10986] + last_layer_output[10987] + last_layer_output[10988] + last_layer_output[10989] + last_layer_output[10990] + last_layer_output[10991] + last_layer_output[10992] + last_layer_output[10993] + last_layer_output[10994] + last_layer_output[10995] + last_layer_output[10996] + last_layer_output[10997] + last_layer_output[10998] + last_layer_output[10999] + last_layer_output[11000] + last_layer_output[11001] + last_layer_output[11002] + last_layer_output[11003] + last_layer_output[11004] + last_layer_output[11005] + last_layer_output[11006] + last_layer_output[11007] + last_layer_output[11008] + last_layer_output[11009] + last_layer_output[11010] + last_layer_output[11011] + last_layer_output[11012] + last_layer_output[11013] + last_layer_output[11014] + last_layer_output[11015] + last_layer_output[11016] + last_layer_output[11017] + last_layer_output[11018] + last_layer_output[11019] + last_layer_output[11020] + last_layer_output[11021] + last_layer_output[11022] + last_layer_output[11023] + last_layer_output[11024] + last_layer_output[11025] + last_layer_output[11026] + last_layer_output[11027] + last_layer_output[11028] + last_layer_output[11029] + last_layer_output[11030] + last_layer_output[11031] + last_layer_output[11032] + last_layer_output[11033] + last_layer_output[11034] + last_layer_output[11035] + last_layer_output[11036] + last_layer_output[11037] + last_layer_output[11038] + last_layer_output[11039] + last_layer_output[11040] + last_layer_output[11041] + last_layer_output[11042] + last_layer_output[11043] + last_layer_output[11044] + last_layer_output[11045] + last_layer_output[11046] + last_layer_output[11047] + last_layer_output[11048] + last_layer_output[11049] + last_layer_output[11050] + last_layer_output[11051] + last_layer_output[11052] + last_layer_output[11053] + last_layer_output[11054] + last_layer_output[11055] + last_layer_output[11056] + last_layer_output[11057] + last_layer_output[11058] + last_layer_output[11059] + last_layer_output[11060] + last_layer_output[11061] + last_layer_output[11062] + last_layer_output[11063] + last_layer_output[11064] + last_layer_output[11065] + last_layer_output[11066] + last_layer_output[11067] + last_layer_output[11068] + last_layer_output[11069] + last_layer_output[11070] + last_layer_output[11071] + last_layer_output[11072] + last_layer_output[11073] + last_layer_output[11074] + last_layer_output[11075] + last_layer_output[11076] + last_layer_output[11077] + last_layer_output[11078] + last_layer_output[11079] + last_layer_output[11080] + last_layer_output[11081] + last_layer_output[11082] + last_layer_output[11083] + last_layer_output[11084] + last_layer_output[11085] + last_layer_output[11086] + last_layer_output[11087] + last_layer_output[11088] + last_layer_output[11089] + last_layer_output[11090] + last_layer_output[11091] + last_layer_output[11092] + last_layer_output[11093] + last_layer_output[11094] + last_layer_output[11095] + last_layer_output[11096] + last_layer_output[11097] + last_layer_output[11098] + last_layer_output[11099] + last_layer_output[11100] + last_layer_output[11101] + last_layer_output[11102] + last_layer_output[11103] + last_layer_output[11104] + last_layer_output[11105] + last_layer_output[11106] + last_layer_output[11107] + last_layer_output[11108] + last_layer_output[11109] + last_layer_output[11110] + last_layer_output[11111] + last_layer_output[11112] + last_layer_output[11113] + last_layer_output[11114] + last_layer_output[11115] + last_layer_output[11116] + last_layer_output[11117] + last_layer_output[11118] + last_layer_output[11119] + last_layer_output[11120] + last_layer_output[11121] + last_layer_output[11122] + last_layer_output[11123] + last_layer_output[11124] + last_layer_output[11125] + last_layer_output[11126] + last_layer_output[11127] + last_layer_output[11128] + last_layer_output[11129] + last_layer_output[11130] + last_layer_output[11131] + last_layer_output[11132] + last_layer_output[11133] + last_layer_output[11134] + last_layer_output[11135] + last_layer_output[11136] + last_layer_output[11137] + last_layer_output[11138] + last_layer_output[11139] + last_layer_output[11140] + last_layer_output[11141] + last_layer_output[11142] + last_layer_output[11143] + last_layer_output[11144] + last_layer_output[11145] + last_layer_output[11146] + last_layer_output[11147] + last_layer_output[11148] + last_layer_output[11149] + last_layer_output[11150] + last_layer_output[11151] + last_layer_output[11152] + last_layer_output[11153] + last_layer_output[11154] + last_layer_output[11155] + last_layer_output[11156] + last_layer_output[11157] + last_layer_output[11158] + last_layer_output[11159] + last_layer_output[11160] + last_layer_output[11161] + last_layer_output[11162] + last_layer_output[11163] + last_layer_output[11164] + last_layer_output[11165] + last_layer_output[11166] + last_layer_output[11167] + last_layer_output[11168] + last_layer_output[11169] + last_layer_output[11170] + last_layer_output[11171] + last_layer_output[11172] + last_layer_output[11173] + last_layer_output[11174] + last_layer_output[11175] + last_layer_output[11176] + last_layer_output[11177] + last_layer_output[11178] + last_layer_output[11179] + last_layer_output[11180] + last_layer_output[11181] + last_layer_output[11182] + last_layer_output[11183] + last_layer_output[11184] + last_layer_output[11185] + last_layer_output[11186] + last_layer_output[11187] + last_layer_output[11188] + last_layer_output[11189] + last_layer_output[11190] + last_layer_output[11191] + last_layer_output[11192] + last_layer_output[11193] + last_layer_output[11194] + last_layer_output[11195] + last_layer_output[11196] + last_layer_output[11197] + last_layer_output[11198] + last_layer_output[11199] + last_layer_output[11200] + last_layer_output[11201] + last_layer_output[11202] + last_layer_output[11203] + last_layer_output[11204] + last_layer_output[11205] + last_layer_output[11206] + last_layer_output[11207] + last_layer_output[11208] + last_layer_output[11209] + last_layer_output[11210] + last_layer_output[11211] + last_layer_output[11212] + last_layer_output[11213] + last_layer_output[11214] + last_layer_output[11215] + last_layer_output[11216] + last_layer_output[11217] + last_layer_output[11218] + last_layer_output[11219] + last_layer_output[11220] + last_layer_output[11221] + last_layer_output[11222] + last_layer_output[11223] + last_layer_output[11224] + last_layer_output[11225] + last_layer_output[11226] + last_layer_output[11227] + last_layer_output[11228] + last_layer_output[11229] + last_layer_output[11230] + last_layer_output[11231] + last_layer_output[11232] + last_layer_output[11233] + last_layer_output[11234] + last_layer_output[11235] + last_layer_output[11236] + last_layer_output[11237] + last_layer_output[11238] + last_layer_output[11239] + last_layer_output[11240] + last_layer_output[11241] + last_layer_output[11242] + last_layer_output[11243] + last_layer_output[11244] + last_layer_output[11245] + last_layer_output[11246] + last_layer_output[11247] + last_layer_output[11248] + last_layer_output[11249] + last_layer_output[11250] + last_layer_output[11251] + last_layer_output[11252] + last_layer_output[11253] + last_layer_output[11254] + last_layer_output[11255] + last_layer_output[11256] + last_layer_output[11257] + last_layer_output[11258] + last_layer_output[11259] + last_layer_output[11260] + last_layer_output[11261] + last_layer_output[11262] + last_layer_output[11263] + last_layer_output[11264] + last_layer_output[11265] + last_layer_output[11266] + last_layer_output[11267] + last_layer_output[11268] + last_layer_output[11269] + last_layer_output[11270] + last_layer_output[11271] + last_layer_output[11272] + last_layer_output[11273] + last_layer_output[11274] + last_layer_output[11275] + last_layer_output[11276] + last_layer_output[11277] + last_layer_output[11278] + last_layer_output[11279] + last_layer_output[11280] + last_layer_output[11281] + last_layer_output[11282] + last_layer_output[11283] + last_layer_output[11284] + last_layer_output[11285] + last_layer_output[11286] + last_layer_output[11287] + last_layer_output[11288] + last_layer_output[11289] + last_layer_output[11290] + last_layer_output[11291] + last_layer_output[11292] + last_layer_output[11293] + last_layer_output[11294] + last_layer_output[11295] + last_layer_output[11296] + last_layer_output[11297] + last_layer_output[11298] + last_layer_output[11299] + last_layer_output[11300] + last_layer_output[11301] + last_layer_output[11302] + last_layer_output[11303] + last_layer_output[11304] + last_layer_output[11305] + last_layer_output[11306] + last_layer_output[11307] + last_layer_output[11308] + last_layer_output[11309] + last_layer_output[11310] + last_layer_output[11311] + last_layer_output[11312] + last_layer_output[11313] + last_layer_output[11314] + last_layer_output[11315] + last_layer_output[11316] + last_layer_output[11317] + last_layer_output[11318] + last_layer_output[11319] + last_layer_output[11320] + last_layer_output[11321] + last_layer_output[11322] + last_layer_output[11323] + last_layer_output[11324] + last_layer_output[11325] + last_layer_output[11326] + last_layer_output[11327] + last_layer_output[11328] + last_layer_output[11329] + last_layer_output[11330] + last_layer_output[11331] + last_layer_output[11332] + last_layer_output[11333] + last_layer_output[11334] + last_layer_output[11335] + last_layer_output[11336] + last_layer_output[11337] + last_layer_output[11338] + last_layer_output[11339] + last_layer_output[11340] + last_layer_output[11341] + last_layer_output[11342] + last_layer_output[11343] + last_layer_output[11344] + last_layer_output[11345] + last_layer_output[11346] + last_layer_output[11347] + last_layer_output[11348] + last_layer_output[11349] + last_layer_output[11350] + last_layer_output[11351] + last_layer_output[11352] + last_layer_output[11353] + last_layer_output[11354] + last_layer_output[11355] + last_layer_output[11356] + last_layer_output[11357] + last_layer_output[11358] + last_layer_output[11359] + last_layer_output[11360] + last_layer_output[11361] + last_layer_output[11362] + last_layer_output[11363] + last_layer_output[11364] + last_layer_output[11365] + last_layer_output[11366] + last_layer_output[11367] + last_layer_output[11368] + last_layer_output[11369] + last_layer_output[11370] + last_layer_output[11371] + last_layer_output[11372] + last_layer_output[11373] + last_layer_output[11374] + last_layer_output[11375] + last_layer_output[11376] + last_layer_output[11377] + last_layer_output[11378] + last_layer_output[11379] + last_layer_output[11380] + last_layer_output[11381] + last_layer_output[11382] + last_layer_output[11383] + last_layer_output[11384] + last_layer_output[11385] + last_layer_output[11386] + last_layer_output[11387] + last_layer_output[11388] + last_layer_output[11389] + last_layer_output[11390] + last_layer_output[11391] + last_layer_output[11392] + last_layer_output[11393] + last_layer_output[11394] + last_layer_output[11395] + last_layer_output[11396] + last_layer_output[11397] + last_layer_output[11398] + last_layer_output[11399] + last_layer_output[11400] + last_layer_output[11401] + last_layer_output[11402] + last_layer_output[11403] + last_layer_output[11404] + last_layer_output[11405] + last_layer_output[11406] + last_layer_output[11407] + last_layer_output[11408] + last_layer_output[11409] + last_layer_output[11410] + last_layer_output[11411] + last_layer_output[11412] + last_layer_output[11413] + last_layer_output[11414] + last_layer_output[11415] + last_layer_output[11416] + last_layer_output[11417] + last_layer_output[11418] + last_layer_output[11419] + last_layer_output[11420] + last_layer_output[11421] + last_layer_output[11422] + last_layer_output[11423] + last_layer_output[11424] + last_layer_output[11425] + last_layer_output[11426] + last_layer_output[11427] + last_layer_output[11428] + last_layer_output[11429] + last_layer_output[11430] + last_layer_output[11431] + last_layer_output[11432] + last_layer_output[11433] + last_layer_output[11434] + last_layer_output[11435] + last_layer_output[11436] + last_layer_output[11437] + last_layer_output[11438] + last_layer_output[11439] + last_layer_output[11440] + last_layer_output[11441] + last_layer_output[11442] + last_layer_output[11443] + last_layer_output[11444] + last_layer_output[11445] + last_layer_output[11446] + last_layer_output[11447] + last_layer_output[11448] + last_layer_output[11449] + last_layer_output[11450] + last_layer_output[11451] + last_layer_output[11452] + last_layer_output[11453] + last_layer_output[11454] + last_layer_output[11455] + last_layer_output[11456] + last_layer_output[11457] + last_layer_output[11458] + last_layer_output[11459] + last_layer_output[11460] + last_layer_output[11461] + last_layer_output[11462] + last_layer_output[11463] + last_layer_output[11464] + last_layer_output[11465] + last_layer_output[11466] + last_layer_output[11467] + last_layer_output[11468] + last_layer_output[11469] + last_layer_output[11470] + last_layer_output[11471] + last_layer_output[11472] + last_layer_output[11473] + last_layer_output[11474] + last_layer_output[11475] + last_layer_output[11476] + last_layer_output[11477] + last_layer_output[11478] + last_layer_output[11479] + last_layer_output[11480] + last_layer_output[11481] + last_layer_output[11482] + last_layer_output[11483] + last_layer_output[11484] + last_layer_output[11485] + last_layer_output[11486] + last_layer_output[11487] + last_layer_output[11488] + last_layer_output[11489] + last_layer_output[11490] + last_layer_output[11491] + last_layer_output[11492] + last_layer_output[11493] + last_layer_output[11494] + last_layer_output[11495] + last_layer_output[11496] + last_layer_output[11497] + last_layer_output[11498] + last_layer_output[11499] + last_layer_output[11500] + last_layer_output[11501] + last_layer_output[11502] + last_layer_output[11503] + last_layer_output[11504] + last_layer_output[11505] + last_layer_output[11506] + last_layer_output[11507] + last_layer_output[11508] + last_layer_output[11509] + last_layer_output[11510] + last_layer_output[11511] + last_layer_output[11512] + last_layer_output[11513] + last_layer_output[11514] + last_layer_output[11515] + last_layer_output[11516] + last_layer_output[11517] + last_layer_output[11518] + last_layer_output[11519] + last_layer_output[11520] + last_layer_output[11521] + last_layer_output[11522] + last_layer_output[11523] + last_layer_output[11524] + last_layer_output[11525] + last_layer_output[11526] + last_layer_output[11527] + last_layer_output[11528] + last_layer_output[11529] + last_layer_output[11530] + last_layer_output[11531] + last_layer_output[11532] + last_layer_output[11533] + last_layer_output[11534] + last_layer_output[11535] + last_layer_output[11536] + last_layer_output[11537] + last_layer_output[11538] + last_layer_output[11539] + last_layer_output[11540] + last_layer_output[11541] + last_layer_output[11542] + last_layer_output[11543] + last_layer_output[11544] + last_layer_output[11545] + last_layer_output[11546] + last_layer_output[11547] + last_layer_output[11548] + last_layer_output[11549] + last_layer_output[11550] + last_layer_output[11551] + last_layer_output[11552] + last_layer_output[11553] + last_layer_output[11554] + last_layer_output[11555] + last_layer_output[11556] + last_layer_output[11557] + last_layer_output[11558] + last_layer_output[11559] + last_layer_output[11560] + last_layer_output[11561] + last_layer_output[11562] + last_layer_output[11563] + last_layer_output[11564] + last_layer_output[11565] + last_layer_output[11566] + last_layer_output[11567] + last_layer_output[11568] + last_layer_output[11569] + last_layer_output[11570] + last_layer_output[11571] + last_layer_output[11572] + last_layer_output[11573] + last_layer_output[11574] + last_layer_output[11575] + last_layer_output[11576] + last_layer_output[11577] + last_layer_output[11578] + last_layer_output[11579] + last_layer_output[11580] + last_layer_output[11581] + last_layer_output[11582] + last_layer_output[11583] + last_layer_output[11584] + last_layer_output[11585] + last_layer_output[11586] + last_layer_output[11587] + last_layer_output[11588] + last_layer_output[11589] + last_layer_output[11590] + last_layer_output[11591] + last_layer_output[11592] + last_layer_output[11593] + last_layer_output[11594] + last_layer_output[11595] + last_layer_output[11596] + last_layer_output[11597] + last_layer_output[11598] + last_layer_output[11599] + last_layer_output[11600] + last_layer_output[11601] + last_layer_output[11602] + last_layer_output[11603] + last_layer_output[11604] + last_layer_output[11605] + last_layer_output[11606] + last_layer_output[11607] + last_layer_output[11608] + last_layer_output[11609] + last_layer_output[11610] + last_layer_output[11611] + last_layer_output[11612] + last_layer_output[11613] + last_layer_output[11614] + last_layer_output[11615] + last_layer_output[11616] + last_layer_output[11617] + last_layer_output[11618] + last_layer_output[11619] + last_layer_output[11620] + last_layer_output[11621] + last_layer_output[11622] + last_layer_output[11623] + last_layer_output[11624] + last_layer_output[11625] + last_layer_output[11626] + last_layer_output[11627] + last_layer_output[11628] + last_layer_output[11629] + last_layer_output[11630] + last_layer_output[11631] + last_layer_output[11632] + last_layer_output[11633] + last_layer_output[11634] + last_layer_output[11635] + last_layer_output[11636] + last_layer_output[11637] + last_layer_output[11638] + last_layer_output[11639] + last_layer_output[11640] + last_layer_output[11641] + last_layer_output[11642] + last_layer_output[11643] + last_layer_output[11644] + last_layer_output[11645] + last_layer_output[11646] + last_layer_output[11647] + last_layer_output[11648] + last_layer_output[11649] + last_layer_output[11650] + last_layer_output[11651] + last_layer_output[11652] + last_layer_output[11653] + last_layer_output[11654] + last_layer_output[11655] + last_layer_output[11656] + last_layer_output[11657] + last_layer_output[11658] + last_layer_output[11659] + last_layer_output[11660] + last_layer_output[11661] + last_layer_output[11662] + last_layer_output[11663] + last_layer_output[11664] + last_layer_output[11665] + last_layer_output[11666] + last_layer_output[11667] + last_layer_output[11668] + last_layer_output[11669] + last_layer_output[11670] + last_layer_output[11671] + last_layer_output[11672] + last_layer_output[11673] + last_layer_output[11674] + last_layer_output[11675] + last_layer_output[11676] + last_layer_output[11677] + last_layer_output[11678] + last_layer_output[11679] + last_layer_output[11680] + last_layer_output[11681] + last_layer_output[11682] + last_layer_output[11683] + last_layer_output[11684] + last_layer_output[11685] + last_layer_output[11686] + last_layer_output[11687] + last_layer_output[11688] + last_layer_output[11689] + last_layer_output[11690] + last_layer_output[11691] + last_layer_output[11692] + last_layer_output[11693] + last_layer_output[11694] + last_layer_output[11695] + last_layer_output[11696] + last_layer_output[11697] + last_layer_output[11698] + last_layer_output[11699] + last_layer_output[11700] + last_layer_output[11701] + last_layer_output[11702] + last_layer_output[11703] + last_layer_output[11704] + last_layer_output[11705] + last_layer_output[11706] + last_layer_output[11707] + last_layer_output[11708] + last_layer_output[11709] + last_layer_output[11710] + last_layer_output[11711] + last_layer_output[11712] + last_layer_output[11713] + last_layer_output[11714] + last_layer_output[11715] + last_layer_output[11716] + last_layer_output[11717] + last_layer_output[11718] + last_layer_output[11719] + last_layer_output[11720] + last_layer_output[11721] + last_layer_output[11722] + last_layer_output[11723] + last_layer_output[11724] + last_layer_output[11725] + last_layer_output[11726] + last_layer_output[11727] + last_layer_output[11728] + last_layer_output[11729] + last_layer_output[11730] + last_layer_output[11731] + last_layer_output[11732] + last_layer_output[11733] + last_layer_output[11734] + last_layer_output[11735] + last_layer_output[11736] + last_layer_output[11737] + last_layer_output[11738] + last_layer_output[11739] + last_layer_output[11740] + last_layer_output[11741] + last_layer_output[11742] + last_layer_output[11743] + last_layer_output[11744] + last_layer_output[11745] + last_layer_output[11746] + last_layer_output[11747] + last_layer_output[11748] + last_layer_output[11749] + last_layer_output[11750] + last_layer_output[11751] + last_layer_output[11752] + last_layer_output[11753] + last_layer_output[11754] + last_layer_output[11755] + last_layer_output[11756] + last_layer_output[11757] + last_layer_output[11758] + last_layer_output[11759] + last_layer_output[11760] + last_layer_output[11761] + last_layer_output[11762] + last_layer_output[11763] + last_layer_output[11764] + last_layer_output[11765] + last_layer_output[11766] + last_layer_output[11767] + last_layer_output[11768] + last_layer_output[11769] + last_layer_output[11770] + last_layer_output[11771] + last_layer_output[11772] + last_layer_output[11773] + last_layer_output[11774] + last_layer_output[11775] + last_layer_output[11776] + last_layer_output[11777] + last_layer_output[11778] + last_layer_output[11779] + last_layer_output[11780] + last_layer_output[11781] + last_layer_output[11782] + last_layer_output[11783] + last_layer_output[11784] + last_layer_output[11785] + last_layer_output[11786] + last_layer_output[11787] + last_layer_output[11788] + last_layer_output[11789] + last_layer_output[11790] + last_layer_output[11791] + last_layer_output[11792] + last_layer_output[11793] + last_layer_output[11794] + last_layer_output[11795] + last_layer_output[11796] + last_layer_output[11797] + last_layer_output[11798] + last_layer_output[11799] + last_layer_output[11800] + last_layer_output[11801] + last_layer_output[11802] + last_layer_output[11803] + last_layer_output[11804] + last_layer_output[11805] + last_layer_output[11806] + last_layer_output[11807] + last_layer_output[11808] + last_layer_output[11809] + last_layer_output[11810] + last_layer_output[11811] + last_layer_output[11812] + last_layer_output[11813] + last_layer_output[11814] + last_layer_output[11815] + last_layer_output[11816] + last_layer_output[11817] + last_layer_output[11818] + last_layer_output[11819] + last_layer_output[11820] + last_layer_output[11821] + last_layer_output[11822] + last_layer_output[11823] + last_layer_output[11824] + last_layer_output[11825] + last_layer_output[11826] + last_layer_output[11827] + last_layer_output[11828] + last_layer_output[11829] + last_layer_output[11830] + last_layer_output[11831] + last_layer_output[11832] + last_layer_output[11833] + last_layer_output[11834] + last_layer_output[11835] + last_layer_output[11836] + last_layer_output[11837] + last_layer_output[11838] + last_layer_output[11839] + last_layer_output[11840] + last_layer_output[11841] + last_layer_output[11842] + last_layer_output[11843] + last_layer_output[11844] + last_layer_output[11845] + last_layer_output[11846] + last_layer_output[11847] + last_layer_output[11848] + last_layer_output[11849] + last_layer_output[11850] + last_layer_output[11851] + last_layer_output[11852] + last_layer_output[11853] + last_layer_output[11854] + last_layer_output[11855] + last_layer_output[11856] + last_layer_output[11857] + last_layer_output[11858] + last_layer_output[11859] + last_layer_output[11860] + last_layer_output[11861] + last_layer_output[11862] + last_layer_output[11863] + last_layer_output[11864] + last_layer_output[11865] + last_layer_output[11866] + last_layer_output[11867] + last_layer_output[11868] + last_layer_output[11869] + last_layer_output[11870] + last_layer_output[11871] + last_layer_output[11872] + last_layer_output[11873] + last_layer_output[11874] + last_layer_output[11875] + last_layer_output[11876] + last_layer_output[11877] + last_layer_output[11878] + last_layer_output[11879] + last_layer_output[11880] + last_layer_output[11881] + last_layer_output[11882] + last_layer_output[11883] + last_layer_output[11884] + last_layer_output[11885] + last_layer_output[11886] + last_layer_output[11887] + last_layer_output[11888] + last_layer_output[11889] + last_layer_output[11890] + last_layer_output[11891] + last_layer_output[11892] + last_layer_output[11893] + last_layer_output[11894] + last_layer_output[11895] + last_layer_output[11896] + last_layer_output[11897] + last_layer_output[11898] + last_layer_output[11899] + last_layer_output[11900] + last_layer_output[11901] + last_layer_output[11902] + last_layer_output[11903] + last_layer_output[11904] + last_layer_output[11905] + last_layer_output[11906] + last_layer_output[11907] + last_layer_output[11908] + last_layer_output[11909] + last_layer_output[11910] + last_layer_output[11911] + last_layer_output[11912] + last_layer_output[11913] + last_layer_output[11914] + last_layer_output[11915] + last_layer_output[11916] + last_layer_output[11917] + last_layer_output[11918] + last_layer_output[11919] + last_layer_output[11920] + last_layer_output[11921] + last_layer_output[11922] + last_layer_output[11923] + last_layer_output[11924] + last_layer_output[11925] + last_layer_output[11926] + last_layer_output[11927] + last_layer_output[11928] + last_layer_output[11929] + last_layer_output[11930] + last_layer_output[11931] + last_layer_output[11932] + last_layer_output[11933] + last_layer_output[11934] + last_layer_output[11935] + last_layer_output[11936] + last_layer_output[11937] + last_layer_output[11938] + last_layer_output[11939] + last_layer_output[11940] + last_layer_output[11941] + last_layer_output[11942] + last_layer_output[11943] + last_layer_output[11944] + last_layer_output[11945] + last_layer_output[11946] + last_layer_output[11947] + last_layer_output[11948] + last_layer_output[11949] + last_layer_output[11950] + last_layer_output[11951] + last_layer_output[11952] + last_layer_output[11953] + last_layer_output[11954] + last_layer_output[11955] + last_layer_output[11956] + last_layer_output[11957] + last_layer_output[11958] + last_layer_output[11959] + last_layer_output[11960] + last_layer_output[11961] + last_layer_output[11962] + last_layer_output[11963] + last_layer_output[11964] + last_layer_output[11965] + last_layer_output[11966] + last_layer_output[11967] + last_layer_output[11968] + last_layer_output[11969] + last_layer_output[11970] + last_layer_output[11971] + last_layer_output[11972] + last_layer_output[11973] + last_layer_output[11974] + last_layer_output[11975] + last_layer_output[11976] + last_layer_output[11977] + last_layer_output[11978] + last_layer_output[11979] + last_layer_output[11980] + last_layer_output[11981] + last_layer_output[11982] + last_layer_output[11983] + last_layer_output[11984] + last_layer_output[11985] + last_layer_output[11986] + last_layer_output[11987] + last_layer_output[11988] + last_layer_output[11989] + last_layer_output[11990] + last_layer_output[11991] + last_layer_output[11992] + last_layer_output[11993] + last_layer_output[11994] + last_layer_output[11995] + last_layer_output[11996] + last_layer_output[11997] + last_layer_output[11998] + last_layer_output[11999];
end
      assign y[109:99]=result[0];
      assign y[98:88]=result[1];
      assign y[87:77]=result[2];
      assign y[76:66]=result[3];
      assign y[65:55]=result[4];
      assign y[54:44]=result[5];
      assign y[43:33]=result[6];
      assign y[32:22]=result[7];
      assign y[21:11]=result[8];
      assign y[10:0]=result[9];
endmodule
