module logic_network (    input wire [399:0] x,
    output wire [99:0] y
);
      wire [7999:0] layer0_out;
      wire [7999:0] layer1_out;
      wire [7999:0] layer2_out;
      wire [7999:0] layer3_out;
      wire [7999:0] layer4_out;
      wire [7999:0] layer5_out;
    assign layer0_out[0] = ~x[19] | x[8];
    assign layer0_out[1] = ~x[153];
    assign layer0_out[2] = ~x[91];
    assign layer0_out[3] = x[367] & x[376];
    assign layer0_out[4] = ~x[308];
    assign layer0_out[5] = x[316];
    assign layer0_out[6] = ~x[64];
    assign layer0_out[7] = ~(x[164] | x[166]);
    assign layer0_out[8] = 1'b0;
    assign layer0_out[9] = x[60] & x[75];
    assign layer0_out[10] = x[170] | x[188];
    assign layer0_out[11] = x[314] | x[321];
    assign layer0_out[12] = x[309];
    assign layer0_out[13] = x[309];
    assign layer0_out[14] = ~x[65];
    assign layer0_out[15] = ~x[152];
    assign layer0_out[16] = x[113] | x[129];
    assign layer0_out[17] = x[314] ^ x[320];
    assign layer0_out[18] = ~(x[381] | x[395]);
    assign layer0_out[19] = ~x[152];
    assign layer0_out[20] = 1'b0;
    assign layer0_out[21] = ~x[323];
    assign layer0_out[22] = x[279] | x[286];
    assign layer0_out[23] = x[105] | x[123];
    assign layer0_out[24] = ~(x[295] | x[297]);
    assign layer0_out[25] = x[320] & x[326];
    assign layer0_out[26] = ~x[130];
    assign layer0_out[27] = x[283] | x[287];
    assign layer0_out[28] = ~(x[126] & x[135]);
    assign layer0_out[29] = 1'b1;
    assign layer0_out[30] = ~(x[1] | x[15]);
    assign layer0_out[31] = ~(x[355] | x[360]);
    assign layer0_out[32] = x[24] | x[36];
    assign layer0_out[33] = x[329] & x[343];
    assign layer0_out[34] = x[8] | x[28];
    assign layer0_out[35] = ~(x[5] | x[23]);
    assign layer0_out[36] = 1'b1;
    assign layer0_out[37] = ~(x[226] & x[231]);
    assign layer0_out[38] = ~x[242];
    assign layer0_out[39] = ~x[108];
    assign layer0_out[40] = ~(x[369] | x[371]);
    assign layer0_out[41] = 1'b0;
    assign layer0_out[42] = x[79] | x[88];
    assign layer0_out[43] = x[46] ^ x[60];
    assign layer0_out[44] = x[287] | x[305];
    assign layer0_out[45] = ~(x[268] ^ x[271]);
    assign layer0_out[46] = ~x[170];
    assign layer0_out[47] = x[249] & ~x[257];
    assign layer0_out[48] = x[84] | x[104];
    assign layer0_out[49] = x[157] & x[167];
    assign layer0_out[50] = ~x[230] | x[217];
    assign layer0_out[51] = ~(x[277] | x[295]);
    assign layer0_out[52] = x[188] ^ x[190];
    assign layer0_out[53] = ~(x[332] & x[346]);
    assign layer0_out[54] = ~(x[5] | x[18]);
    assign layer0_out[55] = 1'b1;
    assign layer0_out[56] = x[25];
    assign layer0_out[57] = x[212];
    assign layer0_out[58] = x[119] | x[126];
    assign layer0_out[59] = ~(x[353] & x[369]);
    assign layer0_out[60] = ~(x[40] ^ x[45]);
    assign layer0_out[61] = x[316];
    assign layer0_out[62] = x[307] & x[327];
    assign layer0_out[63] = x[197];
    assign layer0_out[64] = x[232];
    assign layer0_out[65] = ~x[268];
    assign layer0_out[66] = x[156] ^ x[166];
    assign layer0_out[67] = x[65];
    assign layer0_out[68] = x[95];
    assign layer0_out[69] = x[139] & ~x[119];
    assign layer0_out[70] = x[187];
    assign layer0_out[71] = x[161] | x[163];
    assign layer0_out[72] = ~x[206];
    assign layer0_out[73] = x[216] & x[231];
    assign layer0_out[74] = ~(x[158] & x[177]);
    assign layer0_out[75] = ~x[230];
    assign layer0_out[76] = ~x[249];
    assign layer0_out[77] = ~x[92];
    assign layer0_out[78] = ~(x[360] | x[363]);
    assign layer0_out[79] = ~(x[5] | x[15]);
    assign layer0_out[80] = ~x[258] | x[250];
    assign layer0_out[81] = ~(x[127] | x[146]);
    assign layer0_out[82] = x[244] ^ x[263];
    assign layer0_out[83] = ~(x[276] ^ x[294]);
    assign layer0_out[84] = ~x[330];
    assign layer0_out[85] = ~x[288];
    assign layer0_out[86] = ~(x[386] & x[388]);
    assign layer0_out[87] = ~(x[117] | x[126]);
    assign layer0_out[88] = x[173] | x[179];
    assign layer0_out[89] = ~(x[60] ^ x[70]);
    assign layer0_out[90] = x[145] & x[166];
    assign layer0_out[91] = ~x[120];
    assign layer0_out[92] = x[47];
    assign layer0_out[93] = x[276] & x[279];
    assign layer0_out[94] = x[333] & ~x[313];
    assign layer0_out[95] = x[180] | x[191];
    assign layer0_out[96] = ~x[28] | x[11];
    assign layer0_out[97] = x[192];
    assign layer0_out[98] = ~(x[147] ^ x[156]);
    assign layer0_out[99] = x[159];
    assign layer0_out[100] = ~x[196];
    assign layer0_out[101] = ~x[383];
    assign layer0_out[102] = x[77] | x[98];
    assign layer0_out[103] = ~(x[46] & x[58]);
    assign layer0_out[104] = ~(x[209] & x[214]);
    assign layer0_out[105] = ~x[292] | x[309];
    assign layer0_out[106] = x[23];
    assign layer0_out[107] = ~x[50];
    assign layer0_out[108] = x[21] & ~x[15];
    assign layer0_out[109] = x[314] & ~x[327];
    assign layer0_out[110] = x[173] & ~x[177];
    assign layer0_out[111] = x[142];
    assign layer0_out[112] = ~x[146] | x[138];
    assign layer0_out[113] = x[250] & x[263];
    assign layer0_out[114] = x[56] | x[67];
    assign layer0_out[115] = x[16];
    assign layer0_out[116] = x[136];
    assign layer0_out[117] = ~x[12];
    assign layer0_out[118] = x[53] ^ x[72];
    assign layer0_out[119] = x[270] | x[272];
    assign layer0_out[120] = ~x[206];
    assign layer0_out[121] = ~(x[292] ^ x[312]);
    assign layer0_out[122] = x[126] & ~x[144];
    assign layer0_out[123] = ~(x[164] | x[176]);
    assign layer0_out[124] = x[342];
    assign layer0_out[125] = x[381];
    assign layer0_out[126] = ~x[157] | x[177];
    assign layer0_out[127] = x[23];
    assign layer0_out[128] = ~(x[303] | x[311]);
    assign layer0_out[129] = x[182] | x[197];
    assign layer0_out[130] = ~x[209];
    assign layer0_out[131] = x[395] & x[399];
    assign layer0_out[132] = ~(x[108] & x[129]);
    assign layer0_out[133] = 1'b0;
    assign layer0_out[134] = x[99] & ~x[82];
    assign layer0_out[135] = x[228] & ~x[227];
    assign layer0_out[136] = x[258];
    assign layer0_out[137] = x[353] & x[367];
    assign layer0_out[138] = ~(x[78] | x[86]);
    assign layer0_out[139] = x[176] & ~x[180];
    assign layer0_out[140] = x[303] | x[312];
    assign layer0_out[141] = x[20] | x[31];
    assign layer0_out[142] = x[375];
    assign layer0_out[143] = ~x[268] | x[260];
    assign layer0_out[144] = x[191] & x[209];
    assign layer0_out[145] = ~x[21] | x[8];
    assign layer0_out[146] = x[190] | x[207];
    assign layer0_out[147] = ~(x[376] | x[396]);
    assign layer0_out[148] = 1'b1;
    assign layer0_out[149] = x[100];
    assign layer0_out[150] = x[358] | x[371];
    assign layer0_out[151] = ~x[347];
    assign layer0_out[152] = ~x[63];
    assign layer0_out[153] = x[296] & ~x[305];
    assign layer0_out[154] = x[191] & ~x[179];
    assign layer0_out[155] = x[152] & ~x[144];
    assign layer0_out[156] = ~x[301];
    assign layer0_out[157] = x[337] | x[348];
    assign layer0_out[158] = ~(x[29] | x[41]);
    assign layer0_out[159] = x[238] & ~x[243];
    assign layer0_out[160] = ~(x[371] & x[373]);
    assign layer0_out[161] = x[327] | x[346];
    assign layer0_out[162] = ~(x[89] ^ x[109]);
    assign layer0_out[163] = x[249];
    assign layer0_out[164] = ~x[76] | x[88];
    assign layer0_out[165] = ~x[304] | x[318];
    assign layer0_out[166] = x[356] & ~x[371];
    assign layer0_out[167] = ~(x[80] ^ x[87]);
    assign layer0_out[168] = x[380] | x[395];
    assign layer0_out[169] = ~x[239] | x[223];
    assign layer0_out[170] = ~(x[175] | x[196]);
    assign layer0_out[171] = x[82];
    assign layer0_out[172] = x[309];
    assign layer0_out[173] = ~(x[24] | x[37]);
    assign layer0_out[174] = ~(x[252] | x[254]);
    assign layer0_out[175] = ~x[130] | x[139];
    assign layer0_out[176] = x[344] | x[363];
    assign layer0_out[177] = ~(x[346] & x[354]);
    assign layer0_out[178] = x[343] | x[352];
    assign layer0_out[179] = ~(x[117] | x[138]);
    assign layer0_out[180] = x[355] & x[373];
    assign layer0_out[181] = ~x[288] | x[301];
    assign layer0_out[182] = 1'b1;
    assign layer0_out[183] = ~x[218] | x[234];
    assign layer0_out[184] = ~x[40] | x[39];
    assign layer0_out[185] = ~x[372] | x[360];
    assign layer0_out[186] = x[292] ^ x[298];
    assign layer0_out[187] = ~x[331];
    assign layer0_out[188] = x[285] & ~x[301];
    assign layer0_out[189] = x[87] | x[95];
    assign layer0_out[190] = 1'b0;
    assign layer0_out[191] = ~(x[153] | x[156]);
    assign layer0_out[192] = x[265] | x[281];
    assign layer0_out[193] = 1'b1;
    assign layer0_out[194] = ~(x[325] ^ x[343]);
    assign layer0_out[195] = x[295] | x[303];
    assign layer0_out[196] = ~(x[96] & x[106]);
    assign layer0_out[197] = x[104] | x[120];
    assign layer0_out[198] = x[341] | x[350];
    assign layer0_out[199] = x[164] | x[184];
    assign layer0_out[200] = ~x[239];
    assign layer0_out[201] = x[304] | x[313];
    assign layer0_out[202] = ~(x[60] & x[63]);
    assign layer0_out[203] = x[332];
    assign layer0_out[204] = x[349] | x[364];
    assign layer0_out[205] = x[213] & ~x[225];
    assign layer0_out[206] = x[302] & ~x[314];
    assign layer0_out[207] = x[69] & ~x[56];
    assign layer0_out[208] = x[162] | x[173];
    assign layer0_out[209] = ~(x[205] | x[218]);
    assign layer0_out[210] = x[42] & x[60];
    assign layer0_out[211] = ~(x[187] | x[191]);
    assign layer0_out[212] = x[327];
    assign layer0_out[213] = x[54] ^ x[58];
    assign layer0_out[214] = x[172] & ~x[180];
    assign layer0_out[215] = ~(x[95] | x[99]);
    assign layer0_out[216] = ~(x[350] | x[362]);
    assign layer0_out[217] = ~(x[67] | x[79]);
    assign layer0_out[218] = ~x[53];
    assign layer0_out[219] = ~x[29];
    assign layer0_out[220] = ~x[338] | x[340];
    assign layer0_out[221] = ~x[146];
    assign layer0_out[222] = x[36] ^ x[46];
    assign layer0_out[223] = x[60] ^ x[72];
    assign layer0_out[224] = x[351];
    assign layer0_out[225] = x[147];
    assign layer0_out[226] = x[151] & ~x[145];
    assign layer0_out[227] = x[288] & ~x[274];
    assign layer0_out[228] = x[37] & ~x[40];
    assign layer0_out[229] = x[8] & ~x[0];
    assign layer0_out[230] = 1'b0;
    assign layer0_out[231] = ~(x[18] | x[36]);
    assign layer0_out[232] = ~x[355];
    assign layer0_out[233] = x[49] & x[65];
    assign layer0_out[234] = x[166] | x[167];
    assign layer0_out[235] = x[82] & ~x[71];
    assign layer0_out[236] = 1'b0;
    assign layer0_out[237] = x[171] & ~x[163];
    assign layer0_out[238] = ~(x[91] ^ x[93]);
    assign layer0_out[239] = ~(x[40] ^ x[59]);
    assign layer0_out[240] = x[335] & x[353];
    assign layer0_out[241] = x[118];
    assign layer0_out[242] = ~x[307] | x[315];
    assign layer0_out[243] = ~x[321];
    assign layer0_out[244] = ~(x[203] | x[220]);
    assign layer0_out[245] = x[89] ^ x[107];
    assign layer0_out[246] = x[393];
    assign layer0_out[247] = 1'b0;
    assign layer0_out[248] = x[100] & ~x[86];
    assign layer0_out[249] = ~x[153];
    assign layer0_out[250] = x[52] & ~x[61];
    assign layer0_out[251] = x[193] & ~x[180];
    assign layer0_out[252] = x[372];
    assign layer0_out[253] = x[34] ^ x[54];
    assign layer0_out[254] = ~(x[199] ^ x[215]);
    assign layer0_out[255] = ~x[259];
    assign layer0_out[256] = ~(x[50] | x[60]);
    assign layer0_out[257] = ~(x[302] ^ x[313]);
    assign layer0_out[258] = ~x[377];
    assign layer0_out[259] = 1'b1;
    assign layer0_out[260] = ~(x[37] & x[47]);
    assign layer0_out[261] = ~x[252];
    assign layer0_out[262] = ~x[96];
    assign layer0_out[263] = x[55];
    assign layer0_out[264] = ~x[325];
    assign layer0_out[265] = 1'b0;
    assign layer0_out[266] = x[226] | x[228];
    assign layer0_out[267] = x[269];
    assign layer0_out[268] = ~(x[183] ^ x[196]);
    assign layer0_out[269] = ~(x[204] | x[215]);
    assign layer0_out[270] = ~x[198] | x[201];
    assign layer0_out[271] = x[112];
    assign layer0_out[272] = ~(x[349] | x[351]);
    assign layer0_out[273] = x[334] | x[353];
    assign layer0_out[274] = ~x[127] | x[108];
    assign layer0_out[275] = ~x[30];
    assign layer0_out[276] = ~x[365];
    assign layer0_out[277] = x[253] ^ x[268];
    assign layer0_out[278] = ~x[148];
    assign layer0_out[279] = x[194] & ~x[182];
    assign layer0_out[280] = x[275] | x[279];
    assign layer0_out[281] = 1'b0;
    assign layer0_out[282] = ~x[70];
    assign layer0_out[283] = ~(x[302] & x[312]);
    assign layer0_out[284] = ~(x[150] | x[162]);
    assign layer0_out[285] = x[97] | x[111];
    assign layer0_out[286] = ~(x[38] | x[56]);
    assign layer0_out[287] = ~x[37] | x[53];
    assign layer0_out[288] = ~(x[103] | x[123]);
    assign layer0_out[289] = 1'b0;
    assign layer0_out[290] = x[80];
    assign layer0_out[291] = x[132] | x[153];
    assign layer0_out[292] = ~(x[135] | x[151]);
    assign layer0_out[293] = x[98];
    assign layer0_out[294] = x[143] & ~x[162];
    assign layer0_out[295] = 1'b0;
    assign layer0_out[296] = ~x[320];
    assign layer0_out[297] = x[267] & ~x[255];
    assign layer0_out[298] = ~x[167] | x[154];
    assign layer0_out[299] = ~(x[52] & x[56]);
    assign layer0_out[300] = x[213];
    assign layer0_out[301] = ~x[52];
    assign layer0_out[302] = 1'b0;
    assign layer0_out[303] = x[87] | x[104];
    assign layer0_out[304] = ~x[281];
    assign layer0_out[305] = x[88] | x[98];
    assign layer0_out[306] = ~x[83];
    assign layer0_out[307] = x[96] & x[97];
    assign layer0_out[308] = x[229];
    assign layer0_out[309] = x[230] | x[244];
    assign layer0_out[310] = x[153];
    assign layer0_out[311] = ~x[187];
    assign layer0_out[312] = ~(x[233] ^ x[237]);
    assign layer0_out[313] = ~x[354];
    assign layer0_out[314] = ~x[16];
    assign layer0_out[315] = ~x[10] | x[13];
    assign layer0_out[316] = x[199] ^ x[204];
    assign layer0_out[317] = x[54];
    assign layer0_out[318] = ~(x[352] & x[369]);
    assign layer0_out[319] = ~(x[38] | x[55]);
    assign layer0_out[320] = x[76];
    assign layer0_out[321] = x[228] & x[240];
    assign layer0_out[322] = ~x[52] | x[31];
    assign layer0_out[323] = x[113] & x[119];
    assign layer0_out[324] = ~(x[67] | x[69]);
    assign layer0_out[325] = x[319];
    assign layer0_out[326] = ~(x[77] & x[89]);
    assign layer0_out[327] = ~(x[381] | x[397]);
    assign layer0_out[328] = x[84];
    assign layer0_out[329] = ~x[369];
    assign layer0_out[330] = x[166] & ~x[174];
    assign layer0_out[331] = ~(x[188] | x[201]);
    assign layer0_out[332] = ~(x[109] & x[130]);
    assign layer0_out[333] = ~(x[248] ^ x[263]);
    assign layer0_out[334] = ~(x[71] | x[79]);
    assign layer0_out[335] = x[289];
    assign layer0_out[336] = x[74];
    assign layer0_out[337] = x[69];
    assign layer0_out[338] = x[372] | x[392];
    assign layer0_out[339] = ~(x[267] | x[285]);
    assign layer0_out[340] = x[103];
    assign layer0_out[341] = ~x[267];
    assign layer0_out[342] = x[339];
    assign layer0_out[343] = x[125] & ~x[139];
    assign layer0_out[344] = ~x[334] | x[339];
    assign layer0_out[345] = ~x[231] | x[218];
    assign layer0_out[346] = x[10] | x[29];
    assign layer0_out[347] = x[157];
    assign layer0_out[348] = x[28];
    assign layer0_out[349] = x[62] & ~x[80];
    assign layer0_out[350] = ~(x[356] ^ x[361]);
    assign layer0_out[351] = x[39] & x[56];
    assign layer0_out[352] = x[108] & x[111];
    assign layer0_out[353] = 1'b0;
    assign layer0_out[354] = x[300] | x[317];
    assign layer0_out[355] = ~x[221];
    assign layer0_out[356] = ~(x[57] | x[58]);
    assign layer0_out[357] = 1'b0;
    assign layer0_out[358] = x[150] & ~x[169];
    assign layer0_out[359] = x[329] & ~x[309];
    assign layer0_out[360] = x[360] & ~x[354];
    assign layer0_out[361] = ~(x[122] | x[140]);
    assign layer0_out[362] = ~x[301];
    assign layer0_out[363] = ~(x[328] | x[336]);
    assign layer0_out[364] = x[150];
    assign layer0_out[365] = ~x[84] | x[100];
    assign layer0_out[366] = ~(x[30] & x[34]);
    assign layer0_out[367] = x[138] | x[140];
    assign layer0_out[368] = ~x[213];
    assign layer0_out[369] = ~x[294];
    assign layer0_out[370] = ~x[354] | x[340];
    assign layer0_out[371] = ~(x[162] ^ x[181]);
    assign layer0_out[372] = ~x[56] | x[64];
    assign layer0_out[373] = x[379];
    assign layer0_out[374] = x[30];
    assign layer0_out[375] = ~x[211];
    assign layer0_out[376] = x[335];
    assign layer0_out[377] = x[49] & ~x[55];
    assign layer0_out[378] = x[68];
    assign layer0_out[379] = x[114] | x[118];
    assign layer0_out[380] = ~(x[120] | x[137]);
    assign layer0_out[381] = x[245] & ~x[260];
    assign layer0_out[382] = x[337];
    assign layer0_out[383] = x[42] & ~x[62];
    assign layer0_out[384] = ~(x[154] | x[155]);
    assign layer0_out[385] = x[294] ^ x[303];
    assign layer0_out[386] = ~(x[362] ^ x[373]);
    assign layer0_out[387] = ~x[137];
    assign layer0_out[388] = ~x[151] | x[143];
    assign layer0_out[389] = x[241] | x[261];
    assign layer0_out[390] = x[32] & ~x[13];
    assign layer0_out[391] = x[279] | x[282];
    assign layer0_out[392] = x[302];
    assign layer0_out[393] = x[320];
    assign layer0_out[394] = x[94] | x[95];
    assign layer0_out[395] = ~x[344];
    assign layer0_out[396] = x[202];
    assign layer0_out[397] = x[384] & ~x[366];
    assign layer0_out[398] = x[311] ^ x[315];
    assign layer0_out[399] = ~x[99];
    assign layer0_out[400] = ~(x[382] | x[393]);
    assign layer0_out[401] = 1'b0;
    assign layer0_out[402] = x[101] & ~x[81];
    assign layer0_out[403] = ~(x[252] | x[258]);
    assign layer0_out[404] = x[353] | x[370];
    assign layer0_out[405] = ~(x[336] | x[352]);
    assign layer0_out[406] = x[330] & ~x[311];
    assign layer0_out[407] = ~(x[98] | x[114]);
    assign layer0_out[408] = x[256] ^ x[266];
    assign layer0_out[409] = ~x[94] | x[101];
    assign layer0_out[410] = x[34] ^ x[39];
    assign layer0_out[411] = ~(x[268] ^ x[286]);
    assign layer0_out[412] = x[197];
    assign layer0_out[413] = ~x[22];
    assign layer0_out[414] = x[78] & ~x[92];
    assign layer0_out[415] = x[109];
    assign layer0_out[416] = x[353] | x[365];
    assign layer0_out[417] = 1'b1;
    assign layer0_out[418] = ~x[168];
    assign layer0_out[419] = x[186] & x[191];
    assign layer0_out[420] = ~x[383] | x[387];
    assign layer0_out[421] = x[319] | x[337];
    assign layer0_out[422] = x[173] & ~x[160];
    assign layer0_out[423] = x[199];
    assign layer0_out[424] = x[390] & ~x[384];
    assign layer0_out[425] = ~(x[176] ^ x[189]);
    assign layer0_out[426] = x[270];
    assign layer0_out[427] = ~x[304];
    assign layer0_out[428] = 1'b1;
    assign layer0_out[429] = ~(x[213] | x[233]);
    assign layer0_out[430] = ~x[190];
    assign layer0_out[431] = ~x[129] | x[131];
    assign layer0_out[432] = ~(x[285] | x[302]);
    assign layer0_out[433] = ~x[365];
    assign layer0_out[434] = x[99] & ~x[89];
    assign layer0_out[435] = x[177];
    assign layer0_out[436] = x[165];
    assign layer0_out[437] = 1'b1;
    assign layer0_out[438] = x[291];
    assign layer0_out[439] = x[253];
    assign layer0_out[440] = ~(x[277] | x[292]);
    assign layer0_out[441] = ~x[260] | x[261];
    assign layer0_out[442] = x[8] | x[22];
    assign layer0_out[443] = ~(x[361] & x[373]);
    assign layer0_out[444] = ~x[374];
    assign layer0_out[445] = ~x[65];
    assign layer0_out[446] = x[27] & ~x[18];
    assign layer0_out[447] = x[76] | x[79];
    assign layer0_out[448] = ~x[74];
    assign layer0_out[449] = x[222] | x[233];
    assign layer0_out[450] = 1'b0;
    assign layer0_out[451] = x[383] | x[391];
    assign layer0_out[452] = ~x[125] | x[135];
    assign layer0_out[453] = ~(x[128] ^ x[131]);
    assign layer0_out[454] = x[83] | x[86];
    assign layer0_out[455] = x[187] ^ x[193];
    assign layer0_out[456] = x[337] | x[338];
    assign layer0_out[457] = ~x[265];
    assign layer0_out[458] = ~(x[368] | x[387]);
    assign layer0_out[459] = ~x[11];
    assign layer0_out[460] = x[341];
    assign layer0_out[461] = x[8];
    assign layer0_out[462] = 1'b0;
    assign layer0_out[463] = ~x[388];
    assign layer0_out[464] = x[170] | x[189];
    assign layer0_out[465] = 1'b0;
    assign layer0_out[466] = 1'b0;
    assign layer0_out[467] = x[108] ^ x[125];
    assign layer0_out[468] = ~(x[348] | x[366]);
    assign layer0_out[469] = x[363] & x[375];
    assign layer0_out[470] = ~x[150];
    assign layer0_out[471] = x[133] & ~x[118];
    assign layer0_out[472] = ~(x[318] ^ x[330]);
    assign layer0_out[473] = ~x[386];
    assign layer0_out[474] = ~(x[366] & x[370]);
    assign layer0_out[475] = ~(x[334] & x[341]);
    assign layer0_out[476] = x[160];
    assign layer0_out[477] = x[312] | x[313];
    assign layer0_out[478] = x[339];
    assign layer0_out[479] = x[80];
    assign layer0_out[480] = x[20] | x[23];
    assign layer0_out[481] = ~(x[45] | x[53]);
    assign layer0_out[482] = x[79] | x[97];
    assign layer0_out[483] = ~x[243] | x[234];
    assign layer0_out[484] = ~x[353];
    assign layer0_out[485] = x[269] & ~x[274];
    assign layer0_out[486] = x[24] | x[33];
    assign layer0_out[487] = x[180];
    assign layer0_out[488] = x[394] & ~x[382];
    assign layer0_out[489] = 1'b1;
    assign layer0_out[490] = x[102] | x[122];
    assign layer0_out[491] = ~x[260] | x[257];
    assign layer0_out[492] = ~x[359];
    assign layer0_out[493] = x[111] & ~x[117];
    assign layer0_out[494] = ~x[306] | x[325];
    assign layer0_out[495] = ~x[101] | x[83];
    assign layer0_out[496] = ~x[205] | x[215];
    assign layer0_out[497] = ~(x[252] & x[257]);
    assign layer0_out[498] = ~(x[236] | x[251]);
    assign layer0_out[499] = x[181];
    assign layer0_out[500] = 1'b0;
    assign layer0_out[501] = x[383] & ~x[394];
    assign layer0_out[502] = x[325] | x[336];
    assign layer0_out[503] = ~(x[167] | x[188]);
    assign layer0_out[504] = x[246];
    assign layer0_out[505] = ~x[109] | x[125];
    assign layer0_out[506] = ~x[203];
    assign layer0_out[507] = ~x[118];
    assign layer0_out[508] = x[209] & ~x[213];
    assign layer0_out[509] = ~x[254];
    assign layer0_out[510] = x[386];
    assign layer0_out[511] = x[228] & x[242];
    assign layer0_out[512] = ~x[336] | x[346];
    assign layer0_out[513] = ~(x[255] | x[261]);
    assign layer0_out[514] = x[346];
    assign layer0_out[515] = 1'b1;
    assign layer0_out[516] = x[81] | x[83];
    assign layer0_out[517] = x[277] | x[280];
    assign layer0_out[518] = ~(x[41] | x[55]);
    assign layer0_out[519] = ~x[258];
    assign layer0_out[520] = ~(x[5] | x[24]);
    assign layer0_out[521] = ~(x[201] ^ x[204]);
    assign layer0_out[522] = x[346];
    assign layer0_out[523] = ~x[131];
    assign layer0_out[524] = 1'b0;
    assign layer0_out[525] = ~x[72] | x[55];
    assign layer0_out[526] = x[214] & ~x[230];
    assign layer0_out[527] = ~x[214];
    assign layer0_out[528] = ~(x[160] | x[166]);
    assign layer0_out[529] = ~x[246] | x[260];
    assign layer0_out[530] = ~x[246];
    assign layer0_out[531] = x[165] | x[175];
    assign layer0_out[532] = x[224];
    assign layer0_out[533] = x[268];
    assign layer0_out[534] = x[241] ^ x[254];
    assign layer0_out[535] = x[53];
    assign layer0_out[536] = ~(x[291] | x[302]);
    assign layer0_out[537] = ~x[269] | x[263];
    assign layer0_out[538] = x[239];
    assign layer0_out[539] = x[225] & ~x[229];
    assign layer0_out[540] = x[220] ^ x[224];
    assign layer0_out[541] = 1'b1;
    assign layer0_out[542] = x[267] | x[280];
    assign layer0_out[543] = ~(x[45] & x[48]);
    assign layer0_out[544] = x[222] | x[223];
    assign layer0_out[545] = ~(x[155] | x[172]);
    assign layer0_out[546] = ~x[314];
    assign layer0_out[547] = x[240] | x[256];
    assign layer0_out[548] = x[124] & ~x[110];
    assign layer0_out[549] = x[364] | x[383];
    assign layer0_out[550] = ~x[100] | x[120];
    assign layer0_out[551] = ~x[162];
    assign layer0_out[552] = x[361] | x[372];
    assign layer0_out[553] = x[45] ^ x[63];
    assign layer0_out[554] = x[64];
    assign layer0_out[555] = ~(x[31] & x[37]);
    assign layer0_out[556] = x[48] | x[67];
    assign layer0_out[557] = ~x[289] | x[308];
    assign layer0_out[558] = ~x[227];
    assign layer0_out[559] = ~(x[120] | x[128]);
    assign layer0_out[560] = 1'b1;
    assign layer0_out[561] = x[267] | x[269];
    assign layer0_out[562] = x[291];
    assign layer0_out[563] = x[91];
    assign layer0_out[564] = x[387] | x[388];
    assign layer0_out[565] = x[203] | x[221];
    assign layer0_out[566] = x[116];
    assign layer0_out[567] = x[231] & ~x[251];
    assign layer0_out[568] = 1'b1;
    assign layer0_out[569] = x[101] | x[108];
    assign layer0_out[570] = x[216];
    assign layer0_out[571] = x[189] & x[192];
    assign layer0_out[572] = x[124] ^ x[140];
    assign layer0_out[573] = ~x[72] | x[83];
    assign layer0_out[574] = ~(x[91] ^ x[95]);
    assign layer0_out[575] = 1'b1;
    assign layer0_out[576] = x[198];
    assign layer0_out[577] = x[325] | x[327];
    assign layer0_out[578] = x[32] | x[41];
    assign layer0_out[579] = ~x[241] | x[225];
    assign layer0_out[580] = ~x[324] | x[344];
    assign layer0_out[581] = ~x[190];
    assign layer0_out[582] = x[381];
    assign layer0_out[583] = x[105] | x[124];
    assign layer0_out[584] = x[40] | x[44];
    assign layer0_out[585] = ~(x[100] ^ x[116]);
    assign layer0_out[586] = x[241];
    assign layer0_out[587] = x[76] | x[96];
    assign layer0_out[588] = ~(x[321] ^ x[329]);
    assign layer0_out[589] = x[302] | x[303];
    assign layer0_out[590] = ~x[91];
    assign layer0_out[591] = ~x[33];
    assign layer0_out[592] = ~x[248];
    assign layer0_out[593] = ~(x[387] | x[393]);
    assign layer0_out[594] = ~(x[80] & x[92]);
    assign layer0_out[595] = ~(x[213] | x[222]);
    assign layer0_out[596] = 1'b1;
    assign layer0_out[597] = x[16];
    assign layer0_out[598] = ~(x[165] ^ x[170]);
    assign layer0_out[599] = x[137];
    assign layer0_out[600] = ~x[26];
    assign layer0_out[601] = x[121];
    assign layer0_out[602] = x[175] | x[192];
    assign layer0_out[603] = x[271] | x[275];
    assign layer0_out[604] = x[165];
    assign layer0_out[605] = x[120] | x[122];
    assign layer0_out[606] = x[254] | x[264];
    assign layer0_out[607] = 1'b0;
    assign layer0_out[608] = ~(x[124] | x[144]);
    assign layer0_out[609] = ~x[195] | x[196];
    assign layer0_out[610] = x[135] | x[136];
    assign layer0_out[611] = ~x[221];
    assign layer0_out[612] = x[211] & x[223];
    assign layer0_out[613] = ~x[300];
    assign layer0_out[614] = x[206];
    assign layer0_out[615] = x[220] | x[233];
    assign layer0_out[616] = x[176] & ~x[160];
    assign layer0_out[617] = ~(x[294] | x[307]);
    assign layer0_out[618] = ~(x[256] & x[274]);
    assign layer0_out[619] = x[211];
    assign layer0_out[620] = x[28] | x[33];
    assign layer0_out[621] = ~x[283];
    assign layer0_out[622] = ~(x[226] ^ x[242]);
    assign layer0_out[623] = x[396];
    assign layer0_out[624] = x[3] | x[11];
    assign layer0_out[625] = ~(x[109] | x[129]);
    assign layer0_out[626] = ~(x[23] | x[29]);
    assign layer0_out[627] = x[179];
    assign layer0_out[628] = ~(x[343] | x[351]);
    assign layer0_out[629] = ~(x[359] & x[365]);
    assign layer0_out[630] = x[257];
    assign layer0_out[631] = ~(x[32] | x[44]);
    assign layer0_out[632] = ~x[192] | x[179];
    assign layer0_out[633] = x[244];
    assign layer0_out[634] = ~x[248] | x[251];
    assign layer0_out[635] = ~(x[261] | x[269]);
    assign layer0_out[636] = ~(x[197] & x[213]);
    assign layer0_out[637] = x[2] ^ x[9];
    assign layer0_out[638] = ~x[75] | x[65];
    assign layer0_out[639] = x[324] & x[339];
    assign layer0_out[640] = ~x[341];
    assign layer0_out[641] = ~(x[225] | x[245]);
    assign layer0_out[642] = 1'b0;
    assign layer0_out[643] = x[132] & ~x[126];
    assign layer0_out[644] = ~(x[354] & x[363]);
    assign layer0_out[645] = x[44] | x[56];
    assign layer0_out[646] = x[4] & x[25];
    assign layer0_out[647] = x[147] ^ x[163];
    assign layer0_out[648] = x[253] & x[270];
    assign layer0_out[649] = ~(x[107] | x[108]);
    assign layer0_out[650] = ~(x[6] & x[23]);
    assign layer0_out[651] = ~x[298];
    assign layer0_out[652] = x[59] | x[63];
    assign layer0_out[653] = ~(x[112] ^ x[130]);
    assign layer0_out[654] = 1'b0;
    assign layer0_out[655] = x[352] & ~x[363];
    assign layer0_out[656] = ~x[91];
    assign layer0_out[657] = ~x[268];
    assign layer0_out[658] = ~(x[357] & x[365]);
    assign layer0_out[659] = ~x[224] | x[208];
    assign layer0_out[660] = ~(x[352] | x[355]);
    assign layer0_out[661] = x[22] | x[30];
    assign layer0_out[662] = ~x[374];
    assign layer0_out[663] = ~(x[141] | x[142]);
    assign layer0_out[664] = ~x[188] | x[191];
    assign layer0_out[665] = ~x[96];
    assign layer0_out[666] = ~x[175];
    assign layer0_out[667] = x[31] | x[38];
    assign layer0_out[668] = x[279] & ~x[259];
    assign layer0_out[669] = ~x[59] | x[54];
    assign layer0_out[670] = x[25] | x[39];
    assign layer0_out[671] = ~(x[85] | x[105]);
    assign layer0_out[672] = x[140];
    assign layer0_out[673] = x[78] & ~x[61];
    assign layer0_out[674] = x[202] & x[218];
    assign layer0_out[675] = ~(x[28] & x[35]);
    assign layer0_out[676] = x[102] | x[119];
    assign layer0_out[677] = ~x[260];
    assign layer0_out[678] = x[8];
    assign layer0_out[679] = ~(x[55] & x[71]);
    assign layer0_out[680] = ~x[108];
    assign layer0_out[681] = ~(x[207] ^ x[225]);
    assign layer0_out[682] = ~x[132];
    assign layer0_out[683] = x[379];
    assign layer0_out[684] = ~x[176] | x[186];
    assign layer0_out[685] = x[139] ^ x[152];
    assign layer0_out[686] = 1'b1;
    assign layer0_out[687] = x[118];
    assign layer0_out[688] = ~x[290];
    assign layer0_out[689] = x[204];
    assign layer0_out[690] = x[225] & ~x[217];
    assign layer0_out[691] = ~x[387];
    assign layer0_out[692] = x[147];
    assign layer0_out[693] = 1'b1;
    assign layer0_out[694] = ~(x[124] | x[145]);
    assign layer0_out[695] = x[126] | x[128];
    assign layer0_out[696] = x[18] & x[37];
    assign layer0_out[697] = x[147] | x[165];
    assign layer0_out[698] = 1'b0;
    assign layer0_out[699] = x[329] & x[345];
    assign layer0_out[700] = ~x[174];
    assign layer0_out[701] = ~(x[20] | x[24]);
    assign layer0_out[702] = ~x[268] | x[259];
    assign layer0_out[703] = x[305] | x[313];
    assign layer0_out[704] = ~x[254];
    assign layer0_out[705] = x[230];
    assign layer0_out[706] = x[369];
    assign layer0_out[707] = x[324] & x[328];
    assign layer0_out[708] = x[55] & x[70];
    assign layer0_out[709] = ~x[82] | x[92];
    assign layer0_out[710] = x[87] ^ x[105];
    assign layer0_out[711] = ~(x[299] | x[317]);
    assign layer0_out[712] = ~(x[25] | x[44]);
    assign layer0_out[713] = ~x[57];
    assign layer0_out[714] = x[145] | x[162];
    assign layer0_out[715] = x[337] & ~x[333];
    assign layer0_out[716] = ~(x[218] | x[238]);
    assign layer0_out[717] = x[311] & ~x[291];
    assign layer0_out[718] = x[163] & ~x[149];
    assign layer0_out[719] = x[159];
    assign layer0_out[720] = ~x[138];
    assign layer0_out[721] = 1'b1;
    assign layer0_out[722] = ~x[353];
    assign layer0_out[723] = x[183];
    assign layer0_out[724] = ~(x[381] | x[398]);
    assign layer0_out[725] = ~(x[305] | x[315]);
    assign layer0_out[726] = x[125] | x[146];
    assign layer0_out[727] = x[251] & ~x[270];
    assign layer0_out[728] = ~(x[361] | x[379]);
    assign layer0_out[729] = ~(x[109] ^ x[114]);
    assign layer0_out[730] = x[313] | x[323];
    assign layer0_out[731] = ~(x[80] | x[96]);
    assign layer0_out[732] = x[38];
    assign layer0_out[733] = x[306] & ~x[319];
    assign layer0_out[734] = ~x[109] | x[101];
    assign layer0_out[735] = x[181] ^ x[195];
    assign layer0_out[736] = x[296] ^ x[312];
    assign layer0_out[737] = ~x[86] | x[95];
    assign layer0_out[738] = ~(x[224] & x[229]);
    assign layer0_out[739] = x[334] & ~x[337];
    assign layer0_out[740] = x[159] | x[173];
    assign layer0_out[741] = x[128] & x[132];
    assign layer0_out[742] = x[214];
    assign layer0_out[743] = x[151] ^ x[154];
    assign layer0_out[744] = 1'b0;
    assign layer0_out[745] = ~x[120];
    assign layer0_out[746] = 1'b0;
    assign layer0_out[747] = ~(x[301] & x[310]);
    assign layer0_out[748] = x[119] ^ x[121];
    assign layer0_out[749] = ~x[168];
    assign layer0_out[750] = x[161] ^ x[176];
    assign layer0_out[751] = x[5] & ~x[25];
    assign layer0_out[752] = ~(x[210] | x[227]);
    assign layer0_out[753] = ~(x[331] | x[338]);
    assign layer0_out[754] = x[55] & x[60];
    assign layer0_out[755] = x[264] | x[275];
    assign layer0_out[756] = ~(x[164] | x[185]);
    assign layer0_out[757] = x[39] & ~x[20];
    assign layer0_out[758] = ~(x[382] & x[397]);
    assign layer0_out[759] = x[146];
    assign layer0_out[760] = ~x[149];
    assign layer0_out[761] = x[7] ^ x[19];
    assign layer0_out[762] = ~x[184];
    assign layer0_out[763] = x[185];
    assign layer0_out[764] = ~x[81] | x[79];
    assign layer0_out[765] = ~x[290] | x[301];
    assign layer0_out[766] = x[65];
    assign layer0_out[767] = x[191] & x[194];
    assign layer0_out[768] = x[306];
    assign layer0_out[769] = 1'b1;
    assign layer0_out[770] = ~x[82] | x[100];
    assign layer0_out[771] = x[200] & ~x[189];
    assign layer0_out[772] = x[214] & x[218];
    assign layer0_out[773] = x[162];
    assign layer0_out[774] = ~(x[36] | x[56]);
    assign layer0_out[775] = ~x[321] | x[323];
    assign layer0_out[776] = ~(x[373] | x[382]);
    assign layer0_out[777] = x[47] | x[64];
    assign layer0_out[778] = ~(x[9] | x[12]);
    assign layer0_out[779] = x[257];
    assign layer0_out[780] = x[346] | x[364];
    assign layer0_out[781] = x[155] ^ x[157];
    assign layer0_out[782] = ~x[296];
    assign layer0_out[783] = ~x[251];
    assign layer0_out[784] = ~x[274];
    assign layer0_out[785] = ~(x[395] | x[398]);
    assign layer0_out[786] = x[289] | x[305];
    assign layer0_out[787] = x[79] & x[83];
    assign layer0_out[788] = ~(x[187] ^ x[201]);
    assign layer0_out[789] = x[331];
    assign layer0_out[790] = x[304] & ~x[299];
    assign layer0_out[791] = x[353] & ~x[359];
    assign layer0_out[792] = x[310] ^ x[321];
    assign layer0_out[793] = ~x[272];
    assign layer0_out[794] = ~x[108];
    assign layer0_out[795] = ~x[211] | x[199];
    assign layer0_out[796] = ~x[64];
    assign layer0_out[797] = ~(x[83] & x[90]);
    assign layer0_out[798] = 1'b1;
    assign layer0_out[799] = ~x[234];
    assign layer0_out[800] = ~x[47];
    assign layer0_out[801] = ~(x[155] | x[166]);
    assign layer0_out[802] = x[91];
    assign layer0_out[803] = ~x[171] | x[161];
    assign layer0_out[804] = x[320];
    assign layer0_out[805] = 1'b1;
    assign layer0_out[806] = 1'b1;
    assign layer0_out[807] = x[198] ^ x[218];
    assign layer0_out[808] = x[215];
    assign layer0_out[809] = ~(x[181] | x[193]);
    assign layer0_out[810] = x[140] | x[141];
    assign layer0_out[811] = ~(x[249] ^ x[251]);
    assign layer0_out[812] = x[190] & ~x[203];
    assign layer0_out[813] = x[48] & ~x[43];
    assign layer0_out[814] = ~x[332];
    assign layer0_out[815] = ~x[187] | x[177];
    assign layer0_out[816] = x[344] & x[354];
    assign layer0_out[817] = x[242];
    assign layer0_out[818] = x[88] & ~x[97];
    assign layer0_out[819] = x[1] | x[22];
    assign layer0_out[820] = x[331];
    assign layer0_out[821] = x[54] ^ x[64];
    assign layer0_out[822] = x[65];
    assign layer0_out[823] = ~(x[282] | x[285]);
    assign layer0_out[824] = ~x[250] | x[237];
    assign layer0_out[825] = x[306] & ~x[310];
    assign layer0_out[826] = ~(x[206] ^ x[210]);
    assign layer0_out[827] = 1'b0;
    assign layer0_out[828] = x[280] | x[285];
    assign layer0_out[829] = ~x[391];
    assign layer0_out[830] = x[321] | x[341];
    assign layer0_out[831] = ~x[144];
    assign layer0_out[832] = x[390] | x[392];
    assign layer0_out[833] = ~x[50] | x[63];
    assign layer0_out[834] = x[135];
    assign layer0_out[835] = x[138];
    assign layer0_out[836] = x[179] & ~x[161];
    assign layer0_out[837] = x[268];
    assign layer0_out[838] = ~x[212];
    assign layer0_out[839] = x[70] & x[72];
    assign layer0_out[840] = x[329] | x[349];
    assign layer0_out[841] = ~(x[121] & x[133]);
    assign layer0_out[842] = ~x[4];
    assign layer0_out[843] = ~(x[379] | x[381]);
    assign layer0_out[844] = ~x[142] | x[135];
    assign layer0_out[845] = ~(x[172] & x[187]);
    assign layer0_out[846] = x[313] ^ x[318];
    assign layer0_out[847] = x[290] & x[309];
    assign layer0_out[848] = ~x[141];
    assign layer0_out[849] = ~(x[375] ^ x[394]);
    assign layer0_out[850] = x[149];
    assign layer0_out[851] = x[208];
    assign layer0_out[852] = x[67] & x[82];
    assign layer0_out[853] = x[130];
    assign layer0_out[854] = x[72] & ~x[58];
    assign layer0_out[855] = ~(x[358] | x[374]);
    assign layer0_out[856] = ~x[201] | x[206];
    assign layer0_out[857] = x[304] | x[305];
    assign layer0_out[858] = x[63] | x[84];
    assign layer0_out[859] = ~(x[100] | x[103]);
    assign layer0_out[860] = x[104];
    assign layer0_out[861] = ~x[253];
    assign layer0_out[862] = ~x[122];
    assign layer0_out[863] = ~x[371];
    assign layer0_out[864] = x[327] ^ x[345];
    assign layer0_out[865] = ~x[127];
    assign layer0_out[866] = ~(x[189] | x[191]);
    assign layer0_out[867] = ~x[159] | x[139];
    assign layer0_out[868] = x[60] & x[77];
    assign layer0_out[869] = x[362] & ~x[343];
    assign layer0_out[870] = x[24] | x[25];
    assign layer0_out[871] = ~x[374] | x[355];
    assign layer0_out[872] = ~(x[144] | x[146]);
    assign layer0_out[873] = ~x[88];
    assign layer0_out[874] = ~x[214];
    assign layer0_out[875] = x[134] & ~x[115];
    assign layer0_out[876] = ~x[207];
    assign layer0_out[877] = ~x[274] | x[286];
    assign layer0_out[878] = ~x[108];
    assign layer0_out[879] = x[56] ^ x[71];
    assign layer0_out[880] = 1'b0;
    assign layer0_out[881] = 1'b0;
    assign layer0_out[882] = x[342] & ~x[354];
    assign layer0_out[883] = ~x[364];
    assign layer0_out[884] = ~(x[127] | x[129]);
    assign layer0_out[885] = x[10];
    assign layer0_out[886] = ~x[273];
    assign layer0_out[887] = x[347] & ~x[337];
    assign layer0_out[888] = x[237] | x[248];
    assign layer0_out[889] = ~x[255];
    assign layer0_out[890] = x[147];
    assign layer0_out[891] = x[202] | x[205];
    assign layer0_out[892] = x[280] | x[293];
    assign layer0_out[893] = ~x[187] | x[199];
    assign layer0_out[894] = x[342] | x[346];
    assign layer0_out[895] = ~x[231];
    assign layer0_out[896] = ~x[387];
    assign layer0_out[897] = ~x[87];
    assign layer0_out[898] = x[30];
    assign layer0_out[899] = ~(x[265] & x[284]);
    assign layer0_out[900] = x[315] | x[330];
    assign layer0_out[901] = ~(x[243] | x[246]);
    assign layer0_out[902] = ~(x[366] & x[383]);
    assign layer0_out[903] = x[34] ^ x[45];
    assign layer0_out[904] = ~(x[70] & x[83]);
    assign layer0_out[905] = ~x[219] | x[201];
    assign layer0_out[906] = x[321] ^ x[324];
    assign layer0_out[907] = ~x[20] | x[18];
    assign layer0_out[908] = x[93] & ~x[99];
    assign layer0_out[909] = ~x[236] | x[253];
    assign layer0_out[910] = x[345] | x[359];
    assign layer0_out[911] = ~x[207];
    assign layer0_out[912] = ~(x[52] | x[54]);
    assign layer0_out[913] = ~(x[340] | x[351]);
    assign layer0_out[914] = x[240] ^ x[249];
    assign layer0_out[915] = ~x[307] | x[291];
    assign layer0_out[916] = x[224] | x[227];
    assign layer0_out[917] = ~x[36];
    assign layer0_out[918] = ~x[282] | x[267];
    assign layer0_out[919] = ~(x[35] & x[52]);
    assign layer0_out[920] = x[119];
    assign layer0_out[921] = x[148] & ~x[159];
    assign layer0_out[922] = x[10] | x[26];
    assign layer0_out[923] = x[323] ^ x[338];
    assign layer0_out[924] = x[236] | x[243];
    assign layer0_out[925] = ~(x[239] ^ x[255]);
    assign layer0_out[926] = ~x[156];
    assign layer0_out[927] = x[19];
    assign layer0_out[928] = x[158] ^ x[170];
    assign layer0_out[929] = ~x[378] | x[366];
    assign layer0_out[930] = x[367];
    assign layer0_out[931] = ~x[47];
    assign layer0_out[932] = ~x[288];
    assign layer0_out[933] = ~x[51];
    assign layer0_out[934] = ~x[119] | x[138];
    assign layer0_out[935] = x[250];
    assign layer0_out[936] = x[6] ^ x[21];
    assign layer0_out[937] = x[354] | x[355];
    assign layer0_out[938] = ~x[218];
    assign layer0_out[939] = ~(x[123] | x[124]);
    assign layer0_out[940] = ~(x[17] & x[35]);
    assign layer0_out[941] = ~(x[202] | x[214]);
    assign layer0_out[942] = ~x[297] | x[289];
    assign layer0_out[943] = ~x[248];
    assign layer0_out[944] = ~x[341] | x[351];
    assign layer0_out[945] = x[321];
    assign layer0_out[946] = ~x[47];
    assign layer0_out[947] = ~(x[133] ^ x[136]);
    assign layer0_out[948] = x[240];
    assign layer0_out[949] = x[221] | x[232];
    assign layer0_out[950] = ~(x[166] | x[171]);
    assign layer0_out[951] = x[168] & ~x[157];
    assign layer0_out[952] = x[153] ^ x[155];
    assign layer0_out[953] = x[360];
    assign layer0_out[954] = x[116];
    assign layer0_out[955] = ~(x[61] | x[62]);
    assign layer0_out[956] = ~(x[349] | x[352]);
    assign layer0_out[957] = ~x[356];
    assign layer0_out[958] = 1'b1;
    assign layer0_out[959] = x[180] | x[201];
    assign layer0_out[960] = ~(x[46] | x[56]);
    assign layer0_out[961] = x[356];
    assign layer0_out[962] = ~(x[52] ^ x[55]);
    assign layer0_out[963] = x[366] & ~x[379];
    assign layer0_out[964] = ~(x[281] | x[282]);
    assign layer0_out[965] = ~(x[180] | x[200]);
    assign layer0_out[966] = 1'b0;
    assign layer0_out[967] = x[371];
    assign layer0_out[968] = x[78];
    assign layer0_out[969] = x[119] | x[137];
    assign layer0_out[970] = x[275] | x[280];
    assign layer0_out[971] = x[167] & x[180];
    assign layer0_out[972] = x[103];
    assign layer0_out[973] = ~(x[252] | x[270]);
    assign layer0_out[974] = ~(x[83] | x[102]);
    assign layer0_out[975] = x[172] ^ x[177];
    assign layer0_out[976] = ~x[177];
    assign layer0_out[977] = 1'b1;
    assign layer0_out[978] = 1'b1;
    assign layer0_out[979] = x[165] ^ x[180];
    assign layer0_out[980] = ~(x[136] | x[155]);
    assign layer0_out[981] = ~(x[92] | x[110]);
    assign layer0_out[982] = ~x[386] | x[377];
    assign layer0_out[983] = ~x[29];
    assign layer0_out[984] = ~(x[192] | x[201]);
    assign layer0_out[985] = ~(x[312] | x[323]);
    assign layer0_out[986] = ~x[42] | x[37];
    assign layer0_out[987] = x[124] | x[138];
    assign layer0_out[988] = x[172] & ~x[167];
    assign layer0_out[989] = ~(x[10] | x[31]);
    assign layer0_out[990] = ~(x[307] | x[324]);
    assign layer0_out[991] = ~(x[115] ^ x[130]);
    assign layer0_out[992] = ~x[26] | x[29];
    assign layer0_out[993] = ~(x[349] | x[359]);
    assign layer0_out[994] = x[170];
    assign layer0_out[995] = x[273] & ~x[270];
    assign layer0_out[996] = x[335] & ~x[320];
    assign layer0_out[997] = ~x[334] | x[345];
    assign layer0_out[998] = x[34] & ~x[20];
    assign layer0_out[999] = x[136] | x[157];
    assign layer0_out[1000] = ~(x[222] | x[227]);
    assign layer0_out[1001] = ~(x[260] | x[271]);
    assign layer0_out[1002] = x[313] & x[327];
    assign layer0_out[1003] = x[115];
    assign layer0_out[1004] = ~x[137];
    assign layer0_out[1005] = x[375];
    assign layer0_out[1006] = x[250];
    assign layer0_out[1007] = x[364] & ~x[374];
    assign layer0_out[1008] = ~(x[163] | x[166]);
    assign layer0_out[1009] = ~x[228];
    assign layer0_out[1010] = x[146] & ~x[152];
    assign layer0_out[1011] = ~x[130];
    assign layer0_out[1012] = ~(x[135] | x[146]);
    assign layer0_out[1013] = ~x[360];
    assign layer0_out[1014] = x[72] ^ x[87];
    assign layer0_out[1015] = x[330];
    assign layer0_out[1016] = ~(x[111] ^ x[114]);
    assign layer0_out[1017] = x[122] | x[142];
    assign layer0_out[1018] = x[346] & x[356];
    assign layer0_out[1019] = ~x[9] | x[21];
    assign layer0_out[1020] = x[90] & ~x[104];
    assign layer0_out[1021] = ~(x[60] & x[78]);
    assign layer0_out[1022] = x[190] & x[191];
    assign layer0_out[1023] = ~x[268];
    assign layer0_out[1024] = x[210] ^ x[223];
    assign layer0_out[1025] = 1'b1;
    assign layer0_out[1026] = ~(x[51] ^ x[67]);
    assign layer0_out[1027] = ~(x[156] | x[162]);
    assign layer0_out[1028] = ~x[293];
    assign layer0_out[1029] = x[370] & x[376];
    assign layer0_out[1030] = x[215] & ~x[206];
    assign layer0_out[1031] = ~(x[19] ^ x[23]);
    assign layer0_out[1032] = 1'b1;
    assign layer0_out[1033] = x[61] & ~x[42];
    assign layer0_out[1034] = ~x[97] | x[84];
    assign layer0_out[1035] = x[29] & ~x[36];
    assign layer0_out[1036] = x[141] & x[145];
    assign layer0_out[1037] = ~(x[301] ^ x[318]);
    assign layer0_out[1038] = ~(x[92] | x[94]);
    assign layer0_out[1039] = ~(x[266] ^ x[270]);
    assign layer0_out[1040] = x[81] ^ x[84];
    assign layer0_out[1041] = x[244];
    assign layer0_out[1042] = ~(x[227] ^ x[231]);
    assign layer0_out[1043] = ~x[281] | x[275];
    assign layer0_out[1044] = ~(x[254] | x[261]);
    assign layer0_out[1045] = ~(x[339] | x[359]);
    assign layer0_out[1046] = x[178] | x[179];
    assign layer0_out[1047] = x[254] | x[263];
    assign layer0_out[1048] = ~x[103];
    assign layer0_out[1049] = x[355] | x[366];
    assign layer0_out[1050] = ~(x[55] & x[67]);
    assign layer0_out[1051] = x[287];
    assign layer0_out[1052] = ~x[220];
    assign layer0_out[1053] = 1'b1;
    assign layer0_out[1054] = 1'b1;
    assign layer0_out[1055] = x[326] | x[337];
    assign layer0_out[1056] = x[10] & ~x[20];
    assign layer0_out[1057] = ~x[90];
    assign layer0_out[1058] = ~x[104];
    assign layer0_out[1059] = ~(x[62] & x[63]);
    assign layer0_out[1060] = 1'b1;
    assign layer0_out[1061] = ~x[343] | x[338];
    assign layer0_out[1062] = ~x[366];
    assign layer0_out[1063] = x[307] | x[309];
    assign layer0_out[1064] = 1'b0;
    assign layer0_out[1065] = ~x[329];
    assign layer0_out[1066] = x[387] & x[397];
    assign layer0_out[1067] = x[94] & x[110];
    assign layer0_out[1068] = ~x[263];
    assign layer0_out[1069] = ~(x[120] | x[140]);
    assign layer0_out[1070] = ~x[375] | x[365];
    assign layer0_out[1071] = x[372];
    assign layer0_out[1072] = ~x[363];
    assign layer0_out[1073] = ~(x[99] ^ x[111]);
    assign layer0_out[1074] = ~x[47] | x[26];
    assign layer0_out[1075] = x[178] ^ x[195];
    assign layer0_out[1076] = ~x[96];
    assign layer0_out[1077] = x[62];
    assign layer0_out[1078] = ~(x[161] | x[178]);
    assign layer0_out[1079] = ~(x[107] | x[115]);
    assign layer0_out[1080] = x[169] & x[183];
    assign layer0_out[1081] = ~x[22];
    assign layer0_out[1082] = x[162];
    assign layer0_out[1083] = x[176] & ~x[172];
    assign layer0_out[1084] = x[306] & ~x[320];
    assign layer0_out[1085] = ~(x[92] | x[113]);
    assign layer0_out[1086] = x[267] ^ x[268];
    assign layer0_out[1087] = x[44] | x[45];
    assign layer0_out[1088] = ~(x[201] ^ x[202]);
    assign layer0_out[1089] = x[147] & ~x[143];
    assign layer0_out[1090] = x[70] & x[81];
    assign layer0_out[1091] = ~(x[118] | x[132]);
    assign layer0_out[1092] = x[139];
    assign layer0_out[1093] = 1'b1;
    assign layer0_out[1094] = ~(x[239] ^ x[254]);
    assign layer0_out[1095] = x[65] & x[72];
    assign layer0_out[1096] = ~(x[25] | x[29]);
    assign layer0_out[1097] = ~(x[2] | x[22]);
    assign layer0_out[1098] = x[158] ^ x[171];
    assign layer0_out[1099] = ~x[204] | x[219];
    assign layer0_out[1100] = ~(x[301] ^ x[304]);
    assign layer0_out[1101] = ~x[203];
    assign layer0_out[1102] = ~(x[319] & x[339]);
    assign layer0_out[1103] = x[189] & ~x[180];
    assign layer0_out[1104] = ~x[231];
    assign layer0_out[1105] = ~x[150];
    assign layer0_out[1106] = ~(x[260] ^ x[272]);
    assign layer0_out[1107] = x[45] & ~x[59];
    assign layer0_out[1108] = x[387];
    assign layer0_out[1109] = ~(x[17] | x[21]);
    assign layer0_out[1110] = 1'b0;
    assign layer0_out[1111] = x[288] | x[305];
    assign layer0_out[1112] = x[255] & x[270];
    assign layer0_out[1113] = 1'b0;
    assign layer0_out[1114] = ~x[215] | x[230];
    assign layer0_out[1115] = ~(x[85] | x[97]);
    assign layer0_out[1116] = x[244] & ~x[227];
    assign layer0_out[1117] = ~x[130];
    assign layer0_out[1118] = x[7] & ~x[2];
    assign layer0_out[1119] = ~(x[170] | x[172]);
    assign layer0_out[1120] = x[128];
    assign layer0_out[1121] = x[255] & ~x[248];
    assign layer0_out[1122] = ~(x[331] | x[351]);
    assign layer0_out[1123] = x[255] ^ x[272];
    assign layer0_out[1124] = ~(x[363] ^ x[383]);
    assign layer0_out[1125] = ~x[255] | x[243];
    assign layer0_out[1126] = ~x[287];
    assign layer0_out[1127] = ~(x[211] | x[230]);
    assign layer0_out[1128] = x[295] | x[313];
    assign layer0_out[1129] = ~x[144];
    assign layer0_out[1130] = x[209];
    assign layer0_out[1131] = x[30] & ~x[27];
    assign layer0_out[1132] = ~(x[51] | x[56]);
    assign layer0_out[1133] = x[33];
    assign layer0_out[1134] = x[278] & ~x[294];
    assign layer0_out[1135] = x[296];
    assign layer0_out[1136] = ~x[211];
    assign layer0_out[1137] = x[26] | x[27];
    assign layer0_out[1138] = ~(x[274] | x[284]);
    assign layer0_out[1139] = ~x[174] | x[192];
    assign layer0_out[1140] = ~x[312];
    assign layer0_out[1141] = x[105];
    assign layer0_out[1142] = ~(x[58] ^ x[64]);
    assign layer0_out[1143] = x[76] | x[84];
    assign layer0_out[1144] = ~x[284] | x[289];
    assign layer0_out[1145] = ~(x[317] | x[324]);
    assign layer0_out[1146] = x[185] & ~x[199];
    assign layer0_out[1147] = x[288] & x[292];
    assign layer0_out[1148] = x[327];
    assign layer0_out[1149] = x[272] ^ x[277];
    assign layer0_out[1150] = x[149] & x[170];
    assign layer0_out[1151] = x[25];
    assign layer0_out[1152] = ~x[296] | x[282];
    assign layer0_out[1153] = ~x[288] | x[280];
    assign layer0_out[1154] = ~x[76];
    assign layer0_out[1155] = ~(x[191] | x[205]);
    assign layer0_out[1156] = ~x[247];
    assign layer0_out[1157] = x[291] & x[294];
    assign layer0_out[1158] = ~(x[184] | x[186]);
    assign layer0_out[1159] = ~x[162] | x[182];
    assign layer0_out[1160] = x[286] & x[302];
    assign layer0_out[1161] = x[363];
    assign layer0_out[1162] = ~x[121] | x[102];
    assign layer0_out[1163] = ~(x[271] | x[278]);
    assign layer0_out[1164] = ~x[206] | x[208];
    assign layer0_out[1165] = ~(x[258] ^ x[277]);
    assign layer0_out[1166] = 1'b1;
    assign layer0_out[1167] = x[110];
    assign layer0_out[1168] = x[25] | x[38];
    assign layer0_out[1169] = x[99] & ~x[87];
    assign layer0_out[1170] = x[155] ^ x[161];
    assign layer0_out[1171] = ~(x[136] | x[150]);
    assign layer0_out[1172] = x[116];
    assign layer0_out[1173] = ~(x[145] | x[161]);
    assign layer0_out[1174] = 1'b0;
    assign layer0_out[1175] = ~x[208];
    assign layer0_out[1176] = ~x[356];
    assign layer0_out[1177] = x[153];
    assign layer0_out[1178] = ~(x[370] | x[390]);
    assign layer0_out[1179] = ~x[301] | x[296];
    assign layer0_out[1180] = x[28] | x[44];
    assign layer0_out[1181] = ~x[142];
    assign layer0_out[1182] = x[387];
    assign layer0_out[1183] = x[297] & ~x[294];
    assign layer0_out[1184] = ~x[81];
    assign layer0_out[1185] = x[373] | x[375];
    assign layer0_out[1186] = ~x[30];
    assign layer0_out[1187] = ~x[361];
    assign layer0_out[1188] = ~(x[184] | x[197]);
    assign layer0_out[1189] = ~(x[374] | x[377]);
    assign layer0_out[1190] = x[102] | x[113];
    assign layer0_out[1191] = x[262] ^ x[275];
    assign layer0_out[1192] = x[157];
    assign layer0_out[1193] = x[127] & ~x[120];
    assign layer0_out[1194] = ~x[336] | x[319];
    assign layer0_out[1195] = 1'b0;
    assign layer0_out[1196] = ~(x[115] | x[118]);
    assign layer0_out[1197] = x[290];
    assign layer0_out[1198] = ~x[76] | x[81];
    assign layer0_out[1199] = ~(x[27] ^ x[48]);
    assign layer0_out[1200] = x[9] | x[16];
    assign layer0_out[1201] = x[189] | x[201];
    assign layer0_out[1202] = ~x[119] | x[101];
    assign layer0_out[1203] = x[228];
    assign layer0_out[1204] = ~(x[44] | x[65]);
    assign layer0_out[1205] = ~(x[290] ^ x[306]);
    assign layer0_out[1206] = x[391] & ~x[380];
    assign layer0_out[1207] = ~(x[286] | x[288]);
    assign layer0_out[1208] = x[293] | x[297];
    assign layer0_out[1209] = ~(x[8] | x[24]);
    assign layer0_out[1210] = x[378];
    assign layer0_out[1211] = x[336] & x[338];
    assign layer0_out[1212] = ~(x[350] ^ x[355]);
    assign layer0_out[1213] = ~x[245];
    assign layer0_out[1214] = ~(x[260] | x[263]);
    assign layer0_out[1215] = x[338] & ~x[345];
    assign layer0_out[1216] = x[187] & ~x[196];
    assign layer0_out[1217] = ~(x[23] | x[43]);
    assign layer0_out[1218] = ~(x[331] ^ x[347]);
    assign layer0_out[1219] = ~x[222];
    assign layer0_out[1220] = ~(x[183] & x[186]);
    assign layer0_out[1221] = x[41] & ~x[62];
    assign layer0_out[1222] = x[375];
    assign layer0_out[1223] = x[289] & x[306];
    assign layer0_out[1224] = ~(x[181] | x[200]);
    assign layer0_out[1225] = ~x[6] | x[17];
    assign layer0_out[1226] = ~x[3] | x[15];
    assign layer0_out[1227] = ~x[85] | x[70];
    assign layer0_out[1228] = x[340] | x[345];
    assign layer0_out[1229] = ~x[200];
    assign layer0_out[1230] = x[170];
    assign layer0_out[1231] = x[286] ^ x[304];
    assign layer0_out[1232] = x[130] & ~x[138];
    assign layer0_out[1233] = ~x[267] | x[270];
    assign layer0_out[1234] = x[123];
    assign layer0_out[1235] = 1'b0;
    assign layer0_out[1236] = x[270] & ~x[282];
    assign layer0_out[1237] = ~x[215];
    assign layer0_out[1238] = x[73];
    assign layer0_out[1239] = ~x[168];
    assign layer0_out[1240] = ~x[300] | x[313];
    assign layer0_out[1241] = x[117] | x[128];
    assign layer0_out[1242] = ~x[18];
    assign layer0_out[1243] = x[172] & ~x[184];
    assign layer0_out[1244] = x[222] ^ x[228];
    assign layer0_out[1245] = ~(x[161] ^ x[174]);
    assign layer0_out[1246] = x[284] & x[295];
    assign layer0_out[1247] = ~x[301];
    assign layer0_out[1248] = ~x[47];
    assign layer0_out[1249] = ~(x[75] | x[93]);
    assign layer0_out[1250] = ~x[307] | x[322];
    assign layer0_out[1251] = x[9] & x[17];
    assign layer0_out[1252] = x[113] | x[114];
    assign layer0_out[1253] = 1'b0;
    assign layer0_out[1254] = x[264];
    assign layer0_out[1255] = ~x[85] | x[69];
    assign layer0_out[1256] = ~(x[355] | x[370]);
    assign layer0_out[1257] = x[102] & ~x[85];
    assign layer0_out[1258] = ~(x[43] | x[58]);
    assign layer0_out[1259] = ~x[247] | x[250];
    assign layer0_out[1260] = ~x[73];
    assign layer0_out[1261] = x[297] ^ x[303];
    assign layer0_out[1262] = ~(x[28] & x[45]);
    assign layer0_out[1263] = ~(x[32] ^ x[52]);
    assign layer0_out[1264] = ~(x[152] | x[154]);
    assign layer0_out[1265] = 1'b0;
    assign layer0_out[1266] = ~x[349] | x[340];
    assign layer0_out[1267] = x[139] ^ x[147];
    assign layer0_out[1268] = ~x[388];
    assign layer0_out[1269] = ~(x[340] | x[353]);
    assign layer0_out[1270] = x[151] ^ x[170];
    assign layer0_out[1271] = x[283];
    assign layer0_out[1272] = x[242] & ~x[259];
    assign layer0_out[1273] = x[112];
    assign layer0_out[1274] = ~(x[93] ^ x[95]);
    assign layer0_out[1275] = x[237] | x[247];
    assign layer0_out[1276] = ~(x[169] & x[182]);
    assign layer0_out[1277] = x[21] | x[25];
    assign layer0_out[1278] = x[344];
    assign layer0_out[1279] = 1'b0;
    assign layer0_out[1280] = x[279];
    assign layer0_out[1281] = x[399] & ~x[393];
    assign layer0_out[1282] = ~x[229] | x[236];
    assign layer0_out[1283] = x[261];
    assign layer0_out[1284] = x[85] | x[99];
    assign layer0_out[1285] = x[130];
    assign layer0_out[1286] = ~x[166];
    assign layer0_out[1287] = ~(x[288] & x[290]);
    assign layer0_out[1288] = ~x[235];
    assign layer0_out[1289] = x[181] & x[201];
    assign layer0_out[1290] = ~x[210];
    assign layer0_out[1291] = x[284] & ~x[299];
    assign layer0_out[1292] = x[230];
    assign layer0_out[1293] = x[328];
    assign layer0_out[1294] = x[1] | x[4];
    assign layer0_out[1295] = ~(x[275] | x[276]);
    assign layer0_out[1296] = x[189];
    assign layer0_out[1297] = ~(x[185] ^ x[189]);
    assign layer0_out[1298] = x[313] & x[317];
    assign layer0_out[1299] = x[27] & ~x[19];
    assign layer0_out[1300] = x[122];
    assign layer0_out[1301] = x[55];
    assign layer0_out[1302] = ~(x[232] | x[250]);
    assign layer0_out[1303] = ~(x[311] | x[313]);
    assign layer0_out[1304] = ~x[228];
    assign layer0_out[1305] = x[28] | x[34];
    assign layer0_out[1306] = ~(x[336] & x[354]);
    assign layer0_out[1307] = ~(x[2] | x[3]);
    assign layer0_out[1308] = 1'b0;
    assign layer0_out[1309] = x[377] ^ x[396];
    assign layer0_out[1310] = x[10];
    assign layer0_out[1311] = x[322] & ~x[340];
    assign layer0_out[1312] = x[373] & ~x[384];
    assign layer0_out[1313] = 1'b0;
    assign layer0_out[1314] = ~(x[144] ^ x[147]);
    assign layer0_out[1315] = ~(x[143] & x[163]);
    assign layer0_out[1316] = x[38] | x[43];
    assign layer0_out[1317] = ~(x[298] | x[316]);
    assign layer0_out[1318] = x[205] | x[207];
    assign layer0_out[1319] = ~x[285];
    assign layer0_out[1320] = ~x[246];
    assign layer0_out[1321] = ~x[178];
    assign layer0_out[1322] = x[215] | x[225];
    assign layer0_out[1323] = x[258];
    assign layer0_out[1324] = ~(x[7] | x[20]);
    assign layer0_out[1325] = x[291] & ~x[305];
    assign layer0_out[1326] = x[158];
    assign layer0_out[1327] = ~x[261] | x[268];
    assign layer0_out[1328] = ~x[167] | x[175];
    assign layer0_out[1329] = ~x[390];
    assign layer0_out[1330] = 1'b1;
    assign layer0_out[1331] = x[132];
    assign layer0_out[1332] = ~(x[380] | x[388]);
    assign layer0_out[1333] = ~(x[190] & x[208]);
    assign layer0_out[1334] = x[180] & ~x[199];
    assign layer0_out[1335] = ~(x[63] | x[82]);
    assign layer0_out[1336] = ~(x[129] ^ x[140]);
    assign layer0_out[1337] = x[164] & ~x[174];
    assign layer0_out[1338] = ~x[323] | x[332];
    assign layer0_out[1339] = x[258] | x[268];
    assign layer0_out[1340] = ~(x[353] ^ x[372]);
    assign layer0_out[1341] = ~(x[165] | x[185]);
    assign layer0_out[1342] = x[36] | x[54];
    assign layer0_out[1343] = x[341];
    assign layer0_out[1344] = x[97] ^ x[114];
    assign layer0_out[1345] = x[350];
    assign layer0_out[1346] = ~(x[13] | x[34]);
    assign layer0_out[1347] = x[58];
    assign layer0_out[1348] = ~x[212];
    assign layer0_out[1349] = ~(x[53] & x[64]);
    assign layer0_out[1350] = ~x[381] | x[370];
    assign layer0_out[1351] = x[221] | x[231];
    assign layer0_out[1352] = x[219] | x[232];
    assign layer0_out[1353] = ~(x[167] | x[186]);
    assign layer0_out[1354] = x[133] & x[149];
    assign layer0_out[1355] = ~(x[183] | x[184]);
    assign layer0_out[1356] = ~x[360] | x[367];
    assign layer0_out[1357] = ~x[54] | x[44];
    assign layer0_out[1358] = x[27];
    assign layer0_out[1359] = x[299] & ~x[292];
    assign layer0_out[1360] = ~x[189] | x[172];
    assign layer0_out[1361] = x[263];
    assign layer0_out[1362] = ~x[113];
    assign layer0_out[1363] = x[78] | x[84];
    assign layer0_out[1364] = ~(x[341] | x[343]);
    assign layer0_out[1365] = ~x[102];
    assign layer0_out[1366] = x[77] & ~x[62];
    assign layer0_out[1367] = 1'b1;
    assign layer0_out[1368] = x[142] | x[146];
    assign layer0_out[1369] = ~x[140] | x[157];
    assign layer0_out[1370] = ~(x[322] | x[336]);
    assign layer0_out[1371] = x[6];
    assign layer0_out[1372] = x[246] & ~x[261];
    assign layer0_out[1373] = ~(x[101] | x[116]);
    assign layer0_out[1374] = x[324];
    assign layer0_out[1375] = x[48] | x[66];
    assign layer0_out[1376] = 1'b1;
    assign layer0_out[1377] = ~x[98];
    assign layer0_out[1378] = ~x[323];
    assign layer0_out[1379] = 1'b0;
    assign layer0_out[1380] = ~x[293] | x[274];
    assign layer0_out[1381] = x[262] | x[272];
    assign layer0_out[1382] = x[224] & ~x[243];
    assign layer0_out[1383] = ~(x[332] | x[340]);
    assign layer0_out[1384] = ~(x[54] | x[65]);
    assign layer0_out[1385] = ~x[152];
    assign layer0_out[1386] = ~x[200];
    assign layer0_out[1387] = ~x[215];
    assign layer0_out[1388] = x[319] & ~x[315];
    assign layer0_out[1389] = ~x[45];
    assign layer0_out[1390] = ~x[314];
    assign layer0_out[1391] = x[366];
    assign layer0_out[1392] = ~x[389];
    assign layer0_out[1393] = ~(x[116] ^ x[136]);
    assign layer0_out[1394] = x[264] ^ x[273];
    assign layer0_out[1395] = x[165];
    assign layer0_out[1396] = ~(x[56] & x[60]);
    assign layer0_out[1397] = x[31];
    assign layer0_out[1398] = x[66] ^ x[67];
    assign layer0_out[1399] = x[194] & ~x[204];
    assign layer0_out[1400] = x[143] & x[156];
    assign layer0_out[1401] = x[117];
    assign layer0_out[1402] = ~x[173];
    assign layer0_out[1403] = x[329] | x[346];
    assign layer0_out[1404] = ~(x[29] & x[30]);
    assign layer0_out[1405] = x[317] & x[328];
    assign layer0_out[1406] = ~(x[170] ^ x[190]);
    assign layer0_out[1407] = 1'b0;
    assign layer0_out[1408] = ~x[29] | x[22];
    assign layer0_out[1409] = x[369] | x[372];
    assign layer0_out[1410] = x[69];
    assign layer0_out[1411] = ~x[218];
    assign layer0_out[1412] = ~(x[298] & x[303]);
    assign layer0_out[1413] = ~(x[134] | x[154]);
    assign layer0_out[1414] = ~(x[112] | x[113]);
    assign layer0_out[1415] = x[54] & x[73];
    assign layer0_out[1416] = x[49] & ~x[38];
    assign layer0_out[1417] = ~x[326] | x[313];
    assign layer0_out[1418] = x[326] | x[346];
    assign layer0_out[1419] = ~(x[278] & x[290]);
    assign layer0_out[1420] = ~(x[383] | x[384]);
    assign layer0_out[1421] = x[219];
    assign layer0_out[1422] = ~x[373] | x[388];
    assign layer0_out[1423] = ~x[178] | x[182];
    assign layer0_out[1424] = ~x[174];
    assign layer0_out[1425] = x[262] | x[276];
    assign layer0_out[1426] = x[44] | x[61];
    assign layer0_out[1427] = ~x[308];
    assign layer0_out[1428] = ~(x[39] | x[55]);
    assign layer0_out[1429] = x[189] & ~x[198];
    assign layer0_out[1430] = x[222] | x[226];
    assign layer0_out[1431] = x[221];
    assign layer0_out[1432] = ~x[392] | x[389];
    assign layer0_out[1433] = ~x[236] | x[247];
    assign layer0_out[1434] = 1'b1;
    assign layer0_out[1435] = ~(x[2] | x[12]);
    assign layer0_out[1436] = ~(x[199] ^ x[220]);
    assign layer0_out[1437] = ~x[316];
    assign layer0_out[1438] = x[319] & ~x[325];
    assign layer0_out[1439] = ~x[67] | x[71];
    assign layer0_out[1440] = x[320] & x[338];
    assign layer0_out[1441] = x[46] | x[50];
    assign layer0_out[1442] = x[142] & ~x[151];
    assign layer0_out[1443] = ~(x[297] & x[316]);
    assign layer0_out[1444] = x[365];
    assign layer0_out[1445] = x[177] ^ x[189];
    assign layer0_out[1446] = ~x[108];
    assign layer0_out[1447] = ~x[266];
    assign layer0_out[1448] = x[244] | x[254];
    assign layer0_out[1449] = ~x[217];
    assign layer0_out[1450] = 1'b0;
    assign layer0_out[1451] = x[326] | x[336];
    assign layer0_out[1452] = ~(x[327] & x[328]);
    assign layer0_out[1453] = x[309] & x[318];
    assign layer0_out[1454] = 1'b0;
    assign layer0_out[1455] = x[32];
    assign layer0_out[1456] = x[85] | x[93];
    assign layer0_out[1457] = x[212];
    assign layer0_out[1458] = ~(x[368] & x[379]);
    assign layer0_out[1459] = ~(x[310] | x[312]);
    assign layer0_out[1460] = ~(x[138] | x[155]);
    assign layer0_out[1461] = x[361];
    assign layer0_out[1462] = ~(x[193] ^ x[197]);
    assign layer0_out[1463] = ~(x[235] ^ x[255]);
    assign layer0_out[1464] = x[108];
    assign layer0_out[1465] = ~x[205];
    assign layer0_out[1466] = x[195] ^ x[205];
    assign layer0_out[1467] = ~x[166];
    assign layer0_out[1468] = x[51] ^ x[53];
    assign layer0_out[1469] = ~(x[188] | x[207]);
    assign layer0_out[1470] = x[312] & ~x[332];
    assign layer0_out[1471] = ~(x[67] & x[75]);
    assign layer0_out[1472] = ~x[372] | x[367];
    assign layer0_out[1473] = ~(x[40] & x[41]);
    assign layer0_out[1474] = x[191] ^ x[200];
    assign layer0_out[1475] = x[157] | x[175];
    assign layer0_out[1476] = x[162] & x[177];
    assign layer0_out[1477] = ~(x[116] | x[117]);
    assign layer0_out[1478] = ~(x[46] & x[49]);
    assign layer0_out[1479] = x[125];
    assign layer0_out[1480] = ~x[69] | x[77];
    assign layer0_out[1481] = 1'b1;
    assign layer0_out[1482] = x[371] | x[389];
    assign layer0_out[1483] = ~x[16] | x[5];
    assign layer0_out[1484] = x[296] | x[306];
    assign layer0_out[1485] = x[275] & ~x[292];
    assign layer0_out[1486] = x[180] | x[186];
    assign layer0_out[1487] = ~x[161];
    assign layer0_out[1488] = 1'b1;
    assign layer0_out[1489] = ~x[328] | x[342];
    assign layer0_out[1490] = x[354] & ~x[351];
    assign layer0_out[1491] = ~(x[189] | x[206]);
    assign layer0_out[1492] = ~x[64];
    assign layer0_out[1493] = x[220] | x[238];
    assign layer0_out[1494] = ~x[215] | x[233];
    assign layer0_out[1495] = ~(x[241] | x[248]);
    assign layer0_out[1496] = ~x[221] | x[207];
    assign layer0_out[1497] = 1'b0;
    assign layer0_out[1498] = ~(x[383] ^ x[389]);
    assign layer0_out[1499] = x[273] ^ x[282];
    assign layer0_out[1500] = ~(x[35] ^ x[46]);
    assign layer0_out[1501] = ~(x[55] ^ x[68]);
    assign layer0_out[1502] = ~(x[165] & x[168]);
    assign layer0_out[1503] = x[386] & ~x[368];
    assign layer0_out[1504] = ~(x[104] ^ x[121]);
    assign layer0_out[1505] = ~(x[14] | x[30]);
    assign layer0_out[1506] = ~x[215] | x[229];
    assign layer0_out[1507] = ~x[237] | x[222];
    assign layer0_out[1508] = ~x[210];
    assign layer0_out[1509] = ~(x[381] | x[385]);
    assign layer0_out[1510] = x[205];
    assign layer0_out[1511] = x[49];
    assign layer0_out[1512] = 1'b0;
    assign layer0_out[1513] = ~x[395];
    assign layer0_out[1514] = ~x[95] | x[107];
    assign layer0_out[1515] = ~x[332] | x[329];
    assign layer0_out[1516] = 1'b0;
    assign layer0_out[1517] = x[150];
    assign layer0_out[1518] = ~(x[264] ^ x[267]);
    assign layer0_out[1519] = x[50] ^ x[61];
    assign layer0_out[1520] = ~x[360] | x[359];
    assign layer0_out[1521] = ~x[293] | x[277];
    assign layer0_out[1522] = x[306];
    assign layer0_out[1523] = ~x[356] | x[373];
    assign layer0_out[1524] = x[204] ^ x[209];
    assign layer0_out[1525] = ~(x[80] | x[82]);
    assign layer0_out[1526] = x[158] | x[159];
    assign layer0_out[1527] = x[225];
    assign layer0_out[1528] = ~(x[261] & x[274]);
    assign layer0_out[1529] = x[220] | x[223];
    assign layer0_out[1530] = ~x[173];
    assign layer0_out[1531] = ~(x[18] ^ x[23]);
    assign layer0_out[1532] = ~(x[65] | x[69]);
    assign layer0_out[1533] = x[66] & x[74];
    assign layer0_out[1534] = x[114] ^ x[116];
    assign layer0_out[1535] = x[337] ^ x[339];
    assign layer0_out[1536] = ~x[189];
    assign layer0_out[1537] = x[315] & ~x[310];
    assign layer0_out[1538] = ~(x[148] & x[154]);
    assign layer0_out[1539] = ~(x[301] | x[312]);
    assign layer0_out[1540] = x[51];
    assign layer0_out[1541] = ~(x[55] | x[64]);
    assign layer0_out[1542] = ~x[371];
    assign layer0_out[1543] = x[112];
    assign layer0_out[1544] = x[297] | x[304];
    assign layer0_out[1545] = x[276] & ~x[292];
    assign layer0_out[1546] = ~x[43];
    assign layer0_out[1547] = x[105] | x[115];
    assign layer0_out[1548] = 1'b1;
    assign layer0_out[1549] = ~x[157];
    assign layer0_out[1550] = x[93] & ~x[106];
    assign layer0_out[1551] = ~(x[299] | x[303]);
    assign layer0_out[1552] = ~(x[331] & x[336]);
    assign layer0_out[1553] = ~x[162] | x[174];
    assign layer0_out[1554] = x[350] & x[368];
    assign layer0_out[1555] = x[316];
    assign layer0_out[1556] = ~(x[98] | x[115]);
    assign layer0_out[1557] = x[183];
    assign layer0_out[1558] = 1'b1;
    assign layer0_out[1559] = ~x[324];
    assign layer0_out[1560] = x[237] | x[238];
    assign layer0_out[1561] = x[282];
    assign layer0_out[1562] = ~x[188];
    assign layer0_out[1563] = ~x[358] | x[372];
    assign layer0_out[1564] = x[217] | x[218];
    assign layer0_out[1565] = 1'b0;
    assign layer0_out[1566] = x[191] | x[192];
    assign layer0_out[1567] = ~(x[56] | x[75]);
    assign layer0_out[1568] = ~(x[239] | x[246]);
    assign layer0_out[1569] = x[18] & ~x[15];
    assign layer0_out[1570] = x[118];
    assign layer0_out[1571] = x[192] & ~x[207];
    assign layer0_out[1572] = x[153] & ~x[143];
    assign layer0_out[1573] = ~x[122];
    assign layer0_out[1574] = x[203];
    assign layer0_out[1575] = ~(x[127] ^ x[144]);
    assign layer0_out[1576] = x[368];
    assign layer0_out[1577] = x[131] & ~x[126];
    assign layer0_out[1578] = x[96];
    assign layer0_out[1579] = ~(x[229] ^ x[239]);
    assign layer0_out[1580] = ~x[110];
    assign layer0_out[1581] = ~x[53];
    assign layer0_out[1582] = 1'b1;
    assign layer0_out[1583] = ~(x[245] | x[258]);
    assign layer0_out[1584] = x[178];
    assign layer0_out[1585] = ~(x[139] | x[146]);
    assign layer0_out[1586] = x[100] | x[112];
    assign layer0_out[1587] = x[284] & x[302];
    assign layer0_out[1588] = 1'b1;
    assign layer0_out[1589] = x[303] & ~x[308];
    assign layer0_out[1590] = ~x[343];
    assign layer0_out[1591] = ~(x[35] | x[53]);
    assign layer0_out[1592] = 1'b0;
    assign layer0_out[1593] = 1'b0;
    assign layer0_out[1594] = 1'b1;
    assign layer0_out[1595] = 1'b0;
    assign layer0_out[1596] = x[214] | x[215];
    assign layer0_out[1597] = ~x[255] | x[273];
    assign layer0_out[1598] = x[103] & ~x[114];
    assign layer0_out[1599] = x[248] & ~x[257];
    assign layer0_out[1600] = ~(x[100] | x[115]);
    assign layer0_out[1601] = ~(x[72] | x[74]);
    assign layer0_out[1602] = 1'b1;
    assign layer0_out[1603] = ~(x[130] ^ x[149]);
    assign layer0_out[1604] = x[20];
    assign layer0_out[1605] = x[200] ^ x[205];
    assign layer0_out[1606] = x[155];
    assign layer0_out[1607] = ~x[69] | x[81];
    assign layer0_out[1608] = x[111] & ~x[124];
    assign layer0_out[1609] = x[78] | x[94];
    assign layer0_out[1610] = x[58] | x[59];
    assign layer0_out[1611] = x[35];
    assign layer0_out[1612] = x[110] & x[111];
    assign layer0_out[1613] = x[245] & x[253];
    assign layer0_out[1614] = x[333] & x[336];
    assign layer0_out[1615] = ~x[117] | x[133];
    assign layer0_out[1616] = x[10];
    assign layer0_out[1617] = x[252] & x[272];
    assign layer0_out[1618] = ~x[160];
    assign layer0_out[1619] = ~(x[319] | x[334]);
    assign layer0_out[1620] = x[338];
    assign layer0_out[1621] = 1'b1;
    assign layer0_out[1622] = ~(x[25] & x[41]);
    assign layer0_out[1623] = x[124] & x[131];
    assign layer0_out[1624] = x[293] | x[311];
    assign layer0_out[1625] = ~(x[18] ^ x[38]);
    assign layer0_out[1626] = x[325] | x[339];
    assign layer0_out[1627] = x[193] & x[202];
    assign layer0_out[1628] = ~x[26];
    assign layer0_out[1629] = ~x[263];
    assign layer0_out[1630] = x[328] | x[346];
    assign layer0_out[1631] = x[250] | x[254];
    assign layer0_out[1632] = ~x[274];
    assign layer0_out[1633] = ~(x[286] ^ x[290]);
    assign layer0_out[1634] = ~x[285];
    assign layer0_out[1635] = ~(x[225] ^ x[233]);
    assign layer0_out[1636] = ~x[361] | x[375];
    assign layer0_out[1637] = x[379];
    assign layer0_out[1638] = x[61] & ~x[57];
    assign layer0_out[1639] = x[171];
    assign layer0_out[1640] = ~x[381];
    assign layer0_out[1641] = ~(x[213] ^ x[232]);
    assign layer0_out[1642] = x[255];
    assign layer0_out[1643] = ~(x[59] & x[65]);
    assign layer0_out[1644] = x[32];
    assign layer0_out[1645] = ~(x[338] | x[350]);
    assign layer0_out[1646] = ~x[279];
    assign layer0_out[1647] = ~(x[291] | x[303]);
    assign layer0_out[1648] = ~(x[319] & x[329]);
    assign layer0_out[1649] = ~(x[242] | x[256]);
    assign layer0_out[1650] = ~(x[339] | x[352]);
    assign layer0_out[1651] = ~x[126] | x[139];
    assign layer0_out[1652] = ~(x[121] | x[132]);
    assign layer0_out[1653] = x[228] & ~x[231];
    assign layer0_out[1654] = ~x[150];
    assign layer0_out[1655] = ~x[343];
    assign layer0_out[1656] = x[308] | x[320];
    assign layer0_out[1657] = ~x[91];
    assign layer0_out[1658] = x[329];
    assign layer0_out[1659] = ~x[108];
    assign layer0_out[1660] = x[203];
    assign layer0_out[1661] = x[150] & ~x[146];
    assign layer0_out[1662] = x[81] ^ x[91];
    assign layer0_out[1663] = ~x[168] | x[156];
    assign layer0_out[1664] = ~x[98];
    assign layer0_out[1665] = ~x[32];
    assign layer0_out[1666] = ~x[52] | x[69];
    assign layer0_out[1667] = ~(x[13] | x[33]);
    assign layer0_out[1668] = x[370] | x[374];
    assign layer0_out[1669] = x[215] & ~x[203];
    assign layer0_out[1670] = 1'b0;
    assign layer0_out[1671] = ~x[207] | x[210];
    assign layer0_out[1672] = x[361] & x[377];
    assign layer0_out[1673] = 1'b0;
    assign layer0_out[1674] = x[384] | x[392];
    assign layer0_out[1675] = ~x[144] | x[153];
    assign layer0_out[1676] = x[363];
    assign layer0_out[1677] = ~x[24];
    assign layer0_out[1678] = ~x[138];
    assign layer0_out[1679] = x[274] & x[291];
    assign layer0_out[1680] = ~x[348] | x[341];
    assign layer0_out[1681] = x[374] | x[378];
    assign layer0_out[1682] = ~(x[322] & x[342]);
    assign layer0_out[1683] = x[116] ^ x[124];
    assign layer0_out[1684] = ~(x[58] | x[79]);
    assign layer0_out[1685] = ~x[136];
    assign layer0_out[1686] = ~(x[194] & x[209]);
    assign layer0_out[1687] = ~x[312] | x[294];
    assign layer0_out[1688] = x[81];
    assign layer0_out[1689] = x[181] & ~x[192];
    assign layer0_out[1690] = x[76] & ~x[78];
    assign layer0_out[1691] = x[77] & ~x[65];
    assign layer0_out[1692] = x[258] & ~x[278];
    assign layer0_out[1693] = ~(x[112] | x[116]);
    assign layer0_out[1694] = ~(x[269] ^ x[281]);
    assign layer0_out[1695] = x[199] | x[216];
    assign layer0_out[1696] = ~x[104];
    assign layer0_out[1697] = ~x[98];
    assign layer0_out[1698] = ~(x[341] | x[354]);
    assign layer0_out[1699] = x[78] ^ x[93];
    assign layer0_out[1700] = ~(x[356] ^ x[376]);
    assign layer0_out[1701] = ~x[309] | x[328];
    assign layer0_out[1702] = ~(x[94] | x[115]);
    assign layer0_out[1703] = x[339] ^ x[357];
    assign layer0_out[1704] = ~x[55] | x[34];
    assign layer0_out[1705] = ~x[91];
    assign layer0_out[1706] = x[233] & x[249];
    assign layer0_out[1707] = ~(x[12] | x[29]);
    assign layer0_out[1708] = x[133] | x[147];
    assign layer0_out[1709] = ~x[212] | x[225];
    assign layer0_out[1710] = x[396] & ~x[395];
    assign layer0_out[1711] = x[147];
    assign layer0_out[1712] = ~x[393] | x[378];
    assign layer0_out[1713] = x[44] | x[58];
    assign layer0_out[1714] = x[171] & ~x[191];
    assign layer0_out[1715] = x[367] | x[379];
    assign layer0_out[1716] = ~x[254];
    assign layer0_out[1717] = ~(x[123] | x[144]);
    assign layer0_out[1718] = ~(x[351] & x[369]);
    assign layer0_out[1719] = x[31] | x[47];
    assign layer0_out[1720] = x[309] | x[321];
    assign layer0_out[1721] = ~x[146] | x[159];
    assign layer0_out[1722] = ~x[91] | x[100];
    assign layer0_out[1723] = x[385];
    assign layer0_out[1724] = ~(x[309] | x[315]);
    assign layer0_out[1725] = x[278] ^ x[298];
    assign layer0_out[1726] = x[168] | x[182];
    assign layer0_out[1727] = x[106] & ~x[115];
    assign layer0_out[1728] = x[276];
    assign layer0_out[1729] = ~x[287] | x[300];
    assign layer0_out[1730] = x[315] ^ x[321];
    assign layer0_out[1731] = x[198];
    assign layer0_out[1732] = ~(x[335] & x[342]);
    assign layer0_out[1733] = x[9] & ~x[26];
    assign layer0_out[1734] = ~(x[73] ^ x[78]);
    assign layer0_out[1735] = ~(x[183] | x[199]);
    assign layer0_out[1736] = x[261] | x[264];
    assign layer0_out[1737] = x[209] & x[229];
    assign layer0_out[1738] = ~(x[228] ^ x[245]);
    assign layer0_out[1739] = ~x[72];
    assign layer0_out[1740] = ~(x[134] | x[143]);
    assign layer0_out[1741] = ~(x[209] | x[225]);
    assign layer0_out[1742] = ~x[349] | x[356];
    assign layer0_out[1743] = x[352] ^ x[358];
    assign layer0_out[1744] = ~x[35];
    assign layer0_out[1745] = ~x[302];
    assign layer0_out[1746] = x[148] & ~x[141];
    assign layer0_out[1747] = x[249];
    assign layer0_out[1748] = x[194] ^ x[203];
    assign layer0_out[1749] = 1'b0;
    assign layer0_out[1750] = x[383] & x[388];
    assign layer0_out[1751] = ~x[350];
    assign layer0_out[1752] = ~(x[315] | x[323]);
    assign layer0_out[1753] = x[45] | x[64];
    assign layer0_out[1754] = ~(x[226] ^ x[244]);
    assign layer0_out[1755] = ~(x[381] | x[399]);
    assign layer0_out[1756] = x[71];
    assign layer0_out[1757] = ~x[144];
    assign layer0_out[1758] = ~(x[205] | x[220]);
    assign layer0_out[1759] = x[280];
    assign layer0_out[1760] = ~x[285] | x[279];
    assign layer0_out[1761] = ~x[100];
    assign layer0_out[1762] = 1'b1;
    assign layer0_out[1763] = 1'b0;
    assign layer0_out[1764] = ~(x[278] | x[285]);
    assign layer0_out[1765] = x[327] & x[333];
    assign layer0_out[1766] = x[220] ^ x[239];
    assign layer0_out[1767] = ~(x[127] | x[128]);
    assign layer0_out[1768] = x[236];
    assign layer0_out[1769] = ~x[69];
    assign layer0_out[1770] = ~x[253] | x[244];
    assign layer0_out[1771] = x[247] & ~x[238];
    assign layer0_out[1772] = x[90];
    assign layer0_out[1773] = x[147] & x[153];
    assign layer0_out[1774] = ~x[143];
    assign layer0_out[1775] = 1'b0;
    assign layer0_out[1776] = x[381] & ~x[364];
    assign layer0_out[1777] = x[172];
    assign layer0_out[1778] = ~x[218];
    assign layer0_out[1779] = ~x[157];
    assign layer0_out[1780] = ~(x[227] ^ x[242]);
    assign layer0_out[1781] = x[108] & x[126];
    assign layer0_out[1782] = x[26];
    assign layer0_out[1783] = x[122] ^ x[143];
    assign layer0_out[1784] = ~x[348];
    assign layer0_out[1785] = x[220] & ~x[214];
    assign layer0_out[1786] = ~(x[122] ^ x[124]);
    assign layer0_out[1787] = ~x[259];
    assign layer0_out[1788] = ~(x[359] ^ x[375]);
    assign layer0_out[1789] = ~x[326];
    assign layer0_out[1790] = ~x[61];
    assign layer0_out[1791] = x[293] ^ x[302];
    assign layer0_out[1792] = ~x[157];
    assign layer0_out[1793] = ~(x[72] | x[85]);
    assign layer0_out[1794] = ~(x[217] | x[236]);
    assign layer0_out[1795] = x[111] & ~x[123];
    assign layer0_out[1796] = ~x[206];
    assign layer0_out[1797] = ~x[46] | x[31];
    assign layer0_out[1798] = ~(x[244] | x[261]);
    assign layer0_out[1799] = ~(x[355] | x[368]);
    assign layer0_out[1800] = x[309];
    assign layer0_out[1801] = x[106] & x[113];
    assign layer0_out[1802] = x[58] | x[62];
    assign layer0_out[1803] = ~(x[268] & x[277]);
    assign layer0_out[1804] = x[216];
    assign layer0_out[1805] = x[118] & x[131];
    assign layer0_out[1806] = ~(x[30] | x[44]);
    assign layer0_out[1807] = ~(x[104] | x[123]);
    assign layer0_out[1808] = x[135];
    assign layer0_out[1809] = 1'b1;
    assign layer0_out[1810] = ~(x[360] ^ x[377]);
    assign layer0_out[1811] = ~x[337];
    assign layer0_out[1812] = 1'b1;
    assign layer0_out[1813] = x[163] ^ x[181];
    assign layer0_out[1814] = 1'b0;
    assign layer0_out[1815] = ~x[75] | x[91];
    assign layer0_out[1816] = x[393] & ~x[389];
    assign layer0_out[1817] = x[314] & ~x[328];
    assign layer0_out[1818] = x[255];
    assign layer0_out[1819] = 1'b0;
    assign layer0_out[1820] = 1'b1;
    assign layer0_out[1821] = ~x[145] | x[138];
    assign layer0_out[1822] = ~(x[22] | x[36]);
    assign layer0_out[1823] = ~(x[165] | x[179]);
    assign layer0_out[1824] = x[1] & x[14];
    assign layer0_out[1825] = 1'b0;
    assign layer0_out[1826] = x[140] | x[153];
    assign layer0_out[1827] = x[194];
    assign layer0_out[1828] = x[196];
    assign layer0_out[1829] = x[181] & x[197];
    assign layer0_out[1830] = x[248];
    assign layer0_out[1831] = x[262] & x[273];
    assign layer0_out[1832] = ~(x[335] | x[337]);
    assign layer0_out[1833] = x[53] | x[55];
    assign layer0_out[1834] = ~x[364] | x[344];
    assign layer0_out[1835] = ~x[30];
    assign layer0_out[1836] = x[77] & ~x[81];
    assign layer0_out[1837] = ~x[362] | x[348];
    assign layer0_out[1838] = x[345] ^ x[362];
    assign layer0_out[1839] = 1'b1;
    assign layer0_out[1840] = x[318] & ~x[315];
    assign layer0_out[1841] = x[169];
    assign layer0_out[1842] = x[17];
    assign layer0_out[1843] = x[217] & ~x[208];
    assign layer0_out[1844] = x[132];
    assign layer0_out[1845] = x[217] | x[231];
    assign layer0_out[1846] = x[278] & ~x[273];
    assign layer0_out[1847] = x[379] ^ x[397];
    assign layer0_out[1848] = x[172];
    assign layer0_out[1849] = ~(x[174] ^ x[182]);
    assign layer0_out[1850] = x[48];
    assign layer0_out[1851] = ~x[20];
    assign layer0_out[1852] = ~x[72] | x[63];
    assign layer0_out[1853] = x[72] & ~x[88];
    assign layer0_out[1854] = x[92];
    assign layer0_out[1855] = x[186] & x[204];
    assign layer0_out[1856] = ~x[235] | x[234];
    assign layer0_out[1857] = ~x[229];
    assign layer0_out[1858] = x[27] & ~x[33];
    assign layer0_out[1859] = x[153] | x[174];
    assign layer0_out[1860] = ~x[293];
    assign layer0_out[1861] = 1'b1;
    assign layer0_out[1862] = x[259] | x[270];
    assign layer0_out[1863] = x[61];
    assign layer0_out[1864] = x[270] & x[285];
    assign layer0_out[1865] = x[169] & ~x[156];
    assign layer0_out[1866] = ~x[236];
    assign layer0_out[1867] = x[122] & x[138];
    assign layer0_out[1868] = ~(x[233] | x[235]);
    assign layer0_out[1869] = x[262] & ~x[254];
    assign layer0_out[1870] = ~x[35];
    assign layer0_out[1871] = x[104] ^ x[115];
    assign layer0_out[1872] = x[293] | x[294];
    assign layer0_out[1873] = ~(x[68] & x[88]);
    assign layer0_out[1874] = ~x[28] | x[15];
    assign layer0_out[1875] = ~(x[49] ^ x[69]);
    assign layer0_out[1876] = 1'b0;
    assign layer0_out[1877] = x[43] | x[64];
    assign layer0_out[1878] = ~x[180];
    assign layer0_out[1879] = x[91] & x[99];
    assign layer0_out[1880] = ~(x[54] & x[70]);
    assign layer0_out[1881] = ~x[152];
    assign layer0_out[1882] = ~(x[140] & x[148]);
    assign layer0_out[1883] = ~(x[74] ^ x[78]);
    assign layer0_out[1884] = ~x[219] | x[220];
    assign layer0_out[1885] = x[47] | x[60];
    assign layer0_out[1886] = ~x[344];
    assign layer0_out[1887] = ~(x[330] | x[347]);
    assign layer0_out[1888] = x[72] & ~x[81];
    assign layer0_out[1889] = x[17];
    assign layer0_out[1890] = ~x[170];
    assign layer0_out[1891] = x[166] & ~x[178];
    assign layer0_out[1892] = ~x[213] | x[208];
    assign layer0_out[1893] = x[320];
    assign layer0_out[1894] = ~x[207] | x[227];
    assign layer0_out[1895] = ~x[220];
    assign layer0_out[1896] = ~x[185] | x[174];
    assign layer0_out[1897] = x[260];
    assign layer0_out[1898] = ~(x[174] & x[187]);
    assign layer0_out[1899] = x[260];
    assign layer0_out[1900] = 1'b1;
    assign layer0_out[1901] = ~(x[75] & x[96]);
    assign layer0_out[1902] = x[334] | x[347];
    assign layer0_out[1903] = x[160];
    assign layer0_out[1904] = ~x[314];
    assign layer0_out[1905] = ~(x[183] | x[200]);
    assign layer0_out[1906] = ~(x[23] | x[42]);
    assign layer0_out[1907] = ~x[316];
    assign layer0_out[1908] = ~(x[100] | x[117]);
    assign layer0_out[1909] = x[200];
    assign layer0_out[1910] = x[260] | x[278];
    assign layer0_out[1911] = ~(x[280] | x[283]);
    assign layer0_out[1912] = x[104] & x[116];
    assign layer0_out[1913] = x[188];
    assign layer0_out[1914] = ~(x[60] & x[79]);
    assign layer0_out[1915] = ~x[250] | x[261];
    assign layer0_out[1916] = ~x[41];
    assign layer0_out[1917] = ~(x[6] | x[19]);
    assign layer0_out[1918] = x[238] & ~x[226];
    assign layer0_out[1919] = x[263] & x[274];
    assign layer0_out[1920] = x[245] ^ x[248];
    assign layer0_out[1921] = ~(x[89] ^ x[95]);
    assign layer0_out[1922] = ~x[45];
    assign layer0_out[1923] = x[130];
    assign layer0_out[1924] = ~(x[325] & x[328]);
    assign layer0_out[1925] = ~(x[46] | x[67]);
    assign layer0_out[1926] = x[65] | x[81];
    assign layer0_out[1927] = ~(x[111] | x[115]);
    assign layer0_out[1928] = x[201] & x[209];
    assign layer0_out[1929] = ~(x[341] | x[344]);
    assign layer0_out[1930] = ~(x[115] ^ x[132]);
    assign layer0_out[1931] = ~x[194];
    assign layer0_out[1932] = x[271] & ~x[280];
    assign layer0_out[1933] = x[320] ^ x[333];
    assign layer0_out[1934] = x[33] | x[46];
    assign layer0_out[1935] = ~(x[206] ^ x[220]);
    assign layer0_out[1936] = ~(x[21] | x[23]);
    assign layer0_out[1937] = ~(x[113] | x[115]);
    assign layer0_out[1938] = x[184] | x[185];
    assign layer0_out[1939] = ~(x[34] ^ x[44]);
    assign layer0_out[1940] = ~x[264];
    assign layer0_out[1941] = x[185] | x[198];
    assign layer0_out[1942] = x[29];
    assign layer0_out[1943] = ~(x[273] | x[284]);
    assign layer0_out[1944] = ~(x[238] | x[258]);
    assign layer0_out[1945] = ~(x[254] | x[256]);
    assign layer0_out[1946] = ~x[171];
    assign layer0_out[1947] = x[124] | x[125];
    assign layer0_out[1948] = ~(x[5] | x[19]);
    assign layer0_out[1949] = x[349] | x[369];
    assign layer0_out[1950] = x[278] & ~x[272];
    assign layer0_out[1951] = ~x[71];
    assign layer0_out[1952] = x[25] & ~x[32];
    assign layer0_out[1953] = ~(x[137] & x[156]);
    assign layer0_out[1954] = x[268];
    assign layer0_out[1955] = ~(x[31] ^ x[42]);
    assign layer0_out[1956] = ~(x[141] | x[152]);
    assign layer0_out[1957] = ~(x[33] | x[51]);
    assign layer0_out[1958] = x[345] & x[353];
    assign layer0_out[1959] = x[208];
    assign layer0_out[1960] = x[121] | x[140];
    assign layer0_out[1961] = x[100] | x[104];
    assign layer0_out[1962] = x[390] & ~x[395];
    assign layer0_out[1963] = x[38] & x[54];
    assign layer0_out[1964] = ~x[392];
    assign layer0_out[1965] = ~x[94];
    assign layer0_out[1966] = x[339] & x[341];
    assign layer0_out[1967] = x[171] & ~x[186];
    assign layer0_out[1968] = ~(x[145] | x[146]);
    assign layer0_out[1969] = x[333];
    assign layer0_out[1970] = x[64] | x[79];
    assign layer0_out[1971] = ~(x[49] | x[58]);
    assign layer0_out[1972] = ~x[113];
    assign layer0_out[1973] = x[378] & ~x[373];
    assign layer0_out[1974] = x[92] & ~x[87];
    assign layer0_out[1975] = ~x[375];
    assign layer0_out[1976] = ~(x[17] | x[25]);
    assign layer0_out[1977] = ~x[77] | x[92];
    assign layer0_out[1978] = ~(x[143] ^ x[158]);
    assign layer0_out[1979] = x[345] & ~x[357];
    assign layer0_out[1980] = ~x[249];
    assign layer0_out[1981] = x[334] & x[346];
    assign layer0_out[1982] = x[127] & ~x[109];
    assign layer0_out[1983] = x[221] | x[228];
    assign layer0_out[1984] = x[244];
    assign layer0_out[1985] = ~(x[251] & x[253]);
    assign layer0_out[1986] = x[22] | x[25];
    assign layer0_out[1987] = ~x[37];
    assign layer0_out[1988] = x[126] | x[136];
    assign layer0_out[1989] = 1'b1;
    assign layer0_out[1990] = x[320];
    assign layer0_out[1991] = ~(x[200] | x[216]);
    assign layer0_out[1992] = x[365] | x[378];
    assign layer0_out[1993] = x[307] & ~x[323];
    assign layer0_out[1994] = x[155];
    assign layer0_out[1995] = ~(x[21] | x[37]);
    assign layer0_out[1996] = x[391] | x[394];
    assign layer0_out[1997] = ~(x[249] & x[263]);
    assign layer0_out[1998] = x[9] | x[28];
    assign layer0_out[1999] = ~x[312];
    assign layer0_out[2000] = x[294];
    assign layer0_out[2001] = ~(x[342] | x[345]);
    assign layer0_out[2002] = x[74];
    assign layer0_out[2003] = ~x[133];
    assign layer0_out[2004] = ~(x[216] | x[232]);
    assign layer0_out[2005] = 1'b1;
    assign layer0_out[2006] = x[18] | x[28];
    assign layer0_out[2007] = ~x[256];
    assign layer0_out[2008] = ~x[320];
    assign layer0_out[2009] = ~(x[70] | x[88]);
    assign layer0_out[2010] = ~(x[196] | x[199]);
    assign layer0_out[2011] = 1'b1;
    assign layer0_out[2012] = x[352] | x[360];
    assign layer0_out[2013] = x[24];
    assign layer0_out[2014] = ~x[371];
    assign layer0_out[2015] = x[163] | x[178];
    assign layer0_out[2016] = ~x[120] | x[124];
    assign layer0_out[2017] = ~x[203] | x[206];
    assign layer0_out[2018] = x[106] & ~x[91];
    assign layer0_out[2019] = ~(x[126] | x[129]);
    assign layer0_out[2020] = ~(x[53] & x[67]);
    assign layer0_out[2021] = x[379];
    assign layer0_out[2022] = x[369] | x[370];
    assign layer0_out[2023] = x[238];
    assign layer0_out[2024] = x[91] ^ x[97];
    assign layer0_out[2025] = ~x[197] | x[211];
    assign layer0_out[2026] = x[43] & ~x[34];
    assign layer0_out[2027] = x[35];
    assign layer0_out[2028] = x[42];
    assign layer0_out[2029] = x[191];
    assign layer0_out[2030] = ~x[142];
    assign layer0_out[2031] = x[120] | x[139];
    assign layer0_out[2032] = x[126];
    assign layer0_out[2033] = x[214];
    assign layer0_out[2034] = ~(x[216] ^ x[228]);
    assign layer0_out[2035] = x[225] & ~x[220];
    assign layer0_out[2036] = x[54];
    assign layer0_out[2037] = 1'b0;
    assign layer0_out[2038] = 1'b0;
    assign layer0_out[2039] = 1'b1;
    assign layer0_out[2040] = x[276] & ~x[267];
    assign layer0_out[2041] = x[58];
    assign layer0_out[2042] = ~x[349];
    assign layer0_out[2043] = x[0] & x[1];
    assign layer0_out[2044] = ~(x[286] ^ x[289]);
    assign layer0_out[2045] = ~(x[159] | x[176]);
    assign layer0_out[2046] = ~(x[169] & x[175]);
    assign layer0_out[2047] = ~x[198];
    assign layer0_out[2048] = ~x[193] | x[210];
    assign layer0_out[2049] = x[115] & x[122];
    assign layer0_out[2050] = ~x[86];
    assign layer0_out[2051] = x[320] | x[322];
    assign layer0_out[2052] = ~(x[304] | x[306]);
    assign layer0_out[2053] = ~x[118];
    assign layer0_out[2054] = x[354] & ~x[361];
    assign layer0_out[2055] = ~x[154];
    assign layer0_out[2056] = ~x[372] | x[376];
    assign layer0_out[2057] = x[370] & x[384];
    assign layer0_out[2058] = x[53] & x[71];
    assign layer0_out[2059] = ~(x[155] ^ x[176]);
    assign layer0_out[2060] = x[111] ^ x[113];
    assign layer0_out[2061] = ~x[288];
    assign layer0_out[2062] = x[316] | x[333];
    assign layer0_out[2063] = x[93] | x[98];
    assign layer0_out[2064] = x[73];
    assign layer0_out[2065] = ~(x[198] & x[214]);
    assign layer0_out[2066] = ~(x[132] ^ x[137]);
    assign layer0_out[2067] = ~x[42] | x[34];
    assign layer0_out[2068] = ~(x[348] | x[364]);
    assign layer0_out[2069] = ~(x[272] ^ x[286]);
    assign layer0_out[2070] = 1'b1;
    assign layer0_out[2071] = ~(x[87] & x[98]);
    assign layer0_out[2072] = x[131] & ~x[112];
    assign layer0_out[2073] = ~x[169];
    assign layer0_out[2074] = ~x[377] | x[383];
    assign layer0_out[2075] = ~(x[182] | x[196]);
    assign layer0_out[2076] = ~(x[133] | x[154]);
    assign layer0_out[2077] = ~(x[208] ^ x[223]);
    assign layer0_out[2078] = ~x[245] | x[238];
    assign layer0_out[2079] = ~x[79];
    assign layer0_out[2080] = x[249] | x[268];
    assign layer0_out[2081] = ~x[316];
    assign layer0_out[2082] = ~(x[67] ^ x[84]);
    assign layer0_out[2083] = 1'b0;
    assign layer0_out[2084] = ~(x[158] ^ x[176]);
    assign layer0_out[2085] = ~(x[52] ^ x[73]);
    assign layer0_out[2086] = x[261] & ~x[277];
    assign layer0_out[2087] = x[329] | x[333];
    assign layer0_out[2088] = ~x[367];
    assign layer0_out[2089] = x[27] ^ x[41];
    assign layer0_out[2090] = ~x[101] | x[122];
    assign layer0_out[2091] = ~(x[325] | x[326]);
    assign layer0_out[2092] = x[136] & ~x[120];
    assign layer0_out[2093] = x[237] | x[256];
    assign layer0_out[2094] = x[351] | x[356];
    assign layer0_out[2095] = ~(x[170] | x[176]);
    assign layer0_out[2096] = ~x[40];
    assign layer0_out[2097] = ~(x[169] | x[188]);
    assign layer0_out[2098] = x[11] & ~x[17];
    assign layer0_out[2099] = x[48] ^ x[64];
    assign layer0_out[2100] = ~x[253];
    assign layer0_out[2101] = x[73];
    assign layer0_out[2102] = x[205] ^ x[208];
    assign layer0_out[2103] = x[203];
    assign layer0_out[2104] = x[28];
    assign layer0_out[2105] = ~x[125];
    assign layer0_out[2106] = x[295];
    assign layer0_out[2107] = x[360] & ~x[361];
    assign layer0_out[2108] = ~(x[8] | x[10]);
    assign layer0_out[2109] = ~(x[236] & x[238]);
    assign layer0_out[2110] = x[72] | x[90];
    assign layer0_out[2111] = ~x[348];
    assign layer0_out[2112] = x[355];
    assign layer0_out[2113] = ~(x[300] | x[302]);
    assign layer0_out[2114] = 1'b0;
    assign layer0_out[2115] = x[94];
    assign layer0_out[2116] = x[92];
    assign layer0_out[2117] = ~x[26];
    assign layer0_out[2118] = x[168] ^ x[170];
    assign layer0_out[2119] = ~x[346];
    assign layer0_out[2120] = ~x[44] | x[35];
    assign layer0_out[2121] = x[32];
    assign layer0_out[2122] = ~x[51];
    assign layer0_out[2123] = ~(x[204] ^ x[207]);
    assign layer0_out[2124] = ~x[146];
    assign layer0_out[2125] = x[104] & ~x[99];
    assign layer0_out[2126] = x[202] & x[215];
    assign layer0_out[2127] = x[112] ^ x[120];
    assign layer0_out[2128] = 1'b0;
    assign layer0_out[2129] = x[390] & ~x[397];
    assign layer0_out[2130] = ~(x[77] ^ x[86]);
    assign layer0_out[2131] = ~x[44];
    assign layer0_out[2132] = x[262] | x[266];
    assign layer0_out[2133] = ~x[325];
    assign layer0_out[2134] = x[20] | x[21];
    assign layer0_out[2135] = x[146];
    assign layer0_out[2136] = ~(x[99] ^ x[100]);
    assign layer0_out[2137] = ~x[66];
    assign layer0_out[2138] = ~x[28] | x[12];
    assign layer0_out[2139] = ~(x[67] | x[68]);
    assign layer0_out[2140] = 1'b0;
    assign layer0_out[2141] = x[93] & x[105];
    assign layer0_out[2142] = x[226] & ~x[240];
    assign layer0_out[2143] = ~x[120] | x[132];
    assign layer0_out[2144] = x[339] | x[358];
    assign layer0_out[2145] = x[338];
    assign layer0_out[2146] = ~x[328];
    assign layer0_out[2147] = ~x[380];
    assign layer0_out[2148] = x[219];
    assign layer0_out[2149] = x[288] | x[289];
    assign layer0_out[2150] = 1'b1;
    assign layer0_out[2151] = ~x[91];
    assign layer0_out[2152] = x[259] & ~x[258];
    assign layer0_out[2153] = ~(x[155] | x[164]);
    assign layer0_out[2154] = ~x[164];
    assign layer0_out[2155] = x[348] & ~x[354];
    assign layer0_out[2156] = ~(x[338] | x[355]);
    assign layer0_out[2157] = x[336] ^ x[349];
    assign layer0_out[2158] = x[103] & ~x[85];
    assign layer0_out[2159] = x[41] ^ x[52];
    assign layer0_out[2160] = ~x[94];
    assign layer0_out[2161] = x[296] | x[298];
    assign layer0_out[2162] = ~x[76];
    assign layer0_out[2163] = x[202];
    assign layer0_out[2164] = x[367];
    assign layer0_out[2165] = x[166] ^ x[172];
    assign layer0_out[2166] = ~(x[85] & x[90]);
    assign layer0_out[2167] = ~(x[222] ^ x[230]);
    assign layer0_out[2168] = ~x[317] | x[304];
    assign layer0_out[2169] = x[331] & x[349];
    assign layer0_out[2170] = ~(x[15] & x[16]);
    assign layer0_out[2171] = x[219];
    assign layer0_out[2172] = x[31] | x[50];
    assign layer0_out[2173] = x[293] | x[299];
    assign layer0_out[2174] = ~x[238] | x[222];
    assign layer0_out[2175] = x[125] | x[134];
    assign layer0_out[2176] = x[272];
    assign layer0_out[2177] = ~x[245];
    assign layer0_out[2178] = x[186];
    assign layer0_out[2179] = ~x[75];
    assign layer0_out[2180] = x[355];
    assign layer0_out[2181] = ~(x[211] ^ x[215]);
    assign layer0_out[2182] = ~(x[334] | x[348]);
    assign layer0_out[2183] = x[90];
    assign layer0_out[2184] = ~(x[202] | x[217]);
    assign layer0_out[2185] = x[75] ^ x[79];
    assign layer0_out[2186] = x[132] | x[135];
    assign layer0_out[2187] = ~x[244];
    assign layer0_out[2188] = ~(x[186] ^ x[205]);
    assign layer0_out[2189] = x[184] | x[202];
    assign layer0_out[2190] = x[46] | x[54];
    assign layer0_out[2191] = ~(x[194] & x[205]);
    assign layer0_out[2192] = ~(x[278] ^ x[295]);
    assign layer0_out[2193] = ~(x[7] ^ x[24]);
    assign layer0_out[2194] = ~x[224];
    assign layer0_out[2195] = x[303] | x[322];
    assign layer0_out[2196] = ~(x[46] | x[47]);
    assign layer0_out[2197] = 1'b0;
    assign layer0_out[2198] = ~(x[122] ^ x[125]);
    assign layer0_out[2199] = x[223];
    assign layer0_out[2200] = x[105];
    assign layer0_out[2201] = x[265] & ~x[259];
    assign layer0_out[2202] = ~(x[169] | x[172]);
    assign layer0_out[2203] = x[184];
    assign layer0_out[2204] = x[215] & x[219];
    assign layer0_out[2205] = ~(x[360] | x[365]);
    assign layer0_out[2206] = ~(x[218] | x[236]);
    assign layer0_out[2207] = 1'b1;
    assign layer0_out[2208] = x[378];
    assign layer0_out[2209] = ~(x[267] & x[287]);
    assign layer0_out[2210] = ~(x[4] | x[5]);
    assign layer0_out[2211] = ~(x[365] | x[385]);
    assign layer0_out[2212] = x[399];
    assign layer0_out[2213] = ~(x[247] | x[264]);
    assign layer0_out[2214] = ~x[95];
    assign layer0_out[2215] = x[240];
    assign layer0_out[2216] = 1'b0;
    assign layer0_out[2217] = ~(x[81] | x[99]);
    assign layer0_out[2218] = ~x[321];
    assign layer0_out[2219] = x[221];
    assign layer0_out[2220] = ~x[185];
    assign layer0_out[2221] = ~(x[373] & x[390]);
    assign layer0_out[2222] = ~(x[316] | x[334]);
    assign layer0_out[2223] = 1'b1;
    assign layer0_out[2224] = ~(x[54] ^ x[71]);
    assign layer0_out[2225] = x[67] ^ x[78];
    assign layer0_out[2226] = ~(x[77] ^ x[85]);
    assign layer0_out[2227] = ~(x[121] & x[126]);
    assign layer0_out[2228] = x[329] & x[334];
    assign layer0_out[2229] = x[128];
    assign layer0_out[2230] = ~x[185];
    assign layer0_out[2231] = x[186];
    assign layer0_out[2232] = x[217];
    assign layer0_out[2233] = ~(x[165] | x[171]);
    assign layer0_out[2234] = ~x[105] | x[94];
    assign layer0_out[2235] = x[375] & x[381];
    assign layer0_out[2236] = x[395] & ~x[378];
    assign layer0_out[2237] = ~x[124];
    assign layer0_out[2238] = x[295] | x[315];
    assign layer0_out[2239] = ~(x[144] ^ x[160]);
    assign layer0_out[2240] = ~(x[36] | x[38]);
    assign layer0_out[2241] = ~(x[59] ^ x[76]);
    assign layer0_out[2242] = 1'b1;
    assign layer0_out[2243] = x[151] | x[157];
    assign layer0_out[2244] = x[257] & ~x[242];
    assign layer0_out[2245] = x[301];
    assign layer0_out[2246] = x[326] & ~x[316];
    assign layer0_out[2247] = x[212] | x[213];
    assign layer0_out[2248] = ~(x[375] | x[387]);
    assign layer0_out[2249] = ~(x[264] | x[276]);
    assign layer0_out[2250] = x[244];
    assign layer0_out[2251] = ~(x[380] ^ x[397]);
    assign layer0_out[2252] = x[26];
    assign layer0_out[2253] = x[43] ^ x[63];
    assign layer0_out[2254] = x[264] ^ x[283];
    assign layer0_out[2255] = ~x[265];
    assign layer0_out[2256] = x[62] | x[74];
    assign layer0_out[2257] = x[357] ^ x[375];
    assign layer0_out[2258] = ~x[264];
    assign layer0_out[2259] = 1'b0;
    assign layer0_out[2260] = ~x[95] | x[90];
    assign layer0_out[2261] = x[97] ^ x[100];
    assign layer0_out[2262] = ~(x[34] | x[52]);
    assign layer0_out[2263] = ~(x[242] | x[246]);
    assign layer0_out[2264] = x[244] | x[262];
    assign layer0_out[2265] = x[106] ^ x[125];
    assign layer0_out[2266] = x[12];
    assign layer0_out[2267] = x[136];
    assign layer0_out[2268] = x[355] | x[371];
    assign layer0_out[2269] = x[197];
    assign layer0_out[2270] = 1'b0;
    assign layer0_out[2271] = ~x[142];
    assign layer0_out[2272] = x[365] | x[384];
    assign layer0_out[2273] = x[97] & ~x[109];
    assign layer0_out[2274] = ~x[133];
    assign layer0_out[2275] = ~x[135];
    assign layer0_out[2276] = x[291];
    assign layer0_out[2277] = x[44] & x[48];
    assign layer0_out[2278] = ~(x[323] | x[325]);
    assign layer0_out[2279] = x[308] | x[316];
    assign layer0_out[2280] = ~x[19];
    assign layer0_out[2281] = x[369] & ~x[380];
    assign layer0_out[2282] = x[320] | x[325];
    assign layer0_out[2283] = x[372] | x[379];
    assign layer0_out[2284] = x[112];
    assign layer0_out[2285] = ~x[336] | x[348];
    assign layer0_out[2286] = ~(x[331] & x[340]);
    assign layer0_out[2287] = ~x[61];
    assign layer0_out[2288] = ~x[149];
    assign layer0_out[2289] = ~x[344] | x[335];
    assign layer0_out[2290] = ~x[241] | x[252];
    assign layer0_out[2291] = 1'b0;
    assign layer0_out[2292] = ~(x[220] & x[221]);
    assign layer0_out[2293] = ~x[349];
    assign layer0_out[2294] = ~(x[356] & x[366]);
    assign layer0_out[2295] = ~(x[102] ^ x[117]);
    assign layer0_out[2296] = x[24] & x[27];
    assign layer0_out[2297] = x[143] & x[150];
    assign layer0_out[2298] = x[318] ^ x[337];
    assign layer0_out[2299] = x[161] | x[175];
    assign layer0_out[2300] = x[205];
    assign layer0_out[2301] = ~x[244];
    assign layer0_out[2302] = x[11] & ~x[21];
    assign layer0_out[2303] = x[89];
    assign layer0_out[2304] = x[120] ^ x[138];
    assign layer0_out[2305] = x[13] | x[15];
    assign layer0_out[2306] = x[241] & ~x[257];
    assign layer0_out[2307] = x[90] | x[110];
    assign layer0_out[2308] = ~x[173];
    assign layer0_out[2309] = x[146] | x[148];
    assign layer0_out[2310] = x[39] & ~x[36];
    assign layer0_out[2311] = x[190] | x[205];
    assign layer0_out[2312] = x[364] & ~x[347];
    assign layer0_out[2313] = ~(x[81] & x[88]);
    assign layer0_out[2314] = ~(x[187] | x[204]);
    assign layer0_out[2315] = ~(x[301] | x[321]);
    assign layer0_out[2316] = ~x[213] | x[203];
    assign layer0_out[2317] = x[59];
    assign layer0_out[2318] = ~(x[97] ^ x[104]);
    assign layer0_out[2319] = x[149] & x[150];
    assign layer0_out[2320] = x[209] & ~x[195];
    assign layer0_out[2321] = ~(x[342] | x[358]);
    assign layer0_out[2322] = x[134];
    assign layer0_out[2323] = ~x[269] | x[276];
    assign layer0_out[2324] = ~x[255] | x[252];
    assign layer0_out[2325] = x[109] & x[111];
    assign layer0_out[2326] = x[51] & x[55];
    assign layer0_out[2327] = ~x[309];
    assign layer0_out[2328] = x[207] | x[212];
    assign layer0_out[2329] = x[157];
    assign layer0_out[2330] = ~(x[351] | x[361]);
    assign layer0_out[2331] = ~(x[191] ^ x[195]);
    assign layer0_out[2332] = x[165] & ~x[156];
    assign layer0_out[2333] = 1'b0;
    assign layer0_out[2334] = x[158] ^ x[168];
    assign layer0_out[2335] = ~x[215];
    assign layer0_out[2336] = x[253] & ~x[258];
    assign layer0_out[2337] = x[41] | x[44];
    assign layer0_out[2338] = ~(x[188] & x[189]);
    assign layer0_out[2339] = x[81] | x[87];
    assign layer0_out[2340] = x[358] | x[367];
    assign layer0_out[2341] = x[48] | x[59];
    assign layer0_out[2342] = ~(x[183] | x[202]);
    assign layer0_out[2343] = ~(x[192] ^ x[198]);
    assign layer0_out[2344] = ~x[346];
    assign layer0_out[2345] = ~x[216];
    assign layer0_out[2346] = ~x[269] | x[256];
    assign layer0_out[2347] = x[175];
    assign layer0_out[2348] = 1'b1;
    assign layer0_out[2349] = ~x[49];
    assign layer0_out[2350] = ~(x[42] & x[44]);
    assign layer0_out[2351] = x[391] & x[398];
    assign layer0_out[2352] = ~x[28] | x[14];
    assign layer0_out[2353] = ~(x[226] | x[237]);
    assign layer0_out[2354] = ~x[348];
    assign layer0_out[2355] = x[192];
    assign layer0_out[2356] = x[13] & ~x[14];
    assign layer0_out[2357] = x[392] ^ x[393];
    assign layer0_out[2358] = x[230];
    assign layer0_out[2359] = x[214];
    assign layer0_out[2360] = x[53];
    assign layer0_out[2361] = ~x[333];
    assign layer0_out[2362] = ~x[230];
    assign layer0_out[2363] = x[243] | x[261];
    assign layer0_out[2364] = ~x[331];
    assign layer0_out[2365] = x[308] & x[322];
    assign layer0_out[2366] = x[228] | x[241];
    assign layer0_out[2367] = ~(x[102] | x[111]);
    assign layer0_out[2368] = ~x[101];
    assign layer0_out[2369] = ~x[26];
    assign layer0_out[2370] = ~x[19] | x[1];
    assign layer0_out[2371] = ~x[193] | x[184];
    assign layer0_out[2372] = ~x[42];
    assign layer0_out[2373] = ~(x[315] | x[334]);
    assign layer0_out[2374] = 1'b0;
    assign layer0_out[2375] = x[152] & ~x[137];
    assign layer0_out[2376] = x[73] & ~x[79];
    assign layer0_out[2377] = ~(x[292] ^ x[297]);
    assign layer0_out[2378] = ~x[94] | x[80];
    assign layer0_out[2379] = x[379];
    assign layer0_out[2380] = x[185] & x[206];
    assign layer0_out[2381] = x[376] | x[391];
    assign layer0_out[2382] = ~x[155];
    assign layer0_out[2383] = ~x[183];
    assign layer0_out[2384] = x[122];
    assign layer0_out[2385] = x[371] | x[380];
    assign layer0_out[2386] = x[271] & ~x[251];
    assign layer0_out[2387] = ~(x[68] & x[76]);
    assign layer0_out[2388] = x[179];
    assign layer0_out[2389] = ~(x[149] | x[165]);
    assign layer0_out[2390] = ~x[244];
    assign layer0_out[2391] = ~x[394];
    assign layer0_out[2392] = x[22];
    assign layer0_out[2393] = x[367] & ~x[357];
    assign layer0_out[2394] = x[49] | x[54];
    assign layer0_out[2395] = x[118];
    assign layer0_out[2396] = x[175] | x[195];
    assign layer0_out[2397] = ~x[21] | x[3];
    assign layer0_out[2398] = x[240];
    assign layer0_out[2399] = ~(x[73] & x[90]);
    assign layer0_out[2400] = ~x[332];
    assign layer0_out[2401] = ~x[251];
    assign layer0_out[2402] = x[247] & ~x[233];
    assign layer0_out[2403] = x[97] | x[99];
    assign layer0_out[2404] = ~x[117];
    assign layer0_out[2405] = ~(x[189] | x[207]);
    assign layer0_out[2406] = x[355];
    assign layer0_out[2407] = x[255] & ~x[253];
    assign layer0_out[2408] = 1'b0;
    assign layer0_out[2409] = x[243] & ~x[235];
    assign layer0_out[2410] = x[348] | x[356];
    assign layer0_out[2411] = ~(x[171] ^ x[178]);
    assign layer0_out[2412] = 1'b0;
    assign layer0_out[2413] = x[365];
    assign layer0_out[2414] = ~x[281] | x[270];
    assign layer0_out[2415] = x[330] ^ x[348];
    assign layer0_out[2416] = x[374] ^ x[386];
    assign layer0_out[2417] = 1'b1;
    assign layer0_out[2418] = ~x[137] | x[121];
    assign layer0_out[2419] = ~x[339] | x[354];
    assign layer0_out[2420] = x[21] & x[33];
    assign layer0_out[2421] = ~(x[204] | x[224]);
    assign layer0_out[2422] = x[108];
    assign layer0_out[2423] = x[186];
    assign layer0_out[2424] = x[338] & ~x[352];
    assign layer0_out[2425] = x[25] & ~x[28];
    assign layer0_out[2426] = x[104];
    assign layer0_out[2427] = ~(x[70] | x[82]);
    assign layer0_out[2428] = x[285] & ~x[271];
    assign layer0_out[2429] = ~x[242] | x[252];
    assign layer0_out[2430] = x[107] ^ x[124];
    assign layer0_out[2431] = x[62] & x[83];
    assign layer0_out[2432] = ~x[119];
    assign layer0_out[2433] = 1'b0;
    assign layer0_out[2434] = x[314] & ~x[296];
    assign layer0_out[2435] = ~x[61];
    assign layer0_out[2436] = ~x[167];
    assign layer0_out[2437] = x[66] & x[79];
    assign layer0_out[2438] = 1'b1;
    assign layer0_out[2439] = x[173];
    assign layer0_out[2440] = x[156];
    assign layer0_out[2441] = x[280] & ~x[279];
    assign layer0_out[2442] = ~(x[193] | x[194]);
    assign layer0_out[2443] = 1'b1;
    assign layer0_out[2444] = ~(x[345] | x[365]);
    assign layer0_out[2445] = x[74] ^ x[77];
    assign layer0_out[2446] = 1'b1;
    assign layer0_out[2447] = ~x[303] | x[304];
    assign layer0_out[2448] = x[45] & x[56];
    assign layer0_out[2449] = ~(x[145] & x[156]);
    assign layer0_out[2450] = ~(x[178] | x[197]);
    assign layer0_out[2451] = x[52];
    assign layer0_out[2452] = ~x[68];
    assign layer0_out[2453] = ~(x[16] | x[19]);
    assign layer0_out[2454] = ~x[219];
    assign layer0_out[2455] = ~(x[312] ^ x[317]);
    assign layer0_out[2456] = x[151] & x[167];
    assign layer0_out[2457] = ~x[191] | x[197];
    assign layer0_out[2458] = x[232] & ~x[220];
    assign layer0_out[2459] = x[54] & x[62];
    assign layer0_out[2460] = ~(x[76] & x[92]);
    assign layer0_out[2461] = ~x[281] | x[272];
    assign layer0_out[2462] = ~x[29];
    assign layer0_out[2463] = 1'b0;
    assign layer0_out[2464] = ~(x[246] | x[256]);
    assign layer0_out[2465] = ~(x[265] ^ x[267]);
    assign layer0_out[2466] = ~(x[96] | x[115]);
    assign layer0_out[2467] = ~x[211] | x[220];
    assign layer0_out[2468] = x[165];
    assign layer0_out[2469] = ~x[246];
    assign layer0_out[2470] = x[129] | x[144];
    assign layer0_out[2471] = 1'b0;
    assign layer0_out[2472] = ~(x[173] | x[181]);
    assign layer0_out[2473] = ~x[385] | x[367];
    assign layer0_out[2474] = x[296] & ~x[289];
    assign layer0_out[2475] = ~x[97];
    assign layer0_out[2476] = 1'b1;
    assign layer0_out[2477] = x[306] ^ x[322];
    assign layer0_out[2478] = x[143];
    assign layer0_out[2479] = x[81] & ~x[73];
    assign layer0_out[2480] = x[165];
    assign layer0_out[2481] = ~(x[181] | x[187]);
    assign layer0_out[2482] = 1'b0;
    assign layer0_out[2483] = ~(x[322] | x[331]);
    assign layer0_out[2484] = x[23] & x[33];
    assign layer0_out[2485] = x[59];
    assign layer0_out[2486] = ~x[19];
    assign layer0_out[2487] = x[159] & ~x[138];
    assign layer0_out[2488] = x[295];
    assign layer0_out[2489] = x[374] & ~x[382];
    assign layer0_out[2490] = ~x[229];
    assign layer0_out[2491] = x[43] & x[53];
    assign layer0_out[2492] = ~x[372];
    assign layer0_out[2493] = ~x[379];
    assign layer0_out[2494] = ~x[12];
    assign layer0_out[2495] = x[232] | x[252];
    assign layer0_out[2496] = ~(x[58] ^ x[75]);
    assign layer0_out[2497] = 1'b0;
    assign layer0_out[2498] = x[61];
    assign layer0_out[2499] = x[234] & x[254];
    assign layer0_out[2500] = x[221] & x[236];
    assign layer0_out[2501] = ~(x[74] | x[75]);
    assign layer0_out[2502] = x[222];
    assign layer0_out[2503] = ~(x[74] | x[88]);
    assign layer0_out[2504] = ~x[249] | x[239];
    assign layer0_out[2505] = ~x[232];
    assign layer0_out[2506] = x[310] & ~x[326];
    assign layer0_out[2507] = x[276] | x[293];
    assign layer0_out[2508] = 1'b0;
    assign layer0_out[2509] = x[9] | x[20];
    assign layer0_out[2510] = ~(x[102] | x[110]);
    assign layer0_out[2511] = x[78];
    assign layer0_out[2512] = ~x[240];
    assign layer0_out[2513] = 1'b0;
    assign layer0_out[2514] = x[378] ^ x[384];
    assign layer0_out[2515] = x[350];
    assign layer0_out[2516] = ~x[342] | x[332];
    assign layer0_out[2517] = x[129] | x[149];
    assign layer0_out[2518] = ~x[109];
    assign layer0_out[2519] = 1'b1;
    assign layer0_out[2520] = 1'b0;
    assign layer0_out[2521] = 1'b1;
    assign layer0_out[2522] = ~x[149];
    assign layer0_out[2523] = x[167];
    assign layer0_out[2524] = ~(x[159] | x[167]);
    assign layer0_out[2525] = ~x[18];
    assign layer0_out[2526] = ~(x[92] & x[108]);
    assign layer0_out[2527] = 1'b1;
    assign layer0_out[2528] = x[82];
    assign layer0_out[2529] = x[302];
    assign layer0_out[2530] = x[237] | x[243];
    assign layer0_out[2531] = ~x[186] | x[187];
    assign layer0_out[2532] = x[168] & ~x[147];
    assign layer0_out[2533] = ~x[221];
    assign layer0_out[2534] = ~x[36] | x[52];
    assign layer0_out[2535] = ~(x[22] | x[39]);
    assign layer0_out[2536] = x[27] & ~x[20];
    assign layer0_out[2537] = x[93] ^ x[113];
    assign layer0_out[2538] = x[133] & ~x[119];
    assign layer0_out[2539] = x[238] & ~x[256];
    assign layer0_out[2540] = x[93];
    assign layer0_out[2541] = x[245] | x[246];
    assign layer0_out[2542] = x[19] ^ x[24];
    assign layer0_out[2543] = ~(x[307] ^ x[321]);
    assign layer0_out[2544] = x[50] & x[62];
    assign layer0_out[2545] = x[177];
    assign layer0_out[2546] = ~x[69];
    assign layer0_out[2547] = ~(x[83] | x[94]);
    assign layer0_out[2548] = x[9] & x[13];
    assign layer0_out[2549] = ~x[371];
    assign layer0_out[2550] = x[263];
    assign layer0_out[2551] = x[83] & x[100];
    assign layer0_out[2552] = ~(x[24] | x[28]);
    assign layer0_out[2553] = x[27];
    assign layer0_out[2554] = x[216] | x[219];
    assign layer0_out[2555] = 1'b1;
    assign layer0_out[2556] = x[50];
    assign layer0_out[2557] = x[100] & ~x[89];
    assign layer0_out[2558] = ~x[168] | x[177];
    assign layer0_out[2559] = x[297];
    assign layer0_out[2560] = x[385];
    assign layer0_out[2561] = x[30] ^ x[50];
    assign layer0_out[2562] = ~x[302];
    assign layer0_out[2563] = ~x[84];
    assign layer0_out[2564] = x[222];
    assign layer0_out[2565] = x[57] & ~x[52];
    assign layer0_out[2566] = ~x[169];
    assign layer0_out[2567] = 1'b0;
    assign layer0_out[2568] = x[352] | x[356];
    assign layer0_out[2569] = x[70];
    assign layer0_out[2570] = x[67];
    assign layer0_out[2571] = x[278] & ~x[291];
    assign layer0_out[2572] = x[191] & ~x[196];
    assign layer0_out[2573] = x[88] ^ x[89];
    assign layer0_out[2574] = x[270] ^ x[279];
    assign layer0_out[2575] = ~x[306] | x[293];
    assign layer0_out[2576] = ~x[268];
    assign layer0_out[2577] = ~x[362] | x[380];
    assign layer0_out[2578] = x[235] & ~x[250];
    assign layer0_out[2579] = ~(x[182] | x[185]);
    assign layer0_out[2580] = x[131];
    assign layer0_out[2581] = ~(x[260] | x[277]);
    assign layer0_out[2582] = x[279] & ~x[272];
    assign layer0_out[2583] = x[52];
    assign layer0_out[2584] = ~x[308];
    assign layer0_out[2585] = ~x[168];
    assign layer0_out[2586] = x[82] & x[89];
    assign layer0_out[2587] = ~(x[146] | x[155]);
    assign layer0_out[2588] = x[172];
    assign layer0_out[2589] = x[97] | x[107];
    assign layer0_out[2590] = ~(x[29] ^ x[49]);
    assign layer0_out[2591] = ~(x[362] & x[365]);
    assign layer0_out[2592] = 1'b0;
    assign layer0_out[2593] = ~x[351] | x[353];
    assign layer0_out[2594] = ~(x[153] & x[169]);
    assign layer0_out[2595] = ~x[268];
    assign layer0_out[2596] = x[224];
    assign layer0_out[2597] = ~x[96] | x[100];
    assign layer0_out[2598] = ~(x[45] & x[49]);
    assign layer0_out[2599] = x[384] | x[385];
    assign layer0_out[2600] = ~x[309] | x[316];
    assign layer0_out[2601] = x[319] ^ x[321];
    assign layer0_out[2602] = ~x[128] | x[116];
    assign layer0_out[2603] = ~x[345] | x[356];
    assign layer0_out[2604] = ~x[367] | x[378];
    assign layer0_out[2605] = 1'b0;
    assign layer0_out[2606] = x[121] & ~x[100];
    assign layer0_out[2607] = x[312] | x[329];
    assign layer0_out[2608] = ~(x[33] ^ x[47]);
    assign layer0_out[2609] = 1'b1;
    assign layer0_out[2610] = ~x[272] | x[253];
    assign layer0_out[2611] = x[305] & ~x[298];
    assign layer0_out[2612] = ~(x[355] | x[372]);
    assign layer0_out[2613] = ~x[95];
    assign layer0_out[2614] = ~(x[39] & x[44]);
    assign layer0_out[2615] = ~x[83];
    assign layer0_out[2616] = x[3] & ~x[13];
    assign layer0_out[2617] = x[62];
    assign layer0_out[2618] = ~x[173] | x[164];
    assign layer0_out[2619] = ~x[24];
    assign layer0_out[2620] = ~x[357] | x[343];
    assign layer0_out[2621] = 1'b1;
    assign layer0_out[2622] = x[160] & x[172];
    assign layer0_out[2623] = ~(x[99] ^ x[114]);
    assign layer0_out[2624] = ~(x[217] | x[227]);
    assign layer0_out[2625] = ~(x[75] & x[95]);
    assign layer0_out[2626] = ~x[29] | x[50];
    assign layer0_out[2627] = x[229] | x[249];
    assign layer0_out[2628] = ~x[303];
    assign layer0_out[2629] = ~(x[28] & x[31]);
    assign layer0_out[2630] = x[253] & x[271];
    assign layer0_out[2631] = x[234];
    assign layer0_out[2632] = ~x[368];
    assign layer0_out[2633] = x[358] | x[377];
    assign layer0_out[2634] = ~x[55];
    assign layer0_out[2635] = ~(x[316] | x[329]);
    assign layer0_out[2636] = ~x[283] | x[265];
    assign layer0_out[2637] = x[394] | x[396];
    assign layer0_out[2638] = x[97] | x[113];
    assign layer0_out[2639] = ~(x[202] & x[207]);
    assign layer0_out[2640] = ~x[397];
    assign layer0_out[2641] = x[5] & ~x[26];
    assign layer0_out[2642] = ~(x[85] ^ x[88]);
    assign layer0_out[2643] = x[107];
    assign layer0_out[2644] = x[179];
    assign layer0_out[2645] = x[283] ^ x[293];
    assign layer0_out[2646] = x[279] | x[294];
    assign layer0_out[2647] = x[305] ^ x[323];
    assign layer0_out[2648] = ~x[206];
    assign layer0_out[2649] = ~x[150] | x[139];
    assign layer0_out[2650] = ~x[334];
    assign layer0_out[2651] = x[279];
    assign layer0_out[2652] = ~(x[47] | x[67]);
    assign layer0_out[2653] = ~(x[252] & x[268]);
    assign layer0_out[2654] = ~x[379] | x[385];
    assign layer0_out[2655] = ~x[56];
    assign layer0_out[2656] = ~(x[324] | x[341]);
    assign layer0_out[2657] = x[42] & x[43];
    assign layer0_out[2658] = x[127] | x[143];
    assign layer0_out[2659] = ~x[236];
    assign layer0_out[2660] = ~x[114] | x[121];
    assign layer0_out[2661] = ~x[149];
    assign layer0_out[2662] = ~(x[270] & x[290]);
    assign layer0_out[2663] = 1'b1;
    assign layer0_out[2664] = ~(x[178] & x[180]);
    assign layer0_out[2665] = x[212] | x[227];
    assign layer0_out[2666] = ~x[171] | x[160];
    assign layer0_out[2667] = ~x[309] | x[322];
    assign layer0_out[2668] = x[69] & ~x[86];
    assign layer0_out[2669] = 1'b1;
    assign layer0_out[2670] = x[266] & ~x[254];
    assign layer0_out[2671] = ~x[224];
    assign layer0_out[2672] = ~(x[196] | x[210]);
    assign layer0_out[2673] = ~(x[388] | x[389]);
    assign layer0_out[2674] = x[351];
    assign layer0_out[2675] = ~x[78];
    assign layer0_out[2676] = x[102];
    assign layer0_out[2677] = x[251];
    assign layer0_out[2678] = ~x[138];
    assign layer0_out[2679] = ~(x[9] ^ x[14]);
    assign layer0_out[2680] = 1'b0;
    assign layer0_out[2681] = x[264] ^ x[278];
    assign layer0_out[2682] = ~x[32] | x[17];
    assign layer0_out[2683] = ~x[187];
    assign layer0_out[2684] = ~x[325];
    assign layer0_out[2685] = ~x[88] | x[75];
    assign layer0_out[2686] = x[160];
    assign layer0_out[2687] = x[231];
    assign layer0_out[2688] = ~(x[298] & x[307]);
    assign layer0_out[2689] = x[328] | x[335];
    assign layer0_out[2690] = x[359] ^ x[376];
    assign layer0_out[2691] = ~x[117] | x[113];
    assign layer0_out[2692] = ~x[156];
    assign layer0_out[2693] = x[21];
    assign layer0_out[2694] = x[26];
    assign layer0_out[2695] = ~x[275] | x[282];
    assign layer0_out[2696] = x[381] ^ x[393];
    assign layer0_out[2697] = ~(x[57] | x[68]);
    assign layer0_out[2698] = ~(x[363] ^ x[382]);
    assign layer0_out[2699] = ~x[66];
    assign layer0_out[2700] = x[231] | x[240];
    assign layer0_out[2701] = x[85] & ~x[98];
    assign layer0_out[2702] = x[365];
    assign layer0_out[2703] = ~x[212];
    assign layer0_out[2704] = ~(x[61] | x[80]);
    assign layer0_out[2705] = x[229];
    assign layer0_out[2706] = x[131];
    assign layer0_out[2707] = ~(x[52] | x[72]);
    assign layer0_out[2708] = ~(x[372] | x[387]);
    assign layer0_out[2709] = ~(x[254] & x[273]);
    assign layer0_out[2710] = ~(x[201] | x[222]);
    assign layer0_out[2711] = 1'b0;
    assign layer0_out[2712] = ~(x[40] | x[60]);
    assign layer0_out[2713] = x[302] & x[316];
    assign layer0_out[2714] = x[225];
    assign layer0_out[2715] = ~(x[379] & x[380]);
    assign layer0_out[2716] = ~(x[197] | x[201]);
    assign layer0_out[2717] = x[166];
    assign layer0_out[2718] = ~(x[280] | x[281]);
    assign layer0_out[2719] = ~(x[357] | x[359]);
    assign layer0_out[2720] = ~(x[118] | x[136]);
    assign layer0_out[2721] = ~(x[369] | x[385]);
    assign layer0_out[2722] = 1'b1;
    assign layer0_out[2723] = x[350] & x[352];
    assign layer0_out[2724] = x[386] ^ x[391];
    assign layer0_out[2725] = x[75] | x[81];
    assign layer0_out[2726] = ~(x[287] ^ x[301]);
    assign layer0_out[2727] = ~(x[228] | x[230]);
    assign layer0_out[2728] = 1'b0;
    assign layer0_out[2729] = ~(x[221] ^ x[235]);
    assign layer0_out[2730] = ~(x[227] | x[245]);
    assign layer0_out[2731] = ~(x[225] | x[227]);
    assign layer0_out[2732] = ~(x[95] ^ x[111]);
    assign layer0_out[2733] = ~x[301] | x[298];
    assign layer0_out[2734] = ~x[300] | x[310];
    assign layer0_out[2735] = ~x[246];
    assign layer0_out[2736] = ~x[277];
    assign layer0_out[2737] = x[257] ^ x[272];
    assign layer0_out[2738] = x[38];
    assign layer0_out[2739] = ~x[293];
    assign layer0_out[2740] = ~x[364];
    assign layer0_out[2741] = ~x[272];
    assign layer0_out[2742] = ~x[249];
    assign layer0_out[2743] = x[371] & ~x[359];
    assign layer0_out[2744] = x[231] & x[246];
    assign layer0_out[2745] = ~(x[239] ^ x[256]);
    assign layer0_out[2746] = x[199];
    assign layer0_out[2747] = x[152];
    assign layer0_out[2748] = x[336];
    assign layer0_out[2749] = ~(x[14] | x[16]);
    assign layer0_out[2750] = ~x[169];
    assign layer0_out[2751] = ~x[95];
    assign layer0_out[2752] = x[88];
    assign layer0_out[2753] = ~(x[18] | x[19]);
    assign layer0_out[2754] = ~(x[44] | x[63]);
    assign layer0_out[2755] = x[270] & x[284];
    assign layer0_out[2756] = ~x[287];
    assign layer0_out[2757] = x[77];
    assign layer0_out[2758] = x[291];
    assign layer0_out[2759] = ~x[19];
    assign layer0_out[2760] = ~x[76];
    assign layer0_out[2761] = x[331];
    assign layer0_out[2762] = x[310] | x[316];
    assign layer0_out[2763] = ~(x[128] | x[147]);
    assign layer0_out[2764] = x[50] ^ x[66];
    assign layer0_out[2765] = x[154] ^ x[158];
    assign layer0_out[2766] = ~(x[5] | x[22]);
    assign layer0_out[2767] = ~x[307];
    assign layer0_out[2768] = ~(x[193] | x[208]);
    assign layer0_out[2769] = ~x[107] | x[111];
    assign layer0_out[2770] = x[180];
    assign layer0_out[2771] = x[197] & ~x[212];
    assign layer0_out[2772] = x[127];
    assign layer0_out[2773] = x[146] | x[156];
    assign layer0_out[2774] = x[366] | x[375];
    assign layer0_out[2775] = x[333] ^ x[346];
    assign layer0_out[2776] = x[324] | x[337];
    assign layer0_out[2777] = x[248];
    assign layer0_out[2778] = x[298] ^ x[306];
    assign layer0_out[2779] = x[117] | x[118];
    assign layer0_out[2780] = ~(x[320] | x[340]);
    assign layer0_out[2781] = x[364] | x[376];
    assign layer0_out[2782] = x[223] ^ x[232];
    assign layer0_out[2783] = ~(x[232] | x[237]);
    assign layer0_out[2784] = 1'b0;
    assign layer0_out[2785] = x[139] | x[140];
    assign layer0_out[2786] = 1'b1;
    assign layer0_out[2787] = ~x[370];
    assign layer0_out[2788] = ~x[54] | x[55];
    assign layer0_out[2789] = x[150] | x[152];
    assign layer0_out[2790] = x[262] | x[268];
    assign layer0_out[2791] = 1'b0;
    assign layer0_out[2792] = ~(x[210] | x[230]);
    assign layer0_out[2793] = x[287];
    assign layer0_out[2794] = x[210] | x[217];
    assign layer0_out[2795] = ~(x[171] ^ x[174]);
    assign layer0_out[2796] = x[46] & ~x[34];
    assign layer0_out[2797] = x[368] ^ x[374];
    assign layer0_out[2798] = x[121] | x[141];
    assign layer0_out[2799] = x[294] | x[296];
    assign layer0_out[2800] = x[327] & ~x[310];
    assign layer0_out[2801] = ~x[67] | x[60];
    assign layer0_out[2802] = ~x[248];
    assign layer0_out[2803] = ~(x[188] | x[208]);
    assign layer0_out[2804] = 1'b1;
    assign layer0_out[2805] = x[104] | x[125];
    assign layer0_out[2806] = x[196] & x[205];
    assign layer0_out[2807] = ~x[164];
    assign layer0_out[2808] = x[275];
    assign layer0_out[2809] = x[10] & ~x[19];
    assign layer0_out[2810] = x[37] ^ x[57];
    assign layer0_out[2811] = ~(x[129] | x[130]);
    assign layer0_out[2812] = ~(x[290] & x[294]);
    assign layer0_out[2813] = x[166] | x[182];
    assign layer0_out[2814] = ~(x[24] | x[32]);
    assign layer0_out[2815] = ~x[196];
    assign layer0_out[2816] = ~x[83] | x[67];
    assign layer0_out[2817] = x[39];
    assign layer0_out[2818] = ~(x[345] | x[358]);
    assign layer0_out[2819] = ~(x[346] ^ x[359]);
    assign layer0_out[2820] = 1'b0;
    assign layer0_out[2821] = ~x[288] | x[281];
    assign layer0_out[2822] = x[74];
    assign layer0_out[2823] = ~x[131] | x[148];
    assign layer0_out[2824] = x[267] & ~x[259];
    assign layer0_out[2825] = ~(x[293] & x[308]);
    assign layer0_out[2826] = ~(x[283] | x[302]);
    assign layer0_out[2827] = ~(x[361] ^ x[362]);
    assign layer0_out[2828] = x[381];
    assign layer0_out[2829] = 1'b0;
    assign layer0_out[2830] = x[36] ^ x[48];
    assign layer0_out[2831] = ~(x[51] ^ x[54]);
    assign layer0_out[2832] = ~x[316] | x[328];
    assign layer0_out[2833] = ~x[223];
    assign layer0_out[2834] = ~x[204];
    assign layer0_out[2835] = x[91] & ~x[83];
    assign layer0_out[2836] = x[50] ^ x[64];
    assign layer0_out[2837] = ~(x[200] | x[217]);
    assign layer0_out[2838] = x[362] & ~x[351];
    assign layer0_out[2839] = 1'b1;
    assign layer0_out[2840] = x[97];
    assign layer0_out[2841] = x[256] | x[276];
    assign layer0_out[2842] = ~(x[368] | x[383]);
    assign layer0_out[2843] = x[208];
    assign layer0_out[2844] = x[92];
    assign layer0_out[2845] = x[294] & x[310];
    assign layer0_out[2846] = x[113];
    assign layer0_out[2847] = ~x[165];
    assign layer0_out[2848] = ~x[75];
    assign layer0_out[2849] = x[109] | x[117];
    assign layer0_out[2850] = x[230] & x[235];
    assign layer0_out[2851] = x[85] ^ x[106];
    assign layer0_out[2852] = x[104] & x[110];
    assign layer0_out[2853] = x[241] | x[243];
    assign layer0_out[2854] = x[192] & ~x[188];
    assign layer0_out[2855] = ~x[302];
    assign layer0_out[2856] = ~(x[122] & x[134]);
    assign layer0_out[2857] = ~x[15];
    assign layer0_out[2858] = ~x[365];
    assign layer0_out[2859] = ~x[374] | x[393];
    assign layer0_out[2860] = ~x[152];
    assign layer0_out[2861] = ~x[271];
    assign layer0_out[2862] = ~(x[82] ^ x[95]);
    assign layer0_out[2863] = x[369];
    assign layer0_out[2864] = x[135] & ~x[152];
    assign layer0_out[2865] = x[107] ^ x[123];
    assign layer0_out[2866] = 1'b1;
    assign layer0_out[2867] = ~x[334];
    assign layer0_out[2868] = x[65];
    assign layer0_out[2869] = x[330] | x[339];
    assign layer0_out[2870] = ~x[165];
    assign layer0_out[2871] = x[105] | x[120];
    assign layer0_out[2872] = ~(x[101] | x[114]);
    assign layer0_out[2873] = x[56];
    assign layer0_out[2874] = x[333] | x[335];
    assign layer0_out[2875] = x[33] & ~x[20];
    assign layer0_out[2876] = x[283] & ~x[276];
    assign layer0_out[2877] = ~x[73];
    assign layer0_out[2878] = ~(x[74] | x[89]);
    assign layer0_out[2879] = 1'b0;
    assign layer0_out[2880] = x[265];
    assign layer0_out[2881] = x[366] ^ x[369];
    assign layer0_out[2882] = x[303] | x[313];
    assign layer0_out[2883] = ~(x[33] | x[38]);
    assign layer0_out[2884] = x[200];
    assign layer0_out[2885] = x[304];
    assign layer0_out[2886] = ~(x[226] | x[232]);
    assign layer0_out[2887] = x[345] | x[364];
    assign layer0_out[2888] = x[221];
    assign layer0_out[2889] = ~x[168] | x[185];
    assign layer0_out[2890] = x[82] & ~x[73];
    assign layer0_out[2891] = x[16] & ~x[7];
    assign layer0_out[2892] = x[64] | x[85];
    assign layer0_out[2893] = x[221] & ~x[241];
    assign layer0_out[2894] = ~(x[7] | x[9]);
    assign layer0_out[2895] = ~(x[227] | x[237]);
    assign layer0_out[2896] = ~(x[40] | x[53]);
    assign layer0_out[2897] = ~(x[302] & x[322]);
    assign layer0_out[2898] = ~(x[72] | x[91]);
    assign layer0_out[2899] = ~x[297];
    assign layer0_out[2900] = x[15];
    assign layer0_out[2901] = ~(x[136] | x[156]);
    assign layer0_out[2902] = ~x[47];
    assign layer0_out[2903] = ~(x[140] | x[154]);
    assign layer0_out[2904] = ~(x[116] | x[119]);
    assign layer0_out[2905] = ~(x[337] | x[342]);
    assign layer0_out[2906] = ~(x[140] ^ x[158]);
    assign layer0_out[2907] = x[145] | x[158];
    assign layer0_out[2908] = ~(x[6] | x[15]);
    assign layer0_out[2909] = x[3] & x[8];
    assign layer0_out[2910] = ~(x[245] ^ x[255]);
    assign layer0_out[2911] = x[54];
    assign layer0_out[2912] = ~(x[152] | x[173]);
    assign layer0_out[2913] = ~x[274];
    assign layer0_out[2914] = x[274];
    assign layer0_out[2915] = x[51] & ~x[69];
    assign layer0_out[2916] = x[363] & ~x[367];
    assign layer0_out[2917] = ~(x[9] | x[30]);
    assign layer0_out[2918] = x[150] | x[170];
    assign layer0_out[2919] = ~x[319];
    assign layer0_out[2920] = x[299] & ~x[300];
    assign layer0_out[2921] = 1'b0;
    assign layer0_out[2922] = ~(x[107] ^ x[125]);
    assign layer0_out[2923] = ~(x[336] ^ x[345]);
    assign layer0_out[2924] = 1'b1;
    assign layer0_out[2925] = ~(x[259] ^ x[261]);
    assign layer0_out[2926] = ~(x[26] | x[33]);
    assign layer0_out[2927] = ~(x[201] | x[217]);
    assign layer0_out[2928] = ~x[92];
    assign layer0_out[2929] = ~(x[230] | x[248]);
    assign layer0_out[2930] = x[181] | x[188];
    assign layer0_out[2931] = ~x[370];
    assign layer0_out[2932] = x[165] & x[173];
    assign layer0_out[2933] = ~(x[77] & x[90]);
    assign layer0_out[2934] = x[346] | x[352];
    assign layer0_out[2935] = x[224] | x[231];
    assign layer0_out[2936] = ~x[266] | x[273];
    assign layer0_out[2937] = ~(x[62] & x[71]);
    assign layer0_out[2938] = 1'b0;
    assign layer0_out[2939] = 1'b1;
    assign layer0_out[2940] = ~x[369] | x[350];
    assign layer0_out[2941] = x[48] | x[60];
    assign layer0_out[2942] = x[335];
    assign layer0_out[2943] = 1'b1;
    assign layer0_out[2944] = ~x[219];
    assign layer0_out[2945] = x[15] & x[23];
    assign layer0_out[2946] = 1'b1;
    assign layer0_out[2947] = 1'b1;
    assign layer0_out[2948] = x[184] ^ x[200];
    assign layer0_out[2949] = ~x[74] | x[61];
    assign layer0_out[2950] = x[310] & ~x[314];
    assign layer0_out[2951] = x[232] | x[249];
    assign layer0_out[2952] = x[138];
    assign layer0_out[2953] = x[173];
    assign layer0_out[2954] = ~x[295] | x[301];
    assign layer0_out[2955] = x[28] & x[42];
    assign layer0_out[2956] = x[131] | x[134];
    assign layer0_out[2957] = 1'b1;
    assign layer0_out[2958] = x[386] & ~x[380];
    assign layer0_out[2959] = ~x[172];
    assign layer0_out[2960] = ~(x[192] | x[202]);
    assign layer0_out[2961] = x[179];
    assign layer0_out[2962] = ~x[248] | x[239];
    assign layer0_out[2963] = ~(x[255] | x[259]);
    assign layer0_out[2964] = x[170] ^ x[180];
    assign layer0_out[2965] = x[119] & ~x[98];
    assign layer0_out[2966] = x[168] | x[169];
    assign layer0_out[2967] = ~x[177] | x[164];
    assign layer0_out[2968] = ~x[270];
    assign layer0_out[2969] = x[310] & x[313];
    assign layer0_out[2970] = x[129] ^ x[136];
    assign layer0_out[2971] = x[223];
    assign layer0_out[2972] = ~x[106];
    assign layer0_out[2973] = x[29];
    assign layer0_out[2974] = x[368] & x[370];
    assign layer0_out[2975] = 1'b0;
    assign layer0_out[2976] = x[144] | x[145];
    assign layer0_out[2977] = ~(x[102] ^ x[106]);
    assign layer0_out[2978] = ~x[116];
    assign layer0_out[2979] = x[23];
    assign layer0_out[2980] = x[229];
    assign layer0_out[2981] = ~x[222] | x[211];
    assign layer0_out[2982] = ~(x[126] ^ x[143]);
    assign layer0_out[2983] = ~(x[145] | x[165]);
    assign layer0_out[2984] = 1'b1;
    assign layer0_out[2985] = ~x[25];
    assign layer0_out[2986] = x[220] & x[237];
    assign layer0_out[2987] = x[230] | x[231];
    assign layer0_out[2988] = ~(x[180] | x[197]);
    assign layer0_out[2989] = ~x[142] | x[132];
    assign layer0_out[2990] = ~(x[220] | x[235]);
    assign layer0_out[2991] = ~x[387];
    assign layer0_out[2992] = ~(x[327] | x[347]);
    assign layer0_out[2993] = ~(x[131] | x[150]);
    assign layer0_out[2994] = x[109];
    assign layer0_out[2995] = ~x[212];
    assign layer0_out[2996] = x[137] | x[139];
    assign layer0_out[2997] = x[127] & ~x[107];
    assign layer0_out[2998] = ~x[285] | x[294];
    assign layer0_out[2999] = x[284] | x[303];
    assign layer0_out[3000] = x[220] & ~x[226];
    assign layer0_out[3001] = ~(x[229] | x[242]);
    assign layer0_out[3002] = 1'b1;
    assign layer0_out[3003] = x[41] & x[56];
    assign layer0_out[3004] = ~x[117];
    assign layer0_out[3005] = ~x[267];
    assign layer0_out[3006] = x[363] | x[365];
    assign layer0_out[3007] = x[221] | x[233];
    assign layer0_out[3008] = ~(x[217] & x[235]);
    assign layer0_out[3009] = ~(x[311] | x[314]);
    assign layer0_out[3010] = x[116];
    assign layer0_out[3011] = 1'b1;
    assign layer0_out[3012] = x[216] & ~x[223];
    assign layer0_out[3013] = x[115] ^ x[129];
    assign layer0_out[3014] = ~(x[99] | x[120]);
    assign layer0_out[3015] = x[365];
    assign layer0_out[3016] = 1'b0;
    assign layer0_out[3017] = x[292] ^ x[295];
    assign layer0_out[3018] = x[78] & ~x[62];
    assign layer0_out[3019] = x[231] & x[239];
    assign layer0_out[3020] = x[251];
    assign layer0_out[3021] = x[161];
    assign layer0_out[3022] = ~x[259] | x[276];
    assign layer0_out[3023] = x[150];
    assign layer0_out[3024] = ~x[290];
    assign layer0_out[3025] = ~x[151];
    assign layer0_out[3026] = ~x[143];
    assign layer0_out[3027] = x[291];
    assign layer0_out[3028] = ~x[313];
    assign layer0_out[3029] = 1'b1;
    assign layer0_out[3030] = x[371];
    assign layer0_out[3031] = x[216] | x[218];
    assign layer0_out[3032] = ~(x[238] ^ x[255]);
    assign layer0_out[3033] = ~x[109];
    assign layer0_out[3034] = ~x[286];
    assign layer0_out[3035] = x[169] | x[174];
    assign layer0_out[3036] = x[289];
    assign layer0_out[3037] = ~(x[263] | x[280]);
    assign layer0_out[3038] = ~x[128];
    assign layer0_out[3039] = x[81];
    assign layer0_out[3040] = ~x[68];
    assign layer0_out[3041] = x[16] & ~x[36];
    assign layer0_out[3042] = ~(x[299] | x[308]);
    assign layer0_out[3043] = ~(x[146] | x[162]);
    assign layer0_out[3044] = x[68] | x[83];
    assign layer0_out[3045] = ~x[27];
    assign layer0_out[3046] = x[91];
    assign layer0_out[3047] = x[340] | x[342];
    assign layer0_out[3048] = x[200] ^ x[221];
    assign layer0_out[3049] = x[284];
    assign layer0_out[3050] = x[370];
    assign layer0_out[3051] = x[376] & x[389];
    assign layer0_out[3052] = x[208] & ~x[198];
    assign layer0_out[3053] = x[71] & ~x[85];
    assign layer0_out[3054] = x[383];
    assign layer0_out[3055] = 1'b1;
    assign layer0_out[3056] = 1'b1;
    assign layer0_out[3057] = 1'b1;
    assign layer0_out[3058] = ~(x[203] | x[207]);
    assign layer0_out[3059] = ~x[119];
    assign layer0_out[3060] = x[161];
    assign layer0_out[3061] = x[14] & x[15];
    assign layer0_out[3062] = ~(x[182] | x[201]);
    assign layer0_out[3063] = 1'b1;
    assign layer0_out[3064] = ~(x[266] | x[280]);
    assign layer0_out[3065] = ~x[179] | x[194];
    assign layer0_out[3066] = x[361] | x[376];
    assign layer0_out[3067] = ~(x[304] ^ x[319]);
    assign layer0_out[3068] = x[141] | x[144];
    assign layer0_out[3069] = ~x[266] | x[277];
    assign layer0_out[3070] = x[50] ^ x[56];
    assign layer0_out[3071] = x[220] & ~x[227];
    assign layer0_out[3072] = ~(x[347] | x[353]);
    assign layer0_out[3073] = ~x[87];
    assign layer0_out[3074] = x[145] & x[160];
    assign layer0_out[3075] = x[100] ^ x[105];
    assign layer0_out[3076] = ~(x[42] | x[45]);
    assign layer0_out[3077] = ~(x[261] | x[279]);
    assign layer0_out[3078] = x[362] | x[375];
    assign layer0_out[3079] = x[231];
    assign layer0_out[3080] = x[340] & ~x[343];
    assign layer0_out[3081] = ~x[295];
    assign layer0_out[3082] = ~x[352];
    assign layer0_out[3083] = ~(x[351] | x[371]);
    assign layer0_out[3084] = ~x[8] | x[20];
    assign layer0_out[3085] = ~x[275];
    assign layer0_out[3086] = x[163] | x[180];
    assign layer0_out[3087] = ~(x[107] | x[113]);
    assign layer0_out[3088] = x[121] & ~x[134];
    assign layer0_out[3089] = ~(x[69] | x[70]);
    assign layer0_out[3090] = x[329];
    assign layer0_out[3091] = x[70] & x[87];
    assign layer0_out[3092] = x[358] & ~x[375];
    assign layer0_out[3093] = x[222];
    assign layer0_out[3094] = x[286];
    assign layer0_out[3095] = x[160] & ~x[149];
    assign layer0_out[3096] = x[166] | x[186];
    assign layer0_out[3097] = ~x[364] | x[354];
    assign layer0_out[3098] = ~(x[92] & x[112]);
    assign layer0_out[3099] = ~(x[246] | x[263]);
    assign layer0_out[3100] = ~x[191];
    assign layer0_out[3101] = x[13] | x[27];
    assign layer0_out[3102] = ~x[112];
    assign layer0_out[3103] = x[323] & ~x[330];
    assign layer0_out[3104] = x[225] & ~x[228];
    assign layer0_out[3105] = ~x[136] | x[144];
    assign layer0_out[3106] = x[340] & ~x[358];
    assign layer0_out[3107] = ~x[147] | x[155];
    assign layer0_out[3108] = ~x[338];
    assign layer0_out[3109] = ~(x[306] | x[324]);
    assign layer0_out[3110] = ~x[194];
    assign layer0_out[3111] = x[38];
    assign layer0_out[3112] = x[58];
    assign layer0_out[3113] = x[341] | x[360];
    assign layer0_out[3114] = x[284] ^ x[294];
    assign layer0_out[3115] = ~(x[332] | x[345]);
    assign layer0_out[3116] = ~x[248] | x[232];
    assign layer0_out[3117] = x[353] & x[356];
    assign layer0_out[3118] = x[137] & ~x[150];
    assign layer0_out[3119] = x[103] | x[116];
    assign layer0_out[3120] = x[89] | x[108];
    assign layer0_out[3121] = 1'b1;
    assign layer0_out[3122] = ~x[257] | x[261];
    assign layer0_out[3123] = x[183];
    assign layer0_out[3124] = x[17];
    assign layer0_out[3125] = x[114] | x[115];
    assign layer0_out[3126] = x[315] | x[326];
    assign layer0_out[3127] = x[191] | x[212];
    assign layer0_out[3128] = ~x[135];
    assign layer0_out[3129] = ~x[225];
    assign layer0_out[3130] = x[237] & ~x[251];
    assign layer0_out[3131] = x[234] ^ x[241];
    assign layer0_out[3132] = 1'b0;
    assign layer0_out[3133] = ~(x[122] & x[135]);
    assign layer0_out[3134] = ~(x[8] | x[27]);
    assign layer0_out[3135] = 1'b0;
    assign layer0_out[3136] = x[216];
    assign layer0_out[3137] = x[135] | x[155];
    assign layer0_out[3138] = x[374];
    assign layer0_out[3139] = ~x[250];
    assign layer0_out[3140] = ~(x[65] ^ x[85]);
    assign layer0_out[3141] = ~x[67] | x[87];
    assign layer0_out[3142] = x[239] ^ x[243];
    assign layer0_out[3143] = ~(x[266] ^ x[268]);
    assign layer0_out[3144] = x[214] | x[219];
    assign layer0_out[3145] = x[318];
    assign layer0_out[3146] = ~x[105];
    assign layer0_out[3147] = x[138] | x[141];
    assign layer0_out[3148] = x[164];
    assign layer0_out[3149] = ~(x[183] & x[204]);
    assign layer0_out[3150] = ~x[124];
    assign layer0_out[3151] = ~x[21];
    assign layer0_out[3152] = x[239] & ~x[253];
    assign layer0_out[3153] = ~(x[172] | x[175]);
    assign layer0_out[3154] = x[298] | x[310];
    assign layer0_out[3155] = x[328];
    assign layer0_out[3156] = x[286];
    assign layer0_out[3157] = x[241];
    assign layer0_out[3158] = ~(x[357] | x[371]);
    assign layer0_out[3159] = ~(x[162] | x[164]);
    assign layer0_out[3160] = x[368] | x[388];
    assign layer0_out[3161] = ~(x[216] | x[220]);
    assign layer0_out[3162] = x[132] | x[150];
    assign layer0_out[3163] = ~x[16];
    assign layer0_out[3164] = x[305] & ~x[300];
    assign layer0_out[3165] = 1'b0;
    assign layer0_out[3166] = ~x[67];
    assign layer0_out[3167] = x[307] ^ x[319];
    assign layer0_out[3168] = x[276] ^ x[282];
    assign layer0_out[3169] = x[317] | x[330];
    assign layer0_out[3170] = x[268];
    assign layer0_out[3171] = x[356] | x[359];
    assign layer0_out[3172] = ~x[14] | x[5];
    assign layer0_out[3173] = x[224] & ~x[241];
    assign layer0_out[3174] = ~x[107];
    assign layer0_out[3175] = ~x[48];
    assign layer0_out[3176] = ~x[378] | x[396];
    assign layer0_out[3177] = ~x[127];
    assign layer0_out[3178] = ~x[82] | x[69];
    assign layer0_out[3179] = x[98] & ~x[99];
    assign layer0_out[3180] = ~x[257];
    assign layer0_out[3181] = 1'b0;
    assign layer0_out[3182] = x[261] | x[267];
    assign layer0_out[3183] = x[349];
    assign layer0_out[3184] = ~(x[320] | x[328]);
    assign layer0_out[3185] = ~x[200];
    assign layer0_out[3186] = x[163];
    assign layer0_out[3187] = x[336] & ~x[353];
    assign layer0_out[3188] = ~x[94] | x[75];
    assign layer0_out[3189] = x[37] & ~x[25];
    assign layer0_out[3190] = 1'b0;
    assign layer0_out[3191] = ~(x[344] | x[347]);
    assign layer0_out[3192] = ~x[219];
    assign layer0_out[3193] = ~x[141] | x[158];
    assign layer0_out[3194] = x[316] & ~x[325];
    assign layer0_out[3195] = ~(x[275] | x[278]);
    assign layer0_out[3196] = ~(x[190] ^ x[204]);
    assign layer0_out[3197] = ~(x[41] | x[45]);
    assign layer0_out[3198] = x[296];
    assign layer0_out[3199] = x[15] & ~x[35];
    assign layer0_out[3200] = x[235] | x[238];
    assign layer0_out[3201] = x[219];
    assign layer0_out[3202] = x[193] | x[213];
    assign layer0_out[3203] = ~x[357] | x[342];
    assign layer0_out[3204] = x[289] ^ x[301];
    assign layer0_out[3205] = x[43] ^ x[45];
    assign layer0_out[3206] = x[214] ^ x[225];
    assign layer0_out[3207] = x[59] | x[79];
    assign layer0_out[3208] = ~x[314];
    assign layer0_out[3209] = 1'b1;
    assign layer0_out[3210] = x[368] | x[369];
    assign layer0_out[3211] = ~x[63] | x[66];
    assign layer0_out[3212] = x[46];
    assign layer0_out[3213] = ~x[57];
    assign layer0_out[3214] = ~x[175] | x[170];
    assign layer0_out[3215] = x[28] | x[43];
    assign layer0_out[3216] = x[64];
    assign layer0_out[3217] = ~x[130];
    assign layer0_out[3218] = ~x[391];
    assign layer0_out[3219] = ~(x[192] ^ x[197]);
    assign layer0_out[3220] = ~(x[166] & x[169]);
    assign layer0_out[3221] = x[375] ^ x[383];
    assign layer0_out[3222] = x[72] ^ x[89];
    assign layer0_out[3223] = ~x[347];
    assign layer0_out[3224] = ~(x[385] | x[388]);
    assign layer0_out[3225] = x[102] & x[118];
    assign layer0_out[3226] = ~x[249] | x[260];
    assign layer0_out[3227] = ~(x[325] | x[345]);
    assign layer0_out[3228] = x[373] ^ x[391];
    assign layer0_out[3229] = 1'b0;
    assign layer0_out[3230] = x[69] & x[83];
    assign layer0_out[3231] = x[325];
    assign layer0_out[3232] = x[332];
    assign layer0_out[3233] = x[178] | x[183];
    assign layer0_out[3234] = ~(x[19] ^ x[33]);
    assign layer0_out[3235] = x[15];
    assign layer0_out[3236] = x[23] | x[34];
    assign layer0_out[3237] = ~(x[226] | x[239]);
    assign layer0_out[3238] = ~(x[160] ^ x[163]);
    assign layer0_out[3239] = x[295] | x[312];
    assign layer0_out[3240] = ~(x[142] | x[153]);
    assign layer0_out[3241] = x[314] & x[332];
    assign layer0_out[3242] = x[136] | x[146];
    assign layer0_out[3243] = x[195] ^ x[197];
    assign layer0_out[3244] = ~x[127] | x[117];
    assign layer0_out[3245] = ~x[374];
    assign layer0_out[3246] = ~x[214];
    assign layer0_out[3247] = ~x[33];
    assign layer0_out[3248] = ~x[293];
    assign layer0_out[3249] = ~(x[303] | x[305]);
    assign layer0_out[3250] = ~x[367];
    assign layer0_out[3251] = ~x[379];
    assign layer0_out[3252] = x[334] | x[336];
    assign layer0_out[3253] = x[268];
    assign layer0_out[3254] = ~(x[356] | x[372]);
    assign layer0_out[3255] = x[236];
    assign layer0_out[3256] = ~(x[246] | x[257]);
    assign layer0_out[3257] = x[39];
    assign layer0_out[3258] = ~x[328];
    assign layer0_out[3259] = x[227];
    assign layer0_out[3260] = x[199] & ~x[210];
    assign layer0_out[3261] = x[116] | x[118];
    assign layer0_out[3262] = x[132] | x[141];
    assign layer0_out[3263] = ~(x[101] ^ x[112]);
    assign layer0_out[3264] = ~x[107];
    assign layer0_out[3265] = x[358] | x[359];
    assign layer0_out[3266] = ~x[382];
    assign layer0_out[3267] = x[114];
    assign layer0_out[3268] = x[35] & x[54];
    assign layer0_out[3269] = x[237] | x[257];
    assign layer0_out[3270] = x[282] | x[300];
    assign layer0_out[3271] = x[38] | x[47];
    assign layer0_out[3272] = x[98] & ~x[81];
    assign layer0_out[3273] = x[179] & ~x[197];
    assign layer0_out[3274] = x[191];
    assign layer0_out[3275] = ~(x[215] ^ x[218]);
    assign layer0_out[3276] = x[386] | x[398];
    assign layer0_out[3277] = 1'b1;
    assign layer0_out[3278] = 1'b0;
    assign layer0_out[3279] = ~x[133];
    assign layer0_out[3280] = ~(x[273] & x[292]);
    assign layer0_out[3281] = x[265] ^ x[282];
    assign layer0_out[3282] = x[370] & x[389];
    assign layer0_out[3283] = ~(x[377] | x[384]);
    assign layer0_out[3284] = ~(x[313] & x[319]);
    assign layer0_out[3285] = ~(x[141] | x[161]);
    assign layer0_out[3286] = ~x[207] | x[215];
    assign layer0_out[3287] = x[167];
    assign layer0_out[3288] = x[62] & ~x[60];
    assign layer0_out[3289] = x[49];
    assign layer0_out[3290] = ~x[292];
    assign layer0_out[3291] = x[330] ^ x[345];
    assign layer0_out[3292] = ~x[192];
    assign layer0_out[3293] = 1'b0;
    assign layer0_out[3294] = ~x[119] | x[134];
    assign layer0_out[3295] = x[70] ^ x[86];
    assign layer0_out[3296] = x[207];
    assign layer0_out[3297] = x[173];
    assign layer0_out[3298] = ~x[371] | x[385];
    assign layer0_out[3299] = ~x[117] | x[103];
    assign layer0_out[3300] = ~(x[73] | x[93]);
    assign layer0_out[3301] = x[292];
    assign layer0_out[3302] = x[39] | x[53];
    assign layer0_out[3303] = ~x[94];
    assign layer0_out[3304] = 1'b0;
    assign layer0_out[3305] = ~(x[135] ^ x[139]);
    assign layer0_out[3306] = ~x[246];
    assign layer0_out[3307] = ~x[87];
    assign layer0_out[3308] = ~x[34];
    assign layer0_out[3309] = x[372] | x[377];
    assign layer0_out[3310] = ~(x[234] | x[238]);
    assign layer0_out[3311] = ~(x[278] ^ x[296]);
    assign layer0_out[3312] = x[90] | x[111];
    assign layer0_out[3313] = x[371] ^ x[387];
    assign layer0_out[3314] = x[5] & ~x[2];
    assign layer0_out[3315] = ~x[381] | x[367];
    assign layer0_out[3316] = x[323] & ~x[335];
    assign layer0_out[3317] = ~(x[30] | x[40]);
    assign layer0_out[3318] = ~(x[212] & x[229]);
    assign layer0_out[3319] = ~(x[163] | x[165]);
    assign layer0_out[3320] = ~x[103] | x[86];
    assign layer0_out[3321] = ~(x[299] ^ x[309]);
    assign layer0_out[3322] = x[18] | x[34];
    assign layer0_out[3323] = ~x[303];
    assign layer0_out[3324] = ~x[113];
    assign layer0_out[3325] = ~x[32];
    assign layer0_out[3326] = 1'b1;
    assign layer0_out[3327] = ~x[105];
    assign layer0_out[3328] = x[237] & ~x[224];
    assign layer0_out[3329] = ~x[115] | x[133];
    assign layer0_out[3330] = x[312] | x[314];
    assign layer0_out[3331] = ~x[49];
    assign layer0_out[3332] = x[112] & ~x[126];
    assign layer0_out[3333] = x[393] | x[397];
    assign layer0_out[3334] = x[106] ^ x[123];
    assign layer0_out[3335] = ~x[19] | x[38];
    assign layer0_out[3336] = x[69];
    assign layer0_out[3337] = x[270] ^ x[283];
    assign layer0_out[3338] = ~x[36];
    assign layer0_out[3339] = x[35] & x[51];
    assign layer0_out[3340] = ~x[291] | x[286];
    assign layer0_out[3341] = ~(x[69] ^ x[87]);
    assign layer0_out[3342] = x[348] ^ x[368];
    assign layer0_out[3343] = 1'b1;
    assign layer0_out[3344] = x[105];
    assign layer0_out[3345] = x[346];
    assign layer0_out[3346] = ~(x[0] | x[20]);
    assign layer0_out[3347] = x[130] ^ x[147];
    assign layer0_out[3348] = ~x[169] | x[180];
    assign layer0_out[3349] = ~(x[208] | x[225]);
    assign layer0_out[3350] = x[47] & x[52];
    assign layer0_out[3351] = ~(x[130] & x[132]);
    assign layer0_out[3352] = x[27];
    assign layer0_out[3353] = x[230] & ~x[241];
    assign layer0_out[3354] = x[399] & ~x[392];
    assign layer0_out[3355] = x[221];
    assign layer0_out[3356] = x[49] | x[61];
    assign layer0_out[3357] = x[328] | x[334];
    assign layer0_out[3358] = x[4] | x[11];
    assign layer0_out[3359] = ~(x[323] & x[333]);
    assign layer0_out[3360] = 1'b1;
    assign layer0_out[3361] = x[245] | x[263];
    assign layer0_out[3362] = x[273];
    assign layer0_out[3363] = 1'b0;
    assign layer0_out[3364] = ~(x[363] | x[369]);
    assign layer0_out[3365] = ~(x[181] | x[185]);
    assign layer0_out[3366] = 1'b0;
    assign layer0_out[3367] = ~x[176];
    assign layer0_out[3368] = x[270];
    assign layer0_out[3369] = ~(x[168] | x[189]);
    assign layer0_out[3370] = ~(x[338] | x[342]);
    assign layer0_out[3371] = x[96];
    assign layer0_out[3372] = ~x[323];
    assign layer0_out[3373] = x[354] ^ x[373];
    assign layer0_out[3374] = x[380];
    assign layer0_out[3375] = 1'b0;
    assign layer0_out[3376] = ~x[362];
    assign layer0_out[3377] = x[306];
    assign layer0_out[3378] = x[287];
    assign layer0_out[3379] = x[192];
    assign layer0_out[3380] = ~(x[176] | x[195]);
    assign layer0_out[3381] = x[363];
    assign layer0_out[3382] = ~(x[96] | x[98]);
    assign layer0_out[3383] = x[309];
    assign layer0_out[3384] = x[41] | x[49];
    assign layer0_out[3385] = ~(x[246] | x[249]);
    assign layer0_out[3386] = x[155];
    assign layer0_out[3387] = x[271] & ~x[282];
    assign layer0_out[3388] = ~x[165];
    assign layer0_out[3389] = x[338] ^ x[353];
    assign layer0_out[3390] = ~x[73];
    assign layer0_out[3391] = x[89];
    assign layer0_out[3392] = x[207] | x[214];
    assign layer0_out[3393] = ~x[357] | x[340];
    assign layer0_out[3394] = x[271] | x[279];
    assign layer0_out[3395] = ~x[208] | x[215];
    assign layer0_out[3396] = x[189];
    assign layer0_out[3397] = ~(x[119] | x[123]);
    assign layer0_out[3398] = ~x[191];
    assign layer0_out[3399] = ~x[235];
    assign layer0_out[3400] = x[134] & ~x[137];
    assign layer0_out[3401] = x[297] | x[299];
    assign layer0_out[3402] = x[60] | x[64];
    assign layer0_out[3403] = x[319] | x[335];
    assign layer0_out[3404] = ~(x[43] | x[57]);
    assign layer0_out[3405] = x[111] ^ x[131];
    assign layer0_out[3406] = ~x[237] | x[239];
    assign layer0_out[3407] = x[14] & x[26];
    assign layer0_out[3408] = x[23] | x[36];
    assign layer0_out[3409] = ~(x[224] | x[225]);
    assign layer0_out[3410] = x[348] & ~x[344];
    assign layer0_out[3411] = x[349] & ~x[361];
    assign layer0_out[3412] = ~(x[343] ^ x[360]);
    assign layer0_out[3413] = x[99] | x[108];
    assign layer0_out[3414] = x[17] | x[18];
    assign layer0_out[3415] = 1'b1;
    assign layer0_out[3416] = ~x[14] | x[23];
    assign layer0_out[3417] = ~x[172] | x[168];
    assign layer0_out[3418] = x[318] | x[331];
    assign layer0_out[3419] = ~x[134];
    assign layer0_out[3420] = x[110] | x[119];
    assign layer0_out[3421] = ~x[37];
    assign layer0_out[3422] = ~x[84];
    assign layer0_out[3423] = ~(x[145] ^ x[148]);
    assign layer0_out[3424] = x[5] ^ x[21];
    assign layer0_out[3425] = ~(x[17] | x[20]);
    assign layer0_out[3426] = ~(x[9] | x[29]);
    assign layer0_out[3427] = x[9] & ~x[1];
    assign layer0_out[3428] = x[148] & ~x[151];
    assign layer0_out[3429] = x[345] ^ x[361];
    assign layer0_out[3430] = ~x[94];
    assign layer0_out[3431] = ~(x[206] | x[223]);
    assign layer0_out[3432] = ~x[109] | x[119];
    assign layer0_out[3433] = ~(x[185] ^ x[204]);
    assign layer0_out[3434] = x[42];
    assign layer0_out[3435] = ~(x[64] | x[76]);
    assign layer0_out[3436] = x[373];
    assign layer0_out[3437] = ~x[283] | x[295];
    assign layer0_out[3438] = ~x[175];
    assign layer0_out[3439] = 1'b0;
    assign layer0_out[3440] = ~(x[67] | x[80]);
    assign layer0_out[3441] = x[88];
    assign layer0_out[3442] = ~(x[283] | x[290]);
    assign layer0_out[3443] = x[335];
    assign layer0_out[3444] = ~x[296];
    assign layer0_out[3445] = x[234];
    assign layer0_out[3446] = ~(x[67] | x[77]);
    assign layer0_out[3447] = x[120] | x[135];
    assign layer0_out[3448] = ~(x[277] ^ x[290]);
    assign layer0_out[3449] = x[11];
    assign layer0_out[3450] = ~(x[154] ^ x[171]);
    assign layer0_out[3451] = ~(x[49] ^ x[60]);
    assign layer0_out[3452] = ~(x[265] | x[279]);
    assign layer0_out[3453] = ~x[116];
    assign layer0_out[3454] = x[93] | x[103];
    assign layer0_out[3455] = ~(x[163] | x[182]);
    assign layer0_out[3456] = x[35];
    assign layer0_out[3457] = x[327] & x[330];
    assign layer0_out[3458] = ~(x[175] & x[177]);
    assign layer0_out[3459] = x[241] & ~x[245];
    assign layer0_out[3460] = ~x[8];
    assign layer0_out[3461] = x[49];
    assign layer0_out[3462] = ~x[308] | x[304];
    assign layer0_out[3463] = x[301] & ~x[293];
    assign layer0_out[3464] = x[174] | x[177];
    assign layer0_out[3465] = 1'b1;
    assign layer0_out[3466] = x[192];
    assign layer0_out[3467] = x[390] & ~x[383];
    assign layer0_out[3468] = 1'b1;
    assign layer0_out[3469] = x[180];
    assign layer0_out[3470] = x[38] & ~x[20];
    assign layer0_out[3471] = ~x[138];
    assign layer0_out[3472] = x[55];
    assign layer0_out[3473] = x[17] ^ x[24];
    assign layer0_out[3474] = ~(x[76] | x[94]);
    assign layer0_out[3475] = x[132] | x[139];
    assign layer0_out[3476] = x[60] | x[80];
    assign layer0_out[3477] = ~(x[196] | x[214]);
    assign layer0_out[3478] = 1'b1;
    assign layer0_out[3479] = x[385] | x[390];
    assign layer0_out[3480] = x[244] & x[256];
    assign layer0_out[3481] = ~x[83] | x[64];
    assign layer0_out[3482] = x[235] & ~x[251];
    assign layer0_out[3483] = x[197];
    assign layer0_out[3484] = x[55];
    assign layer0_out[3485] = x[6] & ~x[13];
    assign layer0_out[3486] = x[61];
    assign layer0_out[3487] = 1'b0;
    assign layer0_out[3488] = x[215] | x[217];
    assign layer0_out[3489] = ~(x[83] ^ x[89]);
    assign layer0_out[3490] = x[315] | x[316];
    assign layer0_out[3491] = ~(x[378] | x[397]);
    assign layer0_out[3492] = x[41] ^ x[50];
    assign layer0_out[3493] = ~x[224] | x[226];
    assign layer0_out[3494] = ~x[374];
    assign layer0_out[3495] = ~x[68];
    assign layer0_out[3496] = x[169] | x[190];
    assign layer0_out[3497] = ~x[377];
    assign layer0_out[3498] = ~x[37] | x[23];
    assign layer0_out[3499] = ~(x[287] & x[292]);
    assign layer0_out[3500] = ~(x[71] ^ x[86]);
    assign layer0_out[3501] = ~(x[279] ^ x[281]);
    assign layer0_out[3502] = ~(x[125] ^ x[142]);
    assign layer0_out[3503] = ~x[106] | x[119];
    assign layer0_out[3504] = x[217] & ~x[221];
    assign layer0_out[3505] = ~(x[99] | x[110]);
    assign layer0_out[3506] = x[352] ^ x[364];
    assign layer0_out[3507] = ~x[295] | x[287];
    assign layer0_out[3508] = ~x[85] | x[94];
    assign layer0_out[3509] = x[269] & ~x[277];
    assign layer0_out[3510] = x[190];
    assign layer0_out[3511] = ~(x[233] | x[253]);
    assign layer0_out[3512] = ~(x[346] | x[361]);
    assign layer0_out[3513] = ~(x[255] ^ x[260]);
    assign layer0_out[3514] = ~x[27];
    assign layer0_out[3515] = x[81] ^ x[95];
    assign layer0_out[3516] = x[23] | x[40];
    assign layer0_out[3517] = ~x[267] | x[278];
    assign layer0_out[3518] = x[358] & ~x[349];
    assign layer0_out[3519] = x[91];
    assign layer0_out[3520] = ~x[172] | x[188];
    assign layer0_out[3521] = ~(x[222] | x[236]);
    assign layer0_out[3522] = x[167] ^ x[184];
    assign layer0_out[3523] = ~x[9] | x[8];
    assign layer0_out[3524] = x[368] & ~x[373];
    assign layer0_out[3525] = x[179] | x[182];
    assign layer0_out[3526] = x[114] & ~x[93];
    assign layer0_out[3527] = x[175] | x[193];
    assign layer0_out[3528] = x[191];
    assign layer0_out[3529] = x[111] & x[130];
    assign layer0_out[3530] = x[121] & ~x[142];
    assign layer0_out[3531] = ~x[73] | x[85];
    assign layer0_out[3532] = ~x[230];
    assign layer0_out[3533] = x[273] ^ x[276];
    assign layer0_out[3534] = ~(x[47] & x[48]);
    assign layer0_out[3535] = ~x[283];
    assign layer0_out[3536] = x[361] ^ x[374];
    assign layer0_out[3537] = x[70];
    assign layer0_out[3538] = 1'b1;
    assign layer0_out[3539] = ~x[368];
    assign layer0_out[3540] = x[94] & x[113];
    assign layer0_out[3541] = ~x[68];
    assign layer0_out[3542] = ~(x[345] | x[350]);
    assign layer0_out[3543] = ~(x[308] | x[313]);
    assign layer0_out[3544] = 1'b1;
    assign layer0_out[3545] = ~x[94] | x[73];
    assign layer0_out[3546] = x[43] & ~x[44];
    assign layer0_out[3547] = ~x[172];
    assign layer0_out[3548] = x[137];
    assign layer0_out[3549] = ~x[53];
    assign layer0_out[3550] = ~(x[117] | x[131]);
    assign layer0_out[3551] = ~(x[72] ^ x[76]);
    assign layer0_out[3552] = x[128] & x[137];
    assign layer0_out[3553] = ~(x[6] | x[24]);
    assign layer0_out[3554] = 1'b1;
    assign layer0_out[3555] = ~x[217];
    assign layer0_out[3556] = ~x[86] | x[92];
    assign layer0_out[3557] = x[197] & x[207];
    assign layer0_out[3558] = ~(x[374] | x[394]);
    assign layer0_out[3559] = x[386] | x[397];
    assign layer0_out[3560] = x[174] | x[175];
    assign layer0_out[3561] = x[260];
    assign layer0_out[3562] = ~(x[213] & x[224]);
    assign layer0_out[3563] = x[56] | x[72];
    assign layer0_out[3564] = x[60] & x[65];
    assign layer0_out[3565] = x[249] | x[262];
    assign layer0_out[3566] = x[198];
    assign layer0_out[3567] = x[340];
    assign layer0_out[3568] = x[253] | x[264];
    assign layer0_out[3569] = x[302] | x[306];
    assign layer0_out[3570] = x[169] ^ x[186];
    assign layer0_out[3571] = x[177];
    assign layer0_out[3572] = 1'b0;
    assign layer0_out[3573] = x[245] | x[250];
    assign layer0_out[3574] = ~x[179];
    assign layer0_out[3575] = x[36] ^ x[42];
    assign layer0_out[3576] = ~x[66] | x[53];
    assign layer0_out[3577] = x[99] ^ x[109];
    assign layer0_out[3578] = ~x[167] | x[187];
    assign layer0_out[3579] = 1'b0;
    assign layer0_out[3580] = ~x[89];
    assign layer0_out[3581] = x[393] & x[395];
    assign layer0_out[3582] = 1'b1;
    assign layer0_out[3583] = ~(x[327] ^ x[336]);
    assign layer0_out[3584] = x[258] | x[263];
    assign layer0_out[3585] = ~x[367];
    assign layer0_out[3586] = ~(x[204] & x[211]);
    assign layer0_out[3587] = ~x[40];
    assign layer0_out[3588] = ~x[195];
    assign layer0_out[3589] = x[385];
    assign layer0_out[3590] = ~x[307] | x[308];
    assign layer0_out[3591] = ~(x[290] | x[304]);
    assign layer0_out[3592] = 1'b1;
    assign layer0_out[3593] = 1'b0;
    assign layer0_out[3594] = x[70] & x[76];
    assign layer0_out[3595] = x[228] & x[238];
    assign layer0_out[3596] = ~(x[42] ^ x[46]);
    assign layer0_out[3597] = x[324] | x[332];
    assign layer0_out[3598] = x[236] & x[256];
    assign layer0_out[3599] = x[391];
    assign layer0_out[3600] = x[203] & x[223];
    assign layer0_out[3601] = 1'b0;
    assign layer0_out[3602] = x[24] | x[41];
    assign layer0_out[3603] = x[295] | x[296];
    assign layer0_out[3604] = x[79] & ~x[86];
    assign layer0_out[3605] = ~x[72] | x[51];
    assign layer0_out[3606] = x[243] ^ x[260];
    assign layer0_out[3607] = ~(x[304] & x[322]);
    assign layer0_out[3608] = ~(x[288] & x[291]);
    assign layer0_out[3609] = ~(x[79] & x[95]);
    assign layer0_out[3610] = x[356] & ~x[355];
    assign layer0_out[3611] = ~x[340] | x[324];
    assign layer0_out[3612] = x[282] | x[298];
    assign layer0_out[3613] = ~x[248] | x[262];
    assign layer0_out[3614] = 1'b0;
    assign layer0_out[3615] = ~(x[120] ^ x[130]);
    assign layer0_out[3616] = ~x[302];
    assign layer0_out[3617] = x[312] & ~x[322];
    assign layer0_out[3618] = x[218];
    assign layer0_out[3619] = ~(x[159] ^ x[164]);
    assign layer0_out[3620] = x[219] ^ x[238];
    assign layer0_out[3621] = ~x[61];
    assign layer0_out[3622] = ~(x[314] & x[329]);
    assign layer0_out[3623] = x[296] ^ x[299];
    assign layer0_out[3624] = x[190];
    assign layer0_out[3625] = x[347];
    assign layer0_out[3626] = x[367] & ~x[375];
    assign layer0_out[3627] = x[308];
    assign layer0_out[3628] = x[349];
    assign layer0_out[3629] = x[237];
    assign layer0_out[3630] = x[259] | x[277];
    assign layer0_out[3631] = ~x[245];
    assign layer0_out[3632] = x[367];
    assign layer0_out[3633] = x[136];
    assign layer0_out[3634] = x[179] ^ x[181];
    assign layer0_out[3635] = x[164];
    assign layer0_out[3636] = ~(x[325] | x[331]);
    assign layer0_out[3637] = x[87] ^ x[108];
    assign layer0_out[3638] = x[272];
    assign layer0_out[3639] = x[4] | x[24];
    assign layer0_out[3640] = x[61] ^ x[71];
    assign layer0_out[3641] = x[389];
    assign layer0_out[3642] = x[291] ^ x[308];
    assign layer0_out[3643] = x[166] | x[175];
    assign layer0_out[3644] = ~x[118];
    assign layer0_out[3645] = ~(x[2] | x[21]);
    assign layer0_out[3646] = x[375] | x[395];
    assign layer0_out[3647] = x[245] | x[249];
    assign layer0_out[3648] = ~(x[323] | x[324]);
    assign layer0_out[3649] = x[196] ^ x[209];
    assign layer0_out[3650] = ~x[381];
    assign layer0_out[3651] = x[333] | x[345];
    assign layer0_out[3652] = x[21] ^ x[29];
    assign layer0_out[3653] = ~x[223];
    assign layer0_out[3654] = ~(x[250] ^ x[270]);
    assign layer0_out[3655] = x[178];
    assign layer0_out[3656] = ~x[24];
    assign layer0_out[3657] = ~x[322] | x[319];
    assign layer0_out[3658] = x[24] | x[34];
    assign layer0_out[3659] = ~x[165] | x[161];
    assign layer0_out[3660] = x[176] & ~x[162];
    assign layer0_out[3661] = x[206] & x[224];
    assign layer0_out[3662] = x[125] & ~x[133];
    assign layer0_out[3663] = x[103] ^ x[120];
    assign layer0_out[3664] = x[243] | x[251];
    assign layer0_out[3665] = ~x[21] | x[34];
    assign layer0_out[3666] = ~x[112];
    assign layer0_out[3667] = x[190] & ~x[181];
    assign layer0_out[3668] = ~x[191] | x[206];
    assign layer0_out[3669] = ~(x[149] | x[167]);
    assign layer0_out[3670] = ~(x[173] ^ x[185]);
    assign layer0_out[3671] = ~x[275];
    assign layer0_out[3672] = x[210] & ~x[216];
    assign layer0_out[3673] = x[8] | x[11];
    assign layer0_out[3674] = 1'b1;
    assign layer0_out[3675] = ~(x[72] | x[73]);
    assign layer0_out[3676] = x[266];
    assign layer0_out[3677] = x[48];
    assign layer0_out[3678] = ~x[146] | x[140];
    assign layer0_out[3679] = x[335] & x[354];
    assign layer0_out[3680] = ~x[209] | x[210];
    assign layer0_out[3681] = x[288];
    assign layer0_out[3682] = x[176] | x[194];
    assign layer0_out[3683] = 1'b1;
    assign layer0_out[3684] = x[40] & ~x[48];
    assign layer0_out[3685] = ~x[305];
    assign layer0_out[3686] = x[283] | x[284];
    assign layer0_out[3687] = ~x[276] | x[266];
    assign layer0_out[3688] = ~(x[335] & x[352]);
    assign layer0_out[3689] = ~(x[64] | x[65]);
    assign layer0_out[3690] = x[151] & ~x[141];
    assign layer0_out[3691] = ~(x[311] ^ x[318]);
    assign layer0_out[3692] = x[367];
    assign layer0_out[3693] = 1'b1;
    assign layer0_out[3694] = x[338];
    assign layer0_out[3695] = x[166] ^ x[176];
    assign layer0_out[3696] = ~(x[346] | x[365]);
    assign layer0_out[3697] = ~x[370];
    assign layer0_out[3698] = x[79];
    assign layer0_out[3699] = ~x[64];
    assign layer0_out[3700] = 1'b1;
    assign layer0_out[3701] = x[81] & ~x[102];
    assign layer0_out[3702] = x[346] | x[347];
    assign layer0_out[3703] = ~x[48] | x[53];
    assign layer0_out[3704] = ~(x[62] ^ x[75]);
    assign layer0_out[3705] = x[202] & x[208];
    assign layer0_out[3706] = ~(x[178] ^ x[188]);
    assign layer0_out[3707] = x[294];
    assign layer0_out[3708] = x[24] | x[26];
    assign layer0_out[3709] = x[116] | x[133];
    assign layer0_out[3710] = 1'b1;
    assign layer0_out[3711] = ~x[266];
    assign layer0_out[3712] = x[376] | x[383];
    assign layer0_out[3713] = ~(x[125] ^ x[131]);
    assign layer0_out[3714] = x[201] | x[214];
    assign layer0_out[3715] = ~x[41];
    assign layer0_out[3716] = 1'b1;
    assign layer0_out[3717] = ~x[218];
    assign layer0_out[3718] = ~x[174];
    assign layer0_out[3719] = ~(x[260] | x[275]);
    assign layer0_out[3720] = 1'b0;
    assign layer0_out[3721] = x[88] | x[103];
    assign layer0_out[3722] = ~x[148];
    assign layer0_out[3723] = x[240] & ~x[244];
    assign layer0_out[3724] = ~(x[261] | x[262]);
    assign layer0_out[3725] = x[345] | x[354];
    assign layer0_out[3726] = ~x[364];
    assign layer0_out[3727] = x[321];
    assign layer0_out[3728] = x[112] | x[118];
    assign layer0_out[3729] = x[287] & ~x[306];
    assign layer0_out[3730] = ~x[340];
    assign layer0_out[3731] = x[328] & x[345];
    assign layer0_out[3732] = x[265] & ~x[275];
    assign layer0_out[3733] = ~(x[112] ^ x[119]);
    assign layer0_out[3734] = x[257];
    assign layer0_out[3735] = x[250];
    assign layer0_out[3736] = 1'b1;
    assign layer0_out[3737] = x[185];
    assign layer0_out[3738] = x[54] & x[74];
    assign layer0_out[3739] = x[290];
    assign layer0_out[3740] = ~(x[304] ^ x[315]);
    assign layer0_out[3741] = x[167];
    assign layer0_out[3742] = x[66] | x[77];
    assign layer0_out[3743] = x[363];
    assign layer0_out[3744] = x[255] ^ x[262];
    assign layer0_out[3745] = ~(x[11] & x[29]);
    assign layer0_out[3746] = x[16];
    assign layer0_out[3747] = ~(x[57] ^ x[78]);
    assign layer0_out[3748] = x[85] ^ x[86];
    assign layer0_out[3749] = x[167];
    assign layer0_out[3750] = ~(x[153] & x[168]);
    assign layer0_out[3751] = x[248];
    assign layer0_out[3752] = x[118];
    assign layer0_out[3753] = ~x[268] | x[272];
    assign layer0_out[3754] = 1'b1;
    assign layer0_out[3755] = ~(x[207] ^ x[223]);
    assign layer0_out[3756] = x[6] | x[8];
    assign layer0_out[3757] = x[0];
    assign layer0_out[3758] = x[174];
    assign layer0_out[3759] = ~x[222];
    assign layer0_out[3760] = x[134] | x[141];
    assign layer0_out[3761] = ~(x[40] | x[50]);
    assign layer0_out[3762] = x[91] & ~x[92];
    assign layer0_out[3763] = 1'b0;
    assign layer0_out[3764] = x[90];
    assign layer0_out[3765] = ~(x[113] | x[120]);
    assign layer0_out[3766] = x[73] & x[88];
    assign layer0_out[3767] = ~(x[247] | x[249]);
    assign layer0_out[3768] = ~(x[27] | x[47]);
    assign layer0_out[3769] = x[361] | x[378];
    assign layer0_out[3770] = ~(x[41] & x[58]);
    assign layer0_out[3771] = ~(x[252] & x[266]);
    assign layer0_out[3772] = x[7] & ~x[11];
    assign layer0_out[3773] = ~x[399];
    assign layer0_out[3774] = ~(x[154] & x[173]);
    assign layer0_out[3775] = x[25];
    assign layer0_out[3776] = ~(x[344] | x[346]);
    assign layer0_out[3777] = x[81] ^ x[97];
    assign layer0_out[3778] = x[184] & ~x[174];
    assign layer0_out[3779] = ~x[348] | x[332];
    assign layer0_out[3780] = x[259];
    assign layer0_out[3781] = x[145];
    assign layer0_out[3782] = ~(x[377] ^ x[388]);
    assign layer0_out[3783] = x[313] & ~x[330];
    assign layer0_out[3784] = x[307] ^ x[326];
    assign layer0_out[3785] = x[150] | x[153];
    assign layer0_out[3786] = ~x[24];
    assign layer0_out[3787] = ~(x[199] | x[203]);
    assign layer0_out[3788] = 1'b1;
    assign layer0_out[3789] = x[153];
    assign layer0_out[3790] = ~x[363];
    assign layer0_out[3791] = ~x[56];
    assign layer0_out[3792] = x[172];
    assign layer0_out[3793] = x[55];
    assign layer0_out[3794] = ~(x[180] & x[188]);
    assign layer0_out[3795] = x[300];
    assign layer0_out[3796] = ~(x[156] | x[177]);
    assign layer0_out[3797] = ~(x[375] & x[384]);
    assign layer0_out[3798] = x[297] ^ x[311];
    assign layer0_out[3799] = 1'b0;
    assign layer0_out[3800] = x[374] & x[383];
    assign layer0_out[3801] = x[46] | x[65];
    assign layer0_out[3802] = ~(x[227] & x[241]);
    assign layer0_out[3803] = x[69] ^ x[73];
    assign layer0_out[3804] = 1'b1;
    assign layer0_out[3805] = ~(x[141] ^ x[153]);
    assign layer0_out[3806] = ~(x[340] ^ x[347]);
    assign layer0_out[3807] = x[82];
    assign layer0_out[3808] = ~x[258] | x[267];
    assign layer0_out[3809] = ~(x[341] ^ x[358]);
    assign layer0_out[3810] = x[183] & ~x[195];
    assign layer0_out[3811] = ~(x[326] | x[341]);
    assign layer0_out[3812] = ~x[169] | x[179];
    assign layer0_out[3813] = x[278] & x[283];
    assign layer0_out[3814] = x[44];
    assign layer0_out[3815] = ~(x[239] | x[258]);
    assign layer0_out[3816] = ~(x[299] | x[319]);
    assign layer0_out[3817] = x[218];
    assign layer0_out[3818] = ~x[205];
    assign layer0_out[3819] = ~x[299];
    assign layer0_out[3820] = x[355] | x[358];
    assign layer0_out[3821] = ~x[9];
    assign layer0_out[3822] = ~x[160] | x[153];
    assign layer0_out[3823] = ~(x[83] & x[93]);
    assign layer0_out[3824] = x[83] ^ x[97];
    assign layer0_out[3825] = x[157] | x[159];
    assign layer0_out[3826] = 1'b1;
    assign layer0_out[3827] = x[185] | x[186];
    assign layer0_out[3828] = ~(x[378] | x[379]);
    assign layer0_out[3829] = x[317];
    assign layer0_out[3830] = ~x[340];
    assign layer0_out[3831] = ~(x[168] ^ x[186]);
    assign layer0_out[3832] = ~(x[262] | x[265]);
    assign layer0_out[3833] = ~(x[346] | x[366]);
    assign layer0_out[3834] = x[289] & ~x[276];
    assign layer0_out[3835] = x[260] | x[265];
    assign layer0_out[3836] = ~(x[57] | x[76]);
    assign layer0_out[3837] = x[190];
    assign layer0_out[3838] = ~(x[308] | x[327]);
    assign layer0_out[3839] = x[40] | x[52];
    assign layer0_out[3840] = 1'b1;
    assign layer0_out[3841] = 1'b1;
    assign layer0_out[3842] = ~(x[39] | x[59]);
    assign layer0_out[3843] = x[298];
    assign layer0_out[3844] = x[251] | x[269];
    assign layer0_out[3845] = x[90] & x[92];
    assign layer0_out[3846] = x[88];
    assign layer0_out[3847] = ~(x[281] ^ x[295]);
    assign layer0_out[3848] = x[287];
    assign layer0_out[3849] = x[307] & ~x[311];
    assign layer0_out[3850] = x[283];
    assign layer0_out[3851] = x[74] & x[81];
    assign layer0_out[3852] = x[272] ^ x[290];
    assign layer0_out[3853] = x[385];
    assign layer0_out[3854] = ~(x[140] ^ x[150]);
    assign layer0_out[3855] = 1'b1;
    assign layer0_out[3856] = x[390] & ~x[388];
    assign layer0_out[3857] = x[240];
    assign layer0_out[3858] = ~(x[388] | x[395]);
    assign layer0_out[3859] = ~(x[248] | x[268]);
    assign layer0_out[3860] = ~x[292];
    assign layer0_out[3861] = x[84];
    assign layer0_out[3862] = x[359] ^ x[374];
    assign layer0_out[3863] = ~x[123];
    assign layer0_out[3864] = ~x[386];
    assign layer0_out[3865] = x[383] & ~x[373];
    assign layer0_out[3866] = ~x[267] | x[277];
    assign layer0_out[3867] = ~x[142];
    assign layer0_out[3868] = ~(x[306] | x[307]);
    assign layer0_out[3869] = ~x[183];
    assign layer0_out[3870] = x[216] | x[234];
    assign layer0_out[3871] = x[177];
    assign layer0_out[3872] = ~x[248];
    assign layer0_out[3873] = ~x[77];
    assign layer0_out[3874] = ~x[230];
    assign layer0_out[3875] = x[209] & ~x[220];
    assign layer0_out[3876] = x[125];
    assign layer0_out[3877] = x[123] | x[141];
    assign layer0_out[3878] = ~x[37];
    assign layer0_out[3879] = ~(x[266] ^ x[269]);
    assign layer0_out[3880] = ~x[205];
    assign layer0_out[3881] = x[275];
    assign layer0_out[3882] = ~(x[93] & x[101]);
    assign layer0_out[3883] = ~(x[184] | x[198]);
    assign layer0_out[3884] = x[178] & x[199];
    assign layer0_out[3885] = ~x[230];
    assign layer0_out[3886] = ~(x[338] ^ x[358]);
    assign layer0_out[3887] = x[130] | x[140];
    assign layer0_out[3888] = ~x[338];
    assign layer0_out[3889] = x[333];
    assign layer0_out[3890] = ~(x[223] | x[243]);
    assign layer0_out[3891] = 1'b0;
    assign layer0_out[3892] = ~(x[180] | x[190]);
    assign layer0_out[3893] = ~x[392];
    assign layer0_out[3894] = ~x[61];
    assign layer0_out[3895] = x[173];
    assign layer0_out[3896] = x[177] & ~x[198];
    assign layer0_out[3897] = x[122];
    assign layer0_out[3898] = 1'b1;
    assign layer0_out[3899] = ~x[226] | x[230];
    assign layer0_out[3900] = ~x[71] | x[87];
    assign layer0_out[3901] = ~(x[86] | x[105]);
    assign layer0_out[3902] = ~(x[252] ^ x[256]);
    assign layer0_out[3903] = x[85] | x[96];
    assign layer0_out[3904] = x[18] & ~x[1];
    assign layer0_out[3905] = ~(x[256] | x[257]);
    assign layer0_out[3906] = ~x[240] | x[247];
    assign layer0_out[3907] = x[33] ^ x[41];
    assign layer0_out[3908] = ~x[62];
    assign layer0_out[3909] = ~x[208] | x[211];
    assign layer0_out[3910] = x[223];
    assign layer0_out[3911] = ~(x[209] | x[226]);
    assign layer0_out[3912] = x[184] | x[203];
    assign layer0_out[3913] = ~(x[65] & x[70]);
    assign layer0_out[3914] = x[158] & ~x[163];
    assign layer0_out[3915] = x[98] & x[108];
    assign layer0_out[3916] = x[313] | x[321];
    assign layer0_out[3917] = ~x[231] | x[249];
    assign layer0_out[3918] = 1'b0;
    assign layer0_out[3919] = x[306];
    assign layer0_out[3920] = ~(x[238] | x[239]);
    assign layer0_out[3921] = ~(x[184] | x[199]);
    assign layer0_out[3922] = ~x[288] | x[272];
    assign layer0_out[3923] = x[282] | x[301];
    assign layer0_out[3924] = x[145] & ~x[139];
    assign layer0_out[3925] = x[320];
    assign layer0_out[3926] = x[127] & x[145];
    assign layer0_out[3927] = ~(x[23] ^ x[32]);
    assign layer0_out[3928] = x[347];
    assign layer0_out[3929] = x[126] | x[145];
    assign layer0_out[3930] = ~x[6] | x[0];
    assign layer0_out[3931] = ~x[291];
    assign layer0_out[3932] = x[3] | x[5];
    assign layer0_out[3933] = ~(x[340] & x[350]);
    assign layer0_out[3934] = ~x[281] | x[273];
    assign layer0_out[3935] = x[252] ^ x[261];
    assign layer0_out[3936] = ~(x[88] ^ x[104]);
    assign layer0_out[3937] = ~(x[167] | x[170]);
    assign layer0_out[3938] = ~x[303];
    assign layer0_out[3939] = x[241] ^ x[246];
    assign layer0_out[3940] = 1'b1;
    assign layer0_out[3941] = ~x[288];
    assign layer0_out[3942] = x[258] ^ x[275];
    assign layer0_out[3943] = x[288];
    assign layer0_out[3944] = x[84];
    assign layer0_out[3945] = ~x[343];
    assign layer0_out[3946] = x[47] | x[68];
    assign layer0_out[3947] = ~(x[355] ^ x[357]);
    assign layer0_out[3948] = x[95] | x[114];
    assign layer0_out[3949] = ~x[23];
    assign layer0_out[3950] = x[15] | x[34];
    assign layer0_out[3951] = x[90] & ~x[98];
    assign layer0_out[3952] = ~x[291] | x[290];
    assign layer0_out[3953] = ~x[44] | x[37];
    assign layer0_out[3954] = x[191] & x[210];
    assign layer0_out[3955] = x[337];
    assign layer0_out[3956] = x[154];
    assign layer0_out[3957] = x[237];
    assign layer0_out[3958] = x[91] & ~x[77];
    assign layer0_out[3959] = ~x[369];
    assign layer0_out[3960] = x[86] | x[91];
    assign layer0_out[3961] = ~x[250];
    assign layer0_out[3962] = x[291];
    assign layer0_out[3963] = ~x[290];
    assign layer0_out[3964] = 1'b0;
    assign layer0_out[3965] = ~x[152] | x[153];
    assign layer0_out[3966] = ~x[208];
    assign layer0_out[3967] = ~(x[201] | x[205]);
    assign layer0_out[3968] = x[267] | x[273];
    assign layer0_out[3969] = ~x[115];
    assign layer0_out[3970] = ~x[191] | x[202];
    assign layer0_out[3971] = x[262] | x[281];
    assign layer0_out[3972] = x[252] | x[271];
    assign layer0_out[3973] = ~(x[268] & x[273]);
    assign layer0_out[3974] = ~(x[388] | x[391]);
    assign layer0_out[3975] = x[341];
    assign layer0_out[3976] = x[63];
    assign layer0_out[3977] = ~x[264];
    assign layer0_out[3978] = ~(x[207] | x[226]);
    assign layer0_out[3979] = ~x[142] | x[156];
    assign layer0_out[3980] = x[390];
    assign layer0_out[3981] = x[17];
    assign layer0_out[3982] = x[33] | x[45];
    assign layer0_out[3983] = x[233];
    assign layer0_out[3984] = ~x[398] | x[378];
    assign layer0_out[3985] = ~(x[199] & x[207]);
    assign layer0_out[3986] = x[222] & ~x[209];
    assign layer0_out[3987] = ~(x[135] & x[149]);
    assign layer0_out[3988] = 1'b1;
    assign layer0_out[3989] = ~x[360];
    assign layer0_out[3990] = x[173] & x[183];
    assign layer0_out[3991] = x[298];
    assign layer0_out[3992] = 1'b1;
    assign layer0_out[3993] = x[147] ^ x[161];
    assign layer0_out[3994] = ~x[348];
    assign layer0_out[3995] = ~(x[301] | x[305]);
    assign layer0_out[3996] = x[40] & x[54];
    assign layer0_out[3997] = ~x[372] | x[370];
    assign layer0_out[3998] = x[197] | x[218];
    assign layer0_out[3999] = x[2];
    assign layer0_out[4000] = x[311] ^ x[324];
    assign layer0_out[4001] = x[218] | x[219];
    assign layer0_out[4002] = 1'b1;
    assign layer0_out[4003] = x[164] ^ x[181];
    assign layer0_out[4004] = x[294];
    assign layer0_out[4005] = x[331];
    assign layer0_out[4006] = x[370];
    assign layer0_out[4007] = ~(x[189] | x[194]);
    assign layer0_out[4008] = x[238];
    assign layer0_out[4009] = x[305];
    assign layer0_out[4010] = ~x[247];
    assign layer0_out[4011] = ~x[172] | x[162];
    assign layer0_out[4012] = ~x[14] | x[3];
    assign layer0_out[4013] = x[189] | x[208];
    assign layer0_out[4014] = x[393];
    assign layer0_out[4015] = x[93] ^ x[110];
    assign layer0_out[4016] = x[60] & ~x[44];
    assign layer0_out[4017] = ~x[117] | x[123];
    assign layer0_out[4018] = ~x[309];
    assign layer0_out[4019] = 1'b1;
    assign layer0_out[4020] = x[126];
    assign layer0_out[4021] = ~(x[201] | x[203]);
    assign layer0_out[4022] = 1'b0;
    assign layer0_out[4023] = 1'b1;
    assign layer0_out[4024] = ~(x[318] | x[327]);
    assign layer0_out[4025] = x[92] | x[93];
    assign layer0_out[4026] = ~(x[261] & x[273]);
    assign layer0_out[4027] = ~(x[99] | x[107]);
    assign layer0_out[4028] = ~(x[168] & x[183]);
    assign layer0_out[4029] = x[186] | x[201];
    assign layer0_out[4030] = ~x[249] | x[269];
    assign layer0_out[4031] = x[284];
    assign layer0_out[4032] = x[260];
    assign layer0_out[4033] = ~(x[202] | x[223]);
    assign layer0_out[4034] = x[42];
    assign layer0_out[4035] = x[266] & ~x[279];
    assign layer0_out[4036] = x[38] | x[50];
    assign layer0_out[4037] = x[1] | x[8];
    assign layer0_out[4038] = x[131] & ~x[113];
    assign layer0_out[4039] = 1'b1;
    assign layer0_out[4040] = ~x[0] | x[13];
    assign layer0_out[4041] = ~x[64];
    assign layer0_out[4042] = ~(x[38] & x[52]);
    assign layer0_out[4043] = x[386] & x[396];
    assign layer0_out[4044] = ~(x[332] ^ x[341]);
    assign layer0_out[4045] = x[337];
    assign layer0_out[4046] = ~x[62];
    assign layer0_out[4047] = x[65];
    assign layer0_out[4048] = ~(x[189] ^ x[204]);
    assign layer0_out[4049] = ~(x[379] | x[382]);
    assign layer0_out[4050] = x[294];
    assign layer0_out[4051] = ~x[296] | x[311];
    assign layer0_out[4052] = ~(x[257] | x[273]);
    assign layer0_out[4053] = x[152] | x[164];
    assign layer0_out[4054] = ~(x[330] & x[334]);
    assign layer0_out[4055] = x[37];
    assign layer0_out[4056] = ~x[35];
    assign layer0_out[4057] = ~x[328] | x[340];
    assign layer0_out[4058] = ~x[386] | x[392];
    assign layer0_out[4059] = 1'b1;
    assign layer0_out[4060] = x[99] ^ x[115];
    assign layer0_out[4061] = ~x[101];
    assign layer0_out[4062] = ~x[286] | x[277];
    assign layer0_out[4063] = x[265] & ~x[249];
    assign layer0_out[4064] = ~x[241];
    assign layer0_out[4065] = ~(x[36] | x[55]);
    assign layer0_out[4066] = 1'b1;
    assign layer0_out[4067] = x[396];
    assign layer0_out[4068] = ~x[380] | x[394];
    assign layer0_out[4069] = ~(x[184] | x[188]);
    assign layer0_out[4070] = 1'b1;
    assign layer0_out[4071] = x[35] & ~x[33];
    assign layer0_out[4072] = x[17] & ~x[0];
    assign layer0_out[4073] = ~(x[75] | x[76]);
    assign layer0_out[4074] = ~(x[376] | x[377]);
    assign layer0_out[4075] = x[56];
    assign layer0_out[4076] = ~x[129];
    assign layer0_out[4077] = x[243] ^ x[247];
    assign layer0_out[4078] = 1'b0;
    assign layer0_out[4079] = x[225] | x[232];
    assign layer0_out[4080] = x[63] & ~x[48];
    assign layer0_out[4081] = x[217];
    assign layer0_out[4082] = x[292];
    assign layer0_out[4083] = x[7] | x[10];
    assign layer0_out[4084] = 1'b0;
    assign layer0_out[4085] = ~x[67] | x[62];
    assign layer0_out[4086] = ~x[120];
    assign layer0_out[4087] = x[23];
    assign layer0_out[4088] = x[202] | x[222];
    assign layer0_out[4089] = x[243] & ~x[250];
    assign layer0_out[4090] = x[396] & ~x[382];
    assign layer0_out[4091] = ~x[317];
    assign layer0_out[4092] = x[222] ^ x[229];
    assign layer0_out[4093] = 1'b0;
    assign layer0_out[4094] = ~x[156] | x[167];
    assign layer0_out[4095] = x[316] ^ x[323];
    assign layer0_out[4096] = ~x[222];
    assign layer0_out[4097] = x[7] | x[12];
    assign layer0_out[4098] = x[161] ^ x[169];
    assign layer0_out[4099] = 1'b0;
    assign layer0_out[4100] = ~(x[139] ^ x[155]);
    assign layer0_out[4101] = x[125] & ~x[114];
    assign layer0_out[4102] = ~(x[3] | x[4]);
    assign layer0_out[4103] = x[272] ^ x[289];
    assign layer0_out[4104] = ~x[299];
    assign layer0_out[4105] = x[2];
    assign layer0_out[4106] = ~(x[208] & x[228]);
    assign layer0_out[4107] = ~x[24];
    assign layer0_out[4108] = ~x[26];
    assign layer0_out[4109] = ~x[282];
    assign layer0_out[4110] = 1'b0;
    assign layer0_out[4111] = 1'b0;
    assign layer0_out[4112] = x[131] ^ x[152];
    assign layer0_out[4113] = ~x[204];
    assign layer0_out[4114] = ~x[130];
    assign layer0_out[4115] = x[43];
    assign layer0_out[4116] = ~x[350];
    assign layer0_out[4117] = ~(x[102] | x[114]);
    assign layer0_out[4118] = x[308] ^ x[311];
    assign layer0_out[4119] = ~(x[74] ^ x[94]);
    assign layer0_out[4120] = x[219] & ~x[206];
    assign layer0_out[4121] = ~(x[262] | x[271]);
    assign layer0_out[4122] = x[388] | x[394];
    assign layer0_out[4123] = ~x[207];
    assign layer0_out[4124] = x[190] & x[193];
    assign layer0_out[4125] = x[288] | x[307];
    assign layer0_out[4126] = ~x[146];
    assign layer0_out[4127] = ~x[49];
    assign layer0_out[4128] = x[309] & x[326];
    assign layer0_out[4129] = ~x[69];
    assign layer0_out[4130] = ~x[202];
    assign layer0_out[4131] = ~x[119] | x[128];
    assign layer0_out[4132] = ~x[160] | x[147];
    assign layer0_out[4133] = ~x[242];
    assign layer0_out[4134] = x[307];
    assign layer0_out[4135] = x[106] | x[107];
    assign layer0_out[4136] = ~(x[55] | x[76]);
    assign layer0_out[4137] = ~(x[357] | x[377]);
    assign layer0_out[4138] = ~(x[18] ^ x[29]);
    assign layer0_out[4139] = x[179] & ~x[185];
    assign layer0_out[4140] = ~(x[97] & x[98]);
    assign layer0_out[4141] = ~(x[324] ^ x[326]);
    assign layer0_out[4142] = ~(x[14] | x[33]);
    assign layer0_out[4143] = x[196] | x[216];
    assign layer0_out[4144] = ~x[136] | x[141];
    assign layer0_out[4145] = ~(x[166] ^ x[181]);
    assign layer0_out[4146] = ~(x[59] ^ x[69]);
    assign layer0_out[4147] = x[20];
    assign layer0_out[4148] = 1'b0;
    assign layer0_out[4149] = ~(x[68] | x[82]);
    assign layer0_out[4150] = x[125];
    assign layer0_out[4151] = ~x[269];
    assign layer0_out[4152] = ~(x[46] | x[64]);
    assign layer0_out[4153] = ~x[252] | x[239];
    assign layer0_out[4154] = ~x[56];
    assign layer0_out[4155] = ~x[143];
    assign layer0_out[4156] = ~x[50];
    assign layer0_out[4157] = ~(x[146] ^ x[164]);
    assign layer0_out[4158] = x[148] ^ x[160];
    assign layer0_out[4159] = x[382];
    assign layer0_out[4160] = ~(x[94] ^ x[97]);
    assign layer0_out[4161] = ~x[150];
    assign layer0_out[4162] = ~(x[179] | x[198]);
    assign layer0_out[4163] = x[89] & ~x[81];
    assign layer0_out[4164] = ~x[372];
    assign layer0_out[4165] = x[345] | x[346];
    assign layer0_out[4166] = ~x[263];
    assign layer0_out[4167] = x[84];
    assign layer0_out[4168] = x[101];
    assign layer0_out[4169] = ~(x[193] & x[207]);
    assign layer0_out[4170] = x[240] & x[242];
    assign layer0_out[4171] = ~(x[175] ^ x[178]);
    assign layer0_out[4172] = x[25];
    assign layer0_out[4173] = x[42] & x[55];
    assign layer0_out[4174] = ~x[89];
    assign layer0_out[4175] = x[338];
    assign layer0_out[4176] = x[232];
    assign layer0_out[4177] = ~(x[85] & x[104]);
    assign layer0_out[4178] = ~x[210];
    assign layer0_out[4179] = x[2] | x[4];
    assign layer0_out[4180] = 1'b0;
    assign layer0_out[4181] = x[216] & x[229];
    assign layer0_out[4182] = x[25];
    assign layer0_out[4183] = ~(x[350] ^ x[359]);
    assign layer0_out[4184] = ~(x[22] ^ x[40]);
    assign layer0_out[4185] = x[90];
    assign layer0_out[4186] = 1'b1;
    assign layer0_out[4187] = ~x[310];
    assign layer0_out[4188] = ~x[140];
    assign layer0_out[4189] = 1'b0;
    assign layer0_out[4190] = ~(x[114] ^ x[117]);
    assign layer0_out[4191] = x[251] & ~x[242];
    assign layer0_out[4192] = 1'b0;
    assign layer0_out[4193] = x[230];
    assign layer0_out[4194] = 1'b0;
    assign layer0_out[4195] = x[83] | x[99];
    assign layer0_out[4196] = x[159] | x[174];
    assign layer0_out[4197] = x[323] & x[339];
    assign layer0_out[4198] = ~x[198];
    assign layer0_out[4199] = x[36] & x[53];
    assign layer0_out[4200] = ~x[132] | x[111];
    assign layer0_out[4201] = 1'b1;
    assign layer0_out[4202] = x[133] | x[139];
    assign layer0_out[4203] = x[350] & x[366];
    assign layer0_out[4204] = x[32] ^ x[47];
    assign layer0_out[4205] = x[324] ^ x[338];
    assign layer0_out[4206] = x[104] & ~x[124];
    assign layer0_out[4207] = 1'b1;
    assign layer0_out[4208] = x[162] & ~x[152];
    assign layer0_out[4209] = ~(x[171] | x[189]);
    assign layer0_out[4210] = x[356] | x[358];
    assign layer0_out[4211] = ~x[37] | x[36];
    assign layer0_out[4212] = x[148];
    assign layer0_out[4213] = x[46];
    assign layer0_out[4214] = ~x[36] | x[15];
    assign layer0_out[4215] = x[392];
    assign layer0_out[4216] = ~(x[229] | x[247]);
    assign layer0_out[4217] = x[271];
    assign layer0_out[4218] = x[213];
    assign layer0_out[4219] = x[2];
    assign layer0_out[4220] = x[347] & x[349];
    assign layer0_out[4221] = ~x[314] | x[304];
    assign layer0_out[4222] = ~(x[79] | x[93]);
    assign layer0_out[4223] = ~x[329];
    assign layer0_out[4224] = ~x[366] | x[362];
    assign layer0_out[4225] = ~(x[46] ^ x[66]);
    assign layer0_out[4226] = ~(x[59] ^ x[75]);
    assign layer0_out[4227] = ~x[204];
    assign layer0_out[4228] = ~(x[202] | x[221]);
    assign layer0_out[4229] = ~(x[122] | x[141]);
    assign layer0_out[4230] = x[291] & ~x[271];
    assign layer0_out[4231] = ~(x[115] & x[128]);
    assign layer0_out[4232] = ~(x[241] ^ x[247]);
    assign layer0_out[4233] = x[288] & ~x[303];
    assign layer0_out[4234] = ~(x[271] | x[277]);
    assign layer0_out[4235] = x[153] | x[154];
    assign layer0_out[4236] = ~x[260];
    assign layer0_out[4237] = x[73] & x[77];
    assign layer0_out[4238] = x[8];
    assign layer0_out[4239] = ~(x[276] & x[290]);
    assign layer0_out[4240] = ~(x[177] | x[194]);
    assign layer0_out[4241] = x[154] | x[160];
    assign layer0_out[4242] = x[256] & ~x[245];
    assign layer0_out[4243] = x[80];
    assign layer0_out[4244] = x[165] & ~x[169];
    assign layer0_out[4245] = x[247];
    assign layer0_out[4246] = ~(x[67] ^ x[85]);
    assign layer0_out[4247] = ~x[377];
    assign layer0_out[4248] = x[373] | x[377];
    assign layer0_out[4249] = x[101];
    assign layer0_out[4250] = x[158] & ~x[137];
    assign layer0_out[4251] = x[343] ^ x[348];
    assign layer0_out[4252] = ~(x[21] | x[27]);
    assign layer0_out[4253] = ~x[142];
    assign layer0_out[4254] = ~x[286] | x[292];
    assign layer0_out[4255] = ~(x[352] | x[366]);
    assign layer0_out[4256] = x[88] & ~x[69];
    assign layer0_out[4257] = ~(x[250] | x[268]);
    assign layer0_out[4258] = x[281] | x[297];
    assign layer0_out[4259] = ~x[29];
    assign layer0_out[4260] = x[94] ^ x[111];
    assign layer0_out[4261] = x[31] | x[44];
    assign layer0_out[4262] = x[145];
    assign layer0_out[4263] = x[239] ^ x[259];
    assign layer0_out[4264] = ~(x[182] & x[183]);
    assign layer0_out[4265] = x[392] & ~x[383];
    assign layer0_out[4266] = x[317] | x[336];
    assign layer0_out[4267] = ~(x[197] & x[210]);
    assign layer0_out[4268] = ~x[333];
    assign layer0_out[4269] = ~(x[322] ^ x[325]);
    assign layer0_out[4270] = x[125] | x[140];
    assign layer0_out[4271] = x[234] | x[253];
    assign layer0_out[4272] = x[289] | x[292];
    assign layer0_out[4273] = ~(x[134] | x[151]);
    assign layer0_out[4274] = ~x[257] | x[270];
    assign layer0_out[4275] = x[30] & ~x[36];
    assign layer0_out[4276] = x[109] & ~x[121];
    assign layer0_out[4277] = ~(x[326] | x[328]);
    assign layer0_out[4278] = ~(x[84] | x[96]);
    assign layer0_out[4279] = 1'b0;
    assign layer0_out[4280] = x[224];
    assign layer0_out[4281] = x[61] | x[65];
    assign layer0_out[4282] = x[136];
    assign layer0_out[4283] = x[169] & ~x[160];
    assign layer0_out[4284] = ~x[178] | x[193];
    assign layer0_out[4285] = x[174];
    assign layer0_out[4286] = ~x[340] | x[326];
    assign layer0_out[4287] = x[19] | x[20];
    assign layer0_out[4288] = ~(x[263] | x[268]);
    assign layer0_out[4289] = ~x[196];
    assign layer0_out[4290] = x[129] & ~x[124];
    assign layer0_out[4291] = x[199] & x[200];
    assign layer0_out[4292] = x[140] | x[144];
    assign layer0_out[4293] = x[93] & ~x[111];
    assign layer0_out[4294] = ~x[195];
    assign layer0_out[4295] = ~x[131];
    assign layer0_out[4296] = x[350] | x[370];
    assign layer0_out[4297] = ~(x[336] | x[343]);
    assign layer0_out[4298] = ~x[40];
    assign layer0_out[4299] = x[235];
    assign layer0_out[4300] = ~x[161];
    assign layer0_out[4301] = ~x[356];
    assign layer0_out[4302] = 1'b0;
    assign layer0_out[4303] = ~(x[6] ^ x[20]);
    assign layer0_out[4304] = x[139] & ~x[136];
    assign layer0_out[4305] = x[90] & ~x[79];
    assign layer0_out[4306] = ~(x[217] | x[226]);
    assign layer0_out[4307] = x[127];
    assign layer0_out[4308] = ~(x[66] ^ x[72]);
    assign layer0_out[4309] = ~(x[166] ^ x[173]);
    assign layer0_out[4310] = x[93] & ~x[97];
    assign layer0_out[4311] = ~x[71] | x[52];
    assign layer0_out[4312] = ~x[257];
    assign layer0_out[4313] = ~x[250];
    assign layer0_out[4314] = x[151] | x[160];
    assign layer0_out[4315] = x[46] | x[48];
    assign layer0_out[4316] = x[254] ^ x[258];
    assign layer0_out[4317] = x[379];
    assign layer0_out[4318] = ~(x[92] & x[105]);
    assign layer0_out[4319] = 1'b1;
    assign layer0_out[4320] = x[30] | x[31];
    assign layer0_out[4321] = x[94];
    assign layer0_out[4322] = ~x[201];
    assign layer0_out[4323] = x[161];
    assign layer0_out[4324] = ~(x[37] | x[55]);
    assign layer0_out[4325] = x[271];
    assign layer0_out[4326] = x[300] | x[315];
    assign layer0_out[4327] = x[178] & ~x[173];
    assign layer0_out[4328] = ~x[279] | x[295];
    assign layer0_out[4329] = x[10] ^ x[24];
    assign layer0_out[4330] = ~(x[289] ^ x[300]);
    assign layer0_out[4331] = x[348] & x[361];
    assign layer0_out[4332] = ~(x[266] | x[284]);
    assign layer0_out[4333] = ~x[162];
    assign layer0_out[4334] = x[311];
    assign layer0_out[4335] = x[336] & x[339];
    assign layer0_out[4336] = ~(x[153] | x[170]);
    assign layer0_out[4337] = ~(x[160] | x[162]);
    assign layer0_out[4338] = x[353] ^ x[355];
    assign layer0_out[4339] = x[193] & x[196];
    assign layer0_out[4340] = ~(x[44] ^ x[57]);
    assign layer0_out[4341] = ~(x[348] & x[353]);
    assign layer0_out[4342] = x[286];
    assign layer0_out[4343] = x[11];
    assign layer0_out[4344] = ~x[310] | x[330];
    assign layer0_out[4345] = x[303] & x[318];
    assign layer0_out[4346] = ~x[211];
    assign layer0_out[4347] = ~x[347];
    assign layer0_out[4348] = ~x[266];
    assign layer0_out[4349] = x[131] | x[140];
    assign layer0_out[4350] = ~x[332];
    assign layer0_out[4351] = x[178] | x[194];
    assign layer0_out[4352] = ~(x[213] & x[227]);
    assign layer0_out[4353] = ~x[260] | x[252];
    assign layer0_out[4354] = ~(x[5] | x[8]);
    assign layer0_out[4355] = ~x[378];
    assign layer0_out[4356] = x[62] ^ x[65];
    assign layer0_out[4357] = ~(x[68] | x[85]);
    assign layer0_out[4358] = x[337] | x[354];
    assign layer0_out[4359] = x[67] & ~x[52];
    assign layer0_out[4360] = ~(x[109] | x[110]);
    assign layer0_out[4361] = ~(x[29] & x[46]);
    assign layer0_out[4362] = ~(x[265] | x[269]);
    assign layer0_out[4363] = x[162] ^ x[165];
    assign layer0_out[4364] = x[236] & ~x[252];
    assign layer0_out[4365] = ~(x[343] | x[363]);
    assign layer0_out[4366] = ~x[228];
    assign layer0_out[4367] = ~x[264];
    assign layer0_out[4368] = ~x[346] | x[330];
    assign layer0_out[4369] = x[347];
    assign layer0_out[4370] = ~x[88];
    assign layer0_out[4371] = x[388];
    assign layer0_out[4372] = 1'b0;
    assign layer0_out[4373] = ~(x[380] | x[399]);
    assign layer0_out[4374] = ~x[124];
    assign layer0_out[4375] = x[198] | x[219];
    assign layer0_out[4376] = x[264] ^ x[280];
    assign layer0_out[4377] = ~(x[280] | x[282]);
    assign layer0_out[4378] = ~(x[181] ^ x[183]);
    assign layer0_out[4379] = ~x[384];
    assign layer0_out[4380] = x[29] | x[34];
    assign layer0_out[4381] = ~x[385] | x[399];
    assign layer0_out[4382] = ~(x[35] ^ x[50]);
    assign layer0_out[4383] = ~x[109];
    assign layer0_out[4384] = 1'b1;
    assign layer0_out[4385] = x[182] ^ x[186];
    assign layer0_out[4386] = x[223];
    assign layer0_out[4387] = x[270] | x[276];
    assign layer0_out[4388] = ~x[114] | x[106];
    assign layer0_out[4389] = x[397] | x[399];
    assign layer0_out[4390] = ~x[117];
    assign layer0_out[4391] = x[73] ^ x[76];
    assign layer0_out[4392] = ~x[51];
    assign layer0_out[4393] = ~x[167] | x[160];
    assign layer0_out[4394] = ~x[44] | x[55];
    assign layer0_out[4395] = ~x[106];
    assign layer0_out[4396] = x[175] ^ x[184];
    assign layer0_out[4397] = ~(x[361] & x[380]);
    assign layer0_out[4398] = x[228];
    assign layer0_out[4399] = ~x[269] | x[270];
    assign layer0_out[4400] = ~x[104];
    assign layer0_out[4401] = x[175];
    assign layer0_out[4402] = x[296];
    assign layer0_out[4403] = ~(x[212] | x[216]);
    assign layer0_out[4404] = x[260] & x[280];
    assign layer0_out[4405] = x[299] | x[305];
    assign layer0_out[4406] = x[117] & ~x[115];
    assign layer0_out[4407] = 1'b1;
    assign layer0_out[4408] = x[373];
    assign layer0_out[4409] = ~x[80] | x[93];
    assign layer0_out[4410] = x[1] & x[6];
    assign layer0_out[4411] = x[187];
    assign layer0_out[4412] = ~x[223] | x[228];
    assign layer0_out[4413] = x[213] | x[216];
    assign layer0_out[4414] = x[217];
    assign layer0_out[4415] = ~(x[107] ^ x[120]);
    assign layer0_out[4416] = ~x[387] | x[377];
    assign layer0_out[4417] = x[57] & ~x[46];
    assign layer0_out[4418] = 1'b0;
    assign layer0_out[4419] = x[25] | x[35];
    assign layer0_out[4420] = ~x[390] | x[379];
    assign layer0_out[4421] = ~x[330] | x[338];
    assign layer0_out[4422] = x[162];
    assign layer0_out[4423] = x[343] ^ x[355];
    assign layer0_out[4424] = x[344] & x[355];
    assign layer0_out[4425] = x[349];
    assign layer0_out[4426] = x[44] | x[62];
    assign layer0_out[4427] = x[351] & ~x[365];
    assign layer0_out[4428] = ~x[25] | x[19];
    assign layer0_out[4429] = x[73];
    assign layer0_out[4430] = ~x[371];
    assign layer0_out[4431] = x[89] ^ x[92];
    assign layer0_out[4432] = ~(x[211] & x[218]);
    assign layer0_out[4433] = ~x[166];
    assign layer0_out[4434] = ~x[375];
    assign layer0_out[4435] = 1'b1;
    assign layer0_out[4436] = ~(x[215] | x[222]);
    assign layer0_out[4437] = ~(x[195] | x[200]);
    assign layer0_out[4438] = ~x[293] | x[285];
    assign layer0_out[4439] = ~x[335] | x[318];
    assign layer0_out[4440] = ~(x[205] ^ x[221]);
    assign layer0_out[4441] = ~x[215];
    assign layer0_out[4442] = 1'b0;
    assign layer0_out[4443] = 1'b1;
    assign layer0_out[4444] = ~(x[235] ^ x[237]);
    assign layer0_out[4445] = x[96];
    assign layer0_out[4446] = ~x[36] | x[21];
    assign layer0_out[4447] = ~(x[98] | x[105]);
    assign layer0_out[4448] = x[314];
    assign layer0_out[4449] = x[196];
    assign layer0_out[4450] = ~(x[3] | x[23]);
    assign layer0_out[4451] = x[188] ^ x[202];
    assign layer0_out[4452] = x[328] & ~x[344];
    assign layer0_out[4453] = ~(x[123] ^ x[140]);
    assign layer0_out[4454] = ~(x[6] | x[25]);
    assign layer0_out[4455] = ~x[84];
    assign layer0_out[4456] = x[366];
    assign layer0_out[4457] = x[379];
    assign layer0_out[4458] = x[15] | x[17];
    assign layer0_out[4459] = x[96];
    assign layer0_out[4460] = x[250];
    assign layer0_out[4461] = x[121];
    assign layer0_out[4462] = ~(x[80] | x[100]);
    assign layer0_out[4463] = ~(x[227] ^ x[235]);
    assign layer0_out[4464] = x[86] ^ x[101];
    assign layer0_out[4465] = 1'b1;
    assign layer0_out[4466] = ~(x[228] & x[233]);
    assign layer0_out[4467] = x[94] | x[98];
    assign layer0_out[4468] = ~(x[315] & x[331]);
    assign layer0_out[4469] = x[334] & ~x[314];
    assign layer0_out[4470] = x[369] | x[383];
    assign layer0_out[4471] = ~(x[280] | x[291]);
    assign layer0_out[4472] = ~x[180] | x[159];
    assign layer0_out[4473] = x[210] & ~x[218];
    assign layer0_out[4474] = 1'b0;
    assign layer0_out[4475] = x[366] & ~x[377];
    assign layer0_out[4476] = ~x[260] | x[266];
    assign layer0_out[4477] = ~(x[323] & x[341]);
    assign layer0_out[4478] = ~(x[223] | x[227]);
    assign layer0_out[4479] = x[128];
    assign layer0_out[4480] = x[278] & ~x[292];
    assign layer0_out[4481] = x[214] ^ x[228];
    assign layer0_out[4482] = ~(x[41] | x[48]);
    assign layer0_out[4483] = x[122] & x[123];
    assign layer0_out[4484] = ~(x[208] & x[227]);
    assign layer0_out[4485] = x[204] | x[225];
    assign layer0_out[4486] = x[282] ^ x[295];
    assign layer0_out[4487] = ~x[135] | x[156];
    assign layer0_out[4488] = x[32] | x[53];
    assign layer0_out[4489] = ~(x[251] ^ x[266]);
    assign layer0_out[4490] = x[353] | x[368];
    assign layer0_out[4491] = x[32] | x[51];
    assign layer0_out[4492] = x[164] & ~x[145];
    assign layer0_out[4493] = x[22];
    assign layer0_out[4494] = x[240] & ~x[227];
    assign layer0_out[4495] = 1'b1;
    assign layer0_out[4496] = ~x[19];
    assign layer0_out[4497] = x[180];
    assign layer0_out[4498] = x[1] & ~x[10];
    assign layer0_out[4499] = x[168] | x[171];
    assign layer0_out[4500] = x[68] & x[70];
    assign layer0_out[4501] = x[230] & ~x[223];
    assign layer0_out[4502] = ~x[13] | x[1];
    assign layer0_out[4503] = x[181];
    assign layer0_out[4504] = x[118];
    assign layer0_out[4505] = x[13] & ~x[7];
    assign layer0_out[4506] = x[195] ^ x[216];
    assign layer0_out[4507] = x[30] & ~x[38];
    assign layer0_out[4508] = ~(x[141] | x[156]);
    assign layer0_out[4509] = x[32] ^ x[35];
    assign layer0_out[4510] = x[159] & ~x[140];
    assign layer0_out[4511] = ~x[223];
    assign layer0_out[4512] = x[379] | x[395];
    assign layer0_out[4513] = ~(x[123] | x[126]);
    assign layer0_out[4514] = ~x[208];
    assign layer0_out[4515] = ~x[109] | x[113];
    assign layer0_out[4516] = ~x[193];
    assign layer0_out[4517] = x[273] ^ x[291];
    assign layer0_out[4518] = x[267] & ~x[260];
    assign layer0_out[4519] = x[77] | x[79];
    assign layer0_out[4520] = ~x[108] | x[93];
    assign layer0_out[4521] = ~(x[5] | x[7]);
    assign layer0_out[4522] = ~(x[176] ^ x[184]);
    assign layer0_out[4523] = x[11] & ~x[0];
    assign layer0_out[4524] = ~x[368] | x[359];
    assign layer0_out[4525] = x[308] & ~x[324];
    assign layer0_out[4526] = x[243];
    assign layer0_out[4527] = ~(x[50] | x[59]);
    assign layer0_out[4528] = ~(x[32] & x[36]);
    assign layer0_out[4529] = 1'b0;
    assign layer0_out[4530] = x[70];
    assign layer0_out[4531] = ~(x[280] | x[294]);
    assign layer0_out[4532] = ~x[38];
    assign layer0_out[4533] = x[315] & x[320];
    assign layer0_out[4534] = ~x[33];
    assign layer0_out[4535] = x[83];
    assign layer0_out[4536] = ~x[349] | x[354];
    assign layer0_out[4537] = ~(x[111] | x[119]);
    assign layer0_out[4538] = 1'b1;
    assign layer0_out[4539] = ~x[150];
    assign layer0_out[4540] = ~x[213] | x[198];
    assign layer0_out[4541] = 1'b0;
    assign layer0_out[4542] = ~(x[187] | x[203]);
    assign layer0_out[4543] = ~x[206];
    assign layer0_out[4544] = ~x[39];
    assign layer0_out[4545] = x[161] ^ x[166];
    assign layer0_out[4546] = ~(x[25] & x[46]);
    assign layer0_out[4547] = x[200];
    assign layer0_out[4548] = x[83] & x[87];
    assign layer0_out[4549] = x[166];
    assign layer0_out[4550] = ~x[360] | x[357];
    assign layer0_out[4551] = ~(x[357] | x[376]);
    assign layer0_out[4552] = ~x[302];
    assign layer0_out[4553] = ~(x[117] | x[135]);
    assign layer0_out[4554] = x[280] & ~x[290];
    assign layer0_out[4555] = x[62] | x[70];
    assign layer0_out[4556] = 1'b1;
    assign layer0_out[4557] = ~(x[24] | x[43]);
    assign layer0_out[4558] = ~(x[88] ^ x[95]);
    assign layer0_out[4559] = x[42];
    assign layer0_out[4560] = x[9] | x[11];
    assign layer0_out[4561] = ~(x[256] | x[270]);
    assign layer0_out[4562] = x[272] | x[285];
    assign layer0_out[4563] = ~(x[7] | x[23]);
    assign layer0_out[4564] = ~x[116];
    assign layer0_out[4565] = x[156] ^ x[158];
    assign layer0_out[4566] = x[315];
    assign layer0_out[4567] = ~(x[298] | x[312]);
    assign layer0_out[4568] = x[251];
    assign layer0_out[4569] = x[354] & x[372];
    assign layer0_out[4570] = x[322] & ~x[334];
    assign layer0_out[4571] = ~(x[121] ^ x[135]);
    assign layer0_out[4572] = x[377] & ~x[359];
    assign layer0_out[4573] = 1'b1;
    assign layer0_out[4574] = 1'b0;
    assign layer0_out[4575] = 1'b1;
    assign layer0_out[4576] = ~(x[242] ^ x[254]);
    assign layer0_out[4577] = ~(x[37] ^ x[52]);
    assign layer0_out[4578] = ~(x[182] & x[195]);
    assign layer0_out[4579] = ~(x[148] | x[150]);
    assign layer0_out[4580] = ~x[296] | x[313];
    assign layer0_out[4581] = x[273] ^ x[289];
    assign layer0_out[4582] = ~x[180] | x[164];
    assign layer0_out[4583] = ~(x[66] & x[81]);
    assign layer0_out[4584] = ~x[216] | x[205];
    assign layer0_out[4585] = ~x[284] | x[296];
    assign layer0_out[4586] = ~x[104];
    assign layer0_out[4587] = x[106] & x[124];
    assign layer0_out[4588] = ~x[194];
    assign layer0_out[4589] = ~(x[95] ^ x[96]);
    assign layer0_out[4590] = x[350] | x[354];
    assign layer0_out[4591] = ~x[80];
    assign layer0_out[4592] = x[243] & x[245];
    assign layer0_out[4593] = ~(x[47] | x[54]);
    assign layer0_out[4594] = ~x[337];
    assign layer0_out[4595] = x[194] ^ x[197];
    assign layer0_out[4596] = x[131];
    assign layer0_out[4597] = ~(x[262] | x[263]);
    assign layer0_out[4598] = ~x[367];
    assign layer0_out[4599] = x[59] & ~x[57];
    assign layer0_out[4600] = x[124] | x[142];
    assign layer0_out[4601] = x[215] | x[235];
    assign layer0_out[4602] = x[335] | x[339];
    assign layer0_out[4603] = ~(x[278] & x[287]);
    assign layer0_out[4604] = ~x[139];
    assign layer0_out[4605] = ~(x[140] | x[155]);
    assign layer0_out[4606] = x[285];
    assign layer0_out[4607] = ~(x[373] | x[387]);
    assign layer0_out[4608] = x[381] | x[384];
    assign layer0_out[4609] = ~(x[130] | x[141]);
    assign layer0_out[4610] = x[246] | x[247];
    assign layer0_out[4611] = 1'b0;
    assign layer0_out[4612] = ~x[221];
    assign layer0_out[4613] = x[98] ^ x[106];
    assign layer0_out[4614] = ~(x[58] | x[70]);
    assign layer0_out[4615] = x[87] ^ x[90];
    assign layer0_out[4616] = ~(x[338] ^ x[354]);
    assign layer0_out[4617] = ~x[55];
    assign layer0_out[4618] = ~x[272];
    assign layer0_out[4619] = x[209] & x[216];
    assign layer0_out[4620] = ~x[147];
    assign layer0_out[4621] = x[182] & x[188];
    assign layer0_out[4622] = ~x[191];
    assign layer0_out[4623] = ~x[116] | x[115];
    assign layer0_out[4624] = ~x[364];
    assign layer0_out[4625] = x[251];
    assign layer0_out[4626] = x[74];
    assign layer0_out[4627] = ~x[186] | x[175];
    assign layer0_out[4628] = x[207] & ~x[195];
    assign layer0_out[4629] = x[321] & x[322];
    assign layer0_out[4630] = ~(x[337] & x[341]);
    assign layer0_out[4631] = x[86] ^ x[102];
    assign layer0_out[4632] = x[228] & ~x[248];
    assign layer0_out[4633] = ~(x[152] ^ x[161]);
    assign layer0_out[4634] = ~x[39];
    assign layer0_out[4635] = x[394];
    assign layer0_out[4636] = x[156] ^ x[164];
    assign layer0_out[4637] = x[104] ^ x[117];
    assign layer0_out[4638] = ~x[369];
    assign layer0_out[4639] = ~x[236] | x[241];
    assign layer0_out[4640] = ~(x[303] ^ x[309]);
    assign layer0_out[4641] = x[57] ^ x[60];
    assign layer0_out[4642] = x[263] | x[276];
    assign layer0_out[4643] = x[166];
    assign layer0_out[4644] = x[175] ^ x[180];
    assign layer0_out[4645] = x[53] & ~x[47];
    assign layer0_out[4646] = ~x[288];
    assign layer0_out[4647] = ~(x[137] & x[153]);
    assign layer0_out[4648] = x[142] & x[162];
    assign layer0_out[4649] = x[252];
    assign layer0_out[4650] = ~(x[13] | x[21]);
    assign layer0_out[4651] = ~x[289];
    assign layer0_out[4652] = ~x[192];
    assign layer0_out[4653] = ~x[184];
    assign layer0_out[4654] = ~(x[113] | x[118]);
    assign layer0_out[4655] = x[299];
    assign layer0_out[4656] = ~x[188] | x[197];
    assign layer0_out[4657] = ~x[116];
    assign layer0_out[4658] = x[25] | x[42];
    assign layer0_out[4659] = x[46];
    assign layer0_out[4660] = ~(x[232] | x[240]);
    assign layer0_out[4661] = x[115];
    assign layer0_out[4662] = ~(x[317] | x[319]);
    assign layer0_out[4663] = ~(x[266] | x[267]);
    assign layer0_out[4664] = x[115];
    assign layer0_out[4665] = ~(x[95] | x[106]);
    assign layer0_out[4666] = x[148];
    assign layer0_out[4667] = x[247];
    assign layer0_out[4668] = x[393];
    assign layer0_out[4669] = x[397];
    assign layer0_out[4670] = ~x[179] | x[200];
    assign layer0_out[4671] = ~x[278] | x[262];
    assign layer0_out[4672] = ~(x[251] & x[261]);
    assign layer0_out[4673] = ~x[29];
    assign layer0_out[4674] = ~(x[36] & x[51]);
    assign layer0_out[4675] = x[20] & ~x[4];
    assign layer0_out[4676] = ~x[336] | x[330];
    assign layer0_out[4677] = ~x[178];
    assign layer0_out[4678] = x[84] & ~x[85];
    assign layer0_out[4679] = x[250];
    assign layer0_out[4680] = x[240];
    assign layer0_out[4681] = x[242];
    assign layer0_out[4682] = ~(x[39] & x[57]);
    assign layer0_out[4683] = ~x[50];
    assign layer0_out[4684] = x[53] | x[60];
    assign layer0_out[4685] = x[97];
    assign layer0_out[4686] = ~x[122];
    assign layer0_out[4687] = x[88] & ~x[101];
    assign layer0_out[4688] = x[318] & x[319];
    assign layer0_out[4689] = ~(x[250] | x[266]);
    assign layer0_out[4690] = x[78] & ~x[58];
    assign layer0_out[4691] = x[155] & ~x[148];
    assign layer0_out[4692] = ~x[190] | x[187];
    assign layer0_out[4693] = x[367] | x[370];
    assign layer0_out[4694] = ~x[276];
    assign layer0_out[4695] = x[181];
    assign layer0_out[4696] = ~x[264];
    assign layer0_out[4697] = x[251] & x[262];
    assign layer0_out[4698] = x[345] & x[351];
    assign layer0_out[4699] = x[129] & ~x[116];
    assign layer0_out[4700] = ~(x[90] | x[109]);
    assign layer0_out[4701] = x[191];
    assign layer0_out[4702] = 1'b0;
    assign layer0_out[4703] = ~(x[185] ^ x[202]);
    assign layer0_out[4704] = ~x[194] | x[187];
    assign layer0_out[4705] = x[132] | x[151];
    assign layer0_out[4706] = ~(x[63] & x[65]);
    assign layer0_out[4707] = 1'b1;
    assign layer0_out[4708] = ~x[228] | x[224];
    assign layer0_out[4709] = x[53];
    assign layer0_out[4710] = x[240] ^ x[246];
    assign layer0_out[4711] = x[195] & ~x[189];
    assign layer0_out[4712] = 1'b1;
    assign layer0_out[4713] = x[257] ^ x[276];
    assign layer0_out[4714] = x[38] | x[48];
    assign layer0_out[4715] = 1'b1;
    assign layer0_out[4716] = ~(x[358] | x[366]);
    assign layer0_out[4717] = ~(x[281] ^ x[298]);
    assign layer0_out[4718] = x[148];
    assign layer0_out[4719] = ~(x[24] | x[45]);
    assign layer0_out[4720] = x[345] & ~x[352];
    assign layer0_out[4721] = x[22];
    assign layer0_out[4722] = ~(x[167] | x[169]);
    assign layer0_out[4723] = ~x[386];
    assign layer0_out[4724] = ~(x[288] & x[293]);
    assign layer0_out[4725] = x[322] ^ x[338];
    assign layer0_out[4726] = ~x[171];
    assign layer0_out[4727] = ~x[2] | x[13];
    assign layer0_out[4728] = ~x[207] | x[206];
    assign layer0_out[4729] = x[388] & ~x[397];
    assign layer0_out[4730] = ~x[295];
    assign layer0_out[4731] = ~(x[175] | x[182]);
    assign layer0_out[4732] = x[244] | x[247];
    assign layer0_out[4733] = ~x[151];
    assign layer0_out[4734] = x[103] | x[124];
    assign layer0_out[4735] = ~(x[194] & x[207]);
    assign layer0_out[4736] = ~x[360];
    assign layer0_out[4737] = x[247] & ~x[266];
    assign layer0_out[4738] = x[157] ^ x[174];
    assign layer0_out[4739] = x[157];
    assign layer0_out[4740] = 1'b0;
    assign layer0_out[4741] = ~x[264];
    assign layer0_out[4742] = x[387] ^ x[398];
    assign layer0_out[4743] = ~(x[333] & x[348]);
    assign layer0_out[4744] = x[351] | x[352];
    assign layer0_out[4745] = ~x[89];
    assign layer0_out[4746] = 1'b1;
    assign layer0_out[4747] = ~x[249] | x[258];
    assign layer0_out[4748] = x[350];
    assign layer0_out[4749] = ~(x[217] ^ x[233]);
    assign layer0_out[4750] = ~x[369];
    assign layer0_out[4751] = x[250];
    assign layer0_out[4752] = ~(x[36] | x[57]);
    assign layer0_out[4753] = x[367] & ~x[386];
    assign layer0_out[4754] = ~x[175];
    assign layer0_out[4755] = ~x[240] | x[223];
    assign layer0_out[4756] = x[163] & x[174];
    assign layer0_out[4757] = x[302] & ~x[308];
    assign layer0_out[4758] = x[22] ^ x[41];
    assign layer0_out[4759] = ~(x[313] | x[322]);
    assign layer0_out[4760] = x[371];
    assign layer0_out[4761] = x[310] & x[319];
    assign layer0_out[4762] = x[64] | x[81];
    assign layer0_out[4763] = ~(x[235] & x[242]);
    assign layer0_out[4764] = ~x[390];
    assign layer0_out[4765] = x[112] | x[121];
    assign layer0_out[4766] = ~x[374];
    assign layer0_out[4767] = ~x[168];
    assign layer0_out[4768] = ~(x[98] | x[116]);
    assign layer0_out[4769] = x[116] & x[135];
    assign layer0_out[4770] = 1'b0;
    assign layer0_out[4771] = 1'b0;
    assign layer0_out[4772] = ~x[67];
    assign layer0_out[4773] = x[215] | x[228];
    assign layer0_out[4774] = 1'b1;
    assign layer0_out[4775] = ~x[368];
    assign layer0_out[4776] = ~x[271];
    assign layer0_out[4777] = x[2];
    assign layer0_out[4778] = ~(x[245] | x[265]);
    assign layer0_out[4779] = ~(x[145] | x[159]);
    assign layer0_out[4780] = x[170];
    assign layer0_out[4781] = x[111];
    assign layer0_out[4782] = x[141] & ~x[127];
    assign layer0_out[4783] = ~(x[320] ^ x[332]);
    assign layer0_out[4784] = x[350] ^ x[367];
    assign layer0_out[4785] = x[275] & ~x[288];
    assign layer0_out[4786] = ~(x[178] | x[198]);
    assign layer0_out[4787] = ~(x[166] | x[184]);
    assign layer0_out[4788] = ~(x[76] ^ x[93]);
    assign layer0_out[4789] = x[286] & ~x[305];
    assign layer0_out[4790] = ~(x[143] ^ x[146]);
    assign layer0_out[4791] = ~x[23];
    assign layer0_out[4792] = ~x[146] | x[153];
    assign layer0_out[4793] = x[343];
    assign layer0_out[4794] = x[196] ^ x[217];
    assign layer0_out[4795] = x[214] ^ x[232];
    assign layer0_out[4796] = ~x[382] | x[362];
    assign layer0_out[4797] = 1'b0;
    assign layer0_out[4798] = x[58] | x[63];
    assign layer0_out[4799] = 1'b1;
    assign layer0_out[4800] = x[6] | x[27];
    assign layer0_out[4801] = ~(x[365] | x[381]);
    assign layer0_out[4802] = ~(x[123] | x[133]);
    assign layer0_out[4803] = x[76] & ~x[82];
    assign layer0_out[4804] = ~x[35];
    assign layer0_out[4805] = ~x[58];
    assign layer0_out[4806] = ~x[31] | x[32];
    assign layer0_out[4807] = x[103];
    assign layer0_out[4808] = x[97] & ~x[76];
    assign layer0_out[4809] = x[12] | x[14];
    assign layer0_out[4810] = ~(x[63] | x[80]);
    assign layer0_out[4811] = ~x[241];
    assign layer0_out[4812] = ~(x[82] ^ x[102]);
    assign layer0_out[4813] = ~(x[300] | x[304]);
    assign layer0_out[4814] = ~x[198];
    assign layer0_out[4815] = x[30] | x[49];
    assign layer0_out[4816] = x[129] & x[135];
    assign layer0_out[4817] = x[26] & ~x[37];
    assign layer0_out[4818] = ~(x[0] | x[5]);
    assign layer0_out[4819] = ~x[125];
    assign layer0_out[4820] = x[229] & ~x[223];
    assign layer0_out[4821] = x[79] | x[82];
    assign layer0_out[4822] = ~x[218] | x[213];
    assign layer0_out[4823] = ~x[12] | x[6];
    assign layer0_out[4824] = x[202];
    assign layer0_out[4825] = ~x[357];
    assign layer0_out[4826] = 1'b1;
    assign layer0_out[4827] = x[82] & ~x[66];
    assign layer0_out[4828] = 1'b1;
    assign layer0_out[4829] = x[148] ^ x[158];
    assign layer0_out[4830] = x[311] ^ x[327];
    assign layer0_out[4831] = x[260] & ~x[273];
    assign layer0_out[4832] = ~(x[154] | x[157]);
    assign layer0_out[4833] = ~x[283];
    assign layer0_out[4834] = ~x[128];
    assign layer0_out[4835] = ~(x[100] & x[106]);
    assign layer0_out[4836] = x[232] & ~x[245];
    assign layer0_out[4837] = x[38] | x[59];
    assign layer0_out[4838] = ~(x[99] ^ x[116]);
    assign layer0_out[4839] = ~x[177] | x[159];
    assign layer0_out[4840] = ~x[229];
    assign layer0_out[4841] = ~(x[365] ^ x[376]);
    assign layer0_out[4842] = ~x[204] | x[188];
    assign layer0_out[4843] = ~x[131] | x[119];
    assign layer0_out[4844] = ~x[223];
    assign layer0_out[4845] = x[151] | x[169];
    assign layer0_out[4846] = x[223];
    assign layer0_out[4847] = x[107] | x[126];
    assign layer0_out[4848] = x[31] | x[51];
    assign layer0_out[4849] = x[72];
    assign layer0_out[4850] = x[170] & ~x[178];
    assign layer0_out[4851] = x[137] ^ x[154];
    assign layer0_out[4852] = ~x[314];
    assign layer0_out[4853] = ~x[120] | x[121];
    assign layer0_out[4854] = ~x[290] | x[282];
    assign layer0_out[4855] = 1'b0;
    assign layer0_out[4856] = x[285] | x[296];
    assign layer0_out[4857] = x[321];
    assign layer0_out[4858] = x[386];
    assign layer0_out[4859] = ~(x[174] | x[179]);
    assign layer0_out[4860] = x[318] | x[322];
    assign layer0_out[4861] = ~(x[205] | x[225]);
    assign layer0_out[4862] = x[66] | x[69];
    assign layer0_out[4863] = ~x[333];
    assign layer0_out[4864] = x[75];
    assign layer0_out[4865] = x[222] & ~x[218];
    assign layer0_out[4866] = x[273] | x[285];
    assign layer0_out[4867] = x[300];
    assign layer0_out[4868] = ~(x[94] ^ x[96]);
    assign layer0_out[4869] = ~(x[144] | x[158]);
    assign layer0_out[4870] = x[320];
    assign layer0_out[4871] = ~(x[344] | x[353]);
    assign layer0_out[4872] = x[243] & ~x[227];
    assign layer0_out[4873] = ~x[33];
    assign layer0_out[4874] = ~x[116] | x[130];
    assign layer0_out[4875] = x[342] | x[349];
    assign layer0_out[4876] = ~(x[126] | x[130]);
    assign layer0_out[4877] = x[127] & ~x[133];
    assign layer0_out[4878] = x[135];
    assign layer0_out[4879] = ~x[245] | x[237];
    assign layer0_out[4880] = x[367] & ~x[377];
    assign layer0_out[4881] = ~x[342];
    assign layer0_out[4882] = ~(x[29] & x[42]);
    assign layer0_out[4883] = x[301] | x[303];
    assign layer0_out[4884] = 1'b0;
    assign layer0_out[4885] = ~x[315];
    assign layer0_out[4886] = ~x[256] | x[250];
    assign layer0_out[4887] = ~x[218] | x[220];
    assign layer0_out[4888] = x[216];
    assign layer0_out[4889] = ~x[241] | x[233];
    assign layer0_out[4890] = ~x[255] | x[271];
    assign layer0_out[4891] = x[63] | x[78];
    assign layer0_out[4892] = ~(x[61] & x[82]);
    assign layer0_out[4893] = x[247];
    assign layer0_out[4894] = x[141];
    assign layer0_out[4895] = ~x[202] | x[211];
    assign layer0_out[4896] = ~(x[298] | x[317]);
    assign layer0_out[4897] = ~(x[31] ^ x[48]);
    assign layer0_out[4898] = x[52] | x[62];
    assign layer0_out[4899] = ~(x[150] ^ x[161]);
    assign layer0_out[4900] = 1'b0;
    assign layer0_out[4901] = ~(x[22] | x[43]);
    assign layer0_out[4902] = x[275] & ~x[270];
    assign layer0_out[4903] = ~(x[66] & x[75]);
    assign layer0_out[4904] = x[221] & x[230];
    assign layer0_out[4905] = x[346] | x[351];
    assign layer0_out[4906] = x[115] | x[124];
    assign layer0_out[4907] = ~x[359] | x[340];
    assign layer0_out[4908] = ~(x[210] & x[224]);
    assign layer0_out[4909] = ~(x[120] ^ x[123]);
    assign layer0_out[4910] = ~x[74] | x[65];
    assign layer0_out[4911] = x[158] & ~x[138];
    assign layer0_out[4912] = 1'b0;
    assign layer0_out[4913] = ~x[164];
    assign layer0_out[4914] = x[294];
    assign layer0_out[4915] = ~(x[253] | x[260]);
    assign layer0_out[4916] = x[272] | x[273];
    assign layer0_out[4917] = x[57];
    assign layer0_out[4918] = ~(x[309] | x[319]);
    assign layer0_out[4919] = ~(x[282] ^ x[297]);
    assign layer0_out[4920] = ~x[233];
    assign layer0_out[4921] = x[202] & ~x[213];
    assign layer0_out[4922] = x[311] | x[316];
    assign layer0_out[4923] = x[31] & x[34];
    assign layer0_out[4924] = x[247];
    assign layer0_out[4925] = ~(x[348] | x[367]);
    assign layer0_out[4926] = ~(x[389] ^ x[397]);
    assign layer0_out[4927] = x[113] & ~x[121];
    assign layer0_out[4928] = ~(x[165] | x[167]);
    assign layer0_out[4929] = x[278] & ~x[277];
    assign layer0_out[4930] = 1'b1;
    assign layer0_out[4931] = ~x[316] | x[318];
    assign layer0_out[4932] = x[170] ^ x[184];
    assign layer0_out[4933] = ~x[307] | x[297];
    assign layer0_out[4934] = ~x[159];
    assign layer0_out[4935] = ~(x[271] & x[290]);
    assign layer0_out[4936] = ~(x[157] | x[158]);
    assign layer0_out[4937] = x[110] ^ x[128];
    assign layer0_out[4938] = ~x[306] | x[318];
    assign layer0_out[4939] = x[175];
    assign layer0_out[4940] = ~x[6];
    assign layer0_out[4941] = ~x[274] | x[254];
    assign layer0_out[4942] = x[285];
    assign layer0_out[4943] = x[338];
    assign layer0_out[4944] = ~(x[155] | x[174]);
    assign layer0_out[4945] = ~(x[110] | x[131]);
    assign layer0_out[4946] = ~(x[309] & x[323]);
    assign layer0_out[4947] = ~(x[154] | x[161]);
    assign layer0_out[4948] = x[321];
    assign layer0_out[4949] = x[306] & x[312];
    assign layer0_out[4950] = x[298] ^ x[302];
    assign layer0_out[4951] = x[369];
    assign layer0_out[4952] = ~x[285];
    assign layer0_out[4953] = x[262];
    assign layer0_out[4954] = x[158] & ~x[153];
    assign layer0_out[4955] = ~x[335];
    assign layer0_out[4956] = ~(x[210] | x[228]);
    assign layer0_out[4957] = x[11] & ~x[26];
    assign layer0_out[4958] = ~(x[132] | x[133]);
    assign layer0_out[4959] = ~x[79];
    assign layer0_out[4960] = ~x[333];
    assign layer0_out[4961] = x[5] | x[6];
    assign layer0_out[4962] = ~x[106];
    assign layer0_out[4963] = x[158] | x[178];
    assign layer0_out[4964] = ~(x[368] | x[382]);
    assign layer0_out[4965] = ~(x[109] & x[120]);
    assign layer0_out[4966] = ~(x[353] | x[360]);
    assign layer0_out[4967] = x[290] & ~x[303];
    assign layer0_out[4968] = ~(x[116] | x[137]);
    assign layer0_out[4969] = x[187] & ~x[179];
    assign layer0_out[4970] = ~x[217];
    assign layer0_out[4971] = x[192];
    assign layer0_out[4972] = ~x[352];
    assign layer0_out[4973] = x[172] | x[182];
    assign layer0_out[4974] = x[287];
    assign layer0_out[4975] = 1'b0;
    assign layer0_out[4976] = ~x[383] | x[399];
    assign layer0_out[4977] = ~(x[336] | x[340]);
    assign layer0_out[4978] = ~(x[20] & x[25]);
    assign layer0_out[4979] = x[229] | x[243];
    assign layer0_out[4980] = ~(x[341] & x[342]);
    assign layer0_out[4981] = ~(x[338] | x[349]);
    assign layer0_out[4982] = ~(x[11] | x[31]);
    assign layer0_out[4983] = ~x[100];
    assign layer0_out[4984] = ~x[290];
    assign layer0_out[4985] = x[122] | x[137];
    assign layer0_out[4986] = ~x[335] | x[346];
    assign layer0_out[4987] = ~x[101];
    assign layer0_out[4988] = ~(x[362] | x[376]);
    assign layer0_out[4989] = ~(x[290] | x[299]);
    assign layer0_out[4990] = x[17] & ~x[37];
    assign layer0_out[4991] = x[56];
    assign layer0_out[4992] = x[45] & ~x[47];
    assign layer0_out[4993] = x[245];
    assign layer0_out[4994] = ~(x[308] | x[310]);
    assign layer0_out[4995] = ~(x[276] | x[295]);
    assign layer0_out[4996] = x[114];
    assign layer0_out[4997] = 1'b1;
    assign layer0_out[4998] = x[271] & x[286];
    assign layer0_out[4999] = x[367] ^ x[373];
    assign layer0_out[5000] = ~x[2] | x[11];
    assign layer0_out[5001] = ~x[245] | x[247];
    assign layer0_out[5002] = ~x[344];
    assign layer0_out[5003] = ~x[128] | x[118];
    assign layer0_out[5004] = x[152] ^ x[156];
    assign layer0_out[5005] = x[179] | x[199];
    assign layer0_out[5006] = x[24] & ~x[23];
    assign layer0_out[5007] = x[281] ^ x[290];
    assign layer0_out[5008] = ~x[169];
    assign layer0_out[5009] = ~x[210];
    assign layer0_out[5010] = ~(x[234] ^ x[236]);
    assign layer0_out[5011] = x[377] & ~x[393];
    assign layer0_out[5012] = ~(x[151] & x[159]);
    assign layer0_out[5013] = ~(x[377] | x[397]);
    assign layer0_out[5014] = x[279] & ~x[298];
    assign layer0_out[5015] = x[313];
    assign layer0_out[5016] = x[314] | x[324];
    assign layer0_out[5017] = ~(x[356] | x[360]);
    assign layer0_out[5018] = ~(x[226] & x[229]);
    assign layer0_out[5019] = ~(x[29] & x[47]);
    assign layer0_out[5020] = x[89] & ~x[71];
    assign layer0_out[5021] = ~x[390];
    assign layer0_out[5022] = ~x[329] | x[327];
    assign layer0_out[5023] = x[26] | x[46];
    assign layer0_out[5024] = ~(x[259] | x[264]);
    assign layer0_out[5025] = ~(x[46] | x[62]);
    assign layer0_out[5026] = ~x[68] | x[84];
    assign layer0_out[5027] = 1'b0;
    assign layer0_out[5028] = ~(x[160] | x[181]);
    assign layer0_out[5029] = x[5];
    assign layer0_out[5030] = x[343];
    assign layer0_out[5031] = ~(x[171] | x[173]);
    assign layer0_out[5032] = x[142] | x[158];
    assign layer0_out[5033] = 1'b0;
    assign layer0_out[5034] = ~x[387] | x[379];
    assign layer0_out[5035] = 1'b0;
    assign layer0_out[5036] = x[82] & ~x[98];
    assign layer0_out[5037] = ~(x[3] | x[20]);
    assign layer0_out[5038] = ~(x[27] ^ x[36]);
    assign layer0_out[5039] = ~(x[49] | x[57]);
    assign layer0_out[5040] = x[120] & ~x[126];
    assign layer0_out[5041] = x[194] & x[215];
    assign layer0_out[5042] = ~x[337];
    assign layer0_out[5043] = ~(x[148] ^ x[166]);
    assign layer0_out[5044] = 1'b1;
    assign layer0_out[5045] = ~x[295] | x[298];
    assign layer0_out[5046] = x[335] & ~x[327];
    assign layer0_out[5047] = ~(x[328] | x[331]);
    assign layer0_out[5048] = ~(x[257] & x[275]);
    assign layer0_out[5049] = x[271];
    assign layer0_out[5050] = ~(x[218] | x[233]);
    assign layer0_out[5051] = x[61] ^ x[64];
    assign layer0_out[5052] = ~x[248] | x[250];
    assign layer0_out[5053] = ~(x[348] ^ x[349]);
    assign layer0_out[5054] = x[124] & ~x[128];
    assign layer0_out[5055] = ~x[71];
    assign layer0_out[5056] = x[256] | x[262];
    assign layer0_out[5057] = x[20] | x[40];
    assign layer0_out[5058] = ~x[17];
    assign layer0_out[5059] = ~(x[298] ^ x[300]);
    assign layer0_out[5060] = ~x[291] | x[297];
    assign layer0_out[5061] = ~x[292];
    assign layer0_out[5062] = x[273] | x[275];
    assign layer0_out[5063] = ~(x[51] ^ x[71]);
    assign layer0_out[5064] = ~x[31];
    assign layer0_out[5065] = x[192];
    assign layer0_out[5066] = x[23] & ~x[35];
    assign layer0_out[5067] = x[326] | x[342];
    assign layer0_out[5068] = ~x[261] | x[278];
    assign layer0_out[5069] = ~x[385];
    assign layer0_out[5070] = x[56] | x[66];
    assign layer0_out[5071] = ~x[4];
    assign layer0_out[5072] = x[149] & ~x[159];
    assign layer0_out[5073] = ~(x[376] ^ x[394]);
    assign layer0_out[5074] = ~(x[201] & x[208]);
    assign layer0_out[5075] = ~x[285];
    assign layer0_out[5076] = ~(x[318] | x[338]);
    assign layer0_out[5077] = x[125] | x[126];
    assign layer0_out[5078] = 1'b0;
    assign layer0_out[5079] = x[19] & ~x[17];
    assign layer0_out[5080] = ~x[138];
    assign layer0_out[5081] = x[34] ^ x[36];
    assign layer0_out[5082] = x[377] & ~x[382];
    assign layer0_out[5083] = x[173] | x[193];
    assign layer0_out[5084] = ~(x[144] ^ x[156]);
    assign layer0_out[5085] = x[393] & ~x[398];
    assign layer0_out[5086] = x[193] & x[201];
    assign layer0_out[5087] = ~(x[41] ^ x[43]);
    assign layer0_out[5088] = x[299] ^ x[312];
    assign layer0_out[5089] = 1'b1;
    assign layer0_out[5090] = ~(x[367] | x[387]);
    assign layer0_out[5091] = ~x[58];
    assign layer0_out[5092] = x[128];
    assign layer0_out[5093] = ~x[31];
    assign layer0_out[5094] = ~(x[265] | x[276]);
    assign layer0_out[5095] = x[1] | x[5];
    assign layer0_out[5096] = ~(x[386] | x[399]);
    assign layer0_out[5097] = ~x[169];
    assign layer0_out[5098] = ~x[385] | x[387];
    assign layer0_out[5099] = 1'b0;
    assign layer0_out[5100] = ~(x[243] | x[259]);
    assign layer0_out[5101] = x[180] | x[198];
    assign layer0_out[5102] = ~x[229];
    assign layer0_out[5103] = ~x[61];
    assign layer0_out[5104] = x[186] & x[195];
    assign layer0_out[5105] = x[0] ^ x[10];
    assign layer0_out[5106] = x[144] & ~x[148];
    assign layer0_out[5107] = ~x[183];
    assign layer0_out[5108] = x[220];
    assign layer0_out[5109] = ~x[270];
    assign layer0_out[5110] = x[17];
    assign layer0_out[5111] = ~(x[176] | x[197]);
    assign layer0_out[5112] = ~x[184] | x[187];
    assign layer0_out[5113] = ~x[26];
    assign layer0_out[5114] = ~(x[97] & x[116]);
    assign layer0_out[5115] = x[271] & x[281];
    assign layer0_out[5116] = x[68] | x[87];
    assign layer0_out[5117] = x[8] ^ x[25];
    assign layer0_out[5118] = x[379];
    assign layer0_out[5119] = 1'b1;
    assign layer0_out[5120] = x[162] & ~x[179];
    assign layer0_out[5121] = ~(x[124] & x[127]);
    assign layer0_out[5122] = ~x[82];
    assign layer0_out[5123] = x[105] & ~x[125];
    assign layer0_out[5124] = x[0] & ~x[14];
    assign layer0_out[5125] = x[280];
    assign layer0_out[5126] = ~(x[358] & x[368]);
    assign layer0_out[5127] = ~x[247] | x[256];
    assign layer0_out[5128] = ~x[179];
    assign layer0_out[5129] = x[331] & ~x[341];
    assign layer0_out[5130] = ~x[399] | x[394];
    assign layer0_out[5131] = x[141] & ~x[143];
    assign layer0_out[5132] = x[84];
    assign layer0_out[5133] = x[357];
    assign layer0_out[5134] = x[81] & ~x[67];
    assign layer0_out[5135] = ~(x[316] | x[324]);
    assign layer0_out[5136] = x[41];
    assign layer0_out[5137] = x[56];
    assign layer0_out[5138] = x[54] ^ x[63];
    assign layer0_out[5139] = x[95] | x[104];
    assign layer0_out[5140] = x[260] & ~x[244];
    assign layer0_out[5141] = ~x[43];
    assign layer0_out[5142] = 1'b1;
    assign layer0_out[5143] = ~(x[42] | x[58]);
    assign layer0_out[5144] = x[389];
    assign layer0_out[5145] = ~x[112] | x[108];
    assign layer0_out[5146] = x[81] ^ x[86];
    assign layer0_out[5147] = ~x[238] | x[225];
    assign layer0_out[5148] = ~x[197] | x[196];
    assign layer0_out[5149] = ~x[249] | x[238];
    assign layer0_out[5150] = x[34] & x[48];
    assign layer0_out[5151] = 1'b0;
    assign layer0_out[5152] = x[105] | x[113];
    assign layer0_out[5153] = ~x[202];
    assign layer0_out[5154] = x[237] | x[240];
    assign layer0_out[5155] = ~x[17];
    assign layer0_out[5156] = ~x[281];
    assign layer0_out[5157] = 1'b0;
    assign layer0_out[5158] = ~x[394];
    assign layer0_out[5159] = x[38] & ~x[23];
    assign layer0_out[5160] = ~x[79];
    assign layer0_out[5161] = x[207];
    assign layer0_out[5162] = x[101] & ~x[97];
    assign layer0_out[5163] = 1'b0;
    assign layer0_out[5164] = ~(x[286] | x[301]);
    assign layer0_out[5165] = x[315] & x[332];
    assign layer0_out[5166] = ~(x[33] | x[52]);
    assign layer0_out[5167] = ~(x[330] & x[344]);
    assign layer0_out[5168] = ~x[270];
    assign layer0_out[5169] = ~x[281];
    assign layer0_out[5170] = ~x[125];
    assign layer0_out[5171] = x[102] ^ x[108];
    assign layer0_out[5172] = 1'b1;
    assign layer0_out[5173] = ~(x[257] | x[259]);
    assign layer0_out[5174] = ~(x[218] | x[237]);
    assign layer0_out[5175] = x[303] | x[314];
    assign layer0_out[5176] = x[111] ^ x[126];
    assign layer0_out[5177] = x[30] & ~x[43];
    assign layer0_out[5178] = x[323];
    assign layer0_out[5179] = 1'b1;
    assign layer0_out[5180] = ~(x[287] | x[307]);
    assign layer0_out[5181] = ~x[189] | x[179];
    assign layer0_out[5182] = x[47];
    assign layer0_out[5183] = 1'b1;
    assign layer0_out[5184] = ~x[74];
    assign layer0_out[5185] = ~(x[86] | x[107]);
    assign layer0_out[5186] = x[4];
    assign layer0_out[5187] = ~(x[326] | x[345]);
    assign layer0_out[5188] = x[318] & ~x[299];
    assign layer0_out[5189] = ~x[123];
    assign layer0_out[5190] = x[242] & x[248];
    assign layer0_out[5191] = x[31] | x[49];
    assign layer0_out[5192] = x[253];
    assign layer0_out[5193] = x[316];
    assign layer0_out[5194] = ~x[23];
    assign layer0_out[5195] = x[16] & ~x[13];
    assign layer0_out[5196] = x[182] & ~x[200];
    assign layer0_out[5197] = ~x[153];
    assign layer0_out[5198] = x[218];
    assign layer0_out[5199] = ~x[149];
    assign layer0_out[5200] = x[274] ^ x[276];
    assign layer0_out[5201] = ~x[237] | x[231];
    assign layer0_out[5202] = ~(x[32] ^ x[40]);
    assign layer0_out[5203] = ~(x[9] | x[22]);
    assign layer0_out[5204] = ~(x[45] | x[46]);
    assign layer0_out[5205] = ~x[26] | x[22];
    assign layer0_out[5206] = x[118];
    assign layer0_out[5207] = ~x[44] | x[33];
    assign layer0_out[5208] = x[130] & ~x[117];
    assign layer0_out[5209] = ~(x[362] | x[378]);
    assign layer0_out[5210] = x[177] & x[196];
    assign layer0_out[5211] = x[93] | x[94];
    assign layer0_out[5212] = ~(x[281] | x[300]);
    assign layer0_out[5213] = x[285] ^ x[299];
    assign layer0_out[5214] = ~(x[126] ^ x[142]);
    assign layer0_out[5215] = x[143] ^ x[160];
    assign layer0_out[5216] = ~x[190];
    assign layer0_out[5217] = x[150] | x[158];
    assign layer0_out[5218] = ~(x[284] ^ x[300]);
    assign layer0_out[5219] = ~x[139] | x[134];
    assign layer0_out[5220] = ~x[128] | x[139];
    assign layer0_out[5221] = ~x[107];
    assign layer0_out[5222] = ~x[353];
    assign layer0_out[5223] = x[376];
    assign layer0_out[5224] = 1'b1;
    assign layer0_out[5225] = ~x[206];
    assign layer0_out[5226] = 1'b1;
    assign layer0_out[5227] = 1'b1;
    assign layer0_out[5228] = x[71] & ~x[57];
    assign layer0_out[5229] = x[337];
    assign layer0_out[5230] = ~(x[186] ^ x[189]);
    assign layer0_out[5231] = ~x[170] | x[177];
    assign layer0_out[5232] = x[154];
    assign layer0_out[5233] = ~(x[122] & x[130]);
    assign layer0_out[5234] = x[327];
    assign layer0_out[5235] = x[355] ^ x[367];
    assign layer0_out[5236] = x[330] ^ x[332];
    assign layer0_out[5237] = ~(x[51] | x[57]);
    assign layer0_out[5238] = ~(x[120] | x[141]);
    assign layer0_out[5239] = ~(x[18] ^ x[30]);
    assign layer0_out[5240] = ~(x[311] & x[328]);
    assign layer0_out[5241] = ~(x[366] ^ x[380]);
    assign layer0_out[5242] = x[382];
    assign layer0_out[5243] = x[195] & ~x[193];
    assign layer0_out[5244] = ~(x[337] | x[350]);
    assign layer0_out[5245] = x[159] & x[161];
    assign layer0_out[5246] = x[227];
    assign layer0_out[5247] = ~x[335];
    assign layer0_out[5248] = ~x[312];
    assign layer0_out[5249] = x[339];
    assign layer0_out[5250] = x[79] | x[87];
    assign layer0_out[5251] = ~x[196];
    assign layer0_out[5252] = ~(x[1] | x[11]);
    assign layer0_out[5253] = x[191] & ~x[207];
    assign layer0_out[5254] = ~(x[92] ^ x[99]);
    assign layer0_out[5255] = x[76] & ~x[71];
    assign layer0_out[5256] = ~(x[215] | x[216]);
    assign layer0_out[5257] = x[324] | x[325];
    assign layer0_out[5258] = x[277] | x[294];
    assign layer0_out[5259] = ~(x[133] ^ x[150]);
    assign layer0_out[5260] = ~x[255];
    assign layer0_out[5261] = ~(x[105] ^ x[122]);
    assign layer0_out[5262] = 1'b0;
    assign layer0_out[5263] = ~x[38];
    assign layer0_out[5264] = ~(x[283] ^ x[288]);
    assign layer0_out[5265] = ~x[146];
    assign layer0_out[5266] = 1'b1;
    assign layer0_out[5267] = ~(x[15] | x[20]);
    assign layer0_out[5268] = x[22] | x[31];
    assign layer0_out[5269] = ~x[72];
    assign layer0_out[5270] = x[317] | x[337];
    assign layer0_out[5271] = x[121] & ~x[115];
    assign layer0_out[5272] = ~(x[336] ^ x[337]);
    assign layer0_out[5273] = x[310];
    assign layer0_out[5274] = 1'b0;
    assign layer0_out[5275] = x[248] | x[267];
    assign layer0_out[5276] = ~x[43];
    assign layer0_out[5277] = x[213];
    assign layer0_out[5278] = ~x[67];
    assign layer0_out[5279] = ~x[137] | x[126];
    assign layer0_out[5280] = 1'b1;
    assign layer0_out[5281] = ~x[134] | x[145];
    assign layer0_out[5282] = x[132] ^ x[140];
    assign layer0_out[5283] = x[312] & x[330];
    assign layer0_out[5284] = x[139] | x[156];
    assign layer0_out[5285] = ~x[140] | x[133];
    assign layer0_out[5286] = ~(x[324] ^ x[343]);
    assign layer0_out[5287] = ~(x[166] | x[170]);
    assign layer0_out[5288] = x[22];
    assign layer0_out[5289] = ~(x[33] | x[34]);
    assign layer0_out[5290] = x[356];
    assign layer0_out[5291] = x[30];
    assign layer0_out[5292] = x[208];
    assign layer0_out[5293] = x[360] | x[375];
    assign layer0_out[5294] = x[160] | x[178];
    assign layer0_out[5295] = ~x[37] | x[45];
    assign layer0_out[5296] = ~x[191];
    assign layer0_out[5297] = x[270];
    assign layer0_out[5298] = x[309];
    assign layer0_out[5299] = x[346] | x[350];
    assign layer0_out[5300] = x[94] ^ x[112];
    assign layer0_out[5301] = x[244] ^ x[258];
    assign layer0_out[5302] = x[10] & ~x[3];
    assign layer0_out[5303] = ~x[100];
    assign layer0_out[5304] = x[124];
    assign layer0_out[5305] = x[389] & ~x[395];
    assign layer0_out[5306] = x[99] & ~x[86];
    assign layer0_out[5307] = x[172];
    assign layer0_out[5308] = ~(x[365] | x[379]);
    assign layer0_out[5309] = ~(x[240] | x[245]);
    assign layer0_out[5310] = ~(x[251] & x[265]);
    assign layer0_out[5311] = ~(x[96] ^ x[114]);
    assign layer0_out[5312] = ~x[192];
    assign layer0_out[5313] = ~x[169] | x[176];
    assign layer0_out[5314] = ~(x[32] | x[45]);
    assign layer0_out[5315] = ~(x[209] & x[211]);
    assign layer0_out[5316] = x[109] ^ x[124];
    assign layer0_out[5317] = x[99] | x[112];
    assign layer0_out[5318] = x[51] & ~x[65];
    assign layer0_out[5319] = ~(x[241] | x[260]);
    assign layer0_out[5320] = x[375] | x[376];
    assign layer0_out[5321] = x[226];
    assign layer0_out[5322] = ~(x[48] | x[49]);
    assign layer0_out[5323] = x[135] & ~x[148];
    assign layer0_out[5324] = ~(x[112] ^ x[114]);
    assign layer0_out[5325] = 1'b1;
    assign layer0_out[5326] = x[77] | x[87];
    assign layer0_out[5327] = ~(x[103] | x[105]);
    assign layer0_out[5328] = ~x[24] | x[35];
    assign layer0_out[5329] = ~(x[209] ^ x[230]);
    assign layer0_out[5330] = 1'b0;
    assign layer0_out[5331] = x[89];
    assign layer0_out[5332] = x[169] & ~x[155];
    assign layer0_out[5333] = x[363];
    assign layer0_out[5334] = x[25] | x[33];
    assign layer0_out[5335] = x[300] | x[311];
    assign layer0_out[5336] = ~x[299];
    assign layer0_out[5337] = x[287] & ~x[288];
    assign layer0_out[5338] = ~(x[280] | x[296]);
    assign layer0_out[5339] = ~x[395];
    assign layer0_out[5340] = x[209] & ~x[207];
    assign layer0_out[5341] = ~(x[25] | x[45]);
    assign layer0_out[5342] = ~(x[101] | x[106]);
    assign layer0_out[5343] = ~x[138] | x[156];
    assign layer0_out[5344] = x[392] & ~x[396];
    assign layer0_out[5345] = ~(x[129] ^ x[133]);
    assign layer0_out[5346] = x[315] & x[335];
    assign layer0_out[5347] = x[99];
    assign layer0_out[5348] = x[76] & ~x[83];
    assign layer0_out[5349] = ~x[138];
    assign layer0_out[5350] = ~x[281];
    assign layer0_out[5351] = ~x[163];
    assign layer0_out[5352] = ~x[62] | x[59];
    assign layer0_out[5353] = ~x[149];
    assign layer0_out[5354] = 1'b0;
    assign layer0_out[5355] = ~x[136];
    assign layer0_out[5356] = x[33] & x[49];
    assign layer0_out[5357] = x[131] ^ x[133];
    assign layer0_out[5358] = x[382] & ~x[399];
    assign layer0_out[5359] = ~(x[377] | x[389]);
    assign layer0_out[5360] = ~x[8] | x[12];
    assign layer0_out[5361] = ~(x[176] ^ x[178]);
    assign layer0_out[5362] = ~(x[73] ^ x[75]);
    assign layer0_out[5363] = x[344] | x[356];
    assign layer0_out[5364] = x[324];
    assign layer0_out[5365] = x[14] | x[24];
    assign layer0_out[5366] = x[277] & ~x[273];
    assign layer0_out[5367] = ~(x[382] & x[384]);
    assign layer0_out[5368] = ~(x[84] | x[99]);
    assign layer0_out[5369] = x[19] & ~x[39];
    assign layer0_out[5370] = ~x[135];
    assign layer0_out[5371] = x[199] | x[218];
    assign layer0_out[5372] = ~(x[186] | x[190]);
    assign layer0_out[5373] = ~x[299];
    assign layer0_out[5374] = ~x[300];
    assign layer0_out[5375] = ~x[344];
    assign layer0_out[5376] = x[260];
    assign layer0_out[5377] = ~x[47];
    assign layer0_out[5378] = x[206] & x[218];
    assign layer0_out[5379] = ~(x[100] | x[107]);
    assign layer0_out[5380] = ~x[191] | x[178];
    assign layer0_out[5381] = ~x[271];
    assign layer0_out[5382] = ~(x[350] | x[357]);
    assign layer0_out[5383] = 1'b1;
    assign layer0_out[5384] = ~x[107] | x[93];
    assign layer0_out[5385] = x[369] | x[386];
    assign layer0_out[5386] = x[156];
    assign layer0_out[5387] = x[275] & x[283];
    assign layer0_out[5388] = 1'b0;
    assign layer0_out[5389] = 1'b0;
    assign layer0_out[5390] = x[211];
    assign layer0_out[5391] = ~(x[364] | x[366]);
    assign layer0_out[5392] = x[136] | x[154];
    assign layer0_out[5393] = ~(x[322] | x[341]);
    assign layer0_out[5394] = x[337] | x[345];
    assign layer0_out[5395] = ~x[71] | x[66];
    assign layer0_out[5396] = ~(x[195] | x[202]);
    assign layer0_out[5397] = ~x[89] | x[94];
    assign layer0_out[5398] = ~x[18] | x[33];
    assign layer0_out[5399] = ~x[237];
    assign layer0_out[5400] = x[101];
    assign layer0_out[5401] = ~(x[193] ^ x[198]);
    assign layer0_out[5402] = x[191] & ~x[182];
    assign layer0_out[5403] = x[318] & ~x[298];
    assign layer0_out[5404] = x[343];
    assign layer0_out[5405] = x[335];
    assign layer0_out[5406] = ~(x[369] | x[387]);
    assign layer0_out[5407] = x[257];
    assign layer0_out[5408] = ~(x[77] | x[84]);
    assign layer0_out[5409] = x[217];
    assign layer0_out[5410] = x[21];
    assign layer0_out[5411] = ~x[16] | x[18];
    assign layer0_out[5412] = x[322] & x[333];
    assign layer0_out[5413] = ~x[206];
    assign layer0_out[5414] = x[91] & ~x[79];
    assign layer0_out[5415] = x[134] ^ x[155];
    assign layer0_out[5416] = x[286] & x[296];
    assign layer0_out[5417] = ~(x[307] | x[318]);
    assign layer0_out[5418] = x[366] & ~x[357];
    assign layer0_out[5419] = x[318] | x[320];
    assign layer0_out[5420] = ~(x[192] | x[210]);
    assign layer0_out[5421] = x[172];
    assign layer0_out[5422] = ~(x[7] | x[25]);
    assign layer0_out[5423] = ~(x[200] | x[220]);
    assign layer0_out[5424] = ~(x[150] ^ x[155]);
    assign layer0_out[5425] = ~(x[386] | x[387]);
    assign layer0_out[5426] = x[6] | x[22];
    assign layer0_out[5427] = x[42];
    assign layer0_out[5428] = x[189];
    assign layer0_out[5429] = ~(x[191] | x[203]);
    assign layer0_out[5430] = ~x[345];
    assign layer0_out[5431] = ~x[71];
    assign layer0_out[5432] = ~(x[49] | x[56]);
    assign layer0_out[5433] = x[310] | x[323];
    assign layer0_out[5434] = ~(x[372] & x[382]);
    assign layer0_out[5435] = ~x[298] | x[293];
    assign layer0_out[5436] = ~x[390];
    assign layer0_out[5437] = x[126];
    assign layer0_out[5438] = x[340] | x[341];
    assign layer0_out[5439] = x[194];
    assign layer0_out[5440] = x[161] | x[167];
    assign layer0_out[5441] = x[240] | x[250];
    assign layer0_out[5442] = ~x[72];
    assign layer0_out[5443] = x[131] & ~x[147];
    assign layer0_out[5444] = ~(x[195] & x[214]);
    assign layer0_out[5445] = ~(x[158] | x[175]);
    assign layer0_out[5446] = ~x[129];
    assign layer0_out[5447] = x[33] & ~x[22];
    assign layer0_out[5448] = x[23] & ~x[17];
    assign layer0_out[5449] = x[148] | x[167];
    assign layer0_out[5450] = 1'b0;
    assign layer0_out[5451] = x[97];
    assign layer0_out[5452] = ~x[325];
    assign layer0_out[5453] = x[204] ^ x[206];
    assign layer0_out[5454] = x[66] ^ x[83];
    assign layer0_out[5455] = x[157] & ~x[161];
    assign layer0_out[5456] = x[75] ^ x[89];
    assign layer0_out[5457] = ~x[135] | x[114];
    assign layer0_out[5458] = x[78] & x[87];
    assign layer0_out[5459] = ~x[271] | x[287];
    assign layer0_out[5460] = ~(x[256] | x[272]);
    assign layer0_out[5461] = x[31];
    assign layer0_out[5462] = x[245] | x[262];
    assign layer0_out[5463] = ~(x[293] ^ x[295]);
    assign layer0_out[5464] = ~(x[162] | x[166]);
    assign layer0_out[5465] = ~(x[363] | x[372]);
    assign layer0_out[5466] = x[54];
    assign layer0_out[5467] = x[35] | x[37];
    assign layer0_out[5468] = x[280] & ~x[273];
    assign layer0_out[5469] = ~(x[303] ^ x[316]);
    assign layer0_out[5470] = x[376] & ~x[371];
    assign layer0_out[5471] = x[362] ^ x[363];
    assign layer0_out[5472] = ~x[257];
    assign layer0_out[5473] = ~(x[192] | x[193]);
    assign layer0_out[5474] = ~(x[372] ^ x[380]);
    assign layer0_out[5475] = ~(x[255] | x[263]);
    assign layer0_out[5476] = ~x[151] | x[130];
    assign layer0_out[5477] = ~x[52];
    assign layer0_out[5478] = x[250] & ~x[244];
    assign layer0_out[5479] = ~(x[297] | x[317]);
    assign layer0_out[5480] = ~x[43] | x[31];
    assign layer0_out[5481] = ~(x[264] ^ x[270]);
    assign layer0_out[5482] = ~x[297];
    assign layer0_out[5483] = ~(x[202] ^ x[209]);
    assign layer0_out[5484] = ~x[206];
    assign layer0_out[5485] = ~(x[302] ^ x[315]);
    assign layer0_out[5486] = x[211] | x[212];
    assign layer0_out[5487] = ~(x[248] & x[259]);
    assign layer0_out[5488] = ~x[75];
    assign layer0_out[5489] = ~x[305] | x[317];
    assign layer0_out[5490] = x[149] & ~x[161];
    assign layer0_out[5491] = ~x[392] | x[398];
    assign layer0_out[5492] = ~(x[82] | x[103]);
    assign layer0_out[5493] = x[115];
    assign layer0_out[5494] = x[109];
    assign layer0_out[5495] = x[130] ^ x[137];
    assign layer0_out[5496] = ~(x[233] & x[238]);
    assign layer0_out[5497] = ~(x[51] | x[63]);
    assign layer0_out[5498] = ~(x[135] | x[144]);
    assign layer0_out[5499] = ~x[26];
    assign layer0_out[5500] = ~(x[379] ^ x[394]);
    assign layer0_out[5501] = x[259] ^ x[274];
    assign layer0_out[5502] = x[39] | x[58];
    assign layer0_out[5503] = x[255] & x[274];
    assign layer0_out[5504] = ~x[30] | x[16];
    assign layer0_out[5505] = x[376] & ~x[393];
    assign layer0_out[5506] = x[341] | x[355];
    assign layer0_out[5507] = ~(x[171] | x[180]);
    assign layer0_out[5508] = x[231];
    assign layer0_out[5509] = x[133];
    assign layer0_out[5510] = x[383] | x[398];
    assign layer0_out[5511] = 1'b0;
    assign layer0_out[5512] = ~x[112] | x[129];
    assign layer0_out[5513] = x[363] | x[371];
    assign layer0_out[5514] = x[259] | x[278];
    assign layer0_out[5515] = ~(x[118] | x[135]);
    assign layer0_out[5516] = ~(x[258] & x[262]);
    assign layer0_out[5517] = x[21] & ~x[38];
    assign layer0_out[5518] = x[168] & ~x[159];
    assign layer0_out[5519] = ~x[266] | x[249];
    assign layer0_out[5520] = x[29] | x[48];
    assign layer0_out[5521] = x[32] & ~x[27];
    assign layer0_out[5522] = x[358] & ~x[357];
    assign layer0_out[5523] = x[337] | x[349];
    assign layer0_out[5524] = ~x[314] | x[319];
    assign layer0_out[5525] = ~(x[302] & x[309]);
    assign layer0_out[5526] = ~(x[138] & x[147]);
    assign layer0_out[5527] = ~(x[246] ^ x[252]);
    assign layer0_out[5528] = ~x[203] | x[192];
    assign layer0_out[5529] = ~x[243];
    assign layer0_out[5530] = x[285] | x[287];
    assign layer0_out[5531] = ~x[75];
    assign layer0_out[5532] = ~x[150];
    assign layer0_out[5533] = ~x[374] | x[380];
    assign layer0_out[5534] = ~(x[106] & x[126]);
    assign layer0_out[5535] = 1'b0;
    assign layer0_out[5536] = x[131] ^ x[132];
    assign layer0_out[5537] = x[102];
    assign layer0_out[5538] = ~(x[385] | x[391]);
    assign layer0_out[5539] = x[341] & x[359];
    assign layer0_out[5540] = x[379] & ~x[376];
    assign layer0_out[5541] = x[37] & ~x[41];
    assign layer0_out[5542] = x[282] | x[289];
    assign layer0_out[5543] = x[264];
    assign layer0_out[5544] = ~(x[68] | x[77]);
    assign layer0_out[5545] = 1'b0;
    assign layer0_out[5546] = x[67];
    assign layer0_out[5547] = ~(x[370] | x[388]);
    assign layer0_out[5548] = ~(x[262] ^ x[279]);
    assign layer0_out[5549] = 1'b1;
    assign layer0_out[5550] = x[330] | x[342];
    assign layer0_out[5551] = x[268] & ~x[285];
    assign layer0_out[5552] = ~(x[7] ^ x[27]);
    assign layer0_out[5553] = x[84] ^ x[86];
    assign layer0_out[5554] = ~x[133];
    assign layer0_out[5555] = ~x[380] | x[382];
    assign layer0_out[5556] = x[203];
    assign layer0_out[5557] = ~x[122] | x[110];
    assign layer0_out[5558] = ~(x[98] ^ x[111]);
    assign layer0_out[5559] = x[339] | x[353];
    assign layer0_out[5560] = x[140] & ~x[134];
    assign layer0_out[5561] = ~x[269] | x[260];
    assign layer0_out[5562] = x[106] & ~x[120];
    assign layer0_out[5563] = ~x[381];
    assign layer0_out[5564] = x[51] & ~x[59];
    assign layer0_out[5565] = ~(x[225] ^ x[242]);
    assign layer0_out[5566] = x[152] ^ x[158];
    assign layer0_out[5567] = ~x[229] | x[245];
    assign layer0_out[5568] = x[136];
    assign layer0_out[5569] = ~(x[219] ^ x[226]);
    assign layer0_out[5570] = x[377] & ~x[391];
    assign layer0_out[5571] = x[283] & x[300];
    assign layer0_out[5572] = x[232] ^ x[241];
    assign layer0_out[5573] = ~x[204];
    assign layer0_out[5574] = ~(x[84] | x[93]);
    assign layer0_out[5575] = x[210] | x[226];
    assign layer0_out[5576] = ~(x[332] | x[337]);
    assign layer0_out[5577] = x[68] & ~x[89];
    assign layer0_out[5578] = ~(x[117] | x[134]);
    assign layer0_out[5579] = x[252] | x[259];
    assign layer0_out[5580] = x[85];
    assign layer0_out[5581] = ~x[111];
    assign layer0_out[5582] = ~x[320] | x[330];
    assign layer0_out[5583] = ~(x[128] ^ x[145]);
    assign layer0_out[5584] = x[372] | x[384];
    assign layer0_out[5585] = x[144];
    assign layer0_out[5586] = ~(x[253] | x[269]);
    assign layer0_out[5587] = ~(x[242] ^ x[253]);
    assign layer0_out[5588] = ~(x[146] | x[163]);
    assign layer0_out[5589] = ~(x[111] | x[127]);
    assign layer0_out[5590] = x[151] | x[161];
    assign layer0_out[5591] = x[310] & ~x[291];
    assign layer0_out[5592] = ~(x[339] | x[342]);
    assign layer0_out[5593] = x[5] & x[20];
    assign layer0_out[5594] = ~x[23] | x[22];
    assign layer0_out[5595] = 1'b0;
    assign layer0_out[5596] = ~x[243] | x[228];
    assign layer0_out[5597] = x[23] | x[26];
    assign layer0_out[5598] = ~x[22] | x[10];
    assign layer0_out[5599] = x[203];
    assign layer0_out[5600] = x[1];
    assign layer0_out[5601] = x[80] | x[101];
    assign layer0_out[5602] = ~(x[316] | x[335]);
    assign layer0_out[5603] = ~(x[333] | x[353]);
    assign layer0_out[5604] = x[97] ^ x[105];
    assign layer0_out[5605] = x[317];
    assign layer0_out[5606] = 1'b1;
    assign layer0_out[5607] = x[256] & ~x[258];
    assign layer0_out[5608] = ~(x[208] ^ x[221]);
    assign layer0_out[5609] = ~x[74] | x[93];
    assign layer0_out[5610] = x[258] ^ x[276];
    assign layer0_out[5611] = ~(x[271] | x[273]);
    assign layer0_out[5612] = ~x[286];
    assign layer0_out[5613] = x[92] | x[111];
    assign layer0_out[5614] = ~x[80] | x[77];
    assign layer0_out[5615] = x[188] & ~x[171];
    assign layer0_out[5616] = x[51];
    assign layer0_out[5617] = ~(x[70] | x[74]);
    assign layer0_out[5618] = ~x[198];
    assign layer0_out[5619] = ~(x[35] ^ x[55]);
    assign layer0_out[5620] = x[10] & ~x[12];
    assign layer0_out[5621] = ~x[236] | x[246];
    assign layer0_out[5622] = x[56] | x[62];
    assign layer0_out[5623] = x[278] | x[282];
    assign layer0_out[5624] = x[375] | x[392];
    assign layer0_out[5625] = x[275];
    assign layer0_out[5626] = ~x[192];
    assign layer0_out[5627] = ~(x[4] & x[6]);
    assign layer0_out[5628] = ~x[7];
    assign layer0_out[5629] = x[319] | x[333];
    assign layer0_out[5630] = x[364] & ~x[378];
    assign layer0_out[5631] = ~(x[289] & x[291]);
    assign layer0_out[5632] = x[366] & x[371];
    assign layer0_out[5633] = ~(x[148] | x[165]);
    assign layer0_out[5634] = ~(x[310] & x[320]);
    assign layer0_out[5635] = x[101] & ~x[82];
    assign layer0_out[5636] = ~(x[177] | x[186]);
    assign layer0_out[5637] = ~(x[275] | x[293]);
    assign layer0_out[5638] = x[212] & ~x[223];
    assign layer0_out[5639] = ~(x[1] | x[3]);
    assign layer0_out[5640] = x[367] | x[380];
    assign layer0_out[5641] = x[88] | x[108];
    assign layer0_out[5642] = x[163] & x[167];
    assign layer0_out[5643] = x[388];
    assign layer0_out[5644] = 1'b0;
    assign layer0_out[5645] = x[300] | x[308];
    assign layer0_out[5646] = ~x[55];
    assign layer0_out[5647] = x[194] & x[206];
    assign layer0_out[5648] = x[387] | x[390];
    assign layer0_out[5649] = ~(x[308] ^ x[326]);
    assign layer0_out[5650] = x[331];
    assign layer0_out[5651] = ~x[42];
    assign layer0_out[5652] = x[361] & ~x[343];
    assign layer0_out[5653] = ~(x[286] | x[303]);
    assign layer0_out[5654] = 1'b0;
    assign layer0_out[5655] = x[42] & x[57];
    assign layer0_out[5656] = ~(x[306] | x[309]);
    assign layer0_out[5657] = x[82] & x[93];
    assign layer0_out[5658] = 1'b1;
    assign layer0_out[5659] = x[205] | x[223];
    assign layer0_out[5660] = x[163] & ~x[148];
    assign layer0_out[5661] = x[273];
    assign layer0_out[5662] = ~x[220];
    assign layer0_out[5663] = ~(x[37] & x[39]);
    assign layer0_out[5664] = ~(x[168] & x[175]);
    assign layer0_out[5665] = x[149] ^ x[168];
    assign layer0_out[5666] = ~x[38] | x[35];
    assign layer0_out[5667] = ~x[163] | x[144];
    assign layer0_out[5668] = x[22] | x[42];
    assign layer0_out[5669] = 1'b1;
    assign layer0_out[5670] = ~(x[121] | x[123]);
    assign layer0_out[5671] = x[226] & ~x[213];
    assign layer0_out[5672] = x[151] & ~x[162];
    assign layer0_out[5673] = x[71] | x[80];
    assign layer0_out[5674] = x[191] & ~x[175];
    assign layer0_out[5675] = x[152];
    assign layer0_out[5676] = x[186] & x[192];
    assign layer0_out[5677] = x[124];
    assign layer0_out[5678] = ~(x[195] | x[215]);
    assign layer0_out[5679] = ~x[43];
    assign layer0_out[5680] = ~(x[163] ^ x[183]);
    assign layer0_out[5681] = ~x[267] | x[254];
    assign layer0_out[5682] = ~(x[64] & x[78]);
    assign layer0_out[5683] = x[376] & ~x[388];
    assign layer0_out[5684] = ~(x[205] | x[206]);
    assign layer0_out[5685] = x[143];
    assign layer0_out[5686] = x[59];
    assign layer0_out[5687] = ~x[162];
    assign layer0_out[5688] = ~x[194];
    assign layer0_out[5689] = x[219] ^ x[237];
    assign layer0_out[5690] = ~(x[324] | x[330]);
    assign layer0_out[5691] = x[133] & ~x[153];
    assign layer0_out[5692] = ~(x[115] | x[135]);
    assign layer0_out[5693] = ~(x[336] | x[342]);
    assign layer0_out[5694] = x[230];
    assign layer0_out[5695] = x[208];
    assign layer0_out[5696] = ~(x[322] ^ x[323]);
    assign layer0_out[5697] = x[268] & x[283];
    assign layer0_out[5698] = ~(x[126] & x[147]);
    assign layer0_out[5699] = x[257] ^ x[264];
    assign layer0_out[5700] = x[186] & x[206];
    assign layer0_out[5701] = ~x[331];
    assign layer0_out[5702] = ~x[243];
    assign layer0_out[5703] = x[368];
    assign layer0_out[5704] = ~(x[108] & x[117]);
    assign layer0_out[5705] = x[195] | x[212];
    assign layer0_out[5706] = 1'b1;
    assign layer0_out[5707] = x[60] & ~x[66];
    assign layer0_out[5708] = x[217] & x[223];
    assign layer0_out[5709] = x[98] | x[109];
    assign layer0_out[5710] = ~(x[223] | x[234]);
    assign layer0_out[5711] = x[306];
    assign layer0_out[5712] = x[90] | x[105];
    assign layer0_out[5713] = ~(x[171] ^ x[179]);
    assign layer0_out[5714] = ~x[329];
    assign layer0_out[5715] = ~(x[328] ^ x[348]);
    assign layer0_out[5716] = x[144];
    assign layer0_out[5717] = x[177] & x[195];
    assign layer0_out[5718] = ~x[67];
    assign layer0_out[5719] = ~(x[0] ^ x[3]);
    assign layer0_out[5720] = ~(x[305] & x[319]);
    assign layer0_out[5721] = x[21] ^ x[32];
    assign layer0_out[5722] = ~(x[224] | x[242]);
    assign layer0_out[5723] = ~x[162];
    assign layer0_out[5724] = 1'b0;
    assign layer0_out[5725] = 1'b0;
    assign layer0_out[5726] = ~x[325];
    assign layer0_out[5727] = x[292] | x[303];
    assign layer0_out[5728] = x[244] & ~x[259];
    assign layer0_out[5729] = ~x[71];
    assign layer0_out[5730] = x[12] & ~x[1];
    assign layer0_out[5731] = x[158];
    assign layer0_out[5732] = x[129] | x[139];
    assign layer0_out[5733] = x[277] | x[296];
    assign layer0_out[5734] = ~(x[149] | x[151]);
    assign layer0_out[5735] = 1'b0;
    assign layer0_out[5736] = ~x[313];
    assign layer0_out[5737] = ~x[21] | x[28];
    assign layer0_out[5738] = x[160] ^ x[164];
    assign layer0_out[5739] = ~(x[45] | x[65]);
    assign layer0_out[5740] = x[186] | x[194];
    assign layer0_out[5741] = 1'b0;
    assign layer0_out[5742] = x[287];
    assign layer0_out[5743] = x[65];
    assign layer0_out[5744] = x[87];
    assign layer0_out[5745] = x[27];
    assign layer0_out[5746] = x[75] & ~x[69];
    assign layer0_out[5747] = ~x[93];
    assign layer0_out[5748] = x[70] & ~x[61];
    assign layer0_out[5749] = x[229];
    assign layer0_out[5750] = ~x[58] | x[47];
    assign layer0_out[5751] = x[71] & x[88];
    assign layer0_out[5752] = ~(x[279] & x[287]);
    assign layer0_out[5753] = x[142] & ~x[149];
    assign layer0_out[5754] = ~(x[2] | x[23]);
    assign layer0_out[5755] = x[19];
    assign layer0_out[5756] = ~(x[49] & x[51]);
    assign layer0_out[5757] = x[315] ^ x[325];
    assign layer0_out[5758] = x[121] | x[125];
    assign layer0_out[5759] = 1'b1;
    assign layer0_out[5760] = ~x[232] | x[235];
    assign layer0_out[5761] = ~x[144];
    assign layer0_out[5762] = ~x[27];
    assign layer0_out[5763] = ~x[289];
    assign layer0_out[5764] = 1'b0;
    assign layer0_out[5765] = 1'b0;
    assign layer0_out[5766] = x[269] & ~x[254];
    assign layer0_out[5767] = ~(x[377] | x[379]);
    assign layer0_out[5768] = x[105];
    assign layer0_out[5769] = x[162] | x[163];
    assign layer0_out[5770] = ~(x[89] & x[96]);
    assign layer0_out[5771] = x[130];
    assign layer0_out[5772] = x[15] & ~x[9];
    assign layer0_out[5773] = x[90];
    assign layer0_out[5774] = ~x[38] | x[40];
    assign layer0_out[5775] = x[98];
    assign layer0_out[5776] = x[373] & ~x[386];
    assign layer0_out[5777] = ~x[351] | x[359];
    assign layer0_out[5778] = x[247] & ~x[255];
    assign layer0_out[5779] = x[175] & x[179];
    assign layer0_out[5780] = x[161] | x[164];
    assign layer0_out[5781] = ~x[247];
    assign layer0_out[5782] = ~x[277];
    assign layer0_out[5783] = ~(x[285] ^ x[295]);
    assign layer0_out[5784] = ~x[133] | x[124];
    assign layer0_out[5785] = x[278];
    assign layer0_out[5786] = x[42] | x[50];
    assign layer0_out[5787] = x[240] | x[257];
    assign layer0_out[5788] = ~(x[92] ^ x[95]);
    assign layer0_out[5789] = 1'b1;
    assign layer0_out[5790] = 1'b0;
    assign layer0_out[5791] = ~x[34];
    assign layer0_out[5792] = x[92];
    assign layer0_out[5793] = 1'b0;
    assign layer0_out[5794] = x[67] & ~x[73];
    assign layer0_out[5795] = x[290] | x[310];
    assign layer0_out[5796] = x[380] & ~x[383];
    assign layer0_out[5797] = x[340] | x[360];
    assign layer0_out[5798] = ~x[274];
    assign layer0_out[5799] = x[186] ^ x[193];
    assign layer0_out[5800] = ~x[105] | x[109];
    assign layer0_out[5801] = x[173] | x[180];
    assign layer0_out[5802] = x[363];
    assign layer0_out[5803] = x[198];
    assign layer0_out[5804] = x[333];
    assign layer0_out[5805] = x[150];
    assign layer0_out[5806] = ~x[186] | x[165];
    assign layer0_out[5807] = x[394];
    assign layer0_out[5808] = x[71] & ~x[68];
    assign layer0_out[5809] = ~(x[103] ^ x[108]);
    assign layer0_out[5810] = x[109] & ~x[95];
    assign layer0_out[5811] = ~(x[279] ^ x[297]);
    assign layer0_out[5812] = x[203];
    assign layer0_out[5813] = x[297] | x[314];
    assign layer0_out[5814] = x[195] | x[199];
    assign layer0_out[5815] = x[54] & ~x[41];
    assign layer0_out[5816] = x[21] | x[22];
    assign layer0_out[5817] = x[97] | x[102];
    assign layer0_out[5818] = ~x[340] | x[327];
    assign layer0_out[5819] = 1'b1;
    assign layer0_out[5820] = ~(x[112] | x[117]);
    assign layer0_out[5821] = x[4] & x[10];
    assign layer0_out[5822] = x[151] | x[168];
    assign layer0_out[5823] = x[170];
    assign layer0_out[5824] = ~(x[331] & x[343]);
    assign layer0_out[5825] = ~x[389] | x[373];
    assign layer0_out[5826] = x[61];
    assign layer0_out[5827] = x[23] ^ x[27];
    assign layer0_out[5828] = ~(x[378] | x[392]);
    assign layer0_out[5829] = ~x[236] | x[232];
    assign layer0_out[5830] = ~(x[212] ^ x[228]);
    assign layer0_out[5831] = x[317] | x[329];
    assign layer0_out[5832] = x[254] | x[272];
    assign layer0_out[5833] = x[106];
    assign layer0_out[5834] = ~x[191];
    assign layer0_out[5835] = ~(x[305] | x[322]);
    assign layer0_out[5836] = x[5];
    assign layer0_out[5837] = ~(x[62] | x[81]);
    assign layer0_out[5838] = ~x[321];
    assign layer0_out[5839] = x[278];
    assign layer0_out[5840] = ~x[41];
    assign layer0_out[5841] = ~x[289];
    assign layer0_out[5842] = x[34] | x[49];
    assign layer0_out[5843] = x[106] & x[112];
    assign layer0_out[5844] = x[79] & ~x[85];
    assign layer0_out[5845] = x[51];
    assign layer0_out[5846] = x[319] ^ x[324];
    assign layer0_out[5847] = x[301];
    assign layer0_out[5848] = x[178] ^ x[187];
    assign layer0_out[5849] = x[236];
    assign layer0_out[5850] = x[209] & ~x[199];
    assign layer0_out[5851] = x[237] & x[242];
    assign layer0_out[5852] = ~x[169] | x[177];
    assign layer0_out[5853] = ~x[221] | x[209];
    assign layer0_out[5854] = x[398] & ~x[396];
    assign layer0_out[5855] = x[59] & ~x[55];
    assign layer0_out[5856] = ~(x[322] ^ x[339]);
    assign layer0_out[5857] = ~x[51];
    assign layer0_out[5858] = x[241] | x[253];
    assign layer0_out[5859] = 1'b1;
    assign layer0_out[5860] = x[171];
    assign layer0_out[5861] = 1'b1;
    assign layer0_out[5862] = ~(x[132] ^ x[134]);
    assign layer0_out[5863] = x[7];
    assign layer0_out[5864] = 1'b0;
    assign layer0_out[5865] = x[16] | x[20];
    assign layer0_out[5866] = 1'b0;
    assign layer0_out[5867] = ~x[368] | x[380];
    assign layer0_out[5868] = ~x[22];
    assign layer0_out[5869] = x[50] | x[54];
    assign layer0_out[5870] = ~x[241] | x[226];
    assign layer0_out[5871] = x[18] & x[21];
    assign layer0_out[5872] = ~x[334] | x[320];
    assign layer0_out[5873] = x[347] ^ x[359];
    assign layer0_out[5874] = x[184];
    assign layer0_out[5875] = x[21];
    assign layer0_out[5876] = ~(x[126] | x[141]);
    assign layer0_out[5877] = x[327] & ~x[332];
    assign layer0_out[5878] = ~(x[158] | x[160]);
    assign layer0_out[5879] = ~(x[86] | x[106]);
    assign layer0_out[5880] = ~(x[89] | x[102]);
    assign layer0_out[5881] = x[365];
    assign layer0_out[5882] = ~x[269] | x[278];
    assign layer0_out[5883] = ~x[74] | x[84];
    assign layer0_out[5884] = ~x[41] | x[60];
    assign layer0_out[5885] = ~(x[210] | x[211]);
    assign layer0_out[5886] = x[232] & ~x[238];
    assign layer0_out[5887] = x[334] | x[352];
    assign layer0_out[5888] = x[338] & ~x[329];
    assign layer0_out[5889] = ~x[261];
    assign layer0_out[5890] = ~(x[32] | x[42]);
    assign layer0_out[5891] = 1'b0;
    assign layer0_out[5892] = 1'b0;
    assign layer0_out[5893] = x[223] & ~x[235];
    assign layer0_out[5894] = x[81] & ~x[90];
    assign layer0_out[5895] = ~x[158] | x[165];
    assign layer0_out[5896] = x[14] & ~x[31];
    assign layer0_out[5897] = x[63];
    assign layer0_out[5898] = x[153] | x[167];
    assign layer0_out[5899] = 1'b0;
    assign layer0_out[5900] = ~x[137];
    assign layer0_out[5901] = 1'b0;
    assign layer0_out[5902] = ~x[323];
    assign layer0_out[5903] = x[197] | x[200];
    assign layer0_out[5904] = x[234] ^ x[239];
    assign layer0_out[5905] = x[275] | x[277];
    assign layer0_out[5906] = x[9];
    assign layer0_out[5907] = x[261];
    assign layer0_out[5908] = ~(x[84] & x[103]);
    assign layer0_out[5909] = ~x[85] | x[66];
    assign layer0_out[5910] = ~x[398] | x[380];
    assign layer0_out[5911] = x[368] | x[375];
    assign layer0_out[5912] = ~x[372] | x[378];
    assign layer0_out[5913] = x[376] ^ x[390];
    assign layer0_out[5914] = ~x[6];
    assign layer0_out[5915] = x[69] & ~x[48];
    assign layer0_out[5916] = x[213];
    assign layer0_out[5917] = x[93];
    assign layer0_out[5918] = x[354] ^ x[370];
    assign layer0_out[5919] = ~x[112];
    assign layer0_out[5920] = x[193];
    assign layer0_out[5921] = ~(x[141] & x[162]);
    assign layer0_out[5922] = x[201];
    assign layer0_out[5923] = ~(x[291] | x[304]);
    assign layer0_out[5924] = ~x[254] | x[255];
    assign layer0_out[5925] = ~x[102] | x[107];
    assign layer0_out[5926] = ~(x[83] ^ x[85]);
    assign layer0_out[5927] = ~(x[326] & x[334]);
    assign layer0_out[5928] = x[149] & ~x[136];
    assign layer0_out[5929] = x[396];
    assign layer0_out[5930] = x[117] ^ x[119];
    assign layer0_out[5931] = ~(x[48] & x[62]);
    assign layer0_out[5932] = x[241] & x[250];
    assign layer0_out[5933] = x[282] ^ x[286];
    assign layer0_out[5934] = ~x[334] | x[324];
    assign layer0_out[5935] = x[15] & ~x[31];
    assign layer0_out[5936] = x[12] & ~x[31];
    assign layer0_out[5937] = x[268] | x[282];
    assign layer0_out[5938] = ~(x[221] | x[222]);
    assign layer0_out[5939] = x[26];
    assign layer0_out[5940] = 1'b0;
    assign layer0_out[5941] = x[377] ^ x[395];
    assign layer0_out[5942] = ~(x[184] | x[194]);
    assign layer0_out[5943] = x[13];
    assign layer0_out[5944] = ~x[95];
    assign layer0_out[5945] = ~x[287];
    assign layer0_out[5946] = ~(x[10] & x[28]);
    assign layer0_out[5947] = x[25] | x[34];
    assign layer0_out[5948] = ~x[184];
    assign layer0_out[5949] = ~x[145];
    assign layer0_out[5950] = x[278] | x[280];
    assign layer0_out[5951] = x[320] | x[323];
    assign layer0_out[5952] = ~x[365] | x[349];
    assign layer0_out[5953] = x[252];
    assign layer0_out[5954] = x[185] | x[191];
    assign layer0_out[5955] = 1'b1;
    assign layer0_out[5956] = ~x[349];
    assign layer0_out[5957] = ~x[356];
    assign layer0_out[5958] = x[329];
    assign layer0_out[5959] = ~x[368];
    assign layer0_out[5960] = ~(x[311] | x[320]);
    assign layer0_out[5961] = ~(x[155] & x[158]);
    assign layer0_out[5962] = ~(x[146] | x[147]);
    assign layer0_out[5963] = ~(x[164] & x[168]);
    assign layer0_out[5964] = x[141];
    assign layer0_out[5965] = 1'b0;
    assign layer0_out[5966] = ~x[192] | x[185];
    assign layer0_out[5967] = ~(x[158] | x[167]);
    assign layer0_out[5968] = ~x[253];
    assign layer0_out[5969] = ~x[311] | x[312];
    assign layer0_out[5970] = ~(x[123] | x[137]);
    assign layer0_out[5971] = x[178] & ~x[192];
    assign layer0_out[5972] = ~(x[75] ^ x[90]);
    assign layer0_out[5973] = ~(x[117] | x[137]);
    assign layer0_out[5974] = ~x[386] | x[383];
    assign layer0_out[5975] = x[192] & ~x[204];
    assign layer0_out[5976] = x[226] | x[227];
    assign layer0_out[5977] = ~x[94];
    assign layer0_out[5978] = ~x[237] | x[246];
    assign layer0_out[5979] = ~x[369];
    assign layer0_out[5980] = ~(x[12] & x[33]);
    assign layer0_out[5981] = ~(x[334] | x[350]);
    assign layer0_out[5982] = x[132] & x[152];
    assign layer0_out[5983] = x[282] & x[292];
    assign layer0_out[5984] = ~x[373];
    assign layer0_out[5985] = x[265] | x[273];
    assign layer0_out[5986] = x[163] | x[184];
    assign layer0_out[5987] = ~x[169];
    assign layer0_out[5988] = x[145] & ~x[130];
    assign layer0_out[5989] = x[354];
    assign layer0_out[5990] = ~x[29] | x[38];
    assign layer0_out[5991] = 1'b1;
    assign layer0_out[5992] = x[242];
    assign layer0_out[5993] = x[372];
    assign layer0_out[5994] = 1'b0;
    assign layer0_out[5995] = ~(x[134] ^ x[150]);
    assign layer0_out[5996] = ~x[272] | x[267];
    assign layer0_out[5997] = x[264] | x[271];
    assign layer0_out[5998] = x[72];
    assign layer0_out[5999] = x[82] & ~x[74];
    assign layer0_out[6000] = x[362] & ~x[344];
    assign layer0_out[6001] = x[245] & x[264];
    assign layer0_out[6002] = ~x[309];
    assign layer0_out[6003] = x[200] & x[213];
    assign layer0_out[6004] = ~x[133];
    assign layer0_out[6005] = ~(x[240] | x[259]);
    assign layer0_out[6006] = 1'b0;
    assign layer0_out[6007] = ~x[286];
    assign layer0_out[6008] = x[75] | x[78];
    assign layer0_out[6009] = x[58] | x[76];
    assign layer0_out[6010] = x[73];
    assign layer0_out[6011] = x[68] | x[79];
    assign layer0_out[6012] = ~x[38];
    assign layer0_out[6013] = x[79] | x[96];
    assign layer0_out[6014] = x[17] | x[36];
    assign layer0_out[6015] = x[161] ^ x[181];
    assign layer0_out[6016] = x[321] | x[325];
    assign layer0_out[6017] = x[333] | x[351];
    assign layer0_out[6018] = ~x[102] | x[92];
    assign layer0_out[6019] = x[227] & ~x[233];
    assign layer0_out[6020] = ~x[248];
    assign layer0_out[6021] = x[274];
    assign layer0_out[6022] = x[56] & x[68];
    assign layer0_out[6023] = x[366] | x[382];
    assign layer0_out[6024] = ~(x[157] | x[166]);
    assign layer0_out[6025] = 1'b0;
    assign layer0_out[6026] = 1'b0;
    assign layer0_out[6027] = ~(x[133] | x[143]);
    assign layer0_out[6028] = ~x[123];
    assign layer0_out[6029] = 1'b1;
    assign layer0_out[6030] = x[126] | x[127];
    assign layer0_out[6031] = 1'b0;
    assign layer0_out[6032] = ~(x[129] ^ x[145]);
    assign layer0_out[6033] = ~(x[128] | x[136]);
    assign layer0_out[6034] = x[22];
    assign layer0_out[6035] = ~(x[327] | x[337]);
    assign layer0_out[6036] = ~x[324];
    assign layer0_out[6037] = x[377] & ~x[364];
    assign layer0_out[6038] = x[261] ^ x[263];
    assign layer0_out[6039] = ~x[373];
    assign layer0_out[6040] = ~(x[34] & x[50]);
    assign layer0_out[6041] = x[28] ^ x[46];
    assign layer0_out[6042] = x[103] | x[121];
    assign layer0_out[6043] = ~x[163];
    assign layer0_out[6044] = ~x[129];
    assign layer0_out[6045] = ~(x[292] & x[310]);
    assign layer0_out[6046] = x[357];
    assign layer0_out[6047] = x[372];
    assign layer0_out[6048] = ~(x[281] ^ x[286]);
    assign layer0_out[6049] = ~(x[129] | x[137]);
    assign layer0_out[6050] = x[8];
    assign layer0_out[6051] = x[236] | x[254];
    assign layer0_out[6052] = 1'b0;
    assign layer0_out[6053] = ~(x[26] | x[45]);
    assign layer0_out[6054] = x[227] & ~x[232];
    assign layer0_out[6055] = x[77] ^ x[95];
    assign layer0_out[6056] = ~x[11];
    assign layer0_out[6057] = ~(x[4] | x[18]);
    assign layer0_out[6058] = x[358] | x[376];
    assign layer0_out[6059] = ~x[309] | x[304];
    assign layer0_out[6060] = ~(x[245] & x[257]);
    assign layer0_out[6061] = x[343];
    assign layer0_out[6062] = x[21] ^ x[31];
    assign layer0_out[6063] = ~x[229] | x[235];
    assign layer0_out[6064] = ~(x[59] & x[66]);
    assign layer0_out[6065] = ~(x[326] & x[331]);
    assign layer0_out[6066] = x[393];
    assign layer0_out[6067] = ~(x[326] | x[344]);
    assign layer0_out[6068] = ~x[139];
    assign layer0_out[6069] = ~(x[174] ^ x[176]);
    assign layer0_out[6070] = x[19] & ~x[11];
    assign layer0_out[6071] = x[118] ^ x[129];
    assign layer0_out[6072] = x[3] | x[19];
    assign layer0_out[6073] = ~x[55];
    assign layer0_out[6074] = ~(x[318] | x[332]);
    assign layer0_out[6075] = x[66] | x[86];
    assign layer0_out[6076] = x[199] ^ x[212];
    assign layer0_out[6077] = x[84] | x[105];
    assign layer0_out[6078] = x[128] & x[149];
    assign layer0_out[6079] = ~(x[86] ^ x[89]);
    assign layer0_out[6080] = x[206] | x[226];
    assign layer0_out[6081] = ~(x[76] ^ x[90]);
    assign layer0_out[6082] = ~x[317] | x[333];
    assign layer0_out[6083] = x[199] & ~x[198];
    assign layer0_out[6084] = ~(x[322] | x[327]);
    assign layer0_out[6085] = ~(x[120] ^ x[131]);
    assign layer0_out[6086] = ~x[286];
    assign layer0_out[6087] = x[321] & ~x[302];
    assign layer0_out[6088] = ~(x[68] ^ x[72]);
    assign layer0_out[6089] = ~x[351];
    assign layer0_out[6090] = ~x[16] | x[33];
    assign layer0_out[6091] = ~(x[363] & x[368]);
    assign layer0_out[6092] = ~x[325];
    assign layer0_out[6093] = ~x[353] | x[361];
    assign layer0_out[6094] = x[302] ^ x[319];
    assign layer0_out[6095] = x[35] & x[36];
    assign layer0_out[6096] = ~(x[298] | x[313]);
    assign layer0_out[6097] = ~x[171] | x[176];
    assign layer0_out[6098] = x[14] | x[32];
    assign layer0_out[6099] = 1'b1;
    assign layer0_out[6100] = x[0] | x[12];
    assign layer0_out[6101] = 1'b0;
    assign layer0_out[6102] = ~(x[196] | x[200]);
    assign layer0_out[6103] = x[352] & x[371];
    assign layer0_out[6104] = ~(x[21] | x[30]);
    assign layer0_out[6105] = x[127];
    assign layer0_out[6106] = x[108];
    assign layer0_out[6107] = ~x[196];
    assign layer0_out[6108] = ~(x[218] ^ x[229]);
    assign layer0_out[6109] = x[100] & ~x[85];
    assign layer0_out[6110] = x[320];
    assign layer0_out[6111] = ~x[209] | x[198];
    assign layer0_out[6112] = ~(x[329] & x[348]);
    assign layer0_out[6113] = ~x[7];
    assign layer0_out[6114] = ~(x[236] | x[240]);
    assign layer0_out[6115] = x[102] | x[104];
    assign layer0_out[6116] = ~x[161];
    assign layer0_out[6117] = x[350] | x[353];
    assign layer0_out[6118] = ~x[236];
    assign layer0_out[6119] = ~(x[334] ^ x[342]);
    assign layer0_out[6120] = x[391];
    assign layer0_out[6121] = x[106];
    assign layer0_out[6122] = x[41] & ~x[30];
    assign layer0_out[6123] = x[314] | x[325];
    assign layer0_out[6124] = ~(x[6] | x[16]);
    assign layer0_out[6125] = ~x[183];
    assign layer0_out[6126] = ~x[305] | x[314];
    assign layer0_out[6127] = x[31];
    assign layer0_out[6128] = x[69] & ~x[53];
    assign layer0_out[6129] = ~(x[19] | x[35]);
    assign layer0_out[6130] = x[346] | x[362];
    assign layer0_out[6131] = ~x[368];
    assign layer0_out[6132] = x[389] & ~x[369];
    assign layer0_out[6133] = x[136] | x[140];
    assign layer0_out[6134] = x[391] & ~x[399];
    assign layer0_out[6135] = ~x[106] | x[127];
    assign layer0_out[6136] = x[209];
    assign layer0_out[6137] = 1'b1;
    assign layer0_out[6138] = ~(x[348] ^ x[358]);
    assign layer0_out[6139] = ~x[378] | x[376];
    assign layer0_out[6140] = x[274] | x[275];
    assign layer0_out[6141] = ~x[335];
    assign layer0_out[6142] = ~x[293];
    assign layer0_out[6143] = ~x[187];
    assign layer0_out[6144] = ~x[127];
    assign layer0_out[6145] = ~x[121] | x[111];
    assign layer0_out[6146] = ~(x[50] | x[70]);
    assign layer0_out[6147] = x[367];
    assign layer0_out[6148] = ~(x[312] & x[318]);
    assign layer0_out[6149] = x[324];
    assign layer0_out[6150] = x[49] ^ x[52];
    assign layer0_out[6151] = x[165];
    assign layer0_out[6152] = ~x[144] | x[151];
    assign layer0_out[6153] = ~(x[258] ^ x[261]);
    assign layer0_out[6154] = x[213] | x[229];
    assign layer0_out[6155] = ~(x[373] | x[381]);
    assign layer0_out[6156] = ~x[59];
    assign layer0_out[6157] = x[63] & x[77];
    assign layer0_out[6158] = ~(x[354] ^ x[367]);
    assign layer0_out[6159] = ~(x[261] | x[265]);
    assign layer0_out[6160] = ~(x[366] ^ x[374]);
    assign layer0_out[6161] = ~x[27] | x[46];
    assign layer0_out[6162] = 1'b1;
    assign layer0_out[6163] = ~(x[281] | x[283]);
    assign layer0_out[6164] = x[90];
    assign layer0_out[6165] = x[26];
    assign layer0_out[6166] = x[35] & ~x[14];
    assign layer0_out[6167] = x[235] & x[239];
    assign layer0_out[6168] = x[361];
    assign layer0_out[6169] = x[96] | x[102];
    assign layer0_out[6170] = ~(x[104] | x[118]);
    assign layer0_out[6171] = ~x[178];
    assign layer0_out[6172] = ~x[87] | x[84];
    assign layer0_out[6173] = x[189] & ~x[190];
    assign layer0_out[6174] = x[260] | x[264];
    assign layer0_out[6175] = x[228] & x[232];
    assign layer0_out[6176] = x[225];
    assign layer0_out[6177] = x[277] | x[282];
    assign layer0_out[6178] = x[274];
    assign layer0_out[6179] = x[110];
    assign layer0_out[6180] = ~(x[38] & x[42]);
    assign layer0_out[6181] = ~(x[49] & x[53]);
    assign layer0_out[6182] = ~x[18];
    assign layer0_out[6183] = 1'b0;
    assign layer0_out[6184] = x[234];
    assign layer0_out[6185] = ~(x[275] | x[295]);
    assign layer0_out[6186] = x[236] | x[239];
    assign layer0_out[6187] = x[40];
    assign layer0_out[6188] = x[227];
    assign layer0_out[6189] = ~x[265];
    assign layer0_out[6190] = ~x[352];
    assign layer0_out[6191] = ~(x[144] | x[162]);
    assign layer0_out[6192] = x[57] ^ x[77];
    assign layer0_out[6193] = x[321];
    assign layer0_out[6194] = 1'b0;
    assign layer0_out[6195] = x[297] | x[308];
    assign layer0_out[6196] = x[243] | x[248];
    assign layer0_out[6197] = x[181] | x[186];
    assign layer0_out[6198] = ~(x[81] | x[100]);
    assign layer0_out[6199] = ~x[25];
    assign layer0_out[6200] = ~(x[100] | x[111]);
    assign layer0_out[6201] = ~x[109];
    assign layer0_out[6202] = x[51];
    assign layer0_out[6203] = ~x[169] | x[178];
    assign layer0_out[6204] = ~x[245] | x[236];
    assign layer0_out[6205] = ~(x[232] | x[247]);
    assign layer0_out[6206] = ~x[158] | x[151];
    assign layer0_out[6207] = ~x[49];
    assign layer0_out[6208] = 1'b1;
    assign layer0_out[6209] = x[110] & ~x[123];
    assign layer0_out[6210] = x[325] | x[344];
    assign layer0_out[6211] = x[233] & ~x[232];
    assign layer0_out[6212] = ~(x[294] ^ x[298]);
    assign layer0_out[6213] = x[150];
    assign layer0_out[6214] = x[137];
    assign layer0_out[6215] = 1'b0;
    assign layer0_out[6216] = x[8] & ~x[16];
    assign layer0_out[6217] = x[343] | x[353];
    assign layer0_out[6218] = x[36] & ~x[47];
    assign layer0_out[6219] = ~x[106] | x[118];
    assign layer0_out[6220] = x[234];
    assign layer0_out[6221] = x[69];
    assign layer0_out[6222] = ~(x[126] ^ x[138]);
    assign layer0_out[6223] = ~(x[4] & x[14]);
    assign layer0_out[6224] = x[45] & x[61];
    assign layer0_out[6225] = x[396];
    assign layer0_out[6226] = x[282] & x[284];
    assign layer0_out[6227] = x[218] & ~x[207];
    assign layer0_out[6228] = x[78] ^ x[81];
    assign layer0_out[6229] = 1'b0;
    assign layer0_out[6230] = x[60] & x[76];
    assign layer0_out[6231] = x[276] | x[277];
    assign layer0_out[6232] = ~x[219];
    assign layer0_out[6233] = ~(x[109] ^ x[112]);
    assign layer0_out[6234] = x[185];
    assign layer0_out[6235] = x[339] ^ x[351];
    assign layer0_out[6236] = x[392] | x[397];
    assign layer0_out[6237] = ~x[131];
    assign layer0_out[6238] = x[208] | x[218];
    assign layer0_out[6239] = 1'b0;
    assign layer0_out[6240] = ~(x[150] & x[151]);
    assign layer0_out[6241] = x[297] & x[313];
    assign layer0_out[6242] = ~(x[332] & x[350]);
    assign layer0_out[6243] = x[204] | x[222];
    assign layer0_out[6244] = x[57] & ~x[41];
    assign layer0_out[6245] = x[73];
    assign layer0_out[6246] = ~x[74];
    assign layer0_out[6247] = ~(x[78] & x[80]);
    assign layer0_out[6248] = x[358];
    assign layer0_out[6249] = ~x[111];
    assign layer0_out[6250] = x[237];
    assign layer0_out[6251] = x[182] | x[184];
    assign layer0_out[6252] = ~(x[360] & x[364]);
    assign layer0_out[6253] = ~x[235];
    assign layer0_out[6254] = x[212] & x[215];
    assign layer0_out[6255] = x[262] & x[267];
    assign layer0_out[6256] = ~x[43];
    assign layer0_out[6257] = 1'b1;
    assign layer0_out[6258] = ~(x[116] | x[134]);
    assign layer0_out[6259] = ~x[282];
    assign layer0_out[6260] = 1'b0;
    assign layer0_out[6261] = ~x[235] | x[241];
    assign layer0_out[6262] = x[318] ^ x[326];
    assign layer0_out[6263] = ~(x[384] | x[398]);
    assign layer0_out[6264] = ~(x[280] | x[300]);
    assign layer0_out[6265] = ~(x[24] | x[44]);
    assign layer0_out[6266] = ~(x[155] ^ x[159]);
    assign layer0_out[6267] = ~x[350];
    assign layer0_out[6268] = ~x[253];
    assign layer0_out[6269] = x[282] | x[288];
    assign layer0_out[6270] = x[4];
    assign layer0_out[6271] = x[24];
    assign layer0_out[6272] = ~x[303] | x[285];
    assign layer0_out[6273] = x[299] & ~x[301];
    assign layer0_out[6274] = ~(x[252] & x[267]);
    assign layer0_out[6275] = x[217] | x[219];
    assign layer0_out[6276] = x[190] | x[211];
    assign layer0_out[6277] = x[294];
    assign layer0_out[6278] = ~(x[205] | x[217]);
    assign layer0_out[6279] = ~x[331];
    assign layer0_out[6280] = x[103] & x[119];
    assign layer0_out[6281] = ~(x[291] | x[296]);
    assign layer0_out[6282] = x[359] | x[378];
    assign layer0_out[6283] = ~x[129];
    assign layer0_out[6284] = ~x[311] | x[309];
    assign layer0_out[6285] = x[289] & ~x[285];
    assign layer0_out[6286] = ~(x[226] | x[246]);
    assign layer0_out[6287] = x[85] & x[95];
    assign layer0_out[6288] = ~(x[199] | x[219]);
    assign layer0_out[6289] = ~x[317];
    assign layer0_out[6290] = ~x[148];
    assign layer0_out[6291] = x[32] ^ x[43];
    assign layer0_out[6292] = ~(x[207] | x[220]);
    assign layer0_out[6293] = ~x[5] | x[10];
    assign layer0_out[6294] = x[167] ^ x[183];
    assign layer0_out[6295] = ~(x[26] | x[40]);
    assign layer0_out[6296] = x[318];
    assign layer0_out[6297] = x[75];
    assign layer0_out[6298] = ~(x[260] ^ x[262]);
    assign layer0_out[6299] = ~(x[99] | x[101]);
    assign layer0_out[6300] = x[16];
    assign layer0_out[6301] = ~x[313];
    assign layer0_out[6302] = ~x[215];
    assign layer0_out[6303] = x[208] ^ x[209];
    assign layer0_out[6304] = ~(x[241] & x[256]);
    assign layer0_out[6305] = x[106];
    assign layer0_out[6306] = ~(x[58] ^ x[60]);
    assign layer0_out[6307] = x[73] & ~x[80];
    assign layer0_out[6308] = x[361] | x[364];
    assign layer0_out[6309] = x[196] & ~x[211];
    assign layer0_out[6310] = x[69];
    assign layer0_out[6311] = ~x[193];
    assign layer0_out[6312] = x[136] & ~x[119];
    assign layer0_out[6313] = x[363] ^ x[366];
    assign layer0_out[6314] = x[292] ^ x[296];
    assign layer0_out[6315] = x[275] & x[289];
    assign layer0_out[6316] = x[266];
    assign layer0_out[6317] = x[142];
    assign layer0_out[6318] = ~x[374];
    assign layer0_out[6319] = ~(x[143] | x[148]);
    assign layer0_out[6320] = x[309];
    assign layer0_out[6321] = ~x[131];
    assign layer0_out[6322] = x[378] & x[386];
    assign layer0_out[6323] = x[146];
    assign layer0_out[6324] = x[63] & ~x[55];
    assign layer0_out[6325] = ~x[349];
    assign layer0_out[6326] = ~x[231] | x[234];
    assign layer0_out[6327] = x[39] & ~x[60];
    assign layer0_out[6328] = ~x[230] | x[220];
    assign layer0_out[6329] = ~x[319];
    assign layer0_out[6330] = ~(x[63] | x[83]);
    assign layer0_out[6331] = x[253] & x[273];
    assign layer0_out[6332] = x[191];
    assign layer0_out[6333] = ~x[102];
    assign layer0_out[6334] = ~(x[375] ^ x[386]);
    assign layer0_out[6335] = ~(x[54] ^ x[61]);
    assign layer0_out[6336] = x[116];
    assign layer0_out[6337] = ~x[149];
    assign layer0_out[6338] = ~(x[6] | x[7]);
    assign layer0_out[6339] = ~x[131] | x[121];
    assign layer0_out[6340] = ~(x[8] | x[23]);
    assign layer0_out[6341] = ~(x[108] | x[123]);
    assign layer0_out[6342] = x[198];
    assign layer0_out[6343] = x[58] & ~x[69];
    assign layer0_out[6344] = x[94] | x[103];
    assign layer0_out[6345] = x[304] | x[321];
    assign layer0_out[6346] = ~(x[29] | x[31]);
    assign layer0_out[6347] = 1'b0;
    assign layer0_out[6348] = x[342] & x[362];
    assign layer0_out[6349] = ~(x[110] | x[113]);
    assign layer0_out[6350] = ~x[255] | x[251];
    assign layer0_out[6351] = x[114] | x[120];
    assign layer0_out[6352] = ~x[222] | x[219];
    assign layer0_out[6353] = ~(x[352] | x[357]);
    assign layer0_out[6354] = ~x[77];
    assign layer0_out[6355] = ~(x[342] | x[361]);
    assign layer0_out[6356] = x[67] & ~x[70];
    assign layer0_out[6357] = x[299] ^ x[306];
    assign layer0_out[6358] = ~(x[253] ^ x[256]);
    assign layer0_out[6359] = ~(x[30] ^ x[45]);
    assign layer0_out[6360] = ~x[193];
    assign layer0_out[6361] = ~x[50];
    assign layer0_out[6362] = ~x[12] | x[5];
    assign layer0_out[6363] = x[198];
    assign layer0_out[6364] = x[276];
    assign layer0_out[6365] = ~(x[311] & x[322]);
    assign layer0_out[6366] = ~x[136] | x[132];
    assign layer0_out[6367] = x[380];
    assign layer0_out[6368] = 1'b1;
    assign layer0_out[6369] = x[2] | x[6];
    assign layer0_out[6370] = x[114] & x[127];
    assign layer0_out[6371] = x[199];
    assign layer0_out[6372] = ~x[214];
    assign layer0_out[6373] = ~(x[280] | x[295]);
    assign layer0_out[6374] = x[97] & ~x[95];
    assign layer0_out[6375] = x[342] | x[353];
    assign layer0_out[6376] = x[280];
    assign layer0_out[6377] = x[1] | x[17];
    assign layer0_out[6378] = ~x[119];
    assign layer0_out[6379] = ~(x[268] | x[270]);
    assign layer0_out[6380] = x[186] & ~x[197];
    assign layer0_out[6381] = ~x[192];
    assign layer0_out[6382] = ~(x[361] & x[371]);
    assign layer0_out[6383] = x[224] & x[244];
    assign layer0_out[6384] = x[210];
    assign layer0_out[6385] = 1'b0;
    assign layer0_out[6386] = x[167] | x[178];
    assign layer0_out[6387] = ~x[39] | x[41];
    assign layer0_out[6388] = ~(x[207] | x[222]);
    assign layer0_out[6389] = x[329] & x[335];
    assign layer0_out[6390] = ~(x[340] | x[348]);
    assign layer0_out[6391] = x[96] | x[117];
    assign layer0_out[6392] = x[210] & ~x[195];
    assign layer0_out[6393] = x[377] ^ x[394];
    assign layer0_out[6394] = 1'b1;
    assign layer0_out[6395] = x[382] | x[398];
    assign layer0_out[6396] = ~x[252] | x[243];
    assign layer0_out[6397] = ~x[209] | x[193];
    assign layer0_out[6398] = ~x[88];
    assign layer0_out[6399] = ~x[279] | x[284];
    assign layer0_out[6400] = ~x[370] | x[383];
    assign layer0_out[6401] = x[294] & ~x[302];
    assign layer0_out[6402] = x[71] | x[81];
    assign layer0_out[6403] = x[87];
    assign layer0_out[6404] = ~x[392] | x[379];
    assign layer0_out[6405] = x[34] | x[53];
    assign layer0_out[6406] = ~x[190];
    assign layer0_out[6407] = x[375] ^ x[385];
    assign layer0_out[6408] = x[351] & ~x[342];
    assign layer0_out[6409] = ~(x[347] & x[351]);
    assign layer0_out[6410] = x[133] | x[141];
    assign layer0_out[6411] = x[369] | x[373];
    assign layer0_out[6412] = ~x[159];
    assign layer0_out[6413] = ~x[46];
    assign layer0_out[6414] = x[115];
    assign layer0_out[6415] = x[125] & x[143];
    assign layer0_out[6416] = x[156] & ~x[173];
    assign layer0_out[6417] = x[40] & x[57];
    assign layer0_out[6418] = ~x[213];
    assign layer0_out[6419] = ~x[102];
    assign layer0_out[6420] = ~x[249];
    assign layer0_out[6421] = x[298] | x[304];
    assign layer0_out[6422] = x[159];
    assign layer0_out[6423] = ~x[133];
    assign layer0_out[6424] = ~(x[235] & x[254]);
    assign layer0_out[6425] = 1'b1;
    assign layer0_out[6426] = ~x[131] | x[135];
    assign layer0_out[6427] = ~(x[378] ^ x[380]);
    assign layer0_out[6428] = x[320];
    assign layer0_out[6429] = x[167] ^ x[176];
    assign layer0_out[6430] = ~(x[148] ^ x[153]);
    assign layer0_out[6431] = ~x[218] | x[228];
    assign layer0_out[6432] = ~(x[25] | x[43]);
    assign layer0_out[6433] = ~x[274] | x[273];
    assign layer0_out[6434] = x[136] & ~x[123];
    assign layer0_out[6435] = ~x[355];
    assign layer0_out[6436] = ~(x[213] & x[228]);
    assign layer0_out[6437] = ~x[364] | x[369];
    assign layer0_out[6438] = x[273];
    assign layer0_out[6439] = ~(x[98] | x[100]);
    assign layer0_out[6440] = ~(x[296] | x[316]);
    assign layer0_out[6441] = ~(x[299] | x[316]);
    assign layer0_out[6442] = x[373];
    assign layer0_out[6443] = x[243] | x[254];
    assign layer0_out[6444] = ~x[43];
    assign layer0_out[6445] = x[188] & ~x[193];
    assign layer0_out[6446] = x[239] & x[241];
    assign layer0_out[6447] = ~x[39];
    assign layer0_out[6448] = ~x[109];
    assign layer0_out[6449] = x[332];
    assign layer0_out[6450] = x[4] & ~x[22];
    assign layer0_out[6451] = ~(x[344] | x[359]);
    assign layer0_out[6452] = x[177] & ~x[185];
    assign layer0_out[6453] = x[129] | x[147];
    assign layer0_out[6454] = ~(x[261] ^ x[280]);
    assign layer0_out[6455] = x[283] ^ x[285];
    assign layer0_out[6456] = ~x[274] | x[262];
    assign layer0_out[6457] = ~(x[137] | x[155]);
    assign layer0_out[6458] = ~x[219];
    assign layer0_out[6459] = ~x[110];
    assign layer0_out[6460] = 1'b0;
    assign layer0_out[6461] = x[72];
    assign layer0_out[6462] = ~(x[19] | x[32]);
    assign layer0_out[6463] = ~(x[343] & x[347]);
    assign layer0_out[6464] = x[298];
    assign layer0_out[6465] = x[326] & x[330];
    assign layer0_out[6466] = x[5] ^ x[9];
    assign layer0_out[6467] = x[385] & ~x[397];
    assign layer0_out[6468] = x[382];
    assign layer0_out[6469] = ~x[173];
    assign layer0_out[6470] = ~(x[263] | x[275]);
    assign layer0_out[6471] = x[248] & ~x[231];
    assign layer0_out[6472] = ~(x[43] | x[59]);
    assign layer0_out[6473] = ~x[18];
    assign layer0_out[6474] = ~x[169];
    assign layer0_out[6475] = 1'b0;
    assign layer0_out[6476] = ~(x[162] | x[169]);
    assign layer0_out[6477] = 1'b1;
    assign layer0_out[6478] = x[70] & ~x[51];
    assign layer0_out[6479] = ~(x[215] | x[232]);
    assign layer0_out[6480] = ~(x[38] ^ x[44]);
    assign layer0_out[6481] = x[317] | x[318];
    assign layer0_out[6482] = x[59];
    assign layer0_out[6483] = ~x[170] | x[154];
    assign layer0_out[6484] = ~x[3] | x[16];
    assign layer0_out[6485] = x[265];
    assign layer0_out[6486] = x[304];
    assign layer0_out[6487] = x[197];
    assign layer0_out[6488] = ~(x[347] ^ x[366]);
    assign layer0_out[6489] = x[108];
    assign layer0_out[6490] = x[287] & x[296];
    assign layer0_out[6491] = x[246];
    assign layer0_out[6492] = x[214] | x[229];
    assign layer0_out[6493] = ~(x[40] & x[55]);
    assign layer0_out[6494] = ~(x[217] | x[228]);
    assign layer0_out[6495] = x[314] | x[330];
    assign layer0_out[6496] = x[171];
    assign layer0_out[6497] = ~(x[211] & x[217]);
    assign layer0_out[6498] = ~(x[56] | x[57]);
    assign layer0_out[6499] = ~(x[170] | x[182]);
    assign layer0_out[6500] = x[363] | x[373];
    assign layer0_out[6501] = x[391];
    assign layer0_out[6502] = x[106];
    assign layer0_out[6503] = ~x[122] | x[111];
    assign layer0_out[6504] = ~(x[332] | x[338]);
    assign layer0_out[6505] = ~x[91];
    assign layer0_out[6506] = x[178] ^ x[185];
    assign layer0_out[6507] = x[346];
    assign layer0_out[6508] = x[14] ^ x[34];
    assign layer0_out[6509] = ~x[107] | x[112];
    assign layer0_out[6510] = ~x[159];
    assign layer0_out[6511] = x[140] & ~x[127];
    assign layer0_out[6512] = x[295] & x[311];
    assign layer0_out[6513] = ~x[289];
    assign layer0_out[6514] = x[384] & ~x[374];
    assign layer0_out[6515] = x[308] & ~x[305];
    assign layer0_out[6516] = x[128] | x[144];
    assign layer0_out[6517] = ~(x[27] | x[28]);
    assign layer0_out[6518] = x[30];
    assign layer0_out[6519] = ~x[338];
    assign layer0_out[6520] = ~x[149];
    assign layer0_out[6521] = ~x[259] | x[254];
    assign layer0_out[6522] = 1'b0;
    assign layer0_out[6523] = x[133];
    assign layer0_out[6524] = x[162] & x[178];
    assign layer0_out[6525] = ~(x[30] | x[42]);
    assign layer0_out[6526] = x[377] & x[392];
    assign layer0_out[6527] = ~(x[10] & x[11]);
    assign layer0_out[6528] = 1'b1;
    assign layer0_out[6529] = x[241] | x[244];
    assign layer0_out[6530] = ~(x[177] | x[180]);
    assign layer0_out[6531] = ~x[13] | x[26];
    assign layer0_out[6532] = 1'b1;
    assign layer0_out[6533] = ~(x[75] & x[92]);
    assign layer0_out[6534] = ~(x[203] ^ x[210]);
    assign layer0_out[6535] = ~(x[70] & x[84]);
    assign layer0_out[6536] = x[227];
    assign layer0_out[6537] = 1'b1;
    assign layer0_out[6538] = ~(x[264] | x[277]);
    assign layer0_out[6539] = x[179] & ~x[163];
    assign layer0_out[6540] = x[265] & ~x[254];
    assign layer0_out[6541] = ~(x[45] | x[58]);
    assign layer0_out[6542] = ~x[248];
    assign layer0_out[6543] = ~x[208];
    assign layer0_out[6544] = x[204] ^ x[220];
    assign layer0_out[6545] = ~(x[185] ^ x[190]);
    assign layer0_out[6546] = x[380];
    assign layer0_out[6547] = x[61] | x[75];
    assign layer0_out[6548] = ~(x[28] | x[40]);
    assign layer0_out[6549] = ~x[247];
    assign layer0_out[6550] = 1'b0;
    assign layer0_out[6551] = x[258] ^ x[274];
    assign layer0_out[6552] = ~x[236] | x[226];
    assign layer0_out[6553] = 1'b0;
    assign layer0_out[6554] = ~(x[331] | x[339]);
    assign layer0_out[6555] = 1'b1;
    assign layer0_out[6556] = x[135] ^ x[137];
    assign layer0_out[6557] = 1'b1;
    assign layer0_out[6558] = 1'b0;
    assign layer0_out[6559] = ~(x[173] | x[190]);
    assign layer0_out[6560] = ~x[244];
    assign layer0_out[6561] = x[92] & ~x[71];
    assign layer0_out[6562] = ~x[188];
    assign layer0_out[6563] = ~(x[44] | x[46]);
    assign layer0_out[6564] = x[382] | x[395];
    assign layer0_out[6565] = x[226];
    assign layer0_out[6566] = ~x[149];
    assign layer0_out[6567] = ~x[210] | x[221];
    assign layer0_out[6568] = x[66] & ~x[57];
    assign layer0_out[6569] = ~(x[127] ^ x[138]);
    assign layer0_out[6570] = ~(x[318] | x[325]);
    assign layer0_out[6571] = ~(x[339] ^ x[344]);
    assign layer0_out[6572] = ~(x[142] | x[145]);
    assign layer0_out[6573] = ~x[19] | x[34];
    assign layer0_out[6574] = ~(x[187] ^ x[205]);
    assign layer0_out[6575] = x[101];
    assign layer0_out[6576] = ~x[264];
    assign layer0_out[6577] = x[4];
    assign layer0_out[6578] = x[362];
    assign layer0_out[6579] = x[162] & ~x[148];
    assign layer0_out[6580] = x[78] & ~x[89];
    assign layer0_out[6581] = ~(x[63] ^ x[81]);
    assign layer0_out[6582] = ~x[14];
    assign layer0_out[6583] = ~(x[182] | x[199]);
    assign layer0_out[6584] = ~(x[308] | x[318]);
    assign layer0_out[6585] = x[130];
    assign layer0_out[6586] = ~(x[242] | x[245]);
    assign layer0_out[6587] = ~x[246];
    assign layer0_out[6588] = ~(x[88] ^ x[107]);
    assign layer0_out[6589] = x[103] & ~x[104];
    assign layer0_out[6590] = ~(x[371] | x[391]);
    assign layer0_out[6591] = ~(x[385] | x[386]);
    assign layer0_out[6592] = ~x[261];
    assign layer0_out[6593] = 1'b0;
    assign layer0_out[6594] = x[342] | x[344];
    assign layer0_out[6595] = x[224] & ~x[217];
    assign layer0_out[6596] = ~x[24];
    assign layer0_out[6597] = x[287] ^ x[289];
    assign layer0_out[6598] = x[181] & x[189];
    assign layer0_out[6599] = ~x[125];
    assign layer0_out[6600] = ~x[205] | x[199];
    assign layer0_out[6601] = ~x[107] | x[91];
    assign layer0_out[6602] = x[130] | x[136];
    assign layer0_out[6603] = 1'b0;
    assign layer0_out[6604] = x[125] | x[144];
    assign layer0_out[6605] = x[219];
    assign layer0_out[6606] = ~x[355];
    assign layer0_out[6607] = ~(x[242] | x[244]);
    assign layer0_out[6608] = ~(x[78] & x[82]);
    assign layer0_out[6609] = ~x[258];
    assign layer0_out[6610] = 1'b0;
    assign layer0_out[6611] = x[379] | x[383];
    assign layer0_out[6612] = x[103] ^ x[118];
    assign layer0_out[6613] = ~x[225];
    assign layer0_out[6614] = x[121] | x[127];
    assign layer0_out[6615] = ~(x[155] | x[162]);
    assign layer0_out[6616] = x[371] & ~x[378];
    assign layer0_out[6617] = ~x[290] | x[307];
    assign layer0_out[6618] = x[86];
    assign layer0_out[6619] = x[382] & ~x[385];
    assign layer0_out[6620] = ~(x[351] | x[363]);
    assign layer0_out[6621] = ~x[307];
    assign layer0_out[6622] = ~x[342] | x[331];
    assign layer0_out[6623] = ~(x[259] ^ x[272]);
    assign layer0_out[6624] = ~(x[16] | x[34]);
    assign layer0_out[6625] = ~(x[95] | x[115]);
    assign layer0_out[6626] = x[45];
    assign layer0_out[6627] = ~(x[251] | x[259]);
    assign layer0_out[6628] = x[370];
    assign layer0_out[6629] = x[242] & x[255];
    assign layer0_out[6630] = ~x[77];
    assign layer0_out[6631] = ~(x[228] | x[235]);
    assign layer0_out[6632] = ~x[313];
    assign layer0_out[6633] = x[356] | x[369];
    assign layer0_out[6634] = x[46] | x[53];
    assign layer0_out[6635] = x[114] & ~x[110];
    assign layer0_out[6636] = 1'b1;
    assign layer0_out[6637] = ~(x[303] ^ x[320]);
    assign layer0_out[6638] = ~(x[125] ^ x[127]);
    assign layer0_out[6639] = ~(x[373] ^ x[392]);
    assign layer0_out[6640] = ~x[318];
    assign layer0_out[6641] = x[319];
    assign layer0_out[6642] = x[356];
    assign layer0_out[6643] = ~(x[355] | x[363]);
    assign layer0_out[6644] = x[83] & x[92];
    assign layer0_out[6645] = x[86] ^ x[104];
    assign layer0_out[6646] = ~(x[338] | x[357]);
    assign layer0_out[6647] = ~x[0] | x[15];
    assign layer0_out[6648] = ~(x[260] | x[276]);
    assign layer0_out[6649] = ~(x[195] ^ x[198]);
    assign layer0_out[6650] = ~x[9];
    assign layer0_out[6651] = ~(x[267] ^ x[284]);
    assign layer0_out[6652] = x[242] & ~x[231];
    assign layer0_out[6653] = ~(x[107] | x[118]);
    assign layer0_out[6654] = ~(x[90] ^ x[97]);
    assign layer0_out[6655] = ~(x[238] & x[252]);
    assign layer0_out[6656] = x[125] & x[145];
    assign layer0_out[6657] = ~x[316] | x[306];
    assign layer0_out[6658] = ~x[141];
    assign layer0_out[6659] = x[264] & ~x[263];
    assign layer0_out[6660] = ~(x[318] ^ x[333]);
    assign layer0_out[6661] = ~(x[346] | x[360]);
    assign layer0_out[6662] = x[203] & ~x[186];
    assign layer0_out[6663] = ~(x[83] | x[98]);
    assign layer0_out[6664] = ~(x[117] ^ x[132]);
    assign layer0_out[6665] = ~(x[293] | x[304]);
    assign layer0_out[6666] = ~(x[365] | x[380]);
    assign layer0_out[6667] = x[37];
    assign layer0_out[6668] = x[304] | x[316];
    assign layer0_out[6669] = ~(x[106] | x[117]);
    assign layer0_out[6670] = x[25];
    assign layer0_out[6671] = x[48] ^ x[52];
    assign layer0_out[6672] = ~(x[152] | x[157]);
    assign layer0_out[6673] = x[190] & x[197];
    assign layer0_out[6674] = x[30] & ~x[20];
    assign layer0_out[6675] = ~x[39] | x[23];
    assign layer0_out[6676] = ~(x[264] | x[268]);
    assign layer0_out[6677] = x[24] ^ x[42];
    assign layer0_out[6678] = x[281];
    assign layer0_out[6679] = ~x[88] | x[86];
    assign layer0_out[6680] = ~(x[190] | x[210]);
    assign layer0_out[6681] = ~x[288];
    assign layer0_out[6682] = x[276];
    assign layer0_out[6683] = x[348];
    assign layer0_out[6684] = x[24] & ~x[38];
    assign layer0_out[6685] = ~(x[9] | x[25]);
    assign layer0_out[6686] = ~x[142];
    assign layer0_out[6687] = ~x[188] | x[200];
    assign layer0_out[6688] = ~(x[247] | x[267]);
    assign layer0_out[6689] = ~(x[333] & x[347]);
    assign layer0_out[6690] = x[323];
    assign layer0_out[6691] = ~(x[331] | x[334]);
    assign layer0_out[6692] = x[128] & ~x[146];
    assign layer0_out[6693] = ~x[347];
    assign layer0_out[6694] = ~x[298];
    assign layer0_out[6695] = x[94] | x[108];
    assign layer0_out[6696] = ~(x[157] | x[176]);
    assign layer0_out[6697] = x[250] & ~x[242];
    assign layer0_out[6698] = ~(x[18] ^ x[39]);
    assign layer0_out[6699] = ~x[309] | x[300];
    assign layer0_out[6700] = ~x[203];
    assign layer0_out[6701] = x[105] | x[118];
    assign layer0_out[6702] = x[133];
    assign layer0_out[6703] = ~(x[52] | x[59]);
    assign layer0_out[6704] = x[246] & x[265];
    assign layer0_out[6705] = ~x[308];
    assign layer0_out[6706] = ~(x[50] | x[51]);
    assign layer0_out[6707] = x[202] & ~x[219];
    assign layer0_out[6708] = x[219] | x[224];
    assign layer0_out[6709] = ~x[263];
    assign layer0_out[6710] = x[157];
    assign layer0_out[6711] = x[374];
    assign layer0_out[6712] = x[200] | x[212];
    assign layer0_out[6713] = ~(x[244] & x[251]);
    assign layer0_out[6714] = x[29] & ~x[37];
    assign layer0_out[6715] = ~x[102] | x[91];
    assign layer0_out[6716] = 1'b0;
    assign layer0_out[6717] = x[81] & ~x[85];
    assign layer0_out[6718] = ~(x[45] | x[60]);
    assign layer0_out[6719] = x[384] | x[393];
    assign layer0_out[6720] = x[352];
    assign layer0_out[6721] = ~x[332];
    assign layer0_out[6722] = ~x[394];
    assign layer0_out[6723] = ~x[333];
    assign layer0_out[6724] = x[103];
    assign layer0_out[6725] = x[362] | x[374];
    assign layer0_out[6726] = ~x[81];
    assign layer0_out[6727] = x[61];
    assign layer0_out[6728] = ~(x[313] & x[314]);
    assign layer0_out[6729] = ~x[378];
    assign layer0_out[6730] = x[194] | x[201];
    assign layer0_out[6731] = 1'b0;
    assign layer0_out[6732] = x[309] & ~x[313];
    assign layer0_out[6733] = ~x[211];
    assign layer0_out[6734] = ~x[152] | x[160];
    assign layer0_out[6735] = x[348] & x[350];
    assign layer0_out[6736] = x[353] & x[362];
    assign layer0_out[6737] = ~x[209];
    assign layer0_out[6738] = x[365] ^ x[372];
    assign layer0_out[6739] = ~x[172] | x[161];
    assign layer0_out[6740] = x[203];
    assign layer0_out[6741] = ~x[122];
    assign layer0_out[6742] = x[202] | x[204];
    assign layer0_out[6743] = ~x[31];
    assign layer0_out[6744] = ~x[251];
    assign layer0_out[6745] = ~x[226] | x[233];
    assign layer0_out[6746] = ~(x[46] & x[51]);
    assign layer0_out[6747] = x[246] & ~x[238];
    assign layer0_out[6748] = x[145];
    assign layer0_out[6749] = x[77] | x[93];
    assign layer0_out[6750] = x[198];
    assign layer0_out[6751] = ~x[290];
    assign layer0_out[6752] = x[302];
    assign layer0_out[6753] = x[108];
    assign layer0_out[6754] = ~x[299] | x[302];
    assign layer0_out[6755] = x[118] | x[120];
    assign layer0_out[6756] = ~(x[47] | x[65]);
    assign layer0_out[6757] = x[123] & ~x[112];
    assign layer0_out[6758] = 1'b1;
    assign layer0_out[6759] = ~x[155] | x[168];
    assign layer0_out[6760] = x[326] ^ x[329];
    assign layer0_out[6761] = ~x[10] | x[14];
    assign layer0_out[6762] = ~(x[1] & x[7]);
    assign layer0_out[6763] = ~x[31];
    assign layer0_out[6764] = ~x[26];
    assign layer0_out[6765] = ~x[269];
    assign layer0_out[6766] = x[10] ^ x[16];
    assign layer0_out[6767] = ~x[392];
    assign layer0_out[6768] = x[103] | x[115];
    assign layer0_out[6769] = x[52] & x[68];
    assign layer0_out[6770] = ~(x[341] | x[361]);
    assign layer0_out[6771] = x[309] | x[325];
    assign layer0_out[6772] = x[207] ^ x[213];
    assign layer0_out[6773] = ~x[118];
    assign layer0_out[6774] = ~x[308] | x[288];
    assign layer0_out[6775] = x[164] | x[167];
    assign layer0_out[6776] = x[277] & ~x[262];
    assign layer0_out[6777] = ~x[130];
    assign layer0_out[6778] = ~x[90];
    assign layer0_out[6779] = ~(x[8] ^ x[14]);
    assign layer0_out[6780] = x[348] & x[363];
    assign layer0_out[6781] = ~x[11];
    assign layer0_out[6782] = x[44] & x[59];
    assign layer0_out[6783] = x[257] | x[267];
    assign layer0_out[6784] = x[244] & x[249];
    assign layer0_out[6785] = ~(x[59] ^ x[78]);
    assign layer0_out[6786] = ~(x[47] | x[49]);
    assign layer0_out[6787] = ~(x[303] | x[317]);
    assign layer0_out[6788] = ~x[340];
    assign layer0_out[6789] = 1'b1;
    assign layer0_out[6790] = ~x[342];
    assign layer0_out[6791] = x[167];
    assign layer0_out[6792] = ~x[373];
    assign layer0_out[6793] = ~x[335];
    assign layer0_out[6794] = ~x[269] | x[280];
    assign layer0_out[6795] = ~(x[336] | x[355]);
    assign layer0_out[6796] = x[349] | x[367];
    assign layer0_out[6797] = ~(x[37] | x[56]);
    assign layer0_out[6798] = ~(x[94] | x[99]);
    assign layer0_out[6799] = x[356];
    assign layer0_out[6800] = x[333] | x[341];
    assign layer0_out[6801] = x[302];
    assign layer0_out[6802] = ~(x[319] & x[330]);
    assign layer0_out[6803] = ~(x[244] | x[245]);
    assign layer0_out[6804] = x[347] & ~x[356];
    assign layer0_out[6805] = x[302];
    assign layer0_out[6806] = ~x[67];
    assign layer0_out[6807] = ~x[86];
    assign layer0_out[6808] = ~x[131] | x[145];
    assign layer0_out[6809] = x[53] & x[58];
    assign layer0_out[6810] = ~x[169] | x[149];
    assign layer0_out[6811] = ~(x[223] ^ x[225]);
    assign layer0_out[6812] = ~(x[121] | x[138]);
    assign layer0_out[6813] = x[198] ^ x[206];
    assign layer0_out[6814] = 1'b0;
    assign layer0_out[6815] = ~(x[125] | x[141]);
    assign layer0_out[6816] = x[324] | x[329];
    assign layer0_out[6817] = ~(x[355] & x[365]);
    assign layer0_out[6818] = x[368] & ~x[377];
    assign layer0_out[6819] = x[163] & ~x[155];
    assign layer0_out[6820] = 1'b1;
    assign layer0_out[6821] = ~(x[128] ^ x[141]);
    assign layer0_out[6822] = x[61];
    assign layer0_out[6823] = ~(x[79] | x[92]);
    assign layer0_out[6824] = 1'b0;
    assign layer0_out[6825] = x[78] ^ x[95];
    assign layer0_out[6826] = x[118] | x[121];
    assign layer0_out[6827] = x[151] & ~x[139];
    assign layer0_out[6828] = ~x[129];
    assign layer0_out[6829] = x[376] & ~x[369];
    assign layer0_out[6830] = x[190] | x[200];
    assign layer0_out[6831] = x[384] | x[399];
    assign layer0_out[6832] = x[270];
    assign layer0_out[6833] = ~(x[184] | x[195]);
    assign layer0_out[6834] = x[384] & x[388];
    assign layer0_out[6835] = ~x[263] | x[278];
    assign layer0_out[6836] = ~(x[87] & x[103]);
    assign layer0_out[6837] = ~x[184];
    assign layer0_out[6838] = ~x[169];
    assign layer0_out[6839] = x[28] & x[30];
    assign layer0_out[6840] = ~(x[332] & x[343]);
    assign layer0_out[6841] = ~(x[183] | x[185]);
    assign layer0_out[6842] = x[285] | x[304];
    assign layer0_out[6843] = x[332] ^ x[349];
    assign layer0_out[6844] = ~x[355];
    assign layer0_out[6845] = x[39] & ~x[29];
    assign layer0_out[6846] = x[355] | x[375];
    assign layer0_out[6847] = x[362] & x[372];
    assign layer0_out[6848] = x[206];
    assign layer0_out[6849] = x[56] | x[76];
    assign layer0_out[6850] = ~x[325];
    assign layer0_out[6851] = ~(x[110] & x[121]);
    assign layer0_out[6852] = x[260] & ~x[259];
    assign layer0_out[6853] = ~(x[374] | x[388]);
    assign layer0_out[6854] = ~x[229];
    assign layer0_out[6855] = x[69] | x[78];
    assign layer0_out[6856] = x[387] & ~x[374];
    assign layer0_out[6857] = x[228];
    assign layer0_out[6858] = ~x[322];
    assign layer0_out[6859] = x[328] & x[347];
    assign layer0_out[6860] = 1'b0;
    assign layer0_out[6861] = x[27] & x[45];
    assign layer0_out[6862] = x[148] & ~x[149];
    assign layer0_out[6863] = x[107] | x[119];
    assign layer0_out[6864] = ~x[28];
    assign layer0_out[6865] = x[291] | x[301];
    assign layer0_out[6866] = ~(x[153] | x[157]);
    assign layer0_out[6867] = x[233] & ~x[214];
    assign layer0_out[6868] = ~(x[332] | x[334]);
    assign layer0_out[6869] = x[210] | x[229];
    assign layer0_out[6870] = 1'b0;
    assign layer0_out[6871] = x[379] | x[398];
    assign layer0_out[6872] = x[120] | x[125];
    assign layer0_out[6873] = ~(x[8] | x[26]);
    assign layer0_out[6874] = x[332] & x[335];
    assign layer0_out[6875] = x[190] & ~x[201];
    assign layer0_out[6876] = 1'b1;
    assign layer0_out[6877] = ~(x[266] | x[283]);
    assign layer0_out[6878] = ~x[109] | x[126];
    assign layer0_out[6879] = ~(x[30] | x[37]);
    assign layer0_out[6880] = x[245] & x[254];
    assign layer0_out[6881] = ~(x[236] | x[237]);
    assign layer0_out[6882] = ~x[2] | x[20];
    assign layer0_out[6883] = x[134] | x[135];
    assign layer0_out[6884] = x[224] & ~x[203];
    assign layer0_out[6885] = ~(x[348] & x[352]);
    assign layer0_out[6886] = x[349] & x[366];
    assign layer0_out[6887] = ~x[282];
    assign layer0_out[6888] = ~x[154];
    assign layer0_out[6889] = x[181] & ~x[182];
    assign layer0_out[6890] = x[79] | x[99];
    assign layer0_out[6891] = ~x[283] | x[298];
    assign layer0_out[6892] = ~(x[30] ^ x[39]);
    assign layer0_out[6893] = ~x[278];
    assign layer0_out[6894] = ~x[194];
    assign layer0_out[6895] = ~(x[253] ^ x[259]);
    assign layer0_out[6896] = x[357] | x[363];
    assign layer0_out[6897] = ~(x[317] & x[335]);
    assign layer0_out[6898] = ~x[181];
    assign layer0_out[6899] = ~(x[56] | x[59]);
    assign layer0_out[6900] = x[243];
    assign layer0_out[6901] = x[198] | x[200];
    assign layer0_out[6902] = x[385] & x[389];
    assign layer0_out[6903] = x[144];
    assign layer0_out[6904] = ~x[190] | x[177];
    assign layer0_out[6905] = ~x[168];
    assign layer0_out[6906] = x[114] | x[130];
    assign layer0_out[6907] = x[265] | x[271];
    assign layer0_out[6908] = ~(x[370] & x[373]);
    assign layer0_out[6909] = x[0] & x[21];
    assign layer0_out[6910] = ~(x[257] ^ x[269]);
    assign layer0_out[6911] = x[73] & ~x[60];
    assign layer0_out[6912] = ~x[46] | x[38];
    assign layer0_out[6913] = x[159] ^ x[165];
    assign layer0_out[6914] = ~x[383];
    assign layer0_out[6915] = x[23];
    assign layer0_out[6916] = x[174];
    assign layer0_out[6917] = ~x[39];
    assign layer0_out[6918] = x[36];
    assign layer0_out[6919] = ~x[170];
    assign layer0_out[6920] = 1'b1;
    assign layer0_out[6921] = x[158] & ~x[173];
    assign layer0_out[6922] = ~x[201];
    assign layer0_out[6923] = ~x[386];
    assign layer0_out[6924] = x[154] & ~x[139];
    assign layer0_out[6925] = ~x[293] | x[313];
    assign layer0_out[6926] = x[333] & ~x[342];
    assign layer0_out[6927] = ~(x[174] | x[194]);
    assign layer0_out[6928] = x[303] ^ x[315];
    assign layer0_out[6929] = x[190];
    assign layer0_out[6930] = ~(x[170] | x[171]);
    assign layer0_out[6931] = x[24] & ~x[12];
    assign layer0_out[6932] = ~x[387];
    assign layer0_out[6933] = x[201] & ~x[211];
    assign layer0_out[6934] = ~(x[240] | x[252]);
    assign layer0_out[6935] = ~(x[314] | x[326]);
    assign layer0_out[6936] = x[205] & ~x[193];
    assign layer0_out[6937] = ~(x[172] | x[181]);
    assign layer0_out[6938] = ~(x[116] | x[132]);
    assign layer0_out[6939] = ~(x[280] & x[289]);
    assign layer0_out[6940] = ~x[249];
    assign layer0_out[6941] = x[173];
    assign layer0_out[6942] = x[43];
    assign layer0_out[6943] = ~x[183];
    assign layer0_out[6944] = x[249] | x[259];
    assign layer0_out[6945] = x[311] ^ x[329];
    assign layer0_out[6946] = x[159] | x[160];
    assign layer0_out[6947] = x[300];
    assign layer0_out[6948] = ~(x[105] ^ x[107]);
    assign layer0_out[6949] = ~x[388];
    assign layer0_out[6950] = ~x[201];
    assign layer0_out[6951] = ~(x[246] | x[264]);
    assign layer0_out[6952] = ~(x[303] | x[321]);
    assign layer0_out[6953] = ~x[3] | x[7];
    assign layer0_out[6954] = ~x[268] | x[278];
    assign layer0_out[6955] = x[320] & ~x[329];
    assign layer0_out[6956] = x[372] ^ x[391];
    assign layer0_out[6957] = x[316];
    assign layer0_out[6958] = x[308] ^ x[312];
    assign layer0_out[6959] = x[110] & x[130];
    assign layer0_out[6960] = ~x[123];
    assign layer0_out[6961] = x[28];
    assign layer0_out[6962] = 1'b0;
    assign layer0_out[6963] = x[225] | x[243];
    assign layer0_out[6964] = ~x[306] | x[291];
    assign layer0_out[6965] = ~(x[182] | x[203]);
    assign layer0_out[6966] = ~(x[375] | x[382]);
    assign layer0_out[6967] = ~(x[289] ^ x[290]);
    assign layer0_out[6968] = ~(x[322] | x[332]);
    assign layer0_out[6969] = ~(x[128] & x[142]);
    assign layer0_out[6970] = x[214] | x[234];
    assign layer0_out[6971] = ~(x[342] ^ x[356]);
    assign layer0_out[6972] = ~x[284];
    assign layer0_out[6973] = x[312];
    assign layer0_out[6974] = x[351] | x[370];
    assign layer0_out[6975] = x[303];
    assign layer0_out[6976] = ~x[348];
    assign layer0_out[6977] = x[39];
    assign layer0_out[6978] = ~x[229];
    assign layer0_out[6979] = x[165] ^ x[182];
    assign layer0_out[6980] = x[289];
    assign layer0_out[6981] = x[393] | x[394];
    assign layer0_out[6982] = x[181] & x[196];
    assign layer0_out[6983] = x[370] | x[371];
    assign layer0_out[6984] = ~x[378];
    assign layer0_out[6985] = x[62];
    assign layer0_out[6986] = x[124] ^ x[126];
    assign layer0_out[6987] = ~(x[82] | x[88]);
    assign layer0_out[6988] = ~x[279];
    assign layer0_out[6989] = ~(x[218] | x[224]);
    assign layer0_out[6990] = x[174] | x[180];
    assign layer0_out[6991] = 1'b0;
    assign layer0_out[6992] = ~(x[251] ^ x[257]);
    assign layer0_out[6993] = ~(x[237] ^ x[253]);
    assign layer0_out[6994] = 1'b1;
    assign layer0_out[6995] = x[28];
    assign layer0_out[6996] = ~x[325] | x[340];
    assign layer0_out[6997] = ~(x[349] | x[353]);
    assign layer0_out[6998] = ~x[275];
    assign layer0_out[6999] = ~x[92] | x[73];
    assign layer0_out[7000] = ~x[325];
    assign layer0_out[7001] = ~(x[200] | x[204]);
    assign layer0_out[7002] = ~(x[245] & x[251]);
    assign layer0_out[7003] = ~(x[102] ^ x[105]);
    assign layer0_out[7004] = ~x[347] | x[338];
    assign layer0_out[7005] = x[157] & ~x[163];
    assign layer0_out[7006] = x[352] & x[353];
    assign layer0_out[7007] = ~(x[269] & x[273]);
    assign layer0_out[7008] = ~x[298];
    assign layer0_out[7009] = x[247] & x[252];
    assign layer0_out[7010] = ~x[102] | x[95];
    assign layer0_out[7011] = ~x[122] | x[131];
    assign layer0_out[7012] = ~(x[79] | x[89]);
    assign layer0_out[7013] = ~x[263] | x[279];
    assign layer0_out[7014] = ~x[57];
    assign layer0_out[7015] = x[179] | x[196];
    assign layer0_out[7016] = ~x[86] | x[76];
    assign layer0_out[7017] = ~x[186];
    assign layer0_out[7018] = ~x[117] | x[98];
    assign layer0_out[7019] = x[63] | x[67];
    assign layer0_out[7020] = x[235] | x[252];
    assign layer0_out[7021] = x[344] ^ x[357];
    assign layer0_out[7022] = 1'b0;
    assign layer0_out[7023] = ~(x[229] & x[238]);
    assign layer0_out[7024] = ~x[50] | x[47];
    assign layer0_out[7025] = x[204];
    assign layer0_out[7026] = ~x[324];
    assign layer0_out[7027] = x[60];
    assign layer0_out[7028] = ~(x[215] | x[220]);
    assign layer0_out[7029] = x[297] | x[298];
    assign layer0_out[7030] = x[315];
    assign layer0_out[7031] = ~(x[199] ^ x[206]);
    assign layer0_out[7032] = 1'b1;
    assign layer0_out[7033] = x[265];
    assign layer0_out[7034] = ~(x[253] | x[262]);
    assign layer0_out[7035] = x[390];
    assign layer0_out[7036] = x[200] ^ x[214];
    assign layer0_out[7037] = x[342] | x[343];
    assign layer0_out[7038] = ~x[382];
    assign layer0_out[7039] = x[369] ^ x[378];
    assign layer0_out[7040] = ~x[165];
    assign layer0_out[7041] = x[229] | x[248];
    assign layer0_out[7042] = ~x[57];
    assign layer0_out[7043] = ~x[133];
    assign layer0_out[7044] = x[74] & ~x[57];
    assign layer0_out[7045] = x[36] ^ x[44];
    assign layer0_out[7046] = ~x[75];
    assign layer0_out[7047] = ~(x[120] ^ x[133]);
    assign layer0_out[7048] = ~(x[357] | x[368]);
    assign layer0_out[7049] = 1'b0;
    assign layer0_out[7050] = ~x[187];
    assign layer0_out[7051] = x[243] | x[253];
    assign layer0_out[7052] = ~(x[305] ^ x[307]);
    assign layer0_out[7053] = ~x[319] | x[332];
    assign layer0_out[7054] = ~x[31];
    assign layer0_out[7055] = ~x[221];
    assign layer0_out[7056] = x[58] & x[68];
    assign layer0_out[7057] = x[139] & x[158];
    assign layer0_out[7058] = ~x[322];
    assign layer0_out[7059] = 1'b1;
    assign layer0_out[7060] = x[305] ^ x[318];
    assign layer0_out[7061] = ~x[364] | x[351];
    assign layer0_out[7062] = x[251] & ~x[233];
    assign layer0_out[7063] = ~x[324] | x[318];
    assign layer0_out[7064] = ~x[376];
    assign layer0_out[7065] = x[307];
    assign layer0_out[7066] = ~(x[248] | x[266]);
    assign layer0_out[7067] = ~(x[277] | x[297]);
    assign layer0_out[7068] = ~x[52];
    assign layer0_out[7069] = x[44] ^ x[50];
    assign layer0_out[7070] = x[252] & ~x[248];
    assign layer0_out[7071] = ~x[253];
    assign layer0_out[7072] = ~(x[216] | x[235]);
    assign layer0_out[7073] = ~x[77] | x[71];
    assign layer0_out[7074] = x[195] & ~x[188];
    assign layer0_out[7075] = x[296] & ~x[276];
    assign layer0_out[7076] = 1'b1;
    assign layer0_out[7077] = ~x[172];
    assign layer0_out[7078] = 1'b0;
    assign layer0_out[7079] = ~(x[292] | x[308]);
    assign layer0_out[7080] = x[225] | x[234];
    assign layer0_out[7081] = x[372] ^ x[381];
    assign layer0_out[7082] = ~x[297];
    assign layer0_out[7083] = ~(x[136] | x[151]);
    assign layer0_out[7084] = ~(x[181] | x[198]);
    assign layer0_out[7085] = x[124];
    assign layer0_out[7086] = x[360];
    assign layer0_out[7087] = ~x[288];
    assign layer0_out[7088] = x[355];
    assign layer0_out[7089] = ~(x[127] ^ x[148]);
    assign layer0_out[7090] = ~x[298] | x[291];
    assign layer0_out[7091] = x[32] & ~x[20];
    assign layer0_out[7092] = x[281];
    assign layer0_out[7093] = x[165] | x[183];
    assign layer0_out[7094] = ~(x[42] ^ x[63]);
    assign layer0_out[7095] = ~(x[297] | x[301]);
    assign layer0_out[7096] = ~x[94] | x[88];
    assign layer0_out[7097] = ~(x[323] | x[343]);
    assign layer0_out[7098] = ~(x[305] | x[324]);
    assign layer0_out[7099] = x[89] | x[98];
    assign layer0_out[7100] = x[350] | x[351];
    assign layer0_out[7101] = ~x[152];
    assign layer0_out[7102] = x[34] & ~x[41];
    assign layer0_out[7103] = ~x[167];
    assign layer0_out[7104] = ~x[99];
    assign layer0_out[7105] = x[302] ^ x[317];
    assign layer0_out[7106] = x[331] & x[344];
    assign layer0_out[7107] = ~x[88] | x[91];
    assign layer0_out[7108] = x[324] | x[333];
    assign layer0_out[7109] = x[368];
    assign layer0_out[7110] = ~(x[162] | x[183]);
    assign layer0_out[7111] = ~(x[16] ^ x[28]);
    assign layer0_out[7112] = ~(x[12] | x[32]);
    assign layer0_out[7113] = x[335] | x[336];
    assign layer0_out[7114] = x[263];
    assign layer0_out[7115] = x[279] & ~x[291];
    assign layer0_out[7116] = x[60];
    assign layer0_out[7117] = ~x[47];
    assign layer0_out[7118] = x[114];
    assign layer0_out[7119] = ~x[362];
    assign layer0_out[7120] = x[324];
    assign layer0_out[7121] = ~(x[304] ^ x[307]);
    assign layer0_out[7122] = ~(x[290] & x[292]);
    assign layer0_out[7123] = ~(x[164] & x[175]);
    assign layer0_out[7124] = ~(x[135] ^ x[138]);
    assign layer0_out[7125] = ~x[54] | x[60];
    assign layer0_out[7126] = x[327] & x[339];
    assign layer0_out[7127] = ~(x[308] & x[315]);
    assign layer0_out[7128] = x[142] ^ x[161];
    assign layer0_out[7129] = x[310];
    assign layer0_out[7130] = 1'b1;
    assign layer0_out[7131] = x[284] | x[301];
    assign layer0_out[7132] = x[381] | x[396];
    assign layer0_out[7133] = ~(x[301] ^ x[307]);
    assign layer0_out[7134] = ~(x[45] | x[55]);
    assign layer0_out[7135] = ~x[45];
    assign layer0_out[7136] = ~x[307] | x[295];
    assign layer0_out[7137] = x[162] & ~x[168];
    assign layer0_out[7138] = x[151] ^ x[166];
    assign layer0_out[7139] = ~x[193];
    assign layer0_out[7140] = ~x[113];
    assign layer0_out[7141] = x[172] | x[174];
    assign layer0_out[7142] = x[183] & x[189];
    assign layer0_out[7143] = x[188] ^ x[194];
    assign layer0_out[7144] = ~x[203];
    assign layer0_out[7145] = x[369] ^ x[384];
    assign layer0_out[7146] = ~x[243] | x[231];
    assign layer0_out[7147] = 1'b0;
    assign layer0_out[7148] = ~(x[171] | x[190]);
    assign layer0_out[7149] = x[14] | x[18];
    assign layer0_out[7150] = x[82] | x[83];
    assign layer0_out[7151] = x[101] & ~x[84];
    assign layer0_out[7152] = ~(x[264] ^ x[266]);
    assign layer0_out[7153] = x[102];
    assign layer0_out[7154] = 1'b0;
    assign layer0_out[7155] = x[92] | x[98];
    assign layer0_out[7156] = ~x[17] | x[2];
    assign layer0_out[7157] = ~x[42];
    assign layer0_out[7158] = x[147] ^ x[164];
    assign layer0_out[7159] = x[110] & ~x[125];
    assign layer0_out[7160] = ~x[147];
    assign layer0_out[7161] = ~(x[226] ^ x[243]);
    assign layer0_out[7162] = ~x[355];
    assign layer0_out[7163] = x[97] | x[118];
    assign layer0_out[7164] = x[307] | x[310];
    assign layer0_out[7165] = x[224];
    assign layer0_out[7166] = ~x[105];
    assign layer0_out[7167] = x[121] | x[130];
    assign layer0_out[7168] = x[173];
    assign layer0_out[7169] = ~(x[269] | x[289]);
    assign layer0_out[7170] = ~(x[224] ^ x[236]);
    assign layer0_out[7171] = ~(x[239] | x[245]);
    assign layer0_out[7172] = ~(x[176] ^ x[187]);
    assign layer0_out[7173] = x[333] & ~x[339];
    assign layer0_out[7174] = ~(x[146] & x[161]);
    assign layer0_out[7175] = x[296];
    assign layer0_out[7176] = ~(x[301] & x[315]);
    assign layer0_out[7177] = x[119] & x[122];
    assign layer0_out[7178] = x[238];
    assign layer0_out[7179] = x[70] | x[78];
    assign layer0_out[7180] = x[155] & ~x[152];
    assign layer0_out[7181] = ~(x[269] ^ x[288]);
    assign layer0_out[7182] = x[27] ^ x[29];
    assign layer0_out[7183] = 1'b0;
    assign layer0_out[7184] = ~x[294] | x[295];
    assign layer0_out[7185] = x[234];
    assign layer0_out[7186] = x[368] & ~x[366];
    assign layer0_out[7187] = x[266];
    assign layer0_out[7188] = 1'b1;
    assign layer0_out[7189] = 1'b1;
    assign layer0_out[7190] = ~x[183] | x[190];
    assign layer0_out[7191] = x[100] ^ x[113];
    assign layer0_out[7192] = ~(x[204] ^ x[214]);
    assign layer0_out[7193] = x[269];
    assign layer0_out[7194] = ~x[29];
    assign layer0_out[7195] = x[160];
    assign layer0_out[7196] = ~x[31] | x[17];
    assign layer0_out[7197] = ~(x[281] | x[287]);
    assign layer0_out[7198] = ~(x[373] | x[374]);
    assign layer0_out[7199] = ~x[373];
    assign layer0_out[7200] = 1'b0;
    assign layer0_out[7201] = ~x[0] | x[19];
    assign layer0_out[7202] = ~x[309] | x[317];
    assign layer0_out[7203] = x[358] & ~x[378];
    assign layer0_out[7204] = ~x[97];
    assign layer0_out[7205] = ~x[128];
    assign layer0_out[7206] = x[109];
    assign layer0_out[7207] = ~(x[338] ^ x[348]);
    assign layer0_out[7208] = ~x[198];
    assign layer0_out[7209] = ~(x[384] ^ x[391]);
    assign layer0_out[7210] = ~(x[359] & x[379]);
    assign layer0_out[7211] = x[27];
    assign layer0_out[7212] = ~(x[140] | x[143]);
    assign layer0_out[7213] = ~(x[141] ^ x[146]);
    assign layer0_out[7214] = ~(x[343] | x[354]);
    assign layer0_out[7215] = x[95] ^ x[113];
    assign layer0_out[7216] = ~x[193];
    assign layer0_out[7217] = ~(x[187] | x[188]);
    assign layer0_out[7218] = x[312];
    assign layer0_out[7219] = x[103];
    assign layer0_out[7220] = x[155] & ~x[143];
    assign layer0_out[7221] = x[274];
    assign layer0_out[7222] = 1'b1;
    assign layer0_out[7223] = x[364];
    assign layer0_out[7224] = x[325];
    assign layer0_out[7225] = ~(x[59] | x[61]);
    assign layer0_out[7226] = ~x[161];
    assign layer0_out[7227] = x[170] ^ x[181];
    assign layer0_out[7228] = ~(x[215] & x[221]);
    assign layer0_out[7229] = x[50] & ~x[33];
    assign layer0_out[7230] = 1'b1;
    assign layer0_out[7231] = ~x[330];
    assign layer0_out[7232] = ~x[140] | x[156];
    assign layer0_out[7233] = ~x[83];
    assign layer0_out[7234] = ~(x[135] | x[153]);
    assign layer0_out[7235] = 1'b0;
    assign layer0_out[7236] = x[90] & x[93];
    assign layer0_out[7237] = x[318];
    assign layer0_out[7238] = ~x[146] | x[158];
    assign layer0_out[7239] = ~(x[31] | x[33]);
    assign layer0_out[7240] = 1'b0;
    assign layer0_out[7241] = ~(x[33] | x[53]);
    assign layer0_out[7242] = ~x[300] | x[293];
    assign layer0_out[7243] = x[165];
    assign layer0_out[7244] = x[53];
    assign layer0_out[7245] = ~(x[101] ^ x[120]);
    assign layer0_out[7246] = ~x[116] | x[113];
    assign layer0_out[7247] = x[147] & ~x[154];
    assign layer0_out[7248] = ~x[289] | x[281];
    assign layer0_out[7249] = x[269] & ~x[262];
    assign layer0_out[7250] = ~(x[1] | x[20]);
    assign layer0_out[7251] = ~(x[185] & x[197]);
    assign layer0_out[7252] = ~(x[232] | x[251]);
    assign layer0_out[7253] = ~(x[43] & x[46]);
    assign layer0_out[7254] = ~x[11];
    assign layer0_out[7255] = ~x[205];
    assign layer0_out[7256] = ~x[28];
    assign layer0_out[7257] = x[216] & ~x[233];
    assign layer0_out[7258] = x[50];
    assign layer0_out[7259] = 1'b1;
    assign layer0_out[7260] = ~(x[289] | x[302]);
    assign layer0_out[7261] = 1'b0;
    assign layer0_out[7262] = x[21] | x[39];
    assign layer0_out[7263] = ~x[147];
    assign layer0_out[7264] = ~x[326] | x[312];
    assign layer0_out[7265] = ~x[164];
    assign layer0_out[7266] = ~x[210] | x[208];
    assign layer0_out[7267] = x[347] & ~x[357];
    assign layer0_out[7268] = x[193] & ~x[182];
    assign layer0_out[7269] = ~(x[376] | x[395]);
    assign layer0_out[7270] = x[264] | x[284];
    assign layer0_out[7271] = x[96];
    assign layer0_out[7272] = x[251];
    assign layer0_out[7273] = x[155] | x[160];
    assign layer0_out[7274] = x[129] | x[148];
    assign layer0_out[7275] = ~x[48] | x[61];
    assign layer0_out[7276] = ~(x[378] & x[381]);
    assign layer0_out[7277] = ~x[105] | x[121];
    assign layer0_out[7278] = ~x[215];
    assign layer0_out[7279] = ~(x[174] | x[195]);
    assign layer0_out[7280] = ~x[7];
    assign layer0_out[7281] = ~(x[166] ^ x[183]);
    assign layer0_out[7282] = x[361] ^ x[368];
    assign layer0_out[7283] = x[185] ^ x[187];
    assign layer0_out[7284] = x[121] & ~x[106];
    assign layer0_out[7285] = ~(x[181] ^ x[194]);
    assign layer0_out[7286] = ~x[142];
    assign layer0_out[7287] = x[90] ^ x[107];
    assign layer0_out[7288] = ~x[277];
    assign layer0_out[7289] = ~x[308] | x[306];
    assign layer0_out[7290] = ~x[390] | x[386];
    assign layer0_out[7291] = x[72] | x[80];
    assign layer0_out[7292] = ~(x[93] & x[109]);
    assign layer0_out[7293] = x[11] & ~x[14];
    assign layer0_out[7294] = x[86] | x[87];
    assign layer0_out[7295] = ~x[47];
    assign layer0_out[7296] = 1'b0;
    assign layer0_out[7297] = x[262];
    assign layer0_out[7298] = ~(x[256] | x[260]);
    assign layer0_out[7299] = x[277] | x[284];
    assign layer0_out[7300] = x[230];
    assign layer0_out[7301] = ~x[388];
    assign layer0_out[7302] = x[334] & ~x[333];
    assign layer0_out[7303] = ~(x[329] | x[347]);
    assign layer0_out[7304] = x[285] ^ x[288];
    assign layer0_out[7305] = x[111] & x[116];
    assign layer0_out[7306] = x[101] & ~x[95];
    assign layer0_out[7307] = x[387] & ~x[399];
    assign layer0_out[7308] = x[70] & x[80];
    assign layer0_out[7309] = ~x[240];
    assign layer0_out[7310] = ~(x[13] | x[25]);
    assign layer0_out[7311] = ~(x[363] ^ x[374]);
    assign layer0_out[7312] = x[336] ^ x[356];
    assign layer0_out[7313] = ~(x[211] & x[227]);
    assign layer0_out[7314] = ~x[151] | x[152];
    assign layer0_out[7315] = ~(x[93] | x[96]);
    assign layer0_out[7316] = x[241] & x[249];
    assign layer0_out[7317] = ~(x[209] & x[227]);
    assign layer0_out[7318] = x[269];
    assign layer0_out[7319] = x[123] | x[125];
    assign layer0_out[7320] = x[254];
    assign layer0_out[7321] = x[101] & x[103];
    assign layer0_out[7322] = ~(x[357] | x[372]);
    assign layer0_out[7323] = x[9];
    assign layer0_out[7324] = ~x[326] | x[321];
    assign layer0_out[7325] = x[186];
    assign layer0_out[7326] = x[194];
    assign layer0_out[7327] = ~x[386];
    assign layer0_out[7328] = 1'b1;
    assign layer0_out[7329] = x[128];
    assign layer0_out[7330] = 1'b1;
    assign layer0_out[7331] = x[257] | x[274];
    assign layer0_out[7332] = ~x[265] | x[266];
    assign layer0_out[7333] = ~(x[257] | x[265]);
    assign layer0_out[7334] = ~(x[136] ^ x[142]);
    assign layer0_out[7335] = x[313] & x[328];
    assign layer0_out[7336] = x[289];
    assign layer0_out[7337] = ~x[103] | x[95];
    assign layer0_out[7338] = x[252];
    assign layer0_out[7339] = 1'b1;
    assign layer0_out[7340] = ~(x[131] | x[139]);
    assign layer0_out[7341] = x[151];
    assign layer0_out[7342] = x[244] | x[252];
    assign layer0_out[7343] = x[69];
    assign layer0_out[7344] = ~(x[195] & x[201]);
    assign layer0_out[7345] = ~x[327];
    assign layer0_out[7346] = ~(x[154] | x[156]);
    assign layer0_out[7347] = x[143];
    assign layer0_out[7348] = x[303] ^ x[319];
    assign layer0_out[7349] = ~x[281];
    assign layer0_out[7350] = ~(x[51] ^ x[60]);
    assign layer0_out[7351] = ~(x[136] | x[138]);
    assign layer0_out[7352] = x[145] & ~x[137];
    assign layer0_out[7353] = ~(x[87] | x[106]);
    assign layer0_out[7354] = x[334] | x[338];
    assign layer0_out[7355] = 1'b1;
    assign layer0_out[7356] = ~x[270] | x[262];
    assign layer0_out[7357] = ~x[370];
    assign layer0_out[7358] = x[357] | x[370];
    assign layer0_out[7359] = x[124] & ~x[114];
    assign layer0_out[7360] = ~(x[354] ^ x[359]);
    assign layer0_out[7361] = x[286] & ~x[270];
    assign layer0_out[7362] = ~x[70];
    assign layer0_out[7363] = 1'b0;
    assign layer0_out[7364] = ~x[37];
    assign layer0_out[7365] = ~(x[326] & x[339]);
    assign layer0_out[7366] = ~x[141];
    assign layer0_out[7367] = x[176] & ~x[185];
    assign layer0_out[7368] = 1'b1;
    assign layer0_out[7369] = ~x[40] | x[29];
    assign layer0_out[7370] = x[212] ^ x[232];
    assign layer0_out[7371] = x[190];
    assign layer0_out[7372] = ~(x[351] & x[366]);
    assign layer0_out[7373] = ~(x[244] | x[246]);
    assign layer0_out[7374] = ~(x[294] | x[306]);
    assign layer0_out[7375] = ~x[292] | x[291];
    assign layer0_out[7376] = x[266] ^ x[271];
    assign layer0_out[7377] = x[281] ^ x[294];
    assign layer0_out[7378] = ~x[257];
    assign layer0_out[7379] = x[159];
    assign layer0_out[7380] = ~(x[293] | x[312]);
    assign layer0_out[7381] = x[216] | x[236];
    assign layer0_out[7382] = ~(x[160] | x[170]);
    assign layer0_out[7383] = x[364];
    assign layer0_out[7384] = ~(x[284] | x[298]);
    assign layer0_out[7385] = x[66];
    assign layer0_out[7386] = x[75];
    assign layer0_out[7387] = x[122] | x[136];
    assign layer0_out[7388] = ~x[321];
    assign layer0_out[7389] = 1'b1;
    assign layer0_out[7390] = x[156] ^ x[170];
    assign layer0_out[7391] = ~x[59];
    assign layer0_out[7392] = ~x[95];
    assign layer0_out[7393] = ~(x[317] & x[327]);
    assign layer0_out[7394] = x[345];
    assign layer0_out[7395] = x[57];
    assign layer0_out[7396] = x[47] | x[66];
    assign layer0_out[7397] = ~x[212];
    assign layer0_out[7398] = ~x[171] | x[182];
    assign layer0_out[7399] = ~x[51];
    assign layer0_out[7400] = x[327] & ~x[324];
    assign layer0_out[7401] = ~(x[222] | x[224]);
    assign layer0_out[7402] = x[160];
    assign layer0_out[7403] = ~x[158] | x[149];
    assign layer0_out[7404] = x[97] & ~x[112];
    assign layer0_out[7405] = x[379];
    assign layer0_out[7406] = x[52];
    assign layer0_out[7407] = x[296] & ~x[279];
    assign layer0_out[7408] = x[254];
    assign layer0_out[7409] = ~(x[0] | x[7]);
    assign layer0_out[7410] = ~(x[196] ^ x[201]);
    assign layer0_out[7411] = x[279] & x[299];
    assign layer0_out[7412] = x[185] & ~x[180];
    assign layer0_out[7413] = ~(x[16] | x[31]);
    assign layer0_out[7414] = ~x[122] | x[132];
    assign layer0_out[7415] = ~x[88] | x[100];
    assign layer0_out[7416] = ~x[164];
    assign layer0_out[7417] = x[36];
    assign layer0_out[7418] = ~x[73] | x[91];
    assign layer0_out[7419] = x[79];
    assign layer0_out[7420] = ~x[124];
    assign layer0_out[7421] = x[234];
    assign layer0_out[7422] = x[176];
    assign layer0_out[7423] = ~x[138];
    assign layer0_out[7424] = ~x[303];
    assign layer0_out[7425] = x[93] & ~x[112];
    assign layer0_out[7426] = ~(x[365] | x[374]);
    assign layer0_out[7427] = ~(x[231] | x[241]);
    assign layer0_out[7428] = x[231] & ~x[222];
    assign layer0_out[7429] = x[256];
    assign layer0_out[7430] = ~x[172];
    assign layer0_out[7431] = ~x[81];
    assign layer0_out[7432] = x[96];
    assign layer0_out[7433] = ~x[274];
    assign layer0_out[7434] = x[282] | x[299];
    assign layer0_out[7435] = 1'b1;
    assign layer0_out[7436] = x[12] & x[20];
    assign layer0_out[7437] = x[259] & ~x[241];
    assign layer0_out[7438] = ~(x[302] | x[305]);
    assign layer0_out[7439] = ~x[390];
    assign layer0_out[7440] = ~(x[90] ^ x[108]);
    assign layer0_out[7441] = 1'b1;
    assign layer0_out[7442] = ~x[324];
    assign layer0_out[7443] = ~(x[234] ^ x[250]);
    assign layer0_out[7444] = ~(x[322] ^ x[337]);
    assign layer0_out[7445] = ~x[227];
    assign layer0_out[7446] = x[177];
    assign layer0_out[7447] = 1'b1;
    assign layer0_out[7448] = ~x[286];
    assign layer0_out[7449] = ~x[351];
    assign layer0_out[7450] = x[129] | x[143];
    assign layer0_out[7451] = ~(x[266] | x[285]);
    assign layer0_out[7452] = x[174] & x[193];
    assign layer0_out[7453] = x[392];
    assign layer0_out[7454] = x[164];
    assign layer0_out[7455] = x[178] & x[196];
    assign layer0_out[7456] = ~(x[50] | x[68]);
    assign layer0_out[7457] = x[98] ^ x[112];
    assign layer0_out[7458] = ~x[138];
    assign layer0_out[7459] = ~(x[0] & x[9]);
    assign layer0_out[7460] = ~x[289];
    assign layer0_out[7461] = x[77] & ~x[75];
    assign layer0_out[7462] = x[362] & x[379];
    assign layer0_out[7463] = ~(x[128] | x[148]);
    assign layer0_out[7464] = ~x[365];
    assign layer0_out[7465] = 1'b1;
    assign layer0_out[7466] = 1'b0;
    assign layer0_out[7467] = x[329] & ~x[310];
    assign layer0_out[7468] = ~(x[43] | x[60]);
    assign layer0_out[7469] = x[389] & ~x[378];
    assign layer0_out[7470] = ~(x[138] & x[149]);
    assign layer0_out[7471] = ~(x[85] | x[101]);
    assign layer0_out[7472] = x[354] ^ x[357];
    assign layer0_out[7473] = ~x[317];
    assign layer0_out[7474] = ~(x[221] | x[225]);
    assign layer0_out[7475] = x[287];
    assign layer0_out[7476] = ~(x[93] | x[104]);
    assign layer0_out[7477] = ~x[296];
    assign layer0_out[7478] = ~x[223] | x[209];
    assign layer0_out[7479] = x[47] & ~x[57];
    assign layer0_out[7480] = ~x[355];
    assign layer0_out[7481] = x[304];
    assign layer0_out[7482] = x[225] & ~x[236];
    assign layer0_out[7483] = x[246];
    assign layer0_out[7484] = ~x[206];
    assign layer0_out[7485] = x[144];
    assign layer0_out[7486] = x[71];
    assign layer0_out[7487] = ~(x[105] | x[106]);
    assign layer0_out[7488] = x[81] ^ x[92];
    assign layer0_out[7489] = ~x[30] | x[17];
    assign layer0_out[7490] = x[166] | x[187];
    assign layer0_out[7491] = ~x[364];
    assign layer0_out[7492] = ~(x[145] ^ x[163]);
    assign layer0_out[7493] = 1'b1;
    assign layer0_out[7494] = ~x[170];
    assign layer0_out[7495] = ~(x[294] | x[304]);
    assign layer0_out[7496] = ~(x[185] ^ x[203]);
    assign layer0_out[7497] = ~(x[375] & x[393]);
    assign layer0_out[7498] = ~x[258];
    assign layer0_out[7499] = ~x[361];
    assign layer0_out[7500] = x[195];
    assign layer0_out[7501] = ~x[82];
    assign layer0_out[7502] = ~x[320];
    assign layer0_out[7503] = ~(x[364] ^ x[382]);
    assign layer0_out[7504] = ~x[213] | x[211];
    assign layer0_out[7505] = ~(x[14] | x[21]);
    assign layer0_out[7506] = x[211];
    assign layer0_out[7507] = ~(x[78] | x[88]);
    assign layer0_out[7508] = ~x[375];
    assign layer0_out[7509] = ~(x[185] ^ x[188]);
    assign layer0_out[7510] = x[71] | x[91];
    assign layer0_out[7511] = x[171] ^ x[175];
    assign layer0_out[7512] = ~x[340] | x[335];
    assign layer0_out[7513] = ~(x[314] ^ x[316]);
    assign layer0_out[7514] = ~(x[314] | x[315]);
    assign layer0_out[7515] = x[263] & x[282];
    assign layer0_out[7516] = ~x[233] | x[252];
    assign layer0_out[7517] = ~x[205] | x[211];
    assign layer0_out[7518] = x[27] ^ x[43];
    assign layer0_out[7519] = ~(x[24] | x[40]);
    assign layer0_out[7520] = x[84] ^ x[102];
    assign layer0_out[7521] = 1'b0;
    assign layer0_out[7522] = ~x[30] | x[12];
    assign layer0_out[7523] = x[127];
    assign layer0_out[7524] = ~(x[123] | x[128]);
    assign layer0_out[7525] = ~x[300];
    assign layer0_out[7526] = ~x[264];
    assign layer0_out[7527] = ~x[158] | x[161];
    assign layer0_out[7528] = x[63];
    assign layer0_out[7529] = x[317] & x[322];
    assign layer0_out[7530] = 1'b1;
    assign layer0_out[7531] = x[188] & x[199];
    assign layer0_out[7532] = x[265];
    assign layer0_out[7533] = x[244];
    assign layer0_out[7534] = ~x[103];
    assign layer0_out[7535] = ~x[265];
    assign layer0_out[7536] = x[89] & ~x[93];
    assign layer0_out[7537] = ~(x[230] | x[249]);
    assign layer0_out[7538] = x[19];
    assign layer0_out[7539] = ~(x[64] | x[74]);
    assign layer0_out[7540] = ~x[232] | x[234];
    assign layer0_out[7541] = ~x[197] | x[187];
    assign layer0_out[7542] = ~(x[125] ^ x[137]);
    assign layer0_out[7543] = ~x[363];
    assign layer0_out[7544] = x[189] & ~x[196];
    assign layer0_out[7545] = x[22] & x[34];
    assign layer0_out[7546] = ~x[41];
    assign layer0_out[7547] = x[333];
    assign layer0_out[7548] = ~x[384];
    assign layer0_out[7549] = ~(x[210] | x[222]);
    assign layer0_out[7550] = x[216];
    assign layer0_out[7551] = x[25] | x[31];
    assign layer0_out[7552] = ~(x[202] | x[220]);
    assign layer0_out[7553] = 1'b0;
    assign layer0_out[7554] = x[339] | x[343];
    assign layer0_out[7555] = x[310] & x[318];
    assign layer0_out[7556] = x[21] | x[35];
    assign layer0_out[7557] = x[89];
    assign layer0_out[7558] = ~(x[2] | x[18]);
    assign layer0_out[7559] = 1'b0;
    assign layer0_out[7560] = ~(x[110] & x[115]);
    assign layer0_out[7561] = x[82];
    assign layer0_out[7562] = ~(x[238] ^ x[254]);
    assign layer0_out[7563] = x[102] | x[120];
    assign layer0_out[7564] = x[66] | x[78];
    assign layer0_out[7565] = 1'b1;
    assign layer0_out[7566] = ~x[216] | x[224];
    assign layer0_out[7567] = ~x[53] | x[50];
    assign layer0_out[7568] = x[334] | x[335];
    assign layer0_out[7569] = ~x[100] | x[119];
    assign layer0_out[7570] = ~x[329] | x[337];
    assign layer0_out[7571] = ~x[303];
    assign layer0_out[7572] = ~x[395];
    assign layer0_out[7573] = ~(x[211] | x[229]);
    assign layer0_out[7574] = 1'b1;
    assign layer0_out[7575] = ~x[103] | x[109];
    assign layer0_out[7576] = ~x[396];
    assign layer0_out[7577] = ~(x[322] | x[330]);
    assign layer0_out[7578] = x[189];
    assign layer0_out[7579] = x[335] | x[355];
    assign layer0_out[7580] = ~(x[189] & x[193]);
    assign layer0_out[7581] = ~x[321] | x[339];
    assign layer0_out[7582] = x[291] ^ x[293];
    assign layer0_out[7583] = x[149] ^ x[157];
    assign layer0_out[7584] = ~(x[28] | x[41]);
    assign layer0_out[7585] = ~(x[185] ^ x[201]);
    assign layer0_out[7586] = x[172] & x[173];
    assign layer0_out[7587] = x[238] | x[244];
    assign layer0_out[7588] = ~(x[365] | x[366]);
    assign layer0_out[7589] = ~(x[21] & x[41]);
    assign layer0_out[7590] = ~(x[180] | x[184]);
    assign layer0_out[7591] = x[194] | x[195];
    assign layer0_out[7592] = x[269] ^ x[285];
    assign layer0_out[7593] = x[301];
    assign layer0_out[7594] = ~x[157];
    assign layer0_out[7595] = ~(x[158] | x[174]);
    assign layer0_out[7596] = x[216] | x[217];
    assign layer0_out[7597] = ~x[336] | x[344];
    assign layer0_out[7598] = ~x[246];
    assign layer0_out[7599] = x[371];
    assign layer0_out[7600] = ~x[301];
    assign layer0_out[7601] = ~(x[206] ^ x[213]);
    assign layer0_out[7602] = x[170];
    assign layer0_out[7603] = x[14];
    assign layer0_out[7604] = ~x[44];
    assign layer0_out[7605] = ~x[80];
    assign layer0_out[7606] = ~(x[234] | x[247]);
    assign layer0_out[7607] = ~x[217];
    assign layer0_out[7608] = ~(x[391] | x[392]);
    assign layer0_out[7609] = x[316] & x[327];
    assign layer0_out[7610] = ~(x[45] | x[51]);
    assign layer0_out[7611] = x[161];
    assign layer0_out[7612] = 1'b1;
    assign layer0_out[7613] = x[104] | x[105];
    assign layer0_out[7614] = x[221];
    assign layer0_out[7615] = x[101];
    assign layer0_out[7616] = ~(x[48] & x[58]);
    assign layer0_out[7617] = ~x[274];
    assign layer0_out[7618] = x[350];
    assign layer0_out[7619] = ~(x[139] | x[160]);
    assign layer0_out[7620] = ~x[164];
    assign layer0_out[7621] = ~(x[174] & x[191]);
    assign layer0_out[7622] = x[168] & ~x[188];
    assign layer0_out[7623] = x[139] & ~x[138];
    assign layer0_out[7624] = x[222] | x[234];
    assign layer0_out[7625] = ~(x[19] | x[21]);
    assign layer0_out[7626] = x[271] ^ x[288];
    assign layer0_out[7627] = ~(x[281] | x[293]);
    assign layer0_out[7628] = x[179] & ~x[170];
    assign layer0_out[7629] = ~x[275];
    assign layer0_out[7630] = x[68] | x[75];
    assign layer0_out[7631] = x[334] ^ x[354];
    assign layer0_out[7632] = ~(x[109] | x[123]);
    assign layer0_out[7633] = x[78] | x[98];
    assign layer0_out[7634] = ~(x[66] & x[70]);
    assign layer0_out[7635] = x[200] & ~x[218];
    assign layer0_out[7636] = x[188] & ~x[186];
    assign layer0_out[7637] = ~(x[11] & x[22]);
    assign layer0_out[7638] = ~(x[257] | x[258]);
    assign layer0_out[7639] = x[39] & ~x[54];
    assign layer0_out[7640] = 1'b1;
    assign layer0_out[7641] = ~(x[136] & x[152]);
    assign layer0_out[7642] = ~x[150];
    assign layer0_out[7643] = 1'b0;
    assign layer0_out[7644] = 1'b1;
    assign layer0_out[7645] = 1'b0;
    assign layer0_out[7646] = x[183];
    assign layer0_out[7647] = ~(x[235] ^ x[245]);
    assign layer0_out[7648] = ~x[106];
    assign layer0_out[7649] = x[137];
    assign layer0_out[7650] = ~(x[206] | x[209]);
    assign layer0_out[7651] = 1'b0;
    assign layer0_out[7652] = x[280] & ~x[292];
    assign layer0_out[7653] = x[238] | x[250];
    assign layer0_out[7654] = x[347] ^ x[362];
    assign layer0_out[7655] = x[101] | x[118];
    assign layer0_out[7656] = ~(x[304] & x[310]);
    assign layer0_out[7657] = x[64];
    assign layer0_out[7658] = 1'b1;
    assign layer0_out[7659] = ~(x[314] ^ x[323]);
    assign layer0_out[7660] = ~x[395] | x[385];
    assign layer0_out[7661] = x[313] & x[329];
    assign layer0_out[7662] = x[284];
    assign layer0_out[7663] = x[94] | x[114];
    assign layer0_out[7664] = ~x[218];
    assign layer0_out[7665] = ~x[177] | x[176];
    assign layer0_out[7666] = x[41];
    assign layer0_out[7667] = ~x[385] | x[372];
    assign layer0_out[7668] = x[366] | x[376];
    assign layer0_out[7669] = x[32] & ~x[22];
    assign layer0_out[7670] = x[347] | x[365];
    assign layer0_out[7671] = ~x[73];
    assign layer0_out[7672] = x[184] | x[189];
    assign layer0_out[7673] = ~x[18];
    assign layer0_out[7674] = x[366] | x[367];
    assign layer0_out[7675] = 1'b1;
    assign layer0_out[7676] = x[63];
    assign layer0_out[7677] = ~x[66];
    assign layer0_out[7678] = ~(x[166] ^ x[168]);
    assign layer0_out[7679] = ~x[239];
    assign layer0_out[7680] = ~(x[97] | x[117]);
    assign layer0_out[7681] = ~(x[255] & x[265]);
    assign layer0_out[7682] = x[64] | x[82];
    assign layer0_out[7683] = x[248];
    assign layer0_out[7684] = ~(x[116] & x[123]);
    assign layer0_out[7685] = x[198] | x[207];
    assign layer0_out[7686] = x[101];
    assign layer0_out[7687] = ~x[283];
    assign layer0_out[7688] = ~x[277];
    assign layer0_out[7689] = x[347] ^ x[358];
    assign layer0_out[7690] = ~x[318] | x[321];
    assign layer0_out[7691] = x[337];
    assign layer0_out[7692] = x[64] & ~x[77];
    assign layer0_out[7693] = 1'b1;
    assign layer0_out[7694] = x[96];
    assign layer0_out[7695] = x[245] & ~x[234];
    assign layer0_out[7696] = 1'b1;
    assign layer0_out[7697] = ~(x[100] | x[110]);
    assign layer0_out[7698] = ~(x[154] ^ x[159]);
    assign layer0_out[7699] = x[200] & ~x[202];
    assign layer0_out[7700] = x[85];
    assign layer0_out[7701] = 1'b1;
    assign layer0_out[7702] = x[148];
    assign layer0_out[7703] = ~x[249];
    assign layer0_out[7704] = x[394] & ~x[385];
    assign layer0_out[7705] = x[332];
    assign layer0_out[7706] = ~x[186] | x[199];
    assign layer0_out[7707] = ~(x[179] ^ x[186]);
    assign layer0_out[7708] = ~(x[76] | x[77]);
    assign layer0_out[7709] = ~(x[55] | x[75]);
    assign layer0_out[7710] = 1'b0;
    assign layer0_out[7711] = ~(x[350] ^ x[360]);
    assign layer0_out[7712] = ~(x[80] | x[83]);
    assign layer0_out[7713] = ~(x[147] & x[159]);
    assign layer0_out[7714] = ~x[291];
    assign layer0_out[7715] = x[242] | x[261];
    assign layer0_out[7716] = x[348];
    assign layer0_out[7717] = x[243] ^ x[263];
    assign layer0_out[7718] = ~x[213];
    assign layer0_out[7719] = x[12] | x[18];
    assign layer0_out[7720] = ~x[134] | x[127];
    assign layer0_out[7721] = x[384];
    assign layer0_out[7722] = ~(x[365] | x[373]);
    assign layer0_out[7723] = ~(x[264] & x[282]);
    assign layer0_out[7724] = x[7];
    assign layer0_out[7725] = ~x[383] | x[372];
    assign layer0_out[7726] = x[386] & ~x[384];
    assign layer0_out[7727] = x[73] & ~x[62];
    assign layer0_out[7728] = ~(x[129] | x[141]);
    assign layer0_out[7729] = ~(x[41] | x[59]);
    assign layer0_out[7730] = x[142];
    assign layer0_out[7731] = x[219];
    assign layer0_out[7732] = ~(x[322] | x[324]);
    assign layer0_out[7733] = ~x[277];
    assign layer0_out[7734] = 1'b0;
    assign layer0_out[7735] = ~(x[193] | x[212]);
    assign layer0_out[7736] = x[305] & ~x[290];
    assign layer0_out[7737] = ~x[178];
    assign layer0_out[7738] = ~x[127] | x[119];
    assign layer0_out[7739] = x[209] & ~x[200];
    assign layer0_out[7740] = ~(x[345] & x[347]);
    assign layer0_out[7741] = ~x[346] | x[339];
    assign layer0_out[7742] = x[30];
    assign layer0_out[7743] = ~(x[59] ^ x[77]);
    assign layer0_out[7744] = ~(x[328] | x[343]);
    assign layer0_out[7745] = x[342] | x[360];
    assign layer0_out[7746] = ~x[28];
    assign layer0_out[7747] = x[73];
    assign layer0_out[7748] = x[17] & ~x[13];
    assign layer0_out[7749] = ~x[128];
    assign layer0_out[7750] = x[237];
    assign layer0_out[7751] = x[9] ^ x[18];
    assign layer0_out[7752] = 1'b0;
    assign layer0_out[7753] = x[189] | x[209];
    assign layer0_out[7754] = x[221] ^ x[224];
    assign layer0_out[7755] = x[264] | x[265];
    assign layer0_out[7756] = x[139] & x[142];
    assign layer0_out[7757] = ~(x[256] ^ x[261]);
    assign layer0_out[7758] = x[20] & ~x[13];
    assign layer0_out[7759] = ~x[78] | x[83];
    assign layer0_out[7760] = x[73];
    assign layer0_out[7761] = x[199] & ~x[208];
    assign layer0_out[7762] = x[208] ^ x[214];
    assign layer0_out[7763] = x[56];
    assign layer0_out[7764] = x[154];
    assign layer0_out[7765] = ~(x[311] & x[326]);
    assign layer0_out[7766] = ~x[65] | x[76];
    assign layer0_out[7767] = x[323] | x[342];
    assign layer0_out[7768] = ~x[267] | x[256];
    assign layer0_out[7769] = x[119];
    assign layer0_out[7770] = x[354] & ~x[352];
    assign layer0_out[7771] = 1'b1;
    assign layer0_out[7772] = ~(x[364] | x[365]);
    assign layer0_out[7773] = ~(x[165] & x[184]);
    assign layer0_out[7774] = ~x[22] | x[18];
    assign layer0_out[7775] = x[226] & ~x[208];
    assign layer0_out[7776] = ~x[198] | x[205];
    assign layer0_out[7777] = x[28] | x[48];
    assign layer0_out[7778] = 1'b0;
    assign layer0_out[7779] = x[208];
    assign layer0_out[7780] = x[323] & ~x[337];
    assign layer0_out[7781] = ~x[272];
    assign layer0_out[7782] = x[88] | x[102];
    assign layer0_out[7783] = ~x[324] | x[309];
    assign layer0_out[7784] = x[168] & ~x[178];
    assign layer0_out[7785] = ~(x[200] ^ x[203]);
    assign layer0_out[7786] = ~(x[287] ^ x[291]);
    assign layer0_out[7787] = 1'b1;
    assign layer0_out[7788] = x[36] | x[43];
    assign layer0_out[7789] = x[202] | x[216];
    assign layer0_out[7790] = 1'b1;
    assign layer0_out[7791] = ~(x[228] | x[247]);
    assign layer0_out[7792] = x[28] & ~x[19];
    assign layer0_out[7793] = x[106] ^ x[110];
    assign layer0_out[7794] = x[276] | x[280];
    assign layer0_out[7795] = x[373] & ~x[372];
    assign layer0_out[7796] = ~x[106];
    assign layer0_out[7797] = ~x[263] | x[251];
    assign layer0_out[7798] = ~(x[339] & x[355]);
    assign layer0_out[7799] = x[136] ^ x[153];
    assign layer0_out[7800] = ~(x[70] ^ x[77]);
    assign layer0_out[7801] = x[271] | x[284];
    assign layer0_out[7802] = ~x[162];
    assign layer0_out[7803] = ~x[119] | x[115];
    assign layer0_out[7804] = x[369] & ~x[355];
    assign layer0_out[7805] = ~(x[3] | x[24]);
    assign layer0_out[7806] = ~(x[315] ^ x[322]);
    assign layer0_out[7807] = x[258] & ~x[269];
    assign layer0_out[7808] = ~(x[104] | x[107]);
    assign layer0_out[7809] = ~x[297] | x[283];
    assign layer0_out[7810] = x[263] | x[265];
    assign layer0_out[7811] = x[188] | x[206];
    assign layer0_out[7812] = x[143] | x[145];
    assign layer0_out[7813] = x[272] | x[287];
    assign layer0_out[7814] = x[113] | x[134];
    assign layer0_out[7815] = ~x[355];
    assign layer0_out[7816] = x[195] | x[211];
    assign layer0_out[7817] = x[152];
    assign layer0_out[7818] = ~(x[65] | x[84]);
    assign layer0_out[7819] = ~x[34];
    assign layer0_out[7820] = x[237] & x[249];
    assign layer0_out[7821] = ~(x[53] ^ x[61]);
    assign layer0_out[7822] = ~x[382] | x[370];
    assign layer0_out[7823] = x[266] | x[281];
    assign layer0_out[7824] = ~x[122];
    assign layer0_out[7825] = ~x[236];
    assign layer0_out[7826] = ~(x[54] & x[67]);
    assign layer0_out[7827] = ~x[159];
    assign layer0_out[7828] = ~x[232];
    assign layer0_out[7829] = ~(x[107] | x[128]);
    assign layer0_out[7830] = ~x[318];
    assign layer0_out[7831] = ~x[234];
    assign layer0_out[7832] = ~x[33];
    assign layer0_out[7833] = x[227];
    assign layer0_out[7834] = ~x[168];
    assign layer0_out[7835] = ~(x[324] | x[331]);
    assign layer0_out[7836] = ~x[222];
    assign layer0_out[7837] = x[168] & x[184];
    assign layer0_out[7838] = x[282] | x[283];
    assign layer0_out[7839] = ~x[136];
    assign layer0_out[7840] = ~x[41];
    assign layer0_out[7841] = ~x[336];
    assign layer0_out[7842] = ~(x[142] ^ x[148]);
    assign layer0_out[7843] = ~x[157] | x[160];
    assign layer0_out[7844] = ~(x[301] | x[311]);
    assign layer0_out[7845] = ~(x[180] | x[195]);
    assign layer0_out[7846] = ~(x[112] ^ x[133]);
    assign layer0_out[7847] = ~(x[387] & x[395]);
    assign layer0_out[7848] = ~x[29];
    assign layer0_out[7849] = ~(x[282] | x[302]);
    assign layer0_out[7850] = ~x[143];
    assign layer0_out[7851] = x[107];
    assign layer0_out[7852] = 1'b1;
    assign layer0_out[7853] = 1'b0;
    assign layer0_out[7854] = x[171] & ~x[157];
    assign layer0_out[7855] = ~x[67] | x[88];
    assign layer0_out[7856] = x[254] & x[268];
    assign layer0_out[7857] = x[358];
    assign layer0_out[7858] = x[172];
    assign layer0_out[7859] = ~x[284];
    assign layer0_out[7860] = x[97];
    assign layer0_out[7861] = ~x[134] | x[120];
    assign layer0_out[7862] = ~(x[353] | x[358]);
    assign layer0_out[7863] = ~(x[161] | x[180]);
    assign layer0_out[7864] = x[374] | x[392];
    assign layer0_out[7865] = x[285] & ~x[291];
    assign layer0_out[7866] = x[32];
    assign layer0_out[7867] = x[344] ^ x[358];
    assign layer0_out[7868] = ~(x[177] | x[192]);
    assign layer0_out[7869] = ~(x[318] ^ x[323]);
    assign layer0_out[7870] = x[6] ^ x[11];
    assign layer0_out[7871] = x[322];
    assign layer0_out[7872] = ~x[154] | x[145];
    assign layer0_out[7873] = 1'b0;
    assign layer0_out[7874] = x[369] & ~x[357];
    assign layer0_out[7875] = ~x[335];
    assign layer0_out[7876] = x[172] | x[190];
    assign layer0_out[7877] = x[305];
    assign layer0_out[7878] = x[173] & x[188];
    assign layer0_out[7879] = ~(x[164] ^ x[182]);
    assign layer0_out[7880] = ~x[246];
    assign layer0_out[7881] = ~x[224];
    assign layer0_out[7882] = x[26] & ~x[19];
    assign layer0_out[7883] = ~(x[200] & x[206]);
    assign layer0_out[7884] = x[306] & ~x[300];
    assign layer0_out[7885] = ~(x[264] | x[281]);
    assign layer0_out[7886] = ~x[93] | x[86];
    assign layer0_out[7887] = x[262] ^ x[280];
    assign layer0_out[7888] = x[129] ^ x[146];
    assign layer0_out[7889] = ~x[100] | x[114];
    assign layer0_out[7890] = x[281] ^ x[292];
    assign layer0_out[7891] = ~(x[284] & x[288]);
    assign layer0_out[7892] = ~x[177];
    assign layer0_out[7893] = x[12] & ~x[27];
    assign layer0_out[7894] = x[321];
    assign layer0_out[7895] = x[399];
    assign layer0_out[7896] = x[390];
    assign layer0_out[7897] = ~x[173];
    assign layer0_out[7898] = ~(x[151] & x[153]);
    assign layer0_out[7899] = 1'b1;
    assign layer0_out[7900] = ~x[352] | x[342];
    assign layer0_out[7901] = x[126];
    assign layer0_out[7902] = ~x[223];
    assign layer0_out[7903] = ~x[214];
    assign layer0_out[7904] = ~(x[151] & x[172]);
    assign layer0_out[7905] = ~(x[51] | x[58]);
    assign layer0_out[7906] = x[270] | x[289];
    assign layer0_out[7907] = ~x[38] | x[57];
    assign layer0_out[7908] = x[284] | x[297];
    assign layer0_out[7909] = x[26] & ~x[32];
    assign layer0_out[7910] = 1'b0;
    assign layer0_out[7911] = ~(x[99] ^ x[113]);
    assign layer0_out[7912] = x[264] & ~x[244];
    assign layer0_out[7913] = 1'b1;
    assign layer0_out[7914] = x[327] ^ x[344];
    assign layer0_out[7915] = x[219] & x[231];
    assign layer0_out[7916] = ~x[132];
    assign layer0_out[7917] = x[198];
    assign layer0_out[7918] = ~x[46];
    assign layer0_out[7919] = ~x[289];
    assign layer0_out[7920] = x[181];
    assign layer0_out[7921] = ~x[217] | x[234];
    assign layer0_out[7922] = 1'b0;
    assign layer0_out[7923] = ~x[306];
    assign layer0_out[7924] = ~(x[16] & x[24]);
    assign layer0_out[7925] = x[263] | x[266];
    assign layer0_out[7926] = ~x[369];
    assign layer0_out[7927] = ~x[124];
    assign layer0_out[7928] = ~x[118];
    assign layer0_out[7929] = 1'b1;
    assign layer0_out[7930] = x[4];
    assign layer0_out[7931] = x[118] ^ x[134];
    assign layer0_out[7932] = ~(x[204] & x[216]);
    assign layer0_out[7933] = x[89] & ~x[101];
    assign layer0_out[7934] = ~x[335];
    assign layer0_out[7935] = ~(x[211] | x[225]);
    assign layer0_out[7936] = x[331] | x[350];
    assign layer0_out[7937] = x[364] | x[372];
    assign layer0_out[7938] = 1'b1;
    assign layer0_out[7939] = x[204] | x[205];
    assign layer0_out[7940] = ~(x[227] | x[238]);
    assign layer0_out[7941] = ~x[19];
    assign layer0_out[7942] = ~(x[222] & x[232]);
    assign layer0_out[7943] = ~x[305] | x[297];
    assign layer0_out[7944] = ~(x[364] | x[380]);
    assign layer0_out[7945] = ~(x[53] | x[73]);
    assign layer0_out[7946] = x[171];
    assign layer0_out[7947] = 1'b1;
    assign layer0_out[7948] = x[118] | x[139];
    assign layer0_out[7949] = x[175];
    assign layer0_out[7950] = ~x[226];
    assign layer0_out[7951] = ~(x[281] & x[291]);
    assign layer0_out[7952] = 1'b1;
    assign layer0_out[7953] = x[376];
    assign layer0_out[7954] = ~x[183] | x[172];
    assign layer0_out[7955] = x[281] | x[301];
    assign layer0_out[7956] = x[47];
    assign layer0_out[7957] = x[219] | x[230];
    assign layer0_out[7958] = 1'b0;
    assign layer0_out[7959] = x[192];
    assign layer0_out[7960] = x[293] & ~x[307];
    assign layer0_out[7961] = ~x[15];
    assign layer0_out[7962] = x[143] & x[164];
    assign layer0_out[7963] = x[10] & ~x[17];
    assign layer0_out[7964] = ~(x[108] | x[128]);
    assign layer0_out[7965] = ~(x[156] | x[175]);
    assign layer0_out[7966] = ~x[53];
    assign layer0_out[7967] = x[86] & ~x[90];
    assign layer0_out[7968] = ~x[145];
    assign layer0_out[7969] = ~x[254] | x[240];
    assign layer0_out[7970] = ~(x[11] | x[24]);
    assign layer0_out[7971] = x[148] & ~x[138];
    assign layer0_out[7972] = ~x[319];
    assign layer0_out[7973] = x[290] & x[293];
    assign layer0_out[7974] = x[35];
    assign layer0_out[7975] = x[243] | x[244];
    assign layer0_out[7976] = ~(x[248] | x[249]);
    assign layer0_out[7977] = ~x[358] | x[343];
    assign layer0_out[7978] = x[204] ^ x[221];
    assign layer0_out[7979] = 1'b0;
    assign layer0_out[7980] = ~(x[142] | x[147]);
    assign layer0_out[7981] = ~x[189] | x[203];
    assign layer0_out[7982] = x[72] & x[77];
    assign layer0_out[7983] = ~(x[167] & x[171]);
    assign layer0_out[7984] = ~(x[293] & x[305]);
    assign layer0_out[7985] = x[185] & ~x[167];
    assign layer0_out[7986] = ~x[375] | x[372];
    assign layer0_out[7987] = x[295] & ~x[306];
    assign layer0_out[7988] = ~x[129] | x[119];
    assign layer0_out[7989] = x[391] & x[395];
    assign layer0_out[7990] = ~x[212];
    assign layer0_out[7991] = ~(x[267] | x[286]);
    assign layer0_out[7992] = ~x[99] | x[78];
    assign layer0_out[7993] = ~(x[163] | x[176]);
    assign layer0_out[7994] = ~x[166];
    assign layer0_out[7995] = x[43];
    assign layer0_out[7996] = x[84] & x[90];
    assign layer0_out[7997] = x[269] & ~x[272];
    assign layer0_out[7998] = ~(x[376] | x[380]);
    assign layer0_out[7999] = x[54] | x[57];
    assign layer1_out[0] = layer0_out[7772];
    assign layer1_out[1] = ~layer0_out[4567] | layer0_out[4568];
    assign layer1_out[2] = layer0_out[6876] & layer0_out[6877];
    assign layer1_out[3] = ~layer0_out[2970] | layer0_out[2969];
    assign layer1_out[4] = ~layer0_out[352];
    assign layer1_out[5] = layer0_out[284] & ~layer0_out[285];
    assign layer1_out[6] = ~layer0_out[5512];
    assign layer1_out[7] = layer0_out[1429];
    assign layer1_out[8] = layer0_out[2064];
    assign layer1_out[9] = ~(layer0_out[1453] & layer0_out[1454]);
    assign layer1_out[10] = layer0_out[6960] & layer0_out[6961];
    assign layer1_out[11] = 1'b0;
    assign layer1_out[12] = layer0_out[7536] ^ layer0_out[7537];
    assign layer1_out[13] = layer0_out[6226] ^ layer0_out[6227];
    assign layer1_out[14] = 1'b1;
    assign layer1_out[15] = layer0_out[3143] | layer0_out[3144];
    assign layer1_out[16] = layer0_out[3570] | layer0_out[3571];
    assign layer1_out[17] = ~(layer0_out[789] | layer0_out[790]);
    assign layer1_out[18] = layer0_out[1117] & ~layer0_out[1118];
    assign layer1_out[19] = ~(layer0_out[5246] ^ layer0_out[5247]);
    assign layer1_out[20] = layer0_out[5500] & layer0_out[5501];
    assign layer1_out[21] = layer0_out[4421] | layer0_out[4422];
    assign layer1_out[22] = ~layer0_out[3141] | layer0_out[3140];
    assign layer1_out[23] = layer0_out[4616] & ~layer0_out[4617];
    assign layer1_out[24] = layer0_out[4532] | layer0_out[4533];
    assign layer1_out[25] = layer0_out[3025];
    assign layer1_out[26] = layer0_out[5533];
    assign layer1_out[27] = ~(layer0_out[71] | layer0_out[72]);
    assign layer1_out[28] = layer0_out[943];
    assign layer1_out[29] = ~layer0_out[3314];
    assign layer1_out[30] = layer0_out[6395];
    assign layer1_out[31] = ~(layer0_out[6970] & layer0_out[6971]);
    assign layer1_out[32] = layer0_out[299];
    assign layer1_out[33] = layer0_out[556] & layer0_out[557];
    assign layer1_out[34] = ~layer0_out[3106] | layer0_out[3105];
    assign layer1_out[35] = layer0_out[7496] & ~layer0_out[7495];
    assign layer1_out[36] = layer0_out[1263] | layer0_out[1264];
    assign layer1_out[37] = ~layer0_out[4304];
    assign layer1_out[38] = ~(layer0_out[5225] & layer0_out[5226]);
    assign layer1_out[39] = ~layer0_out[5856];
    assign layer1_out[40] = layer0_out[3805] | layer0_out[3806];
    assign layer1_out[41] = 1'b0;
    assign layer1_out[42] = layer0_out[1076] & ~layer0_out[1077];
    assign layer1_out[43] = ~(layer0_out[1203] | layer0_out[1204]);
    assign layer1_out[44] = ~(layer0_out[7840] & layer0_out[7841]);
    assign layer1_out[45] = ~layer0_out[1667] | layer0_out[1668];
    assign layer1_out[46] = ~layer0_out[5085];
    assign layer1_out[47] = layer0_out[3901];
    assign layer1_out[48] = 1'b1;
    assign layer1_out[49] = layer0_out[1388] & ~layer0_out[1389];
    assign layer1_out[50] = layer0_out[1055];
    assign layer1_out[51] = ~(layer0_out[2302] ^ layer0_out[2303]);
    assign layer1_out[52] = layer0_out[397];
    assign layer1_out[53] = ~layer0_out[1517];
    assign layer1_out[54] = layer0_out[4077];
    assign layer1_out[55] = layer0_out[3690] & ~layer0_out[3689];
    assign layer1_out[56] = layer0_out[7946];
    assign layer1_out[57] = ~(layer0_out[5795] | layer0_out[5796]);
    assign layer1_out[58] = layer0_out[6256];
    assign layer1_out[59] = ~(layer0_out[4214] | layer0_out[4215]);
    assign layer1_out[60] = ~(layer0_out[5267] | layer0_out[5268]);
    assign layer1_out[61] = layer0_out[2893] | layer0_out[2894];
    assign layer1_out[62] = ~layer0_out[3535] | layer0_out[3534];
    assign layer1_out[63] = ~layer0_out[2321] | layer0_out[2322];
    assign layer1_out[64] = 1'b0;
    assign layer1_out[65] = ~(layer0_out[7242] & layer0_out[7243]);
    assign layer1_out[66] = layer0_out[5780];
    assign layer1_out[67] = ~(layer0_out[736] ^ layer0_out[737]);
    assign layer1_out[68] = layer0_out[4576];
    assign layer1_out[69] = layer0_out[1978];
    assign layer1_out[70] = ~(layer0_out[4150] | layer0_out[4151]);
    assign layer1_out[71] = layer0_out[5396];
    assign layer1_out[72] = layer0_out[6427] & ~layer0_out[6426];
    assign layer1_out[73] = ~(layer0_out[5138] | layer0_out[5139]);
    assign layer1_out[74] = layer0_out[3675];
    assign layer1_out[75] = layer0_out[1206] | layer0_out[1207];
    assign layer1_out[76] = ~layer0_out[2450] | layer0_out[2451];
    assign layer1_out[77] = layer0_out[4850];
    assign layer1_out[78] = ~layer0_out[7683];
    assign layer1_out[79] = layer0_out[4128];
    assign layer1_out[80] = 1'b1;
    assign layer1_out[81] = layer0_out[393] ^ layer0_out[394];
    assign layer1_out[82] = ~(layer0_out[1782] & layer0_out[1783]);
    assign layer1_out[83] = ~layer0_out[3205] | layer0_out[3206];
    assign layer1_out[84] = layer0_out[1887] | layer0_out[1888];
    assign layer1_out[85] = ~layer0_out[2170] | layer0_out[2171];
    assign layer1_out[86] = layer0_out[2754] | layer0_out[2755];
    assign layer1_out[87] = layer0_out[7971];
    assign layer1_out[88] = layer0_out[4873] & ~layer0_out[4872];
    assign layer1_out[89] = layer0_out[4310];
    assign layer1_out[90] = layer0_out[5710] & ~layer0_out[5711];
    assign layer1_out[91] = ~(layer0_out[561] ^ layer0_out[562]);
    assign layer1_out[92] = ~layer0_out[6280];
    assign layer1_out[93] = layer0_out[4428];
    assign layer1_out[94] = ~layer0_out[2754];
    assign layer1_out[95] = layer0_out[5424] & ~layer0_out[5425];
    assign layer1_out[96] = ~(layer0_out[2177] ^ layer0_out[2178]);
    assign layer1_out[97] = ~(layer0_out[2185] | layer0_out[2186]);
    assign layer1_out[98] = layer0_out[265];
    assign layer1_out[99] = layer0_out[7576] & layer0_out[7577];
    assign layer1_out[100] = 1'b1;
    assign layer1_out[101] = layer0_out[3620];
    assign layer1_out[102] = layer0_out[6599] | layer0_out[6600];
    assign layer1_out[103] = ~layer0_out[1283];
    assign layer1_out[104] = layer0_out[3033];
    assign layer1_out[105] = ~(layer0_out[2133] | layer0_out[2134]);
    assign layer1_out[106] = layer0_out[6504];
    assign layer1_out[107] = layer0_out[6234] & ~layer0_out[6235];
    assign layer1_out[108] = layer0_out[3652];
    assign layer1_out[109] = ~layer0_out[7843] | layer0_out[7844];
    assign layer1_out[110] = ~(layer0_out[3424] & layer0_out[3425]);
    assign layer1_out[111] = layer0_out[4232] ^ layer0_out[4233];
    assign layer1_out[112] = 1'b0;
    assign layer1_out[113] = layer0_out[7972] & ~layer0_out[7971];
    assign layer1_out[114] = layer0_out[763];
    assign layer1_out[115] = 1'b1;
    assign layer1_out[116] = 1'b0;
    assign layer1_out[117] = ~layer0_out[6735] | layer0_out[6736];
    assign layer1_out[118] = ~layer0_out[865] | layer0_out[866];
    assign layer1_out[119] = layer0_out[7473] & ~layer0_out[7474];
    assign layer1_out[120] = layer0_out[6662];
    assign layer1_out[121] = ~layer0_out[3243];
    assign layer1_out[122] = 1'b1;
    assign layer1_out[123] = layer0_out[7756] & ~layer0_out[7757];
    assign layer1_out[124] = ~(layer0_out[6628] | layer0_out[6629]);
    assign layer1_out[125] = ~layer0_out[1436] | layer0_out[1437];
    assign layer1_out[126] = layer0_out[7029] ^ layer0_out[7030];
    assign layer1_out[127] = ~(layer0_out[7833] ^ layer0_out[7834]);
    assign layer1_out[128] = layer0_out[7682];
    assign layer1_out[129] = layer0_out[2198] & ~layer0_out[2199];
    assign layer1_out[130] = layer0_out[6124] & layer0_out[6125];
    assign layer1_out[131] = layer0_out[127] | layer0_out[128];
    assign layer1_out[132] = 1'b0;
    assign layer1_out[133] = ~layer0_out[1618] | layer0_out[1619];
    assign layer1_out[134] = ~(layer0_out[4059] | layer0_out[4060]);
    assign layer1_out[135] = layer0_out[7436];
    assign layer1_out[136] = layer0_out[7544];
    assign layer1_out[137] = layer0_out[7375] & layer0_out[7376];
    assign layer1_out[138] = 1'b1;
    assign layer1_out[139] = layer0_out[701];
    assign layer1_out[140] = ~(layer0_out[644] & layer0_out[645]);
    assign layer1_out[141] = layer0_out[2601] & ~layer0_out[2602];
    assign layer1_out[142] = 1'b0;
    assign layer1_out[143] = layer0_out[1105] & layer0_out[1106];
    assign layer1_out[144] = ~layer0_out[1132];
    assign layer1_out[145] = layer0_out[2064] & layer0_out[2065];
    assign layer1_out[146] = ~layer0_out[7016] | layer0_out[7015];
    assign layer1_out[147] = ~(layer0_out[6725] ^ layer0_out[6726]);
    assign layer1_out[148] = ~(layer0_out[6129] & layer0_out[6130]);
    assign layer1_out[149] = layer0_out[604] | layer0_out[605];
    assign layer1_out[150] = ~layer0_out[481] | layer0_out[480];
    assign layer1_out[151] = 1'b0;
    assign layer1_out[152] = layer0_out[2377];
    assign layer1_out[153] = ~layer0_out[3526] | layer0_out[3527];
    assign layer1_out[154] = layer0_out[6638] & layer0_out[6639];
    assign layer1_out[155] = layer0_out[517] & ~layer0_out[518];
    assign layer1_out[156] = ~layer0_out[758] | layer0_out[757];
    assign layer1_out[157] = ~(layer0_out[4977] & layer0_out[4978]);
    assign layer1_out[158] = ~(layer0_out[1327] & layer0_out[1328]);
    assign layer1_out[159] = layer0_out[3550];
    assign layer1_out[160] = 1'b1;
    assign layer1_out[161] = ~layer0_out[3726] | layer0_out[3727];
    assign layer1_out[162] = layer0_out[4245] & ~layer0_out[4244];
    assign layer1_out[163] = layer0_out[7291];
    assign layer1_out[164] = layer0_out[3094] & ~layer0_out[3095];
    assign layer1_out[165] = layer0_out[2968];
    assign layer1_out[166] = ~layer0_out[3558];
    assign layer1_out[167] = ~layer0_out[1539] | layer0_out[1538];
    assign layer1_out[168] = ~layer0_out[4030] | layer0_out[4031];
    assign layer1_out[169] = layer0_out[5961];
    assign layer1_out[170] = layer0_out[638] & ~layer0_out[637];
    assign layer1_out[171] = ~layer0_out[3951] | layer0_out[3950];
    assign layer1_out[172] = layer0_out[426];
    assign layer1_out[173] = ~layer0_out[2442];
    assign layer1_out[174] = layer0_out[6516] & ~layer0_out[6515];
    assign layer1_out[175] = ~layer0_out[5752];
    assign layer1_out[176] = layer0_out[4782] | layer0_out[4783];
    assign layer1_out[177] = 1'b0;
    assign layer1_out[178] = layer0_out[5355];
    assign layer1_out[179] = layer0_out[3336];
    assign layer1_out[180] = layer0_out[879];
    assign layer1_out[181] = layer0_out[3862];
    assign layer1_out[182] = ~layer0_out[379] | layer0_out[378];
    assign layer1_out[183] = layer0_out[1565] & layer0_out[1566];
    assign layer1_out[184] = layer0_out[7918];
    assign layer1_out[185] = ~layer0_out[5083];
    assign layer1_out[186] = ~layer0_out[1162];
    assign layer1_out[187] = ~(layer0_out[4758] | layer0_out[4759]);
    assign layer1_out[188] = ~(layer0_out[2918] ^ layer0_out[2919]);
    assign layer1_out[189] = 1'b1;
    assign layer1_out[190] = ~(layer0_out[6386] & layer0_out[6387]);
    assign layer1_out[191] = ~layer0_out[7045];
    assign layer1_out[192] = ~layer0_out[6640];
    assign layer1_out[193] = layer0_out[4943] & layer0_out[4944];
    assign layer1_out[194] = layer0_out[6210] & ~layer0_out[6211];
    assign layer1_out[195] = ~layer0_out[1421];
    assign layer1_out[196] = ~(layer0_out[7067] & layer0_out[7068]);
    assign layer1_out[197] = layer0_out[1754];
    assign layer1_out[198] = ~(layer0_out[5241] | layer0_out[5242]);
    assign layer1_out[199] = ~(layer0_out[5353] | layer0_out[5354]);
    assign layer1_out[200] = ~(layer0_out[4685] & layer0_out[4686]);
    assign layer1_out[201] = ~layer0_out[2009] | layer0_out[2010];
    assign layer1_out[202] = ~layer0_out[3017];
    assign layer1_out[203] = layer0_out[5417] ^ layer0_out[5418];
    assign layer1_out[204] = ~layer0_out[660];
    assign layer1_out[205] = ~layer0_out[5693] | layer0_out[5692];
    assign layer1_out[206] = layer0_out[3980] & ~layer0_out[3981];
    assign layer1_out[207] = 1'b1;
    assign layer1_out[208] = 1'b1;
    assign layer1_out[209] = ~layer0_out[2357] | layer0_out[2358];
    assign layer1_out[210] = ~(layer0_out[4955] ^ layer0_out[4956]);
    assign layer1_out[211] = layer0_out[3706] & ~layer0_out[3705];
    assign layer1_out[212] = layer0_out[7880];
    assign layer1_out[213] = layer0_out[1591];
    assign layer1_out[214] = ~layer0_out[2779];
    assign layer1_out[215] = layer0_out[5677];
    assign layer1_out[216] = ~layer0_out[1428] | layer0_out[1427];
    assign layer1_out[217] = layer0_out[4895] | layer0_out[4896];
    assign layer1_out[218] = layer0_out[3743];
    assign layer1_out[219] = ~layer0_out[2106] | layer0_out[2107];
    assign layer1_out[220] = layer0_out[1250] | layer0_out[1251];
    assign layer1_out[221] = layer0_out[1443] | layer0_out[1444];
    assign layer1_out[222] = ~layer0_out[1804] | layer0_out[1803];
    assign layer1_out[223] = layer0_out[3322];
    assign layer1_out[224] = ~(layer0_out[4429] & layer0_out[4430]);
    assign layer1_out[225] = layer0_out[7679] ^ layer0_out[7680];
    assign layer1_out[226] = layer0_out[1801] ^ layer0_out[1802];
    assign layer1_out[227] = layer0_out[1585] & ~layer0_out[1584];
    assign layer1_out[228] = layer0_out[7289] | layer0_out[7290];
    assign layer1_out[229] = layer0_out[3608] & ~layer0_out[3609];
    assign layer1_out[230] = ~layer0_out[3793];
    assign layer1_out[231] = ~layer0_out[3995] | layer0_out[3994];
    assign layer1_out[232] = layer0_out[46];
    assign layer1_out[233] = 1'b0;
    assign layer1_out[234] = ~(layer0_out[7135] | layer0_out[7136]);
    assign layer1_out[235] = ~layer0_out[4229];
    assign layer1_out[236] = 1'b1;
    assign layer1_out[237] = 1'b1;
    assign layer1_out[238] = layer0_out[2706] ^ layer0_out[2707];
    assign layer1_out[239] = layer0_out[4923];
    assign layer1_out[240] = ~layer0_out[6963];
    assign layer1_out[241] = ~(layer0_out[4643] & layer0_out[4644]);
    assign layer1_out[242] = ~(layer0_out[455] | layer0_out[456]);
    assign layer1_out[243] = ~layer0_out[5819] | layer0_out[5820];
    assign layer1_out[244] = ~(layer0_out[2696] & layer0_out[2697]);
    assign layer1_out[245] = ~(layer0_out[1422] | layer0_out[1423]);
    assign layer1_out[246] = layer0_out[632];
    assign layer1_out[247] = layer0_out[4031] | layer0_out[4032];
    assign layer1_out[248] = ~(layer0_out[2020] & layer0_out[2021]);
    assign layer1_out[249] = ~layer0_out[983];
    assign layer1_out[250] = ~(layer0_out[4174] ^ layer0_out[4175]);
    assign layer1_out[251] = layer0_out[3281] | layer0_out[3282];
    assign layer1_out[252] = 1'b1;
    assign layer1_out[253] = ~(layer0_out[6565] ^ layer0_out[6566]);
    assign layer1_out[254] = layer0_out[3885];
    assign layer1_out[255] = ~(layer0_out[7030] & layer0_out[7031]);
    assign layer1_out[256] = layer0_out[5256] & ~layer0_out[5255];
    assign layer1_out[257] = 1'b0;
    assign layer1_out[258] = ~layer0_out[6567];
    assign layer1_out[259] = ~(layer0_out[4879] | layer0_out[4880]);
    assign layer1_out[260] = ~(layer0_out[4589] & layer0_out[4590]);
    assign layer1_out[261] = ~(layer0_out[2930] | layer0_out[2931]);
    assign layer1_out[262] = layer0_out[5135];
    assign layer1_out[263] = ~layer0_out[311];
    assign layer1_out[264] = layer0_out[7534] & ~layer0_out[7535];
    assign layer1_out[265] = ~layer0_out[828];
    assign layer1_out[266] = ~(layer0_out[297] & layer0_out[298]);
    assign layer1_out[267] = layer0_out[4424];
    assign layer1_out[268] = ~layer0_out[2255];
    assign layer1_out[269] = ~layer0_out[3743] | layer0_out[3744];
    assign layer1_out[270] = ~layer0_out[5771] | layer0_out[5772];
    assign layer1_out[271] = 1'b0;
    assign layer1_out[272] = layer0_out[981] & ~layer0_out[980];
    assign layer1_out[273] = layer0_out[4387] | layer0_out[4388];
    assign layer1_out[274] = layer0_out[2224];
    assign layer1_out[275] = layer0_out[4450] & layer0_out[4451];
    assign layer1_out[276] = layer0_out[2519] & ~layer0_out[2518];
    assign layer1_out[277] = layer0_out[7957];
    assign layer1_out[278] = ~layer0_out[50];
    assign layer1_out[279] = layer0_out[361] & ~layer0_out[362];
    assign layer1_out[280] = layer0_out[7186] & layer0_out[7187];
    assign layer1_out[281] = ~layer0_out[878] | layer0_out[877];
    assign layer1_out[282] = ~layer0_out[4888];
    assign layer1_out[283] = ~(layer0_out[2052] ^ layer0_out[2053]);
    assign layer1_out[284] = layer0_out[152] | layer0_out[153];
    assign layer1_out[285] = layer0_out[4307] & ~layer0_out[4308];
    assign layer1_out[286] = ~(layer0_out[7738] | layer0_out[7739]);
    assign layer1_out[287] = ~layer0_out[6176] | layer0_out[6175];
    assign layer1_out[288] = layer0_out[3594] & ~layer0_out[3595];
    assign layer1_out[289] = ~layer0_out[1326] | layer0_out[1325];
    assign layer1_out[290] = ~layer0_out[2840];
    assign layer1_out[291] = layer0_out[6953] & ~layer0_out[6954];
    assign layer1_out[292] = ~layer0_out[1892] | layer0_out[1893];
    assign layer1_out[293] = ~(layer0_out[707] | layer0_out[708]);
    assign layer1_out[294] = ~(layer0_out[1996] | layer0_out[1997]);
    assign layer1_out[295] = ~(layer0_out[2630] | layer0_out[2631]);
    assign layer1_out[296] = 1'b0;
    assign layer1_out[297] = layer0_out[6335] ^ layer0_out[6336];
    assign layer1_out[298] = 1'b0;
    assign layer1_out[299] = layer0_out[4043] & ~layer0_out[4044];
    assign layer1_out[300] = layer0_out[1908] & ~layer0_out[1909];
    assign layer1_out[301] = ~layer0_out[5833];
    assign layer1_out[302] = layer0_out[7175];
    assign layer1_out[303] = layer0_out[7395] & ~layer0_out[7394];
    assign layer1_out[304] = layer0_out[4551] ^ layer0_out[4552];
    assign layer1_out[305] = ~layer0_out[1502];
    assign layer1_out[306] = ~(layer0_out[1409] | layer0_out[1410]);
    assign layer1_out[307] = ~layer0_out[2139];
    assign layer1_out[308] = layer0_out[3301] & ~layer0_out[3302];
    assign layer1_out[309] = layer0_out[3814] & ~layer0_out[3813];
    assign layer1_out[310] = ~(layer0_out[2574] & layer0_out[2575]);
    assign layer1_out[311] = layer0_out[2474];
    assign layer1_out[312] = layer0_out[418] | layer0_out[419];
    assign layer1_out[313] = ~(layer0_out[6715] | layer0_out[6716]);
    assign layer1_out[314] = layer0_out[5947];
    assign layer1_out[315] = ~layer0_out[1556];
    assign layer1_out[316] = ~layer0_out[1922] | layer0_out[1923];
    assign layer1_out[317] = layer0_out[4670];
    assign layer1_out[318] = layer0_out[2271] & layer0_out[2272];
    assign layer1_out[319] = layer0_out[7223];
    assign layer1_out[320] = layer0_out[2365];
    assign layer1_out[321] = 1'b0;
    assign layer1_out[322] = layer0_out[4219] | layer0_out[4220];
    assign layer1_out[323] = layer0_out[6066] & ~layer0_out[6065];
    assign layer1_out[324] = layer0_out[7295];
    assign layer1_out[325] = layer0_out[1220] & ~layer0_out[1219];
    assign layer1_out[326] = ~layer0_out[6059];
    assign layer1_out[327] = ~layer0_out[5043];
    assign layer1_out[328] = ~layer0_out[4367];
    assign layer1_out[329] = ~layer0_out[5181] | layer0_out[5180];
    assign layer1_out[330] = layer0_out[4560] & ~layer0_out[4559];
    assign layer1_out[331] = layer0_out[2557];
    assign layer1_out[332] = ~layer0_out[146];
    assign layer1_out[333] = 1'b0;
    assign layer1_out[334] = layer0_out[6898] & layer0_out[6899];
    assign layer1_out[335] = layer0_out[5260];
    assign layer1_out[336] = 1'b1;
    assign layer1_out[337] = layer0_out[6542] & layer0_out[6543];
    assign layer1_out[338] = ~layer0_out[3431];
    assign layer1_out[339] = ~(layer0_out[7820] | layer0_out[7821]);
    assign layer1_out[340] = ~layer0_out[6682] | layer0_out[6683];
    assign layer1_out[341] = ~(layer0_out[5925] | layer0_out[5926]);
    assign layer1_out[342] = 1'b1;
    assign layer1_out[343] = layer0_out[1604] | layer0_out[1605];
    assign layer1_out[344] = ~layer0_out[5951];
    assign layer1_out[345] = layer0_out[5364] & ~layer0_out[5363];
    assign layer1_out[346] = layer0_out[6519] & layer0_out[6520];
    assign layer1_out[347] = layer0_out[5812] & ~layer0_out[5811];
    assign layer1_out[348] = ~(layer0_out[4691] & layer0_out[4692]);
    assign layer1_out[349] = layer0_out[2972] & ~layer0_out[2973];
    assign layer1_out[350] = ~layer0_out[6122] | layer0_out[6121];
    assign layer1_out[351] = ~layer0_out[2568] | layer0_out[2567];
    assign layer1_out[352] = ~layer0_out[3660];
    assign layer1_out[353] = layer0_out[493];
    assign layer1_out[354] = 1'b0;
    assign layer1_out[355] = layer0_out[2645] & ~layer0_out[2646];
    assign layer1_out[356] = ~(layer0_out[5698] | layer0_out[5699]);
    assign layer1_out[357] = layer0_out[4738] & ~layer0_out[4737];
    assign layer1_out[358] = ~layer0_out[732];
    assign layer1_out[359] = ~(layer0_out[1735] ^ layer0_out[1736]);
    assign layer1_out[360] = layer0_out[338];
    assign layer1_out[361] = ~layer0_out[7628] | layer0_out[7627];
    assign layer1_out[362] = 1'b1;
    assign layer1_out[363] = ~layer0_out[4786] | layer0_out[4785];
    assign layer1_out[364] = layer0_out[6874];
    assign layer1_out[365] = ~layer0_out[5552];
    assign layer1_out[366] = layer0_out[5906] | layer0_out[5907];
    assign layer1_out[367] = ~layer0_out[4201] | layer0_out[4200];
    assign layer1_out[368] = layer0_out[7758] & ~layer0_out[7757];
    assign layer1_out[369] = layer0_out[5581] & layer0_out[5582];
    assign layer1_out[370] = layer0_out[2396] | layer0_out[2397];
    assign layer1_out[371] = 1'b0;
    assign layer1_out[372] = layer0_out[4213] | layer0_out[4214];
    assign layer1_out[373] = ~layer0_out[6966];
    assign layer1_out[374] = layer0_out[3437];
    assign layer1_out[375] = layer0_out[2029] & ~layer0_out[2030];
    assign layer1_out[376] = 1'b1;
    assign layer1_out[377] = ~layer0_out[1297];
    assign layer1_out[378] = layer0_out[3249] | layer0_out[3250];
    assign layer1_out[379] = ~(layer0_out[1004] | layer0_out[1005]);
    assign layer1_out[380] = layer0_out[7727];
    assign layer1_out[381] = layer0_out[432] & layer0_out[433];
    assign layer1_out[382] = ~layer0_out[735] | layer0_out[734];
    assign layer1_out[383] = layer0_out[1299];
    assign layer1_out[384] = ~layer0_out[5392];
    assign layer1_out[385] = layer0_out[5466] | layer0_out[5467];
    assign layer1_out[386] = ~layer0_out[5044];
    assign layer1_out[387] = layer0_out[3599];
    assign layer1_out[388] = layer0_out[5059] & layer0_out[5060];
    assign layer1_out[389] = layer0_out[1838];
    assign layer1_out[390] = ~layer0_out[533];
    assign layer1_out[391] = layer0_out[6113];
    assign layer1_out[392] = layer0_out[1666];
    assign layer1_out[393] = ~layer0_out[5015];
    assign layer1_out[394] = ~layer0_out[5107] | layer0_out[5108];
    assign layer1_out[395] = ~layer0_out[1382];
    assign layer1_out[396] = layer0_out[7812];
    assign layer1_out[397] = ~(layer0_out[7082] & layer0_out[7083]);
    assign layer1_out[398] = ~(layer0_out[5215] ^ layer0_out[5216]);
    assign layer1_out[399] = layer0_out[3790] & layer0_out[3791];
    assign layer1_out[400] = layer0_out[1689] | layer0_out[1690];
    assign layer1_out[401] = ~layer0_out[7464] | layer0_out[7463];
    assign layer1_out[402] = layer0_out[6878];
    assign layer1_out[403] = ~layer0_out[923] | layer0_out[922];
    assign layer1_out[404] = ~(layer0_out[4845] ^ layer0_out[4846]);
    assign layer1_out[405] = layer0_out[7306] & ~layer0_out[7307];
    assign layer1_out[406] = layer0_out[5639] & ~layer0_out[5638];
    assign layer1_out[407] = ~layer0_out[95] | layer0_out[94];
    assign layer1_out[408] = layer0_out[7440];
    assign layer1_out[409] = layer0_out[4792];
    assign layer1_out[410] = ~(layer0_out[7467] | layer0_out[7468]);
    assign layer1_out[411] = ~layer0_out[847];
    assign layer1_out[412] = layer0_out[3014] & ~layer0_out[3015];
    assign layer1_out[413] = ~layer0_out[3457] | layer0_out[3458];
    assign layer1_out[414] = layer0_out[583] & layer0_out[584];
    assign layer1_out[415] = ~layer0_out[4232];
    assign layer1_out[416] = ~(layer0_out[6512] & layer0_out[6513]);
    assign layer1_out[417] = ~layer0_out[7364];
    assign layer1_out[418] = ~layer0_out[5380] | layer0_out[5379];
    assign layer1_out[419] = layer0_out[639] & ~layer0_out[640];
    assign layer1_out[420] = layer0_out[551] & ~layer0_out[552];
    assign layer1_out[421] = layer0_out[1762] & ~layer0_out[1761];
    assign layer1_out[422] = layer0_out[4249];
    assign layer1_out[423] = layer0_out[2105] & ~layer0_out[2104];
    assign layer1_out[424] = layer0_out[7466] & ~layer0_out[7465];
    assign layer1_out[425] = ~(layer0_out[4889] & layer0_out[4890]);
    assign layer1_out[426] = layer0_out[2166];
    assign layer1_out[427] = layer0_out[3602] ^ layer0_out[3603];
    assign layer1_out[428] = ~(layer0_out[3898] ^ layer0_out[3899]);
    assign layer1_out[429] = ~layer0_out[911] | layer0_out[910];
    assign layer1_out[430] = layer0_out[7000];
    assign layer1_out[431] = ~(layer0_out[2818] & layer0_out[2819]);
    assign layer1_out[432] = layer0_out[2908];
    assign layer1_out[433] = ~(layer0_out[208] | layer0_out[209]);
    assign layer1_out[434] = layer0_out[6893] ^ layer0_out[6894];
    assign layer1_out[435] = ~layer0_out[634] | layer0_out[633];
    assign layer1_out[436] = layer0_out[2468] & layer0_out[2469];
    assign layer1_out[437] = ~layer0_out[1105];
    assign layer1_out[438] = ~layer0_out[2241];
    assign layer1_out[439] = ~(layer0_out[1804] & layer0_out[1805]);
    assign layer1_out[440] = ~layer0_out[1355] | layer0_out[1354];
    assign layer1_out[441] = ~layer0_out[2961] | layer0_out[2960];
    assign layer1_out[442] = ~layer0_out[2520] | layer0_out[2521];
    assign layer1_out[443] = layer0_out[3162] & layer0_out[3163];
    assign layer1_out[444] = layer0_out[1790];
    assign layer1_out[445] = ~layer0_out[2639] | layer0_out[2638];
    assign layer1_out[446] = layer0_out[3899];
    assign layer1_out[447] = layer0_out[461];
    assign layer1_out[448] = layer0_out[1745] & ~layer0_out[1746];
    assign layer1_out[449] = ~layer0_out[2245] | layer0_out[2246];
    assign layer1_out[450] = layer0_out[7351];
    assign layer1_out[451] = ~(layer0_out[6463] ^ layer0_out[6464]);
    assign layer1_out[452] = ~layer0_out[6044];
    assign layer1_out[453] = layer0_out[5063];
    assign layer1_out[454] = layer0_out[7444] ^ layer0_out[7445];
    assign layer1_out[455] = ~layer0_out[6748] | layer0_out[6747];
    assign layer1_out[456] = layer0_out[642];
    assign layer1_out[457] = ~(layer0_out[2815] | layer0_out[2816]);
    assign layer1_out[458] = 1'b1;
    assign layer1_out[459] = layer0_out[3320];
    assign layer1_out[460] = layer0_out[1793] & ~layer0_out[1794];
    assign layer1_out[461] = layer0_out[3577] ^ layer0_out[3578];
    assign layer1_out[462] = layer0_out[645] | layer0_out[646];
    assign layer1_out[463] = ~layer0_out[3389];
    assign layer1_out[464] = ~layer0_out[6187] | layer0_out[6188];
    assign layer1_out[465] = layer0_out[989];
    assign layer1_out[466] = ~(layer0_out[6546] | layer0_out[6547]);
    assign layer1_out[467] = ~layer0_out[7229];
    assign layer1_out[468] = layer0_out[6802] & ~layer0_out[6803];
    assign layer1_out[469] = ~layer0_out[5898];
    assign layer1_out[470] = ~(layer0_out[3976] ^ layer0_out[3977]);
    assign layer1_out[471] = layer0_out[5736] | layer0_out[5737];
    assign layer1_out[472] = ~layer0_out[2995];
    assign layer1_out[473] = layer0_out[4196];
    assign layer1_out[474] = layer0_out[7141];
    assign layer1_out[475] = ~layer0_out[6267] | layer0_out[6268];
    assign layer1_out[476] = layer0_out[2731];
    assign layer1_out[477] = ~(layer0_out[6647] & layer0_out[6648]);
    assign layer1_out[478] = ~layer0_out[7110];
    assign layer1_out[479] = ~layer0_out[2008] | layer0_out[2007];
    assign layer1_out[480] = layer0_out[7212] & layer0_out[7213];
    assign layer1_out[481] = ~layer0_out[6938];
    assign layer1_out[482] = ~layer0_out[7010];
    assign layer1_out[483] = ~(layer0_out[2378] ^ layer0_out[2379]);
    assign layer1_out[484] = ~layer0_out[6127];
    assign layer1_out[485] = layer0_out[649];
    assign layer1_out[486] = ~layer0_out[2228];
    assign layer1_out[487] = ~(layer0_out[1200] & layer0_out[1201]);
    assign layer1_out[488] = layer0_out[4917] & ~layer0_out[4916];
    assign layer1_out[489] = layer0_out[4703];
    assign layer1_out[490] = ~layer0_out[6];
    assign layer1_out[491] = ~layer0_out[5784];
    assign layer1_out[492] = layer0_out[6529];
    assign layer1_out[493] = layer0_out[2101] & layer0_out[2102];
    assign layer1_out[494] = ~(layer0_out[5346] ^ layer0_out[5347]);
    assign layer1_out[495] = layer0_out[5582] & ~layer0_out[5583];
    assign layer1_out[496] = layer0_out[6433] | layer0_out[6434];
    assign layer1_out[497] = layer0_out[1943] & ~layer0_out[1944];
    assign layer1_out[498] = ~layer0_out[1971] | layer0_out[1970];
    assign layer1_out[499] = layer0_out[2211] & ~layer0_out[2212];
    assign layer1_out[500] = ~layer0_out[5757] | layer0_out[5758];
    assign layer1_out[501] = 1'b1;
    assign layer1_out[502] = ~(layer0_out[5030] | layer0_out[5031]);
    assign layer1_out[503] = layer0_out[867] & ~layer0_out[866];
    assign layer1_out[504] = layer0_out[2204];
    assign layer1_out[505] = ~layer0_out[2190] | layer0_out[2189];
    assign layer1_out[506] = ~layer0_out[3655];
    assign layer1_out[507] = ~layer0_out[2413] | layer0_out[2412];
    assign layer1_out[508] = layer0_out[6445] ^ layer0_out[6446];
    assign layer1_out[509] = ~layer0_out[774];
    assign layer1_out[510] = layer0_out[6141];
    assign layer1_out[511] = ~(layer0_out[2174] ^ layer0_out[2175]);
    assign layer1_out[512] = layer0_out[6004] & ~layer0_out[6003];
    assign layer1_out[513] = layer0_out[3291] & ~layer0_out[3292];
    assign layer1_out[514] = layer0_out[2244] & ~layer0_out[2245];
    assign layer1_out[515] = layer0_out[3819] & ~layer0_out[3820];
    assign layer1_out[516] = layer0_out[5530];
    assign layer1_out[517] = layer0_out[1433] | layer0_out[1434];
    assign layer1_out[518] = layer0_out[233] & ~layer0_out[232];
    assign layer1_out[519] = layer0_out[712] & layer0_out[713];
    assign layer1_out[520] = layer0_out[1878] | layer0_out[1879];
    assign layer1_out[521] = layer0_out[234];
    assign layer1_out[522] = layer0_out[4632] & ~layer0_out[4633];
    assign layer1_out[523] = layer0_out[2129];
    assign layer1_out[524] = 1'b0;
    assign layer1_out[525] = ~(layer0_out[5229] ^ layer0_out[5230]);
    assign layer1_out[526] = ~layer0_out[3254];
    assign layer1_out[527] = ~layer0_out[6666] | layer0_out[6667];
    assign layer1_out[528] = layer0_out[1875] & ~layer0_out[1874];
    assign layer1_out[529] = ~(layer0_out[3331] ^ layer0_out[3332]);
    assign layer1_out[530] = ~(layer0_out[3642] | layer0_out[3643]);
    assign layer1_out[531] = ~layer0_out[6023];
    assign layer1_out[532] = ~(layer0_out[2048] | layer0_out[2049]);
    assign layer1_out[533] = ~layer0_out[4117];
    assign layer1_out[534] = ~(layer0_out[4408] ^ layer0_out[4409]);
    assign layer1_out[535] = ~layer0_out[4210];
    assign layer1_out[536] = ~layer0_out[7508] | layer0_out[7507];
    assign layer1_out[537] = layer0_out[871];
    assign layer1_out[538] = layer0_out[2] | layer0_out[3];
    assign layer1_out[539] = ~layer0_out[6890];
    assign layer1_out[540] = ~layer0_out[5069] | layer0_out[5068];
    assign layer1_out[541] = layer0_out[7336];
    assign layer1_out[542] = layer0_out[3213] | layer0_out[3214];
    assign layer1_out[543] = ~layer0_out[2884];
    assign layer1_out[544] = ~(layer0_out[4530] | layer0_out[4531]);
    assign layer1_out[545] = ~(layer0_out[4396] & layer0_out[4397]);
    assign layer1_out[546] = layer0_out[6709] & ~layer0_out[6708];
    assign layer1_out[547] = 1'b0;
    assign layer1_out[548] = 1'b1;
    assign layer1_out[549] = layer0_out[5154];
    assign layer1_out[550] = layer0_out[2790] | layer0_out[2791];
    assign layer1_out[551] = layer0_out[2066];
    assign layer1_out[552] = 1'b0;
    assign layer1_out[553] = ~(layer0_out[6904] & layer0_out[6905]);
    assign layer1_out[554] = layer0_out[3647];
    assign layer1_out[555] = layer0_out[2846] | layer0_out[2847];
    assign layer1_out[556] = ~layer0_out[593];
    assign layer1_out[557] = ~(layer0_out[2963] | layer0_out[2964]);
    assign layer1_out[558] = 1'b1;
    assign layer1_out[559] = ~layer0_out[3642];
    assign layer1_out[560] = layer0_out[5472] ^ layer0_out[5473];
    assign layer1_out[561] = ~layer0_out[5625];
    assign layer1_out[562] = ~layer0_out[3711] | layer0_out[3712];
    assign layer1_out[563] = ~layer0_out[2334];
    assign layer1_out[564] = layer0_out[7697];
    assign layer1_out[565] = layer0_out[2431];
    assign layer1_out[566] = layer0_out[2224];
    assign layer1_out[567] = layer0_out[1694] & ~layer0_out[1695];
    assign layer1_out[568] = ~layer0_out[3494] | layer0_out[3493];
    assign layer1_out[569] = layer0_out[7263];
    assign layer1_out[570] = layer0_out[5007];
    assign layer1_out[571] = layer0_out[6980] & layer0_out[6981];
    assign layer1_out[572] = 1'b1;
    assign layer1_out[573] = ~layer0_out[6928];
    assign layer1_out[574] = layer0_out[6787] & layer0_out[6788];
    assign layer1_out[575] = ~(layer0_out[7488] & layer0_out[7489]);
    assign layer1_out[576] = ~(layer0_out[431] & layer0_out[432]);
    assign layer1_out[577] = layer0_out[4069];
    assign layer1_out[578] = ~layer0_out[3235] | layer0_out[3234];
    assign layer1_out[579] = layer0_out[3822] & ~layer0_out[3821];
    assign layer1_out[580] = 1'b0;
    assign layer1_out[581] = ~(layer0_out[622] | layer0_out[623]);
    assign layer1_out[582] = ~layer0_out[4119];
    assign layer1_out[583] = layer0_out[253] & ~layer0_out[252];
    assign layer1_out[584] = layer0_out[6888];
    assign layer1_out[585] = layer0_out[7349] & ~layer0_out[7350];
    assign layer1_out[586] = ~layer0_out[2823] | layer0_out[2824];
    assign layer1_out[587] = ~(layer0_out[5509] & layer0_out[5510]);
    assign layer1_out[588] = ~layer0_out[6965];
    assign layer1_out[589] = layer0_out[3938] & ~layer0_out[3937];
    assign layer1_out[590] = ~layer0_out[1188];
    assign layer1_out[591] = layer0_out[3831] & layer0_out[3832];
    assign layer1_out[592] = layer0_out[6358];
    assign layer1_out[593] = ~(layer0_out[6244] ^ layer0_out[6245]);
    assign layer1_out[594] = layer0_out[4235] & layer0_out[4236];
    assign layer1_out[595] = ~(layer0_out[7677] ^ layer0_out[7678]);
    assign layer1_out[596] = layer0_out[7217] | layer0_out[7218];
    assign layer1_out[597] = layer0_out[6877];
    assign layer1_out[598] = layer0_out[1229] | layer0_out[1230];
    assign layer1_out[599] = ~(layer0_out[4203] | layer0_out[4204]);
    assign layer1_out[600] = ~layer0_out[4377] | layer0_out[4376];
    assign layer1_out[601] = 1'b1;
    assign layer1_out[602] = layer0_out[3680];
    assign layer1_out[603] = ~layer0_out[1307];
    assign layer1_out[604] = layer0_out[7207] | layer0_out[7208];
    assign layer1_out[605] = ~layer0_out[5392];
    assign layer1_out[606] = ~layer0_out[5924];
    assign layer1_out[607] = ~layer0_out[29];
    assign layer1_out[608] = ~layer0_out[4253];
    assign layer1_out[609] = ~layer0_out[3358];
    assign layer1_out[610] = ~(layer0_out[1237] ^ layer0_out[1238]);
    assign layer1_out[611] = ~(layer0_out[6143] ^ layer0_out[6144]);
    assign layer1_out[612] = ~layer0_out[1656] | layer0_out[1655];
    assign layer1_out[613] = ~(layer0_out[5994] | layer0_out[5995]);
    assign layer1_out[614] = layer0_out[5098] & ~layer0_out[5097];
    assign layer1_out[615] = ~layer0_out[5621];
    assign layer1_out[616] = layer0_out[5387];
    assign layer1_out[617] = layer0_out[7118] ^ layer0_out[7119];
    assign layer1_out[618] = layer0_out[681] & layer0_out[682];
    assign layer1_out[619] = ~(layer0_out[3113] ^ layer0_out[3114]);
    assign layer1_out[620] = ~layer0_out[5465];
    assign layer1_out[621] = ~layer0_out[5768];
    assign layer1_out[622] = ~layer0_out[3090] | layer0_out[3089];
    assign layer1_out[623] = layer0_out[5982] & ~layer0_out[5981];
    assign layer1_out[624] = 1'b1;
    assign layer1_out[625] = ~layer0_out[6777] | layer0_out[6776];
    assign layer1_out[626] = layer0_out[2213];
    assign layer1_out[627] = layer0_out[4588] | layer0_out[4589];
    assign layer1_out[628] = ~(layer0_out[7421] | layer0_out[7422]);
    assign layer1_out[629] = layer0_out[5002] & ~layer0_out[5001];
    assign layer1_out[630] = ~layer0_out[2613];
    assign layer1_out[631] = 1'b1;
    assign layer1_out[632] = ~(layer0_out[1283] | layer0_out[1284]);
    assign layer1_out[633] = ~layer0_out[3553];
    assign layer1_out[634] = layer0_out[3162];
    assign layer1_out[635] = layer0_out[7584] & layer0_out[7585];
    assign layer1_out[636] = layer0_out[2150] & ~layer0_out[2151];
    assign layer1_out[637] = ~layer0_out[6865];
    assign layer1_out[638] = layer0_out[3410];
    assign layer1_out[639] = ~(layer0_out[7600] & layer0_out[7601]);
    assign layer1_out[640] = ~(layer0_out[1386] ^ layer0_out[1387]);
    assign layer1_out[641] = layer0_out[6626];
    assign layer1_out[642] = ~layer0_out[5005] | layer0_out[5006];
    assign layer1_out[643] = 1'b1;
    assign layer1_out[644] = layer0_out[7882] & ~layer0_out[7881];
    assign layer1_out[645] = ~layer0_out[7839] | layer0_out[7840];
    assign layer1_out[646] = ~layer0_out[6294];
    assign layer1_out[647] = layer0_out[4503];
    assign layer1_out[648] = layer0_out[3632] & ~layer0_out[3631];
    assign layer1_out[649] = ~(layer0_out[3893] & layer0_out[3894]);
    assign layer1_out[650] = ~(layer0_out[1544] ^ layer0_out[1545]);
    assign layer1_out[651] = ~layer0_out[1399] | layer0_out[1400];
    assign layer1_out[652] = ~layer0_out[7145];
    assign layer1_out[653] = ~layer0_out[7584] | layer0_out[7583];
    assign layer1_out[654] = ~(layer0_out[2349] & layer0_out[2350]);
    assign layer1_out[655] = layer0_out[6798] & ~layer0_out[6799];
    assign layer1_out[656] = layer0_out[7371] & layer0_out[7372];
    assign layer1_out[657] = ~(layer0_out[7918] ^ layer0_out[7919]);
    assign layer1_out[658] = layer0_out[5258];
    assign layer1_out[659] = ~(layer0_out[1163] & layer0_out[1164]);
    assign layer1_out[660] = layer0_out[38] ^ layer0_out[39];
    assign layer1_out[661] = 1'b1;
    assign layer1_out[662] = ~layer0_out[6508];
    assign layer1_out[663] = 1'b1;
    assign layer1_out[664] = layer0_out[4284];
    assign layer1_out[665] = 1'b1;
    assign layer1_out[666] = ~layer0_out[7802];
    assign layer1_out[667] = layer0_out[4949];
    assign layer1_out[668] = layer0_out[2624] & ~layer0_out[2623];
    assign layer1_out[669] = ~layer0_out[2593] | layer0_out[2594];
    assign layer1_out[670] = layer0_out[1705];
    assign layer1_out[671] = layer0_out[2018];
    assign layer1_out[672] = layer0_out[4198];
    assign layer1_out[673] = ~layer0_out[3784] | layer0_out[3783];
    assign layer1_out[674] = layer0_out[7405] & ~layer0_out[7404];
    assign layer1_out[675] = layer0_out[498] | layer0_out[499];
    assign layer1_out[676] = 1'b1;
    assign layer1_out[677] = ~layer0_out[6272] | layer0_out[6273];
    assign layer1_out[678] = layer0_out[2621] & layer0_out[2622];
    assign layer1_out[679] = layer0_out[3042];
    assign layer1_out[680] = ~layer0_out[4907] | layer0_out[4908];
    assign layer1_out[681] = layer0_out[1830] & layer0_out[1831];
    assign layer1_out[682] = ~layer0_out[5307] | layer0_out[5306];
    assign layer1_out[683] = layer0_out[5201] & ~layer0_out[5200];
    assign layer1_out[684] = 1'b1;
    assign layer1_out[685] = 1'b1;
    assign layer1_out[686] = layer0_out[2862] & ~layer0_out[2861];
    assign layer1_out[687] = ~layer0_out[1130];
    assign layer1_out[688] = ~layer0_out[5233] | layer0_out[5232];
    assign layer1_out[689] = layer0_out[4526] | layer0_out[4527];
    assign layer1_out[690] = layer0_out[5408];
    assign layer1_out[691] = ~layer0_out[697];
    assign layer1_out[692] = ~layer0_out[2505];
    assign layer1_out[693] = layer0_out[4758] & ~layer0_out[4757];
    assign layer1_out[694] = 1'b1;
    assign layer1_out[695] = ~layer0_out[3488];
    assign layer1_out[696] = layer0_out[1377];
    assign layer1_out[697] = layer0_out[3701];
    assign layer1_out[698] = ~layer0_out[449];
    assign layer1_out[699] = ~layer0_out[6439] | layer0_out[6438];
    assign layer1_out[700] = ~layer0_out[7106] | layer0_out[7107];
    assign layer1_out[701] = ~layer0_out[510];
    assign layer1_out[702] = layer0_out[6384] & ~layer0_out[6383];
    assign layer1_out[703] = layer0_out[1705];
    assign layer1_out[704] = ~layer0_out[3970];
    assign layer1_out[705] = ~layer0_out[251];
    assign layer1_out[706] = layer0_out[3753] & ~layer0_out[3752];
    assign layer1_out[707] = layer0_out[4645] & ~layer0_out[4646];
    assign layer1_out[708] = layer0_out[5989] & ~layer0_out[5988];
    assign layer1_out[709] = layer0_out[5077];
    assign layer1_out[710] = layer0_out[2205];
    assign layer1_out[711] = ~layer0_out[1781];
    assign layer1_out[712] = ~layer0_out[3738];
    assign layer1_out[713] = layer0_out[4361] | layer0_out[4362];
    assign layer1_out[714] = layer0_out[3312];
    assign layer1_out[715] = 1'b0;
    assign layer1_out[716] = 1'b0;
    assign layer1_out[717] = ~layer0_out[802];
    assign layer1_out[718] = ~layer0_out[5954];
    assign layer1_out[719] = ~layer0_out[5308];
    assign layer1_out[720] = 1'b1;
    assign layer1_out[721] = ~(layer0_out[2391] & layer0_out[2392]);
    assign layer1_out[722] = ~(layer0_out[3967] & layer0_out[3968]);
    assign layer1_out[723] = ~(layer0_out[3876] | layer0_out[3877]);
    assign layer1_out[724] = ~layer0_out[5673] | layer0_out[5672];
    assign layer1_out[725] = layer0_out[7210] & ~layer0_out[7209];
    assign layer1_out[726] = ~layer0_out[1732];
    assign layer1_out[727] = layer0_out[3317] & ~layer0_out[3316];
    assign layer1_out[728] = ~(layer0_out[5968] & layer0_out[5969]);
    assign layer1_out[729] = ~(layer0_out[4003] ^ layer0_out[4004]);
    assign layer1_out[730] = ~(layer0_out[6027] | layer0_out[6028]);
    assign layer1_out[731] = layer0_out[6613] ^ layer0_out[6614];
    assign layer1_out[732] = layer0_out[2603] | layer0_out[2604];
    assign layer1_out[733] = layer0_out[6185] & ~layer0_out[6186];
    assign layer1_out[734] = ~layer0_out[1678];
    assign layer1_out[735] = layer0_out[2777] & ~layer0_out[2778];
    assign layer1_out[736] = ~layer0_out[1541];
    assign layer1_out[737] = ~layer0_out[5149] | layer0_out[5148];
    assign layer1_out[738] = ~layer0_out[117] | layer0_out[118];
    assign layer1_out[739] = layer0_out[7248];
    assign layer1_out[740] = layer0_out[919];
    assign layer1_out[741] = layer0_out[7540] & ~layer0_out[7541];
    assign layer1_out[742] = layer0_out[453] ^ layer0_out[454];
    assign layer1_out[743] = layer0_out[7278] & ~layer0_out[7277];
    assign layer1_out[744] = layer0_out[2610] & ~layer0_out[2611];
    assign layer1_out[745] = ~(layer0_out[2979] | layer0_out[2980]);
    assign layer1_out[746] = ~layer0_out[4015];
    assign layer1_out[747] = ~layer0_out[6087];
    assign layer1_out[748] = layer0_out[1785];
    assign layer1_out[749] = ~(layer0_out[1958] | layer0_out[1959]);
    assign layer1_out[750] = ~(layer0_out[3088] | layer0_out[3089]);
    assign layer1_out[751] = ~(layer0_out[7787] ^ layer0_out[7788]);
    assign layer1_out[752] = ~layer0_out[7401];
    assign layer1_out[753] = layer0_out[3450] & layer0_out[3451];
    assign layer1_out[754] = ~layer0_out[6033];
    assign layer1_out[755] = layer0_out[1183] | layer0_out[1184];
    assign layer1_out[756] = layer0_out[4919];
    assign layer1_out[757] = ~(layer0_out[2509] ^ layer0_out[2510]);
    assign layer1_out[758] = layer0_out[739] & layer0_out[740];
    assign layer1_out[759] = layer0_out[1401] & ~layer0_out[1402];
    assign layer1_out[760] = ~layer0_out[747] | layer0_out[748];
    assign layer1_out[761] = ~(layer0_out[1096] ^ layer0_out[1097]);
    assign layer1_out[762] = 1'b0;
    assign layer1_out[763] = layer0_out[6131] & ~layer0_out[6132];
    assign layer1_out[764] = ~layer0_out[3122];
    assign layer1_out[765] = layer0_out[4903];
    assign layer1_out[766] = ~layer0_out[556];
    assign layer1_out[767] = ~layer0_out[450] | layer0_out[451];
    assign layer1_out[768] = layer0_out[3615] & ~layer0_out[3616];
    assign layer1_out[769] = ~(layer0_out[2805] ^ layer0_out[2806]);
    assign layer1_out[770] = ~(layer0_out[3996] | layer0_out[3997]);
    assign layer1_out[771] = ~layer0_out[1291];
    assign layer1_out[772] = ~layer0_out[3346] | layer0_out[3347];
    assign layer1_out[773] = ~layer0_out[2260];
    assign layer1_out[774] = layer0_out[4112];
    assign layer1_out[775] = layer0_out[4735] & ~layer0_out[4736];
    assign layer1_out[776] = layer0_out[5548];
    assign layer1_out[777] = layer0_out[824] & ~layer0_out[823];
    assign layer1_out[778] = ~layer0_out[7155];
    assign layer1_out[779] = ~layer0_out[3636];
    assign layer1_out[780] = layer0_out[4013] & ~layer0_out[4012];
    assign layer1_out[781] = layer0_out[7061];
    assign layer1_out[782] = ~layer0_out[5679] | layer0_out[5678];
    assign layer1_out[783] = ~layer0_out[6020] | layer0_out[6019];
    assign layer1_out[784] = ~layer0_out[592] | layer0_out[591];
    assign layer1_out[785] = layer0_out[6090];
    assign layer1_out[786] = ~layer0_out[2770] | layer0_out[2769];
    assign layer1_out[787] = layer0_out[1864] & ~layer0_out[1865];
    assign layer1_out[788] = layer0_out[1810] ^ layer0_out[1811];
    assign layer1_out[789] = 1'b0;
    assign layer1_out[790] = layer0_out[7692] | layer0_out[7693];
    assign layer1_out[791] = layer0_out[846];
    assign layer1_out[792] = ~layer0_out[4029];
    assign layer1_out[793] = layer0_out[4392] | layer0_out[4393];
    assign layer1_out[794] = layer0_out[1692];
    assign layer1_out[795] = ~(layer0_out[5693] & layer0_out[5694]);
    assign layer1_out[796] = layer0_out[7843] & ~layer0_out[7842];
    assign layer1_out[797] = layer0_out[5503] | layer0_out[5504];
    assign layer1_out[798] = layer0_out[7964] & ~layer0_out[7963];
    assign layer1_out[799] = layer0_out[5332];
    assign layer1_out[800] = layer0_out[5513];
    assign layer1_out[801] = ~layer0_out[5987];
    assign layer1_out[802] = ~(layer0_out[5357] & layer0_out[5358]);
    assign layer1_out[803] = ~layer0_out[102];
    assign layer1_out[804] = ~layer0_out[3477] | layer0_out[3476];
    assign layer1_out[805] = layer0_out[3474];
    assign layer1_out[806] = layer0_out[6269] & ~layer0_out[6270];
    assign layer1_out[807] = ~(layer0_out[6606] & layer0_out[6607]);
    assign layer1_out[808] = layer0_out[4135] & ~layer0_out[4134];
    assign layer1_out[809] = layer0_out[1197] | layer0_out[1198];
    assign layer1_out[810] = ~layer0_out[5035];
    assign layer1_out[811] = layer0_out[4177] & ~layer0_out[4176];
    assign layer1_out[812] = layer0_out[7908] | layer0_out[7909];
    assign layer1_out[813] = layer0_out[5244] & ~layer0_out[5243];
    assign layer1_out[814] = ~(layer0_out[4049] & layer0_out[4050]);
    assign layer1_out[815] = 1'b1;
    assign layer1_out[816] = layer0_out[266] | layer0_out[267];
    assign layer1_out[817] = 1'b1;
    assign layer1_out[818] = ~layer0_out[3234] | layer0_out[3233];
    assign layer1_out[819] = layer0_out[3966] | layer0_out[3967];
    assign layer1_out[820] = ~(layer0_out[7163] ^ layer0_out[7164]);
    assign layer1_out[821] = ~(layer0_out[3521] & layer0_out[3522]);
    assign layer1_out[822] = layer0_out[4565];
    assign layer1_out[823] = layer0_out[3580];
    assign layer1_out[824] = 1'b1;
    assign layer1_out[825] = 1'b1;
    assign layer1_out[826] = ~layer0_out[2745];
    assign layer1_out[827] = layer0_out[1141] | layer0_out[1142];
    assign layer1_out[828] = layer0_out[4256] ^ layer0_out[4257];
    assign layer1_out[829] = ~layer0_out[6312];
    assign layer1_out[830] = ~layer0_out[2359];
    assign layer1_out[831] = ~(layer0_out[7936] & layer0_out[7937]);
    assign layer1_out[832] = ~(layer0_out[2718] & layer0_out[2719]);
    assign layer1_out[833] = ~(layer0_out[3385] & layer0_out[3386]);
    assign layer1_out[834] = ~(layer0_out[7100] & layer0_out[7101]);
    assign layer1_out[835] = ~layer0_out[7270];
    assign layer1_out[836] = ~layer0_out[4370];
    assign layer1_out[837] = layer0_out[5506] | layer0_out[5507];
    assign layer1_out[838] = layer0_out[2477];
    assign layer1_out[839] = ~(layer0_out[1866] ^ layer0_out[1867]);
    assign layer1_out[840] = layer0_out[6346] & ~layer0_out[6345];
    assign layer1_out[841] = ~layer0_out[1447] | layer0_out[1448];
    assign layer1_out[842] = ~layer0_out[237];
    assign layer1_out[843] = 1'b0;
    assign layer1_out[844] = layer0_out[4439] & ~layer0_out[4440];
    assign layer1_out[845] = ~layer0_out[314];
    assign layer1_out[846] = layer0_out[3411];
    assign layer1_out[847] = layer0_out[7171];
    assign layer1_out[848] = layer0_out[4192] & ~layer0_out[4191];
    assign layer1_out[849] = ~(layer0_out[6792] & layer0_out[6793]);
    assign layer1_out[850] = ~layer0_out[88] | layer0_out[89];
    assign layer1_out[851] = ~(layer0_out[6949] & layer0_out[6950]);
    assign layer1_out[852] = layer0_out[4187] & layer0_out[4188];
    assign layer1_out[853] = layer0_out[5754] | layer0_out[5755];
    assign layer1_out[854] = layer0_out[12] & layer0_out[13];
    assign layer1_out[855] = layer0_out[143] ^ layer0_out[144];
    assign layer1_out[856] = layer0_out[7864] ^ layer0_out[7865];
    assign layer1_out[857] = layer0_out[5483] & ~layer0_out[5482];
    assign layer1_out[858] = layer0_out[2328] & layer0_out[2329];
    assign layer1_out[859] = ~layer0_out[4195];
    assign layer1_out[860] = layer0_out[3138];
    assign layer1_out[861] = layer0_out[1247];
    assign layer1_out[862] = layer0_out[3553];
    assign layer1_out[863] = layer0_out[1011];
    assign layer1_out[864] = layer0_out[2360] & layer0_out[2361];
    assign layer1_out[865] = ~layer0_out[1293] | layer0_out[1292];
    assign layer1_out[866] = layer0_out[2274] ^ layer0_out[2275];
    assign layer1_out[867] = ~(layer0_out[2952] | layer0_out[2953]);
    assign layer1_out[868] = layer0_out[3559];
    assign layer1_out[869] = layer0_out[762];
    assign layer1_out[870] = ~layer0_out[3809];
    assign layer1_out[871] = layer0_out[7185];
    assign layer1_out[872] = ~(layer0_out[5] | layer0_out[6]);
    assign layer1_out[873] = layer0_out[1272] & ~layer0_out[1273];
    assign layer1_out[874] = layer0_out[6625] & ~layer0_out[6626];
    assign layer1_out[875] = layer0_out[5665] & ~layer0_out[5664];
    assign layer1_out[876] = layer0_out[1742] & ~layer0_out[1743];
    assign layer1_out[877] = layer0_out[7282] & ~layer0_out[7281];
    assign layer1_out[878] = layer0_out[1322] & ~layer0_out[1321];
    assign layer1_out[879] = ~(layer0_out[276] | layer0_out[277]);
    assign layer1_out[880] = ~layer0_out[722];
    assign layer1_out[881] = layer0_out[112] | layer0_out[113];
    assign layer1_out[882] = ~layer0_out[7205];
    assign layer1_out[883] = ~layer0_out[5884];
    assign layer1_out[884] = ~layer0_out[4898];
    assign layer1_out[885] = layer0_out[6679];
    assign layer1_out[886] = ~(layer0_out[2035] ^ layer0_out[2036]);
    assign layer1_out[887] = layer0_out[5505] | layer0_out[5506];
    assign layer1_out[888] = layer0_out[6990];
    assign layer1_out[889] = ~layer0_out[7896] | layer0_out[7895];
    assign layer1_out[890] = layer0_out[339];
    assign layer1_out[891] = layer0_out[2486] & ~layer0_out[2485];
    assign layer1_out[892] = layer0_out[6535] & ~layer0_out[6534];
    assign layer1_out[893] = layer0_out[6920] & ~layer0_out[6919];
    assign layer1_out[894] = layer0_out[1474] | layer0_out[1475];
    assign layer1_out[895] = layer0_out[6930];
    assign layer1_out[896] = layer0_out[1191] ^ layer0_out[1192];
    assign layer1_out[897] = layer0_out[3062];
    assign layer1_out[898] = ~(layer0_out[3380] & layer0_out[3381]);
    assign layer1_out[899] = ~(layer0_out[6985] | layer0_out[6986]);
    assign layer1_out[900] = ~(layer0_out[6616] & layer0_out[6617]);
    assign layer1_out[901] = layer0_out[2354];
    assign layer1_out[902] = 1'b0;
    assign layer1_out[903] = ~(layer0_out[4352] & layer0_out[4353]);
    assign layer1_out[904] = layer0_out[576];
    assign layer1_out[905] = layer0_out[5265];
    assign layer1_out[906] = ~layer0_out[6735];
    assign layer1_out[907] = ~layer0_out[3385];
    assign layer1_out[908] = 1'b1;
    assign layer1_out[909] = ~(layer0_out[4974] & layer0_out[4975]);
    assign layer1_out[910] = layer0_out[7439] & ~layer0_out[7438];
    assign layer1_out[911] = layer0_out[3335] & ~layer0_out[3334];
    assign layer1_out[912] = layer0_out[3839];
    assign layer1_out[913] = 1'b1;
    assign layer1_out[914] = ~layer0_out[2561];
    assign layer1_out[915] = ~(layer0_out[2129] & layer0_out[2130]);
    assign layer1_out[916] = ~(layer0_out[1347] | layer0_out[1348]);
    assign layer1_out[917] = ~layer0_out[2399] | layer0_out[2400];
    assign layer1_out[918] = ~layer0_out[4959];
    assign layer1_out[919] = layer0_out[2113];
    assign layer1_out[920] = ~(layer0_out[2240] ^ layer0_out[2241]);
    assign layer1_out[921] = layer0_out[5147] | layer0_out[5148];
    assign layer1_out[922] = ~(layer0_out[4190] | layer0_out[4191]);
    assign layer1_out[923] = layer0_out[6740] & ~layer0_out[6741];
    assign layer1_out[924] = layer0_out[939];
    assign layer1_out[925] = layer0_out[3732] & layer0_out[3733];
    assign layer1_out[926] = layer0_out[6986] ^ layer0_out[6987];
    assign layer1_out[927] = ~(layer0_out[5935] | layer0_out[5936]);
    assign layer1_out[928] = layer0_out[7356] & ~layer0_out[7357];
    assign layer1_out[929] = ~layer0_out[5381] | layer0_out[5380];
    assign layer1_out[930] = 1'b1;
    assign layer1_out[931] = layer0_out[495] & ~layer0_out[494];
    assign layer1_out[932] = ~layer0_out[6754] | layer0_out[6753];
    assign layer1_out[933] = ~layer0_out[1998];
    assign layer1_out[934] = 1'b1;
    assign layer1_out[935] = ~layer0_out[2352] | layer0_out[2353];
    assign layer1_out[936] = ~(layer0_out[5015] | layer0_out[5016]);
    assign layer1_out[937] = ~(layer0_out[7366] & layer0_out[7367]);
    assign layer1_out[938] = ~layer0_out[1586];
    assign layer1_out[939] = layer0_out[2564] & ~layer0_out[2563];
    assign layer1_out[940] = layer0_out[3952] & ~layer0_out[3953];
    assign layer1_out[941] = layer0_out[4167] | layer0_out[4168];
    assign layer1_out[942] = ~layer0_out[7924] | layer0_out[7925];
    assign layer1_out[943] = layer0_out[263] | layer0_out[264];
    assign layer1_out[944] = ~(layer0_out[1903] ^ layer0_out[1904]);
    assign layer1_out[945] = ~(layer0_out[3413] ^ layer0_out[3414]);
    assign layer1_out[946] = layer0_out[5091] | layer0_out[5092];
    assign layer1_out[947] = ~layer0_out[7357] | layer0_out[7358];
    assign layer1_out[948] = layer0_out[3047] ^ layer0_out[3048];
    assign layer1_out[949] = ~layer0_out[1617];
    assign layer1_out[950] = ~layer0_out[7535] | layer0_out[7536];
    assign layer1_out[951] = ~(layer0_out[7405] | layer0_out[7406]);
    assign layer1_out[952] = 1'b0;
    assign layer1_out[953] = ~layer0_out[2109];
    assign layer1_out[954] = layer0_out[3150] ^ layer0_out[3151];
    assign layer1_out[955] = ~(layer0_out[1549] & layer0_out[1550]);
    assign layer1_out[956] = ~layer0_out[5225];
    assign layer1_out[957] = layer0_out[4227];
    assign layer1_out[958] = layer0_out[598] & ~layer0_out[597];
    assign layer1_out[959] = layer0_out[5343];
    assign layer1_out[960] = ~layer0_out[3202] | layer0_out[3201];
    assign layer1_out[961] = ~(layer0_out[3307] | layer0_out[3308]);
    assign layer1_out[962] = ~(layer0_out[7780] | layer0_out[7781]);
    assign layer1_out[963] = ~(layer0_out[535] | layer0_out[536]);
    assign layer1_out[964] = ~layer0_out[7397] | layer0_out[7396];
    assign layer1_out[965] = ~layer0_out[90];
    assign layer1_out[966] = layer0_out[4829];
    assign layer1_out[967] = layer0_out[1471] | layer0_out[1472];
    assign layer1_out[968] = layer0_out[5200];
    assign layer1_out[969] = ~layer0_out[3936];
    assign layer1_out[970] = layer0_out[5883] & ~layer0_out[5882];
    assign layer1_out[971] = layer0_out[1897] ^ layer0_out[1898];
    assign layer1_out[972] = ~layer0_out[3032] | layer0_out[3031];
    assign layer1_out[973] = layer0_out[2090] & ~layer0_out[2091];
    assign layer1_out[974] = layer0_out[6643] & ~layer0_out[6642];
    assign layer1_out[975] = layer0_out[3370];
    assign layer1_out[976] = layer0_out[6556];
    assign layer1_out[977] = layer0_out[3117] & ~layer0_out[3116];
    assign layer1_out[978] = layer0_out[924] & layer0_out[925];
    assign layer1_out[979] = ~(layer0_out[5269] | layer0_out[5270]);
    assign layer1_out[980] = ~layer0_out[3266] | layer0_out[3265];
    assign layer1_out[981] = ~layer0_out[771];
    assign layer1_out[982] = ~layer0_out[1698];
    assign layer1_out[983] = ~layer0_out[1657] | layer0_out[1658];
    assign layer1_out[984] = layer0_out[3889] & ~layer0_out[3888];
    assign layer1_out[985] = layer0_out[4847] & ~layer0_out[4846];
    assign layer1_out[986] = ~layer0_out[1319] | layer0_out[1318];
    assign layer1_out[987] = ~layer0_out[3517];
    assign layer1_out[988] = ~(layer0_out[2075] & layer0_out[2076]);
    assign layer1_out[989] = ~(layer0_out[7009] ^ layer0_out[7010]);
    assign layer1_out[990] = layer0_out[4351] & ~layer0_out[4352];
    assign layer1_out[991] = ~layer0_out[4900];
    assign layer1_out[992] = 1'b1;
    assign layer1_out[993] = ~layer0_out[6671] | layer0_out[6670];
    assign layer1_out[994] = layer0_out[86] & layer0_out[87];
    assign layer1_out[995] = layer0_out[1363];
    assign layer1_out[996] = layer0_out[3798];
    assign layer1_out[997] = ~(layer0_out[1971] ^ layer0_out[1972]);
    assign layer1_out[998] = ~layer0_out[942] | layer0_out[941];
    assign layer1_out[999] = layer0_out[1313];
    assign layer1_out[1000] = ~(layer0_out[7422] & layer0_out[7423]);
    assign layer1_out[1001] = layer0_out[6733] & ~layer0_out[6732];
    assign layer1_out[1002] = layer0_out[5112] & ~layer0_out[5113];
    assign layer1_out[1003] = ~(layer0_out[7377] ^ layer0_out[7378]);
    assign layer1_out[1004] = layer0_out[764] | layer0_out[765];
    assign layer1_out[1005] = ~layer0_out[1469];
    assign layer1_out[1006] = layer0_out[7258] | layer0_out[7259];
    assign layer1_out[1007] = layer0_out[1232] & layer0_out[1233];
    assign layer1_out[1008] = ~layer0_out[6386];
    assign layer1_out[1009] = layer0_out[998] ^ layer0_out[999];
    assign layer1_out[1010] = ~(layer0_out[6950] ^ layer0_out[6951]);
    assign layer1_out[1011] = ~layer0_out[3622];
    assign layer1_out[1012] = ~layer0_out[2234];
    assign layer1_out[1013] = ~layer0_out[4631];
    assign layer1_out[1014] = ~layer0_out[2989] | layer0_out[2988];
    assign layer1_out[1015] = ~(layer0_out[1834] & layer0_out[1835]);
    assign layer1_out[1016] = layer0_out[6408] & ~layer0_out[6409];
    assign layer1_out[1017] = layer0_out[181];
    assign layer1_out[1018] = ~layer0_out[6238] | layer0_out[6237];
    assign layer1_out[1019] = ~layer0_out[1738] | layer0_out[1737];
    assign layer1_out[1020] = layer0_out[1708];
    assign layer1_out[1021] = layer0_out[5787] & ~layer0_out[5788];
    assign layer1_out[1022] = ~(layer0_out[6164] ^ layer0_out[6165]);
    assign layer1_out[1023] = layer0_out[4456];
    assign layer1_out[1024] = ~(layer0_out[75] & layer0_out[76]);
    assign layer1_out[1025] = layer0_out[97] | layer0_out[98];
    assign layer1_out[1026] = 1'b0;
    assign layer1_out[1027] = ~(layer0_out[4908] ^ layer0_out[4909]);
    assign layer1_out[1028] = ~layer0_out[813];
    assign layer1_out[1029] = ~(layer0_out[2086] | layer0_out[2087]);
    assign layer1_out[1030] = ~(layer0_out[1257] ^ layer0_out[1258]);
    assign layer1_out[1031] = ~layer0_out[3275];
    assign layer1_out[1032] = 1'b1;
    assign layer1_out[1033] = 1'b1;
    assign layer1_out[1034] = ~layer0_out[6816];
    assign layer1_out[1035] = ~layer0_out[2990] | layer0_out[2989];
    assign layer1_out[1036] = layer0_out[7460] & layer0_out[7461];
    assign layer1_out[1037] = 1'b1;
    assign layer1_out[1038] = layer0_out[872];
    assign layer1_out[1039] = ~layer0_out[5272];
    assign layer1_out[1040] = ~(layer0_out[2871] ^ layer0_out[2872]);
    assign layer1_out[1041] = ~layer0_out[6527];
    assign layer1_out[1042] = layer0_out[7258];
    assign layer1_out[1043] = ~layer0_out[19] | layer0_out[18];
    assign layer1_out[1044] = ~(layer0_out[6714] ^ layer0_out[6715]);
    assign layer1_out[1045] = layer0_out[3377] | layer0_out[3378];
    assign layer1_out[1046] = layer0_out[3792] & ~layer0_out[3791];
    assign layer1_out[1047] = ~layer0_out[6944];
    assign layer1_out[1048] = layer0_out[6113] & layer0_out[6114];
    assign layer1_out[1049] = layer0_out[3440];
    assign layer1_out[1050] = layer0_out[4278];
    assign layer1_out[1051] = 1'b0;
    assign layer1_out[1052] = ~(layer0_out[1018] | layer0_out[1019]);
    assign layer1_out[1053] = layer0_out[6029] & layer0_out[6030];
    assign layer1_out[1054] = ~(layer0_out[6456] ^ layer0_out[6457]);
    assign layer1_out[1055] = ~layer0_out[2876];
    assign layer1_out[1056] = ~layer0_out[4299] | layer0_out[4300];
    assign layer1_out[1057] = ~layer0_out[6538];
    assign layer1_out[1058] = ~layer0_out[2767];
    assign layer1_out[1059] = layer0_out[6120] & ~layer0_out[6121];
    assign layer1_out[1060] = layer0_out[778];
    assign layer1_out[1061] = ~(layer0_out[5937] | layer0_out[5938]);
    assign layer1_out[1062] = ~layer0_out[1889] | layer0_out[1890];
    assign layer1_out[1063] = layer0_out[1851] ^ layer0_out[1852];
    assign layer1_out[1064] = layer0_out[115] | layer0_out[116];
    assign layer1_out[1065] = 1'b0;
    assign layer1_out[1066] = ~layer0_out[4509] | layer0_out[4510];
    assign layer1_out[1067] = ~(layer0_out[6840] & layer0_out[6841]);
    assign layer1_out[1068] = layer0_out[77];
    assign layer1_out[1069] = layer0_out[2159] & ~layer0_out[2158];
    assign layer1_out[1070] = ~layer0_out[5278];
    assign layer1_out[1071] = ~(layer0_out[6570] & layer0_out[6571]);
    assign layer1_out[1072] = layer0_out[7816] | layer0_out[7817];
    assign layer1_out[1073] = ~layer0_out[176];
    assign layer1_out[1074] = ~(layer0_out[4295] | layer0_out[4296]);
    assign layer1_out[1075] = ~(layer0_out[31] & layer0_out[32]);
    assign layer1_out[1076] = layer0_out[5170] & layer0_out[5171];
    assign layer1_out[1077] = ~layer0_out[5666];
    assign layer1_out[1078] = ~layer0_out[6554] | layer0_out[6553];
    assign layer1_out[1079] = 1'b0;
    assign layer1_out[1080] = layer0_out[3663] & ~layer0_out[3664];
    assign layer1_out[1081] = layer0_out[5401] | layer0_out[5402];
    assign layer1_out[1082] = ~(layer0_out[3485] | layer0_out[3486]);
    assign layer1_out[1083] = ~(layer0_out[1048] & layer0_out[1049]);
    assign layer1_out[1084] = ~layer0_out[4636] | layer0_out[4635];
    assign layer1_out[1085] = layer0_out[1025] ^ layer0_out[1026];
    assign layer1_out[1086] = ~(layer0_out[487] | layer0_out[488]);
    assign layer1_out[1087] = layer0_out[7107] ^ layer0_out[7108];
    assign layer1_out[1088] = layer0_out[7454] & ~layer0_out[7455];
    assign layer1_out[1089] = 1'b1;
    assign layer1_out[1090] = layer0_out[3687] & ~layer0_out[3686];
    assign layer1_out[1091] = layer0_out[5915];
    assign layer1_out[1092] = layer0_out[7148] & layer0_out[7149];
    assign layer1_out[1093] = ~(layer0_out[7054] ^ layer0_out[7055]);
    assign layer1_out[1094] = layer0_out[6814] | layer0_out[6815];
    assign layer1_out[1095] = ~layer0_out[7567];
    assign layer1_out[1096] = 1'b1;
    assign layer1_out[1097] = ~layer0_out[4963];
    assign layer1_out[1098] = layer0_out[6974] ^ layer0_out[6975];
    assign layer1_out[1099] = ~(layer0_out[1928] | layer0_out[1929]);
    assign layer1_out[1100] = layer0_out[332] | layer0_out[333];
    assign layer1_out[1101] = layer0_out[5746] | layer0_out[5747];
    assign layer1_out[1102] = ~layer0_out[5673];
    assign layer1_out[1103] = layer0_out[5761] ^ layer0_out[5762];
    assign layer1_out[1104] = ~(layer0_out[7622] | layer0_out[7623]);
    assign layer1_out[1105] = layer0_out[5860] & layer0_out[5861];
    assign layer1_out[1106] = layer0_out[1387];
    assign layer1_out[1107] = ~layer0_out[111] | layer0_out[110];
    assign layer1_out[1108] = 1'b1;
    assign layer1_out[1109] = ~(layer0_out[1277] & layer0_out[1278]);
    assign layer1_out[1110] = layer0_out[3110] & ~layer0_out[3109];
    assign layer1_out[1111] = layer0_out[2052] & ~layer0_out[2051];
    assign layer1_out[1112] = ~layer0_out[1818];
    assign layer1_out[1113] = ~layer0_out[7957] | layer0_out[7956];
    assign layer1_out[1114] = ~layer0_out[6608];
    assign layer1_out[1115] = ~(layer0_out[4051] & layer0_out[4052]);
    assign layer1_out[1116] = layer0_out[6096] | layer0_out[6097];
    assign layer1_out[1117] = ~layer0_out[2315] | layer0_out[2314];
    assign layer1_out[1118] = layer0_out[74] & ~layer0_out[73];
    assign layer1_out[1119] = ~(layer0_out[4657] | layer0_out[4658]);
    assign layer1_out[1120] = ~layer0_out[4166];
    assign layer1_out[1121] = ~(layer0_out[4821] | layer0_out[4822]);
    assign layer1_out[1122] = layer0_out[2658];
    assign layer1_out[1123] = layer0_out[7234];
    assign layer1_out[1124] = layer0_out[5907];
    assign layer1_out[1125] = layer0_out[1610] ^ layer0_out[1611];
    assign layer1_out[1126] = layer0_out[3184] & ~layer0_out[3183];
    assign layer1_out[1127] = ~(layer0_out[4483] & layer0_out[4484]);
    assign layer1_out[1128] = layer0_out[6475] | layer0_out[6476];
    assign layer1_out[1129] = layer0_out[1915] & layer0_out[1916];
    assign layer1_out[1130] = 1'b1;
    assign layer1_out[1131] = layer0_out[1307] ^ layer0_out[1308];
    assign layer1_out[1132] = ~layer0_out[7289] | layer0_out[7288];
    assign layer1_out[1133] = layer0_out[1566];
    assign layer1_out[1134] = ~(layer0_out[174] ^ layer0_out[175]);
    assign layer1_out[1135] = layer0_out[7681] | layer0_out[7682];
    assign layer1_out[1136] = ~layer0_out[4381];
    assign layer1_out[1137] = layer0_out[203];
    assign layer1_out[1138] = ~(layer0_out[5813] | layer0_out[5814]);
    assign layer1_out[1139] = layer0_out[167];
    assign layer1_out[1140] = layer0_out[4895] & ~layer0_out[4894];
    assign layer1_out[1141] = ~(layer0_out[4494] & layer0_out[4495]);
    assign layer1_out[1142] = ~layer0_out[375];
    assign layer1_out[1143] = layer0_out[5651] & ~layer0_out[5652];
    assign layer1_out[1144] = layer0_out[5091] & ~layer0_out[5090];
    assign layer1_out[1145] = ~layer0_out[188] | layer0_out[189];
    assign layer1_out[1146] = layer0_out[4524];
    assign layer1_out[1147] = ~(layer0_out[5808] ^ layer0_out[5809]);
    assign layer1_out[1148] = ~(layer0_out[7611] & layer0_out[7612]);
    assign layer1_out[1149] = layer0_out[2983] ^ layer0_out[2984];
    assign layer1_out[1150] = layer0_out[851] & ~layer0_out[852];
    assign layer1_out[1151] = ~(layer0_out[2488] ^ layer0_out[2489]);
    assign layer1_out[1152] = layer0_out[3492] & layer0_out[3493];
    assign layer1_out[1153] = layer0_out[2579];
    assign layer1_out[1154] = layer0_out[381];
    assign layer1_out[1155] = ~(layer0_out[6951] & layer0_out[6952]);
    assign layer1_out[1156] = layer0_out[200];
    assign layer1_out[1157] = 1'b1;
    assign layer1_out[1158] = ~layer0_out[2198];
    assign layer1_out[1159] = 1'b0;
    assign layer1_out[1160] = ~layer0_out[5647];
    assign layer1_out[1161] = layer0_out[2329] & ~layer0_out[2330];
    assign layer1_out[1162] = layer0_out[4407] | layer0_out[4408];
    assign layer1_out[1163] = ~(layer0_out[2466] & layer0_out[2467]);
    assign layer1_out[1164] = layer0_out[507] ^ layer0_out[508];
    assign layer1_out[1165] = layer0_out[3035];
    assign layer1_out[1166] = ~layer0_out[7378];
    assign layer1_out[1167] = ~(layer0_out[20] & layer0_out[21]);
    assign layer1_out[1168] = ~layer0_out[6594];
    assign layer1_out[1169] = layer0_out[4105];
    assign layer1_out[1170] = ~(layer0_out[890] ^ layer0_out[891]);
    assign layer1_out[1171] = layer0_out[11];
    assign layer1_out[1172] = layer0_out[5046] & ~layer0_out[5045];
    assign layer1_out[1173] = layer0_out[1559] | layer0_out[1560];
    assign layer1_out[1174] = layer0_out[7904] ^ layer0_out[7905];
    assign layer1_out[1175] = layer0_out[725] & layer0_out[726];
    assign layer1_out[1176] = layer0_out[2661] & layer0_out[2662];
    assign layer1_out[1177] = layer0_out[7232] & layer0_out[7233];
    assign layer1_out[1178] = layer0_out[7786];
    assign layer1_out[1179] = 1'b0;
    assign layer1_out[1180] = layer0_out[2671];
    assign layer1_out[1181] = layer0_out[2585] ^ layer0_out[2586];
    assign layer1_out[1182] = ~(layer0_out[2852] ^ layer0_out[2853]);
    assign layer1_out[1183] = layer0_out[383] & ~layer0_out[382];
    assign layer1_out[1184] = ~layer0_out[7485] | layer0_out[7486];
    assign layer1_out[1185] = layer0_out[7767] & ~layer0_out[7768];
    assign layer1_out[1186] = layer0_out[6770] & ~layer0_out[6771];
    assign layer1_out[1187] = ~(layer0_out[3573] & layer0_out[3574]);
    assign layer1_out[1188] = layer0_out[6240];
    assign layer1_out[1189] = ~(layer0_out[2787] | layer0_out[2788]);
    assign layer1_out[1190] = layer0_out[4211] & layer0_out[4212];
    assign layer1_out[1191] = ~layer0_out[7931] | layer0_out[7930];
    assign layer1_out[1192] = ~layer0_out[1174] | layer0_out[1173];
    assign layer1_out[1193] = layer0_out[1564] & ~layer0_out[1563];
    assign layer1_out[1194] = ~layer0_out[7202];
    assign layer1_out[1195] = layer0_out[1660] | layer0_out[1661];
    assign layer1_out[1196] = layer0_out[3666] & ~layer0_out[3667];
    assign layer1_out[1197] = ~layer0_out[1349] | layer0_out[1348];
    assign layer1_out[1198] = ~layer0_out[4948] | layer0_out[4949];
    assign layer1_out[1199] = layer0_out[3888];
    assign layer1_out[1200] = ~layer0_out[7491];
    assign layer1_out[1201] = layer0_out[2590];
    assign layer1_out[1202] = ~layer0_out[7560];
    assign layer1_out[1203] = ~layer0_out[250];
    assign layer1_out[1204] = ~(layer0_out[686] | layer0_out[687]);
    assign layer1_out[1205] = ~layer0_out[4809];
    assign layer1_out[1206] = ~(layer0_out[2510] | layer0_out[2511]);
    assign layer1_out[1207] = layer0_out[7891] & ~layer0_out[7890];
    assign layer1_out[1208] = ~(layer0_out[2400] | layer0_out[2401]);
    assign layer1_out[1209] = ~layer0_out[7253] | layer0_out[7254];
    assign layer1_out[1210] = layer0_out[4769];
    assign layer1_out[1211] = ~(layer0_out[1562] & layer0_out[1563]);
    assign layer1_out[1212] = ~layer0_out[5282] | layer0_out[5281];
    assign layer1_out[1213] = ~(layer0_out[856] & layer0_out[857]);
    assign layer1_out[1214] = layer0_out[7042] & layer0_out[7043];
    assign layer1_out[1215] = layer0_out[68];
    assign layer1_out[1216] = ~layer0_out[2763];
    assign layer1_out[1217] = layer0_out[1441];
    assign layer1_out[1218] = ~layer0_out[6381] | layer0_out[6382];
    assign layer1_out[1219] = ~layer0_out[4116] | layer0_out[4115];
    assign layer1_out[1220] = layer0_out[4638] & layer0_out[4639];
    assign layer1_out[1221] = ~(layer0_out[6745] ^ layer0_out[6746]);
    assign layer1_out[1222] = layer0_out[4061] & ~layer0_out[4060];
    assign layer1_out[1223] = ~layer0_out[5895] | layer0_out[5896];
    assign layer1_out[1224] = layer0_out[3067] & ~layer0_out[3066];
    assign layer1_out[1225] = ~(layer0_out[7001] & layer0_out[7002]);
    assign layer1_out[1226] = layer0_out[2182];
    assign layer1_out[1227] = ~layer0_out[1676] | layer0_out[1675];
    assign layer1_out[1228] = layer0_out[6811] & layer0_out[6812];
    assign layer1_out[1229] = ~layer0_out[5397] | layer0_out[5398];
    assign layer1_out[1230] = ~layer0_out[363];
    assign layer1_out[1231] = layer0_out[4470];
    assign layer1_out[1232] = 1'b1;
    assign layer1_out[1233] = ~layer0_out[5765];
    assign layer1_out[1234] = layer0_out[5448] ^ layer0_out[5449];
    assign layer1_out[1235] = ~layer0_out[3579] | layer0_out[3578];
    assign layer1_out[1236] = ~layer0_out[7772];
    assign layer1_out[1237] = layer0_out[1071];
    assign layer1_out[1238] = ~(layer0_out[1638] | layer0_out[1639]);
    assign layer1_out[1239] = ~layer0_out[6850] | layer0_out[6849];
    assign layer1_out[1240] = ~(layer0_out[4360] | layer0_out[4361]);
    assign layer1_out[1241] = layer0_out[5801];
    assign layer1_out[1242] = ~layer0_out[438];
    assign layer1_out[1243] = layer0_out[4540];
    assign layer1_out[1244] = layer0_out[759] & layer0_out[760];
    assign layer1_out[1245] = layer0_out[5716] | layer0_out[5717];
    assign layer1_out[1246] = ~layer0_out[3185] | layer0_out[3186];
    assign layer1_out[1247] = ~(layer0_out[1213] & layer0_out[1214]);
    assign layer1_out[1248] = ~layer0_out[3887];
    assign layer1_out[1249] = ~layer0_out[7117] | layer0_out[7118];
    assign layer1_out[1250] = ~(layer0_out[4165] | layer0_out[4166]);
    assign layer1_out[1251] = layer0_out[4046];
    assign layer1_out[1252] = ~layer0_out[6039] | layer0_out[6038];
    assign layer1_out[1253] = ~layer0_out[6693] | layer0_out[6694];
    assign layer1_out[1254] = ~layer0_out[631];
    assign layer1_out[1255] = ~layer0_out[725] | layer0_out[724];
    assign layer1_out[1256] = layer0_out[5105];
    assign layer1_out[1257] = layer0_out[5998];
    assign layer1_out[1258] = layer0_out[723] ^ layer0_out[724];
    assign layer1_out[1259] = 1'b0;
    assign layer1_out[1260] = ~layer0_out[7751];
    assign layer1_out[1261] = ~layer0_out[814];
    assign layer1_out[1262] = layer0_out[5026] & ~layer0_out[5025];
    assign layer1_out[1263] = layer0_out[5422];
    assign layer1_out[1264] = layer0_out[7233] & ~layer0_out[7234];
    assign layer1_out[1265] = ~(layer0_out[5980] & layer0_out[5981]);
    assign layer1_out[1266] = layer0_out[2293] ^ layer0_out[2294];
    assign layer1_out[1267] = ~layer0_out[7367];
    assign layer1_out[1268] = layer0_out[5231] & layer0_out[5232];
    assign layer1_out[1269] = layer0_out[1964];
    assign layer1_out[1270] = layer0_out[5211];
    assign layer1_out[1271] = layer0_out[5963] & layer0_out[5964];
    assign layer1_out[1272] = layer0_out[7203] & ~layer0_out[7202];
    assign layer1_out[1273] = ~layer0_out[6244];
    assign layer1_out[1274] = ~(layer0_out[6733] & layer0_out[6734]);
    assign layer1_out[1275] = 1'b1;
    assign layer1_out[1276] = layer0_out[6762] & ~layer0_out[6761];
    assign layer1_out[1277] = layer0_out[706] | layer0_out[707];
    assign layer1_out[1278] = layer0_out[2271];
    assign layer1_out[1279] = ~layer0_out[6050] | layer0_out[6049];
    assign layer1_out[1280] = ~layer0_out[837] | layer0_out[836];
    assign layer1_out[1281] = layer0_out[6595];
    assign layer1_out[1282] = ~(layer0_out[5161] | layer0_out[5162]);
    assign layer1_out[1283] = layer0_out[2447];
    assign layer1_out[1284] = layer0_out[7552];
    assign layer1_out[1285] = layer0_out[4189] & ~layer0_out[4188];
    assign layer1_out[1286] = layer0_out[2945] & layer0_out[2946];
    assign layer1_out[1287] = ~layer0_out[3464];
    assign layer1_out[1288] = ~(layer0_out[4766] & layer0_out[4767]);
    assign layer1_out[1289] = layer0_out[5790] & ~layer0_out[5789];
    assign layer1_out[1290] = 1'b1;
    assign layer1_out[1291] = ~(layer0_out[7461] ^ layer0_out[7462]);
    assign layer1_out[1292] = layer0_out[5858];
    assign layer1_out[1293] = layer0_out[595];
    assign layer1_out[1294] = ~layer0_out[7759];
    assign layer1_out[1295] = layer0_out[4663];
    assign layer1_out[1296] = layer0_out[6189];
    assign layer1_out[1297] = layer0_out[688] & ~layer0_out[689];
    assign layer1_out[1298] = layer0_out[691];
    assign layer1_out[1299] = layer0_out[4590] & layer0_out[4591];
    assign layer1_out[1300] = layer0_out[2108];
    assign layer1_out[1301] = ~layer0_out[407] | layer0_out[408];
    assign layer1_out[1302] = layer0_out[2318] & layer0_out[2319];
    assign layer1_out[1303] = ~layer0_out[1597] | layer0_out[1596];
    assign layer1_out[1304] = ~(layer0_out[2138] ^ layer0_out[2139]);
    assign layer1_out[1305] = layer0_out[6810] & ~layer0_out[6811];
    assign layer1_out[1306] = ~layer0_out[7607] | layer0_out[7608];
    assign layer1_out[1307] = ~(layer0_out[4928] & layer0_out[4929]);
    assign layer1_out[1308] = layer0_out[2655] & layer0_out[2656];
    assign layer1_out[1309] = 1'b0;
    assign layer1_out[1310] = ~(layer0_out[2764] | layer0_out[2765]);
    assign layer1_out[1311] = ~layer0_out[5211];
    assign layer1_out[1312] = ~layer0_out[1056] | layer0_out[1057];
    assign layer1_out[1313] = ~(layer0_out[1097] | layer0_out[1098]);
    assign layer1_out[1314] = layer0_out[1682] & ~layer0_out[1681];
    assign layer1_out[1315] = layer0_out[2217];
    assign layer1_out[1316] = layer0_out[971] & ~layer0_out[970];
    assign layer1_out[1317] = ~layer0_out[2971] | layer0_out[2972];
    assign layer1_out[1318] = layer0_out[3547];
    assign layer1_out[1319] = layer0_out[1755] & layer0_out[1756];
    assign layer1_out[1320] = ~layer0_out[2524] | layer0_out[2523];
    assign layer1_out[1321] = layer0_out[1966] & ~layer0_out[1965];
    assign layer1_out[1322] = ~(layer0_out[2812] & layer0_out[2813]);
    assign layer1_out[1323] = layer0_out[7086] & layer0_out[7087];
    assign layer1_out[1324] = ~layer0_out[4162] | layer0_out[4163];
    assign layer1_out[1325] = layer0_out[1877] ^ layer0_out[1878];
    assign layer1_out[1326] = ~layer0_out[940] | layer0_out[939];
    assign layer1_out[1327] = 1'b1;
    assign layer1_out[1328] = layer0_out[3297];
    assign layer1_out[1329] = layer0_out[7237] & ~layer0_out[7236];
    assign layer1_out[1330] = layer0_out[7807] & layer0_out[7808];
    assign layer1_out[1331] = ~(layer0_out[242] | layer0_out[243]);
    assign layer1_out[1332] = layer0_out[4080] & ~layer0_out[4079];
    assign layer1_out[1333] = layer0_out[3151];
    assign layer1_out[1334] = layer0_out[3483] & ~layer0_out[3482];
    assign layer1_out[1335] = layer0_out[1134] | layer0_out[1135];
    assign layer1_out[1336] = layer0_out[6519] & ~layer0_out[6518];
    assign layer1_out[1337] = 1'b1;
    assign layer1_out[1338] = layer0_out[1975] & ~layer0_out[1974];
    assign layer1_out[1339] = layer0_out[7652];
    assign layer1_out[1340] = layer0_out[1987] & layer0_out[1988];
    assign layer1_out[1341] = ~layer0_out[195];
    assign layer1_out[1342] = 1'b0;
    assign layer1_out[1343] = 1'b0;
    assign layer1_out[1344] = ~layer0_out[3058];
    assign layer1_out[1345] = ~layer0_out[3402];
    assign layer1_out[1346] = layer0_out[6342];
    assign layer1_out[1347] = ~(layer0_out[1792] | layer0_out[1793]);
    assign layer1_out[1348] = ~layer0_out[2608];
    assign layer1_out[1349] = ~layer0_out[4006];
    assign layer1_out[1350] = layer0_out[6303] & ~layer0_out[6304];
    assign layer1_out[1351] = layer0_out[3173];
    assign layer1_out[1352] = 1'b0;
    assign layer1_out[1353] = ~(layer0_out[7139] | layer0_out[7140]);
    assign layer1_out[1354] = layer0_out[2868] | layer0_out[2869];
    assign layer1_out[1355] = layer0_out[973] & ~layer0_out[972];
    assign layer1_out[1356] = ~(layer0_out[4113] ^ layer0_out[4114]);
    assign layer1_out[1357] = ~layer0_out[1995];
    assign layer1_out[1358] = ~(layer0_out[7020] ^ layer0_out[7021]);
    assign layer1_out[1359] = layer0_out[921];
    assign layer1_out[1360] = 1'b0;
    assign layer1_out[1361] = layer0_out[4336];
    assign layer1_out[1362] = 1'b1;
    assign layer1_out[1363] = 1'b0;
    assign layer1_out[1364] = layer0_out[3391] & layer0_out[3392];
    assign layer1_out[1365] = ~layer0_out[1254];
    assign layer1_out[1366] = layer0_out[992] | layer0_out[993];
    assign layer1_out[1367] = layer0_out[6524];
    assign layer1_out[1368] = ~layer0_out[210];
    assign layer1_out[1369] = layer0_out[7115] & layer0_out[7116];
    assign layer1_out[1370] = layer0_out[1008] & ~layer0_out[1009];
    assign layer1_out[1371] = ~(layer0_out[2015] & layer0_out[2016]);
    assign layer1_out[1372] = layer0_out[726] & ~layer0_out[727];
    assign layer1_out[1373] = layer0_out[1921];
    assign layer1_out[1374] = layer0_out[2053] & ~layer0_out[2054];
    assign layer1_out[1375] = layer0_out[1528] & layer0_out[1529];
    assign layer1_out[1376] = ~(layer0_out[6198] | layer0_out[6199]);
    assign layer1_out[1377] = ~layer0_out[4823];
    assign layer1_out[1378] = layer0_out[4810];
    assign layer1_out[1379] = layer0_out[7862] & layer0_out[7863];
    assign layer1_out[1380] = layer0_out[5205] & ~layer0_out[5206];
    assign layer1_out[1381] = ~layer0_out[2756];
    assign layer1_out[1382] = ~layer0_out[1040];
    assign layer1_out[1383] = ~(layer0_out[6050] ^ layer0_out[6051]);
    assign layer1_out[1384] = ~layer0_out[10];
    assign layer1_out[1385] = 1'b1;
    assign layer1_out[1386] = ~layer0_out[2530];
    assign layer1_out[1387] = layer0_out[5732] | layer0_out[5733];
    assign layer1_out[1388] = ~layer0_out[3548] | layer0_out[3549];
    assign layer1_out[1389] = ~layer0_out[5779];
    assign layer1_out[1390] = ~(layer0_out[7411] | layer0_out[7412]);
    assign layer1_out[1391] = ~layer0_out[7935];
    assign layer1_out[1392] = 1'b1;
    assign layer1_out[1393] = ~layer0_out[7061] | layer0_out[7060];
    assign layer1_out[1394] = ~layer0_out[6945];
    assign layer1_out[1395] = layer0_out[7279];
    assign layer1_out[1396] = layer0_out[7342] | layer0_out[7343];
    assign layer1_out[1397] = layer0_out[3920];
    assign layer1_out[1398] = layer0_out[1744];
    assign layer1_out[1399] = ~layer0_out[100] | layer0_out[101];
    assign layer1_out[1400] = layer0_out[808] & layer0_out[809];
    assign layer1_out[1401] = layer0_out[7601];
    assign layer1_out[1402] = ~layer0_out[4403];
    assign layer1_out[1403] = ~layer0_out[7469];
    assign layer1_out[1404] = ~layer0_out[638] | layer0_out[639];
    assign layer1_out[1405] = ~layer0_out[482];
    assign layer1_out[1406] = layer0_out[2046] ^ layer0_out[2047];
    assign layer1_out[1407] = ~layer0_out[6174];
    assign layer1_out[1408] = ~layer0_out[2753];
    assign layer1_out[1409] = ~(layer0_out[2484] ^ layer0_out[2485]);
    assign layer1_out[1410] = layer0_out[1102] & ~layer0_out[1103];
    assign layer1_out[1411] = ~layer0_out[6696];
    assign layer1_out[1412] = ~layer0_out[7093];
    assign layer1_out[1413] = ~layer0_out[7192] | layer0_out[7191];
    assign layer1_out[1414] = layer0_out[3495];
    assign layer1_out[1415] = ~layer0_out[1352];
    assign layer1_out[1416] = layer0_out[3022] & ~layer0_out[3023];
    assign layer1_out[1417] = 1'b0;
    assign layer1_out[1418] = 1'b1;
    assign layer1_out[1419] = ~layer0_out[4282];
    assign layer1_out[1420] = layer0_out[2376];
    assign layer1_out[1421] = layer0_out[80] & ~layer0_out[79];
    assign layer1_out[1422] = layer0_out[3866] & ~layer0_out[3865];
    assign layer1_out[1423] = layer0_out[7614] | layer0_out[7615];
    assign layer1_out[1424] = layer0_out[4117] & ~layer0_out[4116];
    assign layer1_out[1425] = layer0_out[6353];
    assign layer1_out[1426] = ~layer0_out[2908] | layer0_out[2909];
    assign layer1_out[1427] = ~layer0_out[6857];
    assign layer1_out[1428] = layer0_out[4836] & ~layer0_out[4835];
    assign layer1_out[1429] = layer0_out[1500] & layer0_out[1501];
    assign layer1_out[1430] = ~layer0_out[6035];
    assign layer1_out[1431] = ~(layer0_out[4096] & layer0_out[4097]);
    assign layer1_out[1432] = layer0_out[4111] & ~layer0_out[4112];
    assign layer1_out[1433] = layer0_out[449] & ~layer0_out[448];
    assign layer1_out[1434] = ~layer0_out[6200];
    assign layer1_out[1435] = ~layer0_out[4806] | layer0_out[4805];
    assign layer1_out[1436] = layer0_out[585];
    assign layer1_out[1437] = ~layer0_out[1920] | layer0_out[1919];
    assign layer1_out[1438] = ~layer0_out[5537];
    assign layer1_out[1439] = ~(layer0_out[2180] | layer0_out[2181]);
    assign layer1_out[1440] = layer0_out[1449] & ~layer0_out[1450];
    assign layer1_out[1441] = layer0_out[3059];
    assign layer1_out[1442] = layer0_out[5131];
    assign layer1_out[1443] = layer0_out[470];
    assign layer1_out[1444] = ~layer0_out[2309];
    assign layer1_out[1445] = layer0_out[6102];
    assign layer1_out[1446] = ~(layer0_out[718] | layer0_out[719]);
    assign layer1_out[1447] = ~(layer0_out[1940] ^ layer0_out[1941]);
    assign layer1_out[1448] = layer0_out[4662];
    assign layer1_out[1449] = layer0_out[2059] ^ layer0_out[2060];
    assign layer1_out[1450] = layer0_out[386] & ~layer0_out[385];
    assign layer1_out[1451] = ~layer0_out[7377];
    assign layer1_out[1452] = ~(layer0_out[1133] | layer0_out[1134]);
    assign layer1_out[1453] = layer0_out[995] & ~layer0_out[996];
    assign layer1_out[1454] = ~layer0_out[7064] | layer0_out[7065];
    assign layer1_out[1455] = ~layer0_out[6163];
    assign layer1_out[1456] = ~layer0_out[3648];
    assign layer1_out[1457] = ~layer0_out[5536];
    assign layer1_out[1458] = ~layer0_out[5415];
    assign layer1_out[1459] = ~(layer0_out[7537] | layer0_out[7538]);
    assign layer1_out[1460] = 1'b0;
    assign layer1_out[1461] = ~(layer0_out[4242] | layer0_out[4243]);
    assign layer1_out[1462] = layer0_out[2859] | layer0_out[2860];
    assign layer1_out[1463] = layer0_out[3486];
    assign layer1_out[1464] = layer0_out[3951];
    assign layer1_out[1465] = ~layer0_out[6227];
    assign layer1_out[1466] = ~layer0_out[5187];
    assign layer1_out[1467] = ~layer0_out[6369];
    assign layer1_out[1468] = layer0_out[1508];
    assign layer1_out[1469] = ~layer0_out[2196];
    assign layer1_out[1470] = 1'b0;
    assign layer1_out[1471] = layer0_out[6067];
    assign layer1_out[1472] = ~layer0_out[7869];
    assign layer1_out[1473] = layer0_out[3014];
    assign layer1_out[1474] = layer0_out[4478] & ~layer0_out[4479];
    assign layer1_out[1475] = ~layer0_out[7936];
    assign layer1_out[1476] = 1'b1;
    assign layer1_out[1477] = layer0_out[1121] ^ layer0_out[1122];
    assign layer1_out[1478] = layer0_out[1920];
    assign layer1_out[1479] = layer0_out[5503];
    assign layer1_out[1480] = layer0_out[7993];
    assign layer1_out[1481] = ~layer0_out[1034];
    assign layer1_out[1482] = layer0_out[7944] & ~layer0_out[7943];
    assign layer1_out[1483] = ~layer0_out[6621];
    assign layer1_out[1484] = layer0_out[1360] & ~layer0_out[1359];
    assign layer1_out[1485] = ~layer0_out[1643] | layer0_out[1642];
    assign layer1_out[1486] = layer0_out[1703] & ~layer0_out[1704];
    assign layer1_out[1487] = layer0_out[6340] & ~layer0_out[6339];
    assign layer1_out[1488] = layer0_out[85] & ~layer0_out[84];
    assign layer1_out[1489] = layer0_out[7380] | layer0_out[7381];
    assign layer1_out[1490] = layer0_out[4127];
    assign layer1_out[1491] = layer0_out[2154] & layer0_out[2155];
    assign layer1_out[1492] = layer0_out[2072] & ~layer0_out[2071];
    assign layer1_out[1493] = ~layer0_out[5897];
    assign layer1_out[1494] = layer0_out[6285] & ~layer0_out[6286];
    assign layer1_out[1495] = layer0_out[6159];
    assign layer1_out[1496] = layer0_out[6349] & layer0_out[6350];
    assign layer1_out[1497] = 1'b0;
    assign layer1_out[1498] = ~(layer0_out[2439] ^ layer0_out[2440]);
    assign layer1_out[1499] = ~layer0_out[2556];
    assign layer1_out[1500] = layer0_out[7779];
    assign layer1_out[1501] = ~layer0_out[7331];
    assign layer1_out[1502] = layer0_out[979] & layer0_out[980];
    assign layer1_out[1503] = layer0_out[6655] & ~layer0_out[6654];
    assign layer1_out[1504] = ~(layer0_out[4542] & layer0_out[4543]);
    assign layer1_out[1505] = layer0_out[1273];
    assign layer1_out[1506] = layer0_out[2041] | layer0_out[2042];
    assign layer1_out[1507] = layer0_out[2318] & ~layer0_out[2317];
    assign layer1_out[1508] = ~(layer0_out[2458] | layer0_out[2459]);
    assign layer1_out[1509] = layer0_out[5713];
    assign layer1_out[1510] = layer0_out[1435];
    assign layer1_out[1511] = layer0_out[4524] ^ layer0_out[4525];
    assign layer1_out[1512] = layer0_out[6333];
    assign layer1_out[1513] = ~layer0_out[3794] | layer0_out[3793];
    assign layer1_out[1514] = ~layer0_out[642] | layer0_out[643];
    assign layer1_out[1515] = layer0_out[6188] & ~layer0_out[6189];
    assign layer1_out[1516] = layer0_out[1582] & ~layer0_out[1581];
    assign layer1_out[1517] = ~layer0_out[1397];
    assign layer1_out[1518] = layer0_out[6623] & ~layer0_out[6624];
    assign layer1_out[1519] = 1'b1;
    assign layer1_out[1520] = ~(layer0_out[1305] & layer0_out[1306]);
    assign layer1_out[1521] = layer0_out[5308] | layer0_out[5309];
    assign layer1_out[1522] = 1'b0;
    assign layer1_out[1523] = layer0_out[1078];
    assign layer1_out[1524] = ~layer0_out[1831] | layer0_out[1832];
    assign layer1_out[1525] = layer0_out[1630] & ~layer0_out[1629];
    assign layer1_out[1526] = ~(layer0_out[3713] | layer0_out[3714]);
    assign layer1_out[1527] = layer0_out[858];
    assign layer1_out[1528] = ~layer0_out[2107] | layer0_out[2108];
    assign layer1_out[1529] = ~layer0_out[2057];
    assign layer1_out[1530] = layer0_out[3628] | layer0_out[3629];
    assign layer1_out[1531] = layer0_out[3867] & ~layer0_out[3868];
    assign layer1_out[1532] = layer0_out[982];
    assign layer1_out[1533] = layer0_out[825] | layer0_out[826];
    assign layer1_out[1534] = ~(layer0_out[3120] & layer0_out[3121]);
    assign layer1_out[1535] = layer0_out[2646] | layer0_out[2647];
    assign layer1_out[1536] = layer0_out[5339];
    assign layer1_out[1537] = ~(layer0_out[1639] ^ layer0_out[1640]);
    assign layer1_out[1538] = ~layer0_out[4482];
    assign layer1_out[1539] = ~layer0_out[2878];
    assign layer1_out[1540] = layer0_out[7041];
    assign layer1_out[1541] = layer0_out[5938] & layer0_out[5939];
    assign layer1_out[1542] = ~layer0_out[2040];
    assign layer1_out[1543] = layer0_out[492] & ~layer0_out[491];
    assign layer1_out[1544] = layer0_out[3802] & ~layer0_out[3801];
    assign layer1_out[1545] = layer0_out[3785];
    assign layer1_out[1546] = layer0_out[3747] & ~layer0_out[3748];
    assign layer1_out[1547] = ~layer0_out[3709];
    assign layer1_out[1548] = ~layer0_out[666] | layer0_out[665];
    assign layer1_out[1549] = layer0_out[6163] | layer0_out[6164];
    assign layer1_out[1550] = layer0_out[2628] ^ layer0_out[2629];
    assign layer1_out[1551] = layer0_out[2942] & layer0_out[2943];
    assign layer1_out[1552] = ~(layer0_out[3707] | layer0_out[3708]);
    assign layer1_out[1553] = ~layer0_out[6261] | layer0_out[6260];
    assign layer1_out[1554] = ~layer0_out[2117] | layer0_out[2116];
    assign layer1_out[1555] = ~layer0_out[7724] | layer0_out[7723];
    assign layer1_out[1556] = layer0_out[7619] & ~layer0_out[7618];
    assign layer1_out[1557] = layer0_out[6800] & ~layer0_out[6799];
    assign layer1_out[1558] = layer0_out[1366];
    assign layer1_out[1559] = ~(layer0_out[4548] ^ layer0_out[4549]);
    assign layer1_out[1560] = ~layer0_out[2332];
    assign layer1_out[1561] = ~layer0_out[609] | layer0_out[608];
    assign layer1_out[1562] = ~layer0_out[4531];
    assign layer1_out[1563] = layer0_out[5846] | layer0_out[5847];
    assign layer1_out[1564] = ~(layer0_out[3230] ^ layer0_out[3231]);
    assign layer1_out[1565] = layer0_out[4637] | layer0_out[4638];
    assign layer1_out[1566] = layer0_out[6493];
    assign layer1_out[1567] = layer0_out[2175] & ~layer0_out[2176];
    assign layer1_out[1568] = layer0_out[6618];
    assign layer1_out[1569] = layer0_out[7914] | layer0_out[7915];
    assign layer1_out[1570] = layer0_out[794] | layer0_out[795];
    assign layer1_out[1571] = layer0_out[2785];
    assign layer1_out[1572] = layer0_out[5108] & layer0_out[5109];
    assign layer1_out[1573] = layer0_out[6838];
    assign layer1_out[1574] = 1'b0;
    assign layer1_out[1575] = layer0_out[4391] & ~layer0_out[4390];
    assign layer1_out[1576] = layer0_out[7181];
    assign layer1_out[1577] = layer0_out[2540];
    assign layer1_out[1578] = layer0_out[4444] & ~layer0_out[4445];
    assign layer1_out[1579] = 1'b1;
    assign layer1_out[1580] = ~layer0_out[2927] | layer0_out[2926];
    assign layer1_out[1581] = ~(layer0_out[6176] & layer0_out[6177]);
    assign layer1_out[1582] = layer0_out[5023];
    assign layer1_out[1583] = layer0_out[7729] ^ layer0_out[7730];
    assign layer1_out[1584] = 1'b0;
    assign layer1_out[1585] = layer0_out[6588];
    assign layer1_out[1586] = layer0_out[151] | layer0_out[152];
    assign layer1_out[1587] = ~layer0_out[331];
    assign layer1_out[1588] = layer0_out[1489] & layer0_out[1490];
    assign layer1_out[1589] = 1'b0;
    assign layer1_out[1590] = ~layer0_out[4760];
    assign layer1_out[1591] = layer0_out[1345];
    assign layer1_out[1592] = layer0_out[3186] & ~layer0_out[3187];
    assign layer1_out[1593] = ~layer0_out[2419];
    assign layer1_out[1594] = ~(layer0_out[2310] & layer0_out[2311]);
    assign layer1_out[1595] = 1'b0;
    assign layer1_out[1596] = layer0_out[4750];
    assign layer1_out[1597] = ~(layer0_out[2031] | layer0_out[2032]);
    assign layer1_out[1598] = ~(layer0_out[6320] | layer0_out[6321]);
    assign layer1_out[1599] = ~(layer0_out[5642] | layer0_out[5643]);
    assign layer1_out[1600] = ~layer0_out[4693];
    assign layer1_out[1601] = layer0_out[6967];
    assign layer1_out[1602] = ~(layer0_out[7765] | layer0_out[7766]);
    assign layer1_out[1603] = layer0_out[66];
    assign layer1_out[1604] = ~(layer0_out[4047] ^ layer0_out[4048]);
    assign layer1_out[1605] = layer0_out[954] ^ layer0_out[955];
    assign layer1_out[1606] = ~layer0_out[1442];
    assign layer1_out[1607] = ~layer0_out[3689] | layer0_out[3688];
    assign layer1_out[1608] = layer0_out[5494] | layer0_out[5495];
    assign layer1_out[1609] = ~layer0_out[1116] | layer0_out[1117];
    assign layer1_out[1610] = layer0_out[3076] & ~layer0_out[3077];
    assign layer1_out[1611] = ~layer0_out[222];
    assign layer1_out[1612] = ~(layer0_out[7704] & layer0_out[7705]);
    assign layer1_out[1613] = ~layer0_out[2299];
    assign layer1_out[1614] = ~layer0_out[540];
    assign layer1_out[1615] = ~layer0_out[1136];
    assign layer1_out[1616] = ~layer0_out[765];
    assign layer1_out[1617] = ~layer0_out[2103] | layer0_out[2104];
    assign layer1_out[1618] = layer0_out[6923];
    assign layer1_out[1619] = ~(layer0_out[4512] | layer0_out[4513]);
    assign layer1_out[1620] = ~(layer0_out[3432] ^ layer0_out[3433]);
    assign layer1_out[1621] = ~layer0_out[5316];
    assign layer1_out[1622] = ~layer0_out[3413];
    assign layer1_out[1623] = layer0_out[3795] | layer0_out[3796];
    assign layer1_out[1624] = layer0_out[1215] ^ layer0_out[1216];
    assign layer1_out[1625] = layer0_out[7742];
    assign layer1_out[1626] = layer0_out[522];
    assign layer1_out[1627] = layer0_out[5198] & layer0_out[5199];
    assign layer1_out[1628] = layer0_out[2951] & ~layer0_out[2950];
    assign layer1_out[1629] = ~(layer0_out[6968] ^ layer0_out[6969]);
    assign layer1_out[1630] = 1'b0;
    assign layer1_out[1631] = ~layer0_out[1445];
    assign layer1_out[1632] = ~layer0_out[4496];
    assign layer1_out[1633] = ~layer0_out[1383] | layer0_out[1384];
    assign layer1_out[1634] = layer0_out[5885] & ~layer0_out[5884];
    assign layer1_out[1635] = layer0_out[5296] | layer0_out[5297];
    assign layer1_out[1636] = ~layer0_out[2821];
    assign layer1_out[1637] = ~layer0_out[6975];
    assign layer1_out[1638] = layer0_out[6355];
    assign layer1_out[1639] = ~layer0_out[6372] | layer0_out[6373];
    assign layer1_out[1640] = ~layer0_out[3993];
    assign layer1_out[1641] = layer0_out[690];
    assign layer1_out[1642] = layer0_out[5032];
    assign layer1_out[1643] = ~(layer0_out[5087] | layer0_out[5088]);
    assign layer1_out[1644] = layer0_out[6484] & ~layer0_out[6483];
    assign layer1_out[1645] = layer0_out[2424] & ~layer0_out[2423];
    assign layer1_out[1646] = ~(layer0_out[857] & layer0_out[858]);
    assign layer1_out[1647] = ~layer0_out[6249] | layer0_out[6250];
    assign layer1_out[1648] = ~layer0_out[2820];
    assign layer1_out[1649] = layer0_out[7732] & ~layer0_out[7733];
    assign layer1_out[1650] = ~layer0_out[4700] | layer0_out[4699];
    assign layer1_out[1651] = layer0_out[422] & ~layer0_out[421];
    assign layer1_out[1652] = ~(layer0_out[7967] ^ layer0_out[7968]);
    assign layer1_out[1653] = ~layer0_out[2456] | layer0_out[2455];
    assign layer1_out[1654] = ~layer0_out[7033];
    assign layer1_out[1655] = layer0_out[7650];
    assign layer1_out[1656] = ~(layer0_out[4726] | layer0_out[4727]);
    assign layer1_out[1657] = ~layer0_out[2698] | layer0_out[2697];
    assign layer1_out[1658] = layer0_out[7748];
    assign layer1_out[1659] = layer0_out[2799] & ~layer0_out[2798];
    assign layer1_out[1660] = layer0_out[4765];
    assign layer1_out[1661] = 1'b0;
    assign layer1_out[1662] = layer0_out[1967] & layer0_out[1968];
    assign layer1_out[1663] = layer0_out[6405];
    assign layer1_out[1664] = ~layer0_out[1895];
    assign layer1_out[1665] = ~(layer0_out[7472] | layer0_out[7473]);
    assign layer1_out[1666] = 1'b1;
    assign layer1_out[1667] = ~layer0_out[4553];
    assign layer1_out[1668] = layer0_out[4464];
    assign layer1_out[1669] = ~(layer0_out[4944] | layer0_out[4945]);
    assign layer1_out[1670] = layer0_out[4806] & layer0_out[4807];
    assign layer1_out[1671] = layer0_out[901];
    assign layer1_out[1672] = ~(layer0_out[2512] | layer0_out[2513]);
    assign layer1_out[1673] = layer0_out[1936] & ~layer0_out[1935];
    assign layer1_out[1674] = ~(layer0_out[4641] ^ layer0_out[4642]);
    assign layer1_out[1675] = layer0_out[2547] & ~layer0_out[2548];
    assign layer1_out[1676] = layer0_out[2718];
    assign layer1_out[1677] = layer0_out[3849] ^ layer0_out[3850];
    assign layer1_out[1678] = layer0_out[3812] | layer0_out[3813];
    assign layer1_out[1679] = ~(layer0_out[7305] | layer0_out[7306]);
    assign layer1_out[1680] = layer0_out[6448];
    assign layer1_out[1681] = ~(layer0_out[519] & layer0_out[520]);
    assign layer1_out[1682] = layer0_out[2503];
    assign layer1_out[1683] = layer0_out[5098];
    assign layer1_out[1684] = ~layer0_out[5189];
    assign layer1_out[1685] = layer0_out[4297] & layer0_out[4298];
    assign layer1_out[1686] = ~layer0_out[2887];
    assign layer1_out[1687] = layer0_out[943];
    assign layer1_out[1688] = layer0_out[6903] | layer0_out[6904];
    assign layer1_out[1689] = ~(layer0_out[2346] | layer0_out[2347]);
    assign layer1_out[1690] = ~(layer0_out[5222] | layer0_out[5223]);
    assign layer1_out[1691] = ~layer0_out[886] | layer0_out[887];
    assign layer1_out[1692] = ~layer0_out[7088];
    assign layer1_out[1693] = layer0_out[7573];
    assign layer1_out[1694] = ~(layer0_out[625] ^ layer0_out[626]);
    assign layer1_out[1695] = layer0_out[899] & layer0_out[900];
    assign layer1_out[1696] = layer0_out[4447] & ~layer0_out[4446];
    assign layer1_out[1697] = layer0_out[4612];
    assign layer1_out[1698] = layer0_out[4481];
    assign layer1_out[1699] = layer0_out[194] ^ layer0_out[195];
    assign layer1_out[1700] = 1'b0;
    assign layer1_out[1701] = 1'b1;
    assign layer1_out[1702] = layer0_out[3418] & ~layer0_out[3419];
    assign layer1_out[1703] = layer0_out[3255] | layer0_out[3256];
    assign layer1_out[1704] = layer0_out[376];
    assign layer1_out[1705] = 1'b0;
    assign layer1_out[1706] = 1'b0;
    assign layer1_out[1707] = layer0_out[1731] & ~layer0_out[1730];
    assign layer1_out[1708] = ~layer0_out[161];
    assign layer1_out[1709] = ~layer0_out[7407];
    assign layer1_out[1710] = 1'b1;
    assign layer1_out[1711] = ~(layer0_out[991] & layer0_out[992]);
    assign layer1_out[1712] = 1'b0;
    assign layer1_out[1713] = ~layer0_out[3434] | layer0_out[3435];
    assign layer1_out[1714] = ~layer0_out[1063];
    assign layer1_out[1715] = layer0_out[6849] & ~layer0_out[6848];
    assign layer1_out[1716] = ~layer0_out[6730] | layer0_out[6729];
    assign layer1_out[1717] = ~(layer0_out[7215] & layer0_out[7216]);
    assign layer1_out[1718] = ~(layer0_out[1762] | layer0_out[1763]);
    assign layer1_out[1719] = ~layer0_out[2616] | layer0_out[2615];
    assign layer1_out[1720] = ~(layer0_out[658] & layer0_out[659]);
    assign layer1_out[1721] = layer0_out[4534];
    assign layer1_out[1722] = layer0_out[3141] & layer0_out[3142];
    assign layer1_out[1723] = ~layer0_out[7679];
    assign layer1_out[1724] = ~layer0_out[6317] | layer0_out[6318];
    assign layer1_out[1725] = ~layer0_out[2672];
    assign layer1_out[1726] = ~layer0_out[2036] | layer0_out[2037];
    assign layer1_out[1727] = ~layer0_out[5417];
    assign layer1_out[1728] = ~layer0_out[3256] | layer0_out[3257];
    assign layer1_out[1729] = layer0_out[4665];
    assign layer1_out[1730] = 1'b1;
    assign layer1_out[1731] = ~(layer0_out[582] ^ layer0_out[583]);
    assign layer1_out[1732] = ~layer0_out[5084] | layer0_out[5083];
    assign layer1_out[1733] = layer0_out[7937];
    assign layer1_out[1734] = ~layer0_out[7208];
    assign layer1_out[1735] = ~layer0_out[3047] | layer0_out[3046];
    assign layer1_out[1736] = ~layer0_out[4743];
    assign layer1_out[1737] = ~layer0_out[4864];
    assign layer1_out[1738] = ~(layer0_out[680] | layer0_out[681]);
    assign layer1_out[1739] = ~(layer0_out[4272] & layer0_out[4273]);
    assign layer1_out[1740] = layer0_out[880] & layer0_out[881];
    assign layer1_out[1741] = 1'b0;
    assign layer1_out[1742] = layer0_out[3975] | layer0_out[3976];
    assign layer1_out[1743] = ~layer0_out[783] | layer0_out[782];
    assign layer1_out[1744] = layer0_out[6843] & layer0_out[6844];
    assign layer1_out[1745] = ~(layer0_out[489] | layer0_out[490]);
    assign layer1_out[1746] = layer0_out[987] | layer0_out[988];
    assign layer1_out[1747] = ~layer0_out[908];
    assign layer1_out[1748] = ~layer0_out[2727];
    assign layer1_out[1749] = 1'b0;
    assign layer1_out[1750] = ~layer0_out[3842];
    assign layer1_out[1751] = layer0_out[1063];
    assign layer1_out[1752] = ~(layer0_out[2112] ^ layer0_out[2113]);
    assign layer1_out[1753] = layer0_out[4902] & ~layer0_out[4901];
    assign layer1_out[1754] = layer0_out[4554];
    assign layer1_out[1755] = ~layer0_out[5829];
    assign layer1_out[1756] = ~(layer0_out[2829] & layer0_out[2830]);
    assign layer1_out[1757] = ~layer0_out[7075] | layer0_out[7076];
    assign layer1_out[1758] = ~(layer0_out[5146] & layer0_out[5147]);
    assign layer1_out[1759] = ~layer0_out[4304] | layer0_out[4303];
    assign layer1_out[1760] = layer0_out[6150];
    assign layer1_out[1761] = layer0_out[1810];
    assign layer1_out[1762] = ~layer0_out[5890];
    assign layer1_out[1763] = ~(layer0_out[6398] & layer0_out[6399]);
    assign layer1_out[1764] = layer0_out[4125] & ~layer0_out[4124];
    assign layer1_out[1765] = 1'b1;
    assign layer1_out[1766] = 1'b1;
    assign layer1_out[1767] = ~layer0_out[6228];
    assign layer1_out[1768] = layer0_out[5818] ^ layer0_out[5819];
    assign layer1_out[1769] = layer0_out[1537] | layer0_out[1538];
    assign layer1_out[1770] = layer0_out[5703] & layer0_out[5704];
    assign layer1_out[1771] = ~layer0_out[7340];
    assign layer1_out[1772] = ~layer0_out[4557];
    assign layer1_out[1773] = layer0_out[6896];
    assign layer1_out[1774] = ~layer0_out[5568];
    assign layer1_out[1775] = layer0_out[6361] & ~layer0_out[6360];
    assign layer1_out[1776] = ~(layer0_out[107] | layer0_out[108]);
    assign layer1_out[1777] = layer0_out[3261] | layer0_out[3262];
    assign layer1_out[1778] = layer0_out[3074] & ~layer0_out[3075];
    assign layer1_out[1779] = 1'b0;
    assign layer1_out[1780] = ~layer0_out[4868];
    assign layer1_out[1781] = 1'b0;
    assign layer1_out[1782] = layer0_out[2686] ^ layer0_out[2687];
    assign layer1_out[1783] = ~(layer0_out[5688] | layer0_out[5689]);
    assign layer1_out[1784] = layer0_out[132];
    assign layer1_out[1785] = layer0_out[6992];
    assign layer1_out[1786] = 1'b1;
    assign layer1_out[1787] = ~layer0_out[5727];
    assign layer1_out[1788] = ~layer0_out[7666];
    assign layer1_out[1789] = ~layer0_out[6429];
    assign layer1_out[1790] = layer0_out[1455] & layer0_out[1456];
    assign layer1_out[1791] = ~layer0_out[6465] | layer0_out[6466];
    assign layer1_out[1792] = ~layer0_out[2675] | layer0_out[2676];
    assign layer1_out[1793] = ~layer0_out[574];
    assign layer1_out[1794] = layer0_out[2335];
    assign layer1_out[1795] = layer0_out[5023] & layer0_out[5024];
    assign layer1_out[1796] = ~layer0_out[7388];
    assign layer1_out[1797] = layer0_out[7909];
    assign layer1_out[1798] = layer0_out[3807];
    assign layer1_out[1799] = 1'b1;
    assign layer1_out[1800] = ~layer0_out[4913];
    assign layer1_out[1801] = layer0_out[6507] & ~layer0_out[6506];
    assign layer1_out[1802] = layer0_out[5993] & ~layer0_out[5994];
    assign layer1_out[1803] = ~layer0_out[5587] | layer0_out[5586];
    assign layer1_out[1804] = ~(layer0_out[5667] & layer0_out[5668]);
    assign layer1_out[1805] = ~layer0_out[5521] | layer0_out[5520];
    assign layer1_out[1806] = ~(layer0_out[7445] & layer0_out[7446]);
    assign layer1_out[1807] = layer0_out[3892];
    assign layer1_out[1808] = layer0_out[6829];
    assign layer1_out[1809] = ~(layer0_out[3376] & layer0_out[3377]);
    assign layer1_out[1810] = ~layer0_out[2084];
    assign layer1_out[1811] = layer0_out[312];
    assign layer1_out[1812] = layer0_out[6853];
    assign layer1_out[1813] = ~(layer0_out[3857] ^ layer0_out[3858]);
    assign layer1_out[1814] = layer0_out[3767];
    assign layer1_out[1815] = layer0_out[3957] & layer0_out[3958];
    assign layer1_out[1816] = ~(layer0_out[2327] & layer0_out[2328]);
    assign layer1_out[1817] = 1'b1;
    assign layer1_out[1818] = layer0_out[1226] & ~layer0_out[1225];
    assign layer1_out[1819] = ~layer0_out[6040];
    assign layer1_out[1820] = ~(layer0_out[3909] & layer0_out[3910]);
    assign layer1_out[1821] = ~layer0_out[475];
    assign layer1_out[1822] = layer0_out[1142] ^ layer0_out[1143];
    assign layer1_out[1823] = ~layer0_out[1167];
    assign layer1_out[1824] = ~(layer0_out[3415] & layer0_out[3416]);
    assign layer1_out[1825] = ~layer0_out[2032] | layer0_out[2033];
    assign layer1_out[1826] = 1'b0;
    assign layer1_out[1827] = layer0_out[786] & ~layer0_out[785];
    assign layer1_out[1828] = ~(layer0_out[149] | layer0_out[150]);
    assign layer1_out[1829] = 1'b0;
    assign layer1_out[1830] = layer0_out[6074];
    assign layer1_out[1831] = ~(layer0_out[7763] | layer0_out[7764]);
    assign layer1_out[1832] = ~layer0_out[7914];
    assign layer1_out[1833] = 1'b0;
    assign layer1_out[1834] = layer0_out[7994] & ~layer0_out[7995];
    assign layer1_out[1835] = ~layer0_out[1112];
    assign layer1_out[1836] = layer0_out[902] & ~layer0_out[903];
    assign layer1_out[1837] = ~layer0_out[6961];
    assign layer1_out[1838] = layer0_out[2809];
    assign layer1_out[1839] = layer0_out[4098];
    assign layer1_out[1840] = ~layer0_out[4402];
    assign layer1_out[1841] = layer0_out[2882];
    assign layer1_out[1842] = layer0_out[6258];
    assign layer1_out[1843] = layer0_out[4080];
    assign layer1_out[1844] = ~(layer0_out[7069] & layer0_out[7070]);
    assign layer1_out[1845] = ~(layer0_out[5558] & layer0_out[5559]);
    assign layer1_out[1846] = ~layer0_out[3833];
    assign layer1_out[1847] = layer0_out[3815];
    assign layer1_out[1848] = ~(layer0_out[6536] & layer0_out[6537]);
    assign layer1_out[1849] = ~(layer0_out[5866] ^ layer0_out[5867]);
    assign layer1_out[1850] = 1'b1;
    assign layer1_out[1851] = layer0_out[7483] ^ layer0_out[7484];
    assign layer1_out[1852] = layer0_out[6602];
    assign layer1_out[1853] = layer0_out[1881] ^ layer0_out[1882];
    assign layer1_out[1854] = ~layer0_out[6122] | layer0_out[6123];
    assign layer1_out[1855] = ~layer0_out[6019];
    assign layer1_out[1856] = ~(layer0_out[277] | layer0_out[278]);
    assign layer1_out[1857] = ~layer0_out[7701] | layer0_out[7702];
    assign layer1_out[1858] = ~layer0_out[853];
    assign layer1_out[1859] = layer0_out[4017];
    assign layer1_out[1860] = ~(layer0_out[162] | layer0_out[163]);
    assign layer1_out[1861] = layer0_out[586];
    assign layer1_out[1862] = ~(layer0_out[2255] & layer0_out[2256]);
    assign layer1_out[1863] = ~(layer0_out[7858] | layer0_out[7859]);
    assign layer1_out[1864] = layer0_out[4488] & layer0_out[4489];
    assign layer1_out[1865] = ~layer0_out[1728];
    assign layer1_out[1866] = layer0_out[7882];
    assign layer1_out[1867] = ~(layer0_out[7046] ^ layer0_out[7047]);
    assign layer1_out[1868] = ~layer0_out[5809];
    assign layer1_out[1869] = layer0_out[6601] | layer0_out[6602];
    assign layer1_out[1870] = ~layer0_out[4041] | layer0_out[4042];
    assign layer1_out[1871] = layer0_out[495] & layer0_out[496];
    assign layer1_out[1872] = ~layer0_out[5841];
    assign layer1_out[1873] = ~(layer0_out[4397] | layer0_out[4398]);
    assign layer1_out[1874] = ~layer0_out[2496] | layer0_out[2495];
    assign layer1_out[1875] = ~(layer0_out[2778] | layer0_out[2779]);
    assign layer1_out[1876] = ~layer0_out[7026] | layer0_out[7025];
    assign layer1_out[1877] = layer0_out[6575] | layer0_out[6576];
    assign layer1_out[1878] = layer0_out[2428] ^ layer0_out[2429];
    assign layer1_out[1879] = ~(layer0_out[392] ^ layer0_out[393]);
    assign layer1_out[1880] = layer0_out[1668] & ~layer0_out[1669];
    assign layer1_out[1881] = ~layer0_out[3878] | layer0_out[3879];
    assign layer1_out[1882] = layer0_out[4104] & layer0_out[4105];
    assign layer1_out[1883] = layer0_out[1607] | layer0_out[1608];
    assign layer1_out[1884] = layer0_out[4597] ^ layer0_out[4598];
    assign layer1_out[1885] = ~layer0_out[669] | layer0_out[668];
    assign layer1_out[1886] = ~layer0_out[1151] | layer0_out[1152];
    assign layer1_out[1887] = layer0_out[1602] & ~layer0_out[1603];
    assign layer1_out[1888] = layer0_out[2202];
    assign layer1_out[1889] = 1'b1;
    assign layer1_out[1890] = 1'b0;
    assign layer1_out[1891] = layer0_out[2415];
    assign layer1_out[1892] = ~layer0_out[1464];
    assign layer1_out[1893] = ~(layer0_out[5701] | layer0_out[5702]);
    assign layer1_out[1894] = layer0_out[6827];
    assign layer1_out[1895] = ~(layer0_out[85] | layer0_out[86]);
    assign layer1_out[1896] = ~(layer0_out[6897] & layer0_out[6898]);
    assign layer1_out[1897] = ~layer0_out[2058] | layer0_out[2057];
    assign layer1_out[1898] = ~(layer0_out[6779] | layer0_out[6780]);
    assign layer1_out[1899] = layer0_out[5036] & layer0_out[5037];
    assign layer1_out[1900] = ~layer0_out[5304];
    assign layer1_out[1901] = ~layer0_out[1362];
    assign layer1_out[1902] = layer0_out[815] & ~layer0_out[814];
    assign layer1_out[1903] = layer0_out[1615];
    assign layer1_out[1904] = ~(layer0_out[1862] ^ layer0_out[1863]);
    assign layer1_out[1905] = layer0_out[1514] & layer0_out[1515];
    assign layer1_out[1906] = ~layer0_out[172];
    assign layer1_out[1907] = ~layer0_out[286] | layer0_out[285];
    assign layer1_out[1908] = layer0_out[514] & ~layer0_out[515];
    assign layer1_out[1909] = ~layer0_out[4876] | layer0_out[4877];
    assign layer1_out[1910] = layer0_out[6995] & ~layer0_out[6996];
    assign layer1_out[1911] = ~layer0_out[7801] | layer0_out[7800];
    assign layer1_out[1912] = layer0_out[5303];
    assign layer1_out[1913] = layer0_out[163] & layer0_out[164];
    assign layer1_out[1914] = layer0_out[484] & ~layer0_out[485];
    assign layer1_out[1915] = ~(layer0_out[434] | layer0_out[435]);
    assign layer1_out[1916] = 1'b1;
    assign layer1_out[1917] = ~layer0_out[1252];
    assign layer1_out[1918] = layer0_out[504] & layer0_out[505];
    assign layer1_out[1919] = ~layer0_out[3606];
    assign layer1_out[1920] = ~(layer0_out[7590] & layer0_out[7591]);
    assign layer1_out[1921] = layer0_out[6771];
    assign layer1_out[1922] = 1'b0;
    assign layer1_out[1923] = layer0_out[5173] | layer0_out[5174];
    assign layer1_out[1924] = ~layer0_out[2865] | layer0_out[2864];
    assign layer1_out[1925] = 1'b0;
    assign layer1_out[1926] = ~layer0_out[7832];
    assign layer1_out[1927] = layer0_out[4718];
    assign layer1_out[1928] = 1'b1;
    assign layer1_out[1929] = layer0_out[5920];
    assign layer1_out[1930] = ~layer0_out[5555] | layer0_out[5554];
    assign layer1_out[1931] = ~layer0_out[619];
    assign layer1_out[1932] = ~layer0_out[2324] | layer0_out[2323];
    assign layer1_out[1933] = ~(layer0_out[1795] | layer0_out[1796]);
    assign layer1_out[1934] = ~(layer0_out[6629] & layer0_out[6630]);
    assign layer1_out[1935] = layer0_out[81];
    assign layer1_out[1936] = 1'b1;
    assign layer1_out[1937] = layer0_out[6236] & ~layer0_out[6235];
    assign layer1_out[1938] = layer0_out[2418] | layer0_out[2419];
    assign layer1_out[1939] = ~layer0_out[3246];
    assign layer1_out[1940] = layer0_out[6794];
    assign layer1_out[1941] = ~layer0_out[7694] | layer0_out[7695];
    assign layer1_out[1942] = ~layer0_out[410];
    assign layer1_out[1943] = layer0_out[4625];
    assign layer1_out[1944] = layer0_out[2858] & layer0_out[2859];
    assign layer1_out[1945] = 1'b1;
    assign layer1_out[1946] = layer0_out[7558] & ~layer0_out[7557];
    assign layer1_out[1947] = ~layer0_out[6136] | layer0_out[6135];
    assign layer1_out[1948] = layer0_out[5495];
    assign layer1_out[1949] = layer0_out[3144] | layer0_out[3145];
    assign layer1_out[1950] = ~layer0_out[2552] | layer0_out[2553];
    assign layer1_out[1951] = layer0_out[4323] & ~layer0_out[4322];
    assign layer1_out[1952] = layer0_out[4980] & ~layer0_out[4981];
    assign layer1_out[1953] = ~(layer0_out[6564] | layer0_out[6565]);
    assign layer1_out[1954] = layer0_out[4722];
    assign layer1_out[1955] = ~layer0_out[2703];
    assign layer1_out[1956] = ~layer0_out[629] | layer0_out[628];
    assign layer1_out[1957] = ~(layer0_out[7648] & layer0_out[7649]);
    assign layer1_out[1958] = ~(layer0_out[4513] ^ layer0_out[4514]);
    assign layer1_out[1959] = layer0_out[3724] & ~layer0_out[3723];
    assign layer1_out[1960] = layer0_out[7160] | layer0_out[7161];
    assign layer1_out[1961] = ~(layer0_out[1861] & layer0_out[1862]);
    assign layer1_out[1962] = layer0_out[4543];
    assign layer1_out[1963] = layer0_out[5565];
    assign layer1_out[1964] = ~layer0_out[6656];
    assign layer1_out[1965] = ~layer0_out[3993];
    assign layer1_out[1966] = ~layer0_out[993];
    assign layer1_out[1967] = layer0_out[4937];
    assign layer1_out[1968] = ~(layer0_out[245] | layer0_out[246]);
    assign layer1_out[1969] = ~(layer0_out[1870] ^ layer0_out[1871]);
    assign layer1_out[1970] = layer0_out[6297];
    assign layer1_out[1971] = ~(layer0_out[2449] & layer0_out[2450]);
    assign layer1_out[1972] = ~layer0_out[1510] | layer0_out[1511];
    assign layer1_out[1973] = ~(layer0_out[1246] ^ layer0_out[1247]);
    assign layer1_out[1974] = layer0_out[5040] | layer0_out[5041];
    assign layer1_out[1975] = ~layer0_out[1391] | layer0_out[1392];
    assign layer1_out[1976] = layer0_out[3904];
    assign layer1_out[1977] = ~(layer0_out[4462] | layer0_out[4463]);
    assign layer1_out[1978] = layer0_out[2870] & ~layer0_out[2871];
    assign layer1_out[1979] = layer0_out[7481] & ~layer0_out[7482];
    assign layer1_out[1980] = layer0_out[3699];
    assign layer1_out[1981] = ~layer0_out[4241];
    assign layer1_out[1982] = layer0_out[6391] | layer0_out[6392];
    assign layer1_out[1983] = ~layer0_out[743];
    assign layer1_out[1984] = layer0_out[4493];
    assign layer1_out[1985] = ~(layer0_out[1127] ^ layer0_out[1128]);
    assign layer1_out[1986] = layer0_out[6809];
    assign layer1_out[1987] = layer0_out[2889];
    assign layer1_out[1988] = layer0_out[3421];
    assign layer1_out[1989] = ~layer0_out[7716] | layer0_out[7717];
    assign layer1_out[1990] = ~(layer0_out[6229] & layer0_out[6230]);
    assign layer1_out[1991] = ~layer0_out[7097];
    assign layer1_out[1992] = ~layer0_out[3021] | layer0_out[3022];
    assign layer1_out[1993] = ~layer0_out[2922];
    assign layer1_out[1994] = layer0_out[4420] ^ layer0_out[4421];
    assign layer1_out[1995] = 1'b0;
    assign layer1_out[1996] = ~layer0_out[1053] | layer0_out[1052];
    assign layer1_out[1997] = layer0_out[6100];
    assign layer1_out[1998] = ~layer0_out[7487];
    assign layer1_out[1999] = layer0_out[397] | layer0_out[398];
    assign layer1_out[2000] = ~(layer0_out[3131] | layer0_out[3132]);
    assign layer1_out[2001] = ~(layer0_out[1917] ^ layer0_out[1918]);
    assign layer1_out[2002] = ~(layer0_out[2534] & layer0_out[2535]);
    assign layer1_out[2003] = layer0_out[5177] & ~layer0_out[5176];
    assign layer1_out[2004] = ~layer0_out[7847] | layer0_out[7846];
    assign layer1_out[2005] = layer0_out[7410];
    assign layer1_out[2006] = layer0_out[749];
    assign layer1_out[2007] = ~layer0_out[4049] | layer0_out[4048];
    assign layer1_out[2008] = layer0_out[3111];
    assign layer1_out[2009] = ~(layer0_out[7314] & layer0_out[7315]);
    assign layer1_out[2010] = layer0_out[3539];
    assign layer1_out[2011] = layer0_out[4422] & ~layer0_out[4423];
    assign layer1_out[2012] = ~(layer0_out[4873] | layer0_out[4874]);
    assign layer1_out[2013] = 1'b0;
    assign layer1_out[2014] = layer0_out[7300];
    assign layer1_out[2015] = ~layer0_out[7294];
    assign layer1_out[2016] = layer0_out[1949] | layer0_out[1950];
    assign layer1_out[2017] = layer0_out[6585] ^ layer0_out[6586];
    assign layer1_out[2018] = ~(layer0_out[1248] & layer0_out[1249]);
    assign layer1_out[2019] = ~layer0_out[1380];
    assign layer1_out[2020] = layer0_out[5713] & ~layer0_out[5714];
    assign layer1_out[2021] = layer0_out[1853] | layer0_out[1854];
    assign layer1_out[2022] = 1'b1;
    assign layer1_out[2023] = layer0_out[7784] ^ layer0_out[7785];
    assign layer1_out[2024] = ~layer0_out[4493];
    assign layer1_out[2025] = ~layer0_out[3177];
    assign layer1_out[2026] = ~(layer0_out[4545] & layer0_out[4546]);
    assign layer1_out[2027] = layer0_out[664];
    assign layer1_out[2028] = ~layer0_out[3400] | layer0_out[3399];
    assign layer1_out[2029] = layer0_out[5619] & ~layer0_out[5618];
    assign layer1_out[2030] = layer0_out[4090] & ~layer0_out[4091];
    assign layer1_out[2031] = layer0_out[5791];
    assign layer1_out[2032] = ~layer0_out[4546] | layer0_out[4547];
    assign layer1_out[2033] = layer0_out[4691];
    assign layer1_out[2034] = layer0_out[2710];
    assign layer1_out[2035] = layer0_out[3998] & ~layer0_out[3997];
    assign layer1_out[2036] = ~layer0_out[6401];
    assign layer1_out[2037] = layer0_out[2006];
    assign layer1_out[2038] = ~(layer0_out[6479] & layer0_out[6480]);
    assign layer1_out[2039] = layer0_out[6485] | layer0_out[6486];
    assign layer1_out[2040] = ~(layer0_out[3617] | layer0_out[3618]);
    assign layer1_out[2041] = layer0_out[6577];
    assign layer1_out[2042] = ~(layer0_out[7084] ^ layer0_out[7085]);
    assign layer1_out[2043] = ~layer0_out[5772] | layer0_out[5773];
    assign layer1_out[2044] = layer0_out[6069];
    assign layer1_out[2045] = ~layer0_out[2178] | layer0_out[2179];
    assign layer1_out[2046] = ~layer0_out[5449];
    assign layer1_out[2047] = 1'b0;
    assign layer1_out[2048] = ~(layer0_out[5762] & layer0_out[5763]);
    assign layer1_out[2049] = ~layer0_out[5115];
    assign layer1_out[2050] = layer0_out[7808] & layer0_out[7809];
    assign layer1_out[2051] = layer0_out[4340];
    assign layer1_out[2052] = layer0_out[7391] & ~layer0_out[7390];
    assign layer1_out[2053] = layer0_out[7413];
    assign layer1_out[2054] = 1'b0;
    assign layer1_out[2055] = ~layer0_out[2653] | layer0_out[2654];
    assign layer1_out[2056] = layer0_out[7835];
    assign layer1_out[2057] = 1'b1;
    assign layer1_out[2058] = ~layer0_out[6111] | layer0_out[6112];
    assign layer1_out[2059] = layer0_out[5192];
    assign layer1_out[2060] = layer0_out[1123] & layer0_out[1124];
    assign layer1_out[2061] = ~layer0_out[6809];
    assign layer1_out[2062] = layer0_out[7190];
    assign layer1_out[2063] = ~layer0_out[280] | layer0_out[281];
    assign layer1_out[2064] = ~layer0_out[5135] | layer0_out[5136];
    assign layer1_out[2065] = 1'b1;
    assign layer1_out[2066] = ~layer0_out[7503];
    assign layer1_out[2067] = layer0_out[3009] | layer0_out[3010];
    assign layer1_out[2068] = layer0_out[1520] ^ layer0_out[1521];
    assign layer1_out[2069] = ~layer0_out[5333] | layer0_out[5334];
    assign layer1_out[2070] = layer0_out[7304];
    assign layer1_out[2071] = layer0_out[6964] & layer0_out[6965];
    assign layer1_out[2072] = ~layer0_out[7356];
    assign layer1_out[2073] = layer0_out[5624] & ~layer0_out[5623];
    assign layer1_out[2074] = layer0_out[3558];
    assign layer1_out[2075] = ~layer0_out[2023];
    assign layer1_out[2076] = ~layer0_out[4739];
    assign layer1_out[2077] = ~(layer0_out[3807] & layer0_out[3808]);
    assign layer1_out[2078] = layer0_out[7916] & ~layer0_out[7915];
    assign layer1_out[2079] = ~layer0_out[4800];
    assign layer1_out[2080] = layer0_out[7155] & layer0_out[7156];
    assign layer1_out[2081] = 1'b0;
    assign layer1_out[2082] = ~(layer0_out[490] ^ layer0_out[491]);
    assign layer1_out[2083] = layer0_out[3503];
    assign layer1_out[2084] = layer0_out[3779] & layer0_out[3780];
    assign layer1_out[2085] = layer0_out[3485] & ~layer0_out[3484];
    assign layer1_out[2086] = ~(layer0_out[3904] | layer0_out[3905]);
    assign layer1_out[2087] = layer0_out[2565] | layer0_out[2566];
    assign layer1_out[2088] = ~layer0_out[2130];
    assign layer1_out[2089] = ~(layer0_out[4984] | layer0_out[4985]);
    assign layer1_out[2090] = ~layer0_out[3739] | layer0_out[3740];
    assign layer1_out[2091] = layer0_out[5003] ^ layer0_out[5004];
    assign layer1_out[2092] = ~(layer0_out[7582] & layer0_out[7583]);
    assign layer1_out[2093] = ~layer0_out[7539] | layer0_out[7538];
    assign layer1_out[2094] = layer0_out[1372] | layer0_out[1373];
    assign layer1_out[2095] = ~(layer0_out[7428] | layer0_out[7429]);
    assign layer1_out[2096] = layer0_out[1022] ^ layer0_out[1023];
    assign layer1_out[2097] = layer0_out[3075] | layer0_out[3076];
    assign layer1_out[2098] = layer0_out[1365];
    assign layer1_out[2099] = layer0_out[7642];
    assign layer1_out[2100] = ~layer0_out[7462];
    assign layer1_out[2101] = layer0_out[2602] & ~layer0_out[2603];
    assign layer1_out[2102] = layer0_out[6777] & layer0_out[6778];
    assign layer1_out[2103] = ~(layer0_out[7379] | layer0_out[7380]);
    assign layer1_out[2104] = ~layer0_out[7028] | layer0_out[7027];
    assign layer1_out[2105] = ~(layer0_out[5484] ^ layer0_out[5485]);
    assign layer1_out[2106] = ~layer0_out[3365];
    assign layer1_out[2107] = ~(layer0_out[5631] ^ layer0_out[5632]);
    assign layer1_out[2108] = ~(layer0_out[2824] | layer0_out[2825]);
    assign layer1_out[2109] = ~(layer0_out[4751] & layer0_out[4752]);
    assign layer1_out[2110] = ~layer0_out[5152];
    assign layer1_out[2111] = ~layer0_out[4931];
    assign layer1_out[2112] = layer0_out[6008] & layer0_out[6009];
    assign layer1_out[2113] = ~layer0_out[1451] | layer0_out[1452];
    assign layer1_out[2114] = 1'b1;
    assign layer1_out[2115] = 1'b1;
    assign layer1_out[2116] = layer0_out[3348] ^ layer0_out[3349];
    assign layer1_out[2117] = ~layer0_out[2739] | layer0_out[2738];
    assign layer1_out[2118] = layer0_out[3902] & ~layer0_out[3903];
    assign layer1_out[2119] = ~layer0_out[5835];
    assign layer1_out[2120] = layer0_out[2199] | layer0_out[2200];
    assign layer1_out[2121] = layer0_out[669] & layer0_out[670];
    assign layer1_out[2122] = layer0_out[2569] & layer0_out[2570];
    assign layer1_out[2123] = ~(layer0_out[5418] | layer0_out[5419]);
    assign layer1_out[2124] = layer0_out[7625] & ~layer0_out[7626];
    assign layer1_out[2125] = ~layer0_out[673] | layer0_out[674];
    assign layer1_out[2126] = layer0_out[5377];
    assign layer1_out[2127] = layer0_out[2536];
    assign layer1_out[2128] = ~(layer0_out[3020] & layer0_out[3021]);
    assign layer1_out[2129] = ~layer0_out[6804];
    assign layer1_out[2130] = ~layer0_out[5074] | layer0_out[5075];
    assign layer1_out[2131] = layer0_out[5474] & ~layer0_out[5475];
    assign layer1_out[2132] = ~layer0_out[67];
    assign layer1_out[2133] = layer0_out[5596] & layer0_out[5597];
    assign layer1_out[2134] = 1'b0;
    assign layer1_out[2135] = layer0_out[6524] | layer0_out[6525];
    assign layer1_out[2136] = ~layer0_out[6110];
    assign layer1_out[2137] = ~layer0_out[5626];
    assign layer1_out[2138] = layer0_out[6033];
    assign layer1_out[2139] = ~layer0_out[5933];
    assign layer1_out[2140] = layer0_out[394] & layer0_out[395];
    assign layer1_out[2141] = ~(layer0_out[4181] | layer0_out[4182]);
    assign layer1_out[2142] = ~(layer0_out[728] & layer0_out[729]);
    assign layer1_out[2143] = layer0_out[3398] & ~layer0_out[3397];
    assign layer1_out[2144] = layer0_out[7965] ^ layer0_out[7966];
    assign layer1_out[2145] = layer0_out[4875] & layer0_out[4876];
    assign layer1_out[2146] = ~layer0_out[3229] | layer0_out[3228];
    assign layer1_out[2147] = ~layer0_out[6883];
    assign layer1_out[2148] = ~(layer0_out[224] & layer0_out[225]);
    assign layer1_out[2149] = 1'b1;
    assign layer1_out[2150] = layer0_out[6816] & layer0_out[6817];
    assign layer1_out[2151] = ~layer0_out[5629];
    assign layer1_out[2152] = ~layer0_out[7978];
    assign layer1_out[2153] = ~(layer0_out[4107] | layer0_out[4108]);
    assign layer1_out[2154] = 1'b1;
    assign layer1_out[2155] = layer0_out[3854] & layer0_out[3855];
    assign layer1_out[2156] = layer0_out[3603];
    assign layer1_out[2157] = 1'b1;
    assign layer1_out[2158] = layer0_out[5793] | layer0_out[5794];
    assign layer1_out[2159] = ~(layer0_out[3868] | layer0_out[3869]);
    assign layer1_out[2160] = ~(layer0_out[3926] & layer0_out[3927]);
    assign layer1_out[2161] = layer0_out[2307] & layer0_out[2308];
    assign layer1_out[2162] = layer0_out[7036] & ~layer0_out[7037];
    assign layer1_out[2163] = layer0_out[7382] | layer0_out[7383];
    assign layer1_out[2164] = layer0_out[4840] ^ layer0_out[4841];
    assign layer1_out[2165] = layer0_out[1249];
    assign layer1_out[2166] = layer0_out[2265] & ~layer0_out[2266];
    assign layer1_out[2167] = layer0_out[2058];
    assign layer1_out[2168] = layer0_out[1913];
    assign layer1_out[2169] = layer0_out[2995];
    assign layer1_out[2170] = layer0_out[1997] | layer0_out[1998];
    assign layer1_out[2171] = layer0_out[5413] & ~layer0_out[5414];
    assign layer1_out[2172] = ~(layer0_out[2925] & layer0_out[2926]);
    assign layer1_out[2173] = layer0_out[2368] & ~layer0_out[2369];
    assign layer1_out[2174] = ~layer0_out[7426] | layer0_out[7425];
    assign layer1_out[2175] = ~layer0_out[5546];
    assign layer1_out[2176] = 1'b1;
    assign layer1_out[2177] = layer0_out[215] & ~layer0_out[214];
    assign layer1_out[2178] = ~layer0_out[2705];
    assign layer1_out[2179] = layer0_out[6020] | layer0_out[6021];
    assign layer1_out[2180] = ~layer0_out[4404] | layer0_out[4405];
    assign layer1_out[2181] = ~layer0_out[562] | layer0_out[563];
    assign layer1_out[2182] = ~(layer0_out[4458] | layer0_out[4459]);
    assign layer1_out[2183] = layer0_out[5840] & ~layer0_out[5839];
    assign layer1_out[2184] = layer0_out[3114];
    assign layer1_out[2185] = ~(layer0_out[567] | layer0_out[568]);
    assign layer1_out[2186] = ~layer0_out[7021];
    assign layer1_out[2187] = ~layer0_out[7227] | layer0_out[7226];
    assign layer1_out[2188] = layer0_out[5944] & ~layer0_out[5945];
    assign layer1_out[2189] = ~layer0_out[6328];
    assign layer1_out[2190] = ~layer0_out[1830];
    assign layer1_out[2191] = ~layer0_out[1386] | layer0_out[1385];
    assign layer1_out[2192] = 1'b0;
    assign layer1_out[2193] = layer0_out[3101] | layer0_out[3102];
    assign layer1_out[2194] = layer0_out[1962] & layer0_out[1963];
    assign layer1_out[2195] = ~layer0_out[5633];
    assign layer1_out[2196] = ~layer0_out[4003];
    assign layer1_out[2197] = layer0_out[4200] & ~layer0_out[4199];
    assign layer1_out[2198] = layer0_out[5230] & layer0_out[5231];
    assign layer1_out[2199] = layer0_out[6393] | layer0_out[6394];
    assign layer1_out[2200] = ~layer0_out[4713] | layer0_out[4712];
    assign layer1_out[2201] = ~layer0_out[5546] | layer0_out[5547];
    assign layer1_out[2202] = ~(layer0_out[4040] | layer0_out[4041]);
    assign layer1_out[2203] = ~layer0_out[2684];
    assign layer1_out[2204] = layer0_out[3197] & ~layer0_out[3198];
    assign layer1_out[2205] = layer0_out[93] & ~layer0_out[92];
    assign layer1_out[2206] = layer0_out[7362];
    assign layer1_out[2207] = ~layer0_out[4174];
    assign layer1_out[2208] = layer0_out[622] & ~layer0_out[621];
    assign layer1_out[2209] = layer0_out[3351] & ~layer0_out[3350];
    assign layer1_out[2210] = ~layer0_out[6177];
    assign layer1_out[2211] = layer0_out[3944] ^ layer0_out[3945];
    assign layer1_out[2212] = layer0_out[4000] | layer0_out[4001];
    assign layer1_out[2213] = layer0_out[1461] & ~layer0_out[1460];
    assign layer1_out[2214] = layer0_out[4672] & ~layer0_out[4671];
    assign layer1_out[2215] = ~layer0_out[3644];
    assign layer1_out[2216] = layer0_out[1210];
    assign layer1_out[2217] = ~layer0_out[7604];
    assign layer1_out[2218] = ~layer0_out[4635];
    assign layer1_out[2219] = layer0_out[6832] & ~layer0_out[6831];
    assign layer1_out[2220] = ~layer0_out[7159];
    assign layer1_out[2221] = ~layer0_out[4145];
    assign layer1_out[2222] = ~layer0_out[3658];
    assign layer1_out[2223] = 1'b0;
    assign layer1_out[2224] = ~(layer0_out[3922] | layer0_out[3923]);
    assign layer1_out[2225] = ~layer0_out[7851] | layer0_out[7850];
    assign layer1_out[2226] = ~layer0_out[5905];
    assign layer1_out[2227] = 1'b0;
    assign layer1_out[2228] = ~(layer0_out[5216] ^ layer0_out[5217]);
    assign layer1_out[2229] = ~layer0_out[5866];
    assign layer1_out[2230] = ~(layer0_out[7397] & layer0_out[7398]);
    assign layer1_out[2231] = layer0_out[2093] & ~layer0_out[2094];
    assign layer1_out[2232] = ~layer0_out[4431];
    assign layer1_out[2233] = layer0_out[1843] & ~layer0_out[1844];
    assign layer1_out[2234] = layer0_out[1760] | layer0_out[1761];
    assign layer1_out[2235] = layer0_out[7302] & ~layer0_out[7303];
    assign layer1_out[2236] = layer0_out[2087] ^ layer0_out[2088];
    assign layer1_out[2237] = layer0_out[5305];
    assign layer1_out[2238] = layer0_out[4259] & ~layer0_out[4258];
    assign layer1_out[2239] = ~layer0_out[2677] | layer0_out[2676];
    assign layer1_out[2240] = ~(layer0_out[5268] ^ layer0_out[5269]);
    assign layer1_out[2241] = ~layer0_out[1183] | layer0_out[1182];
    assign layer1_out[2242] = ~layer0_out[7231];
    assign layer1_out[2243] = ~(layer0_out[4565] | layer0_out[4566]);
    assign layer1_out[2244] = layer0_out[7219] | layer0_out[7220];
    assign layer1_out[2245] = layer0_out[4053];
    assign layer1_out[2246] = 1'b1;
    assign layer1_out[2247] = ~layer0_out[5868] | layer0_out[5869];
    assign layer1_out[2248] = layer0_out[1985] & layer0_out[1986];
    assign layer1_out[2249] = layer0_out[3650] ^ layer0_out[3651];
    assign layer1_out[2250] = ~layer0_out[2452];
    assign layer1_out[2251] = layer0_out[7040];
    assign layer1_out[2252] = ~layer0_out[3569];
    assign layer1_out[2253] = layer0_out[472] & ~layer0_out[471];
    assign layer1_out[2254] = ~layer0_out[516];
    assign layer1_out[2255] = 1'b1;
    assign layer1_out[2256] = layer0_out[6775] & ~layer0_out[6776];
    assign layer1_out[2257] = layer0_out[165] | layer0_out[166];
    assign layer1_out[2258] = layer0_out[1909] | layer0_out[1910];
    assign layer1_out[2259] = ~layer0_out[5753];
    assign layer1_out[2260] = layer0_out[5553];
    assign layer1_out[2261] = layer0_out[2194] ^ layer0_out[2195];
    assign layer1_out[2262] = ~layer0_out[5178];
    assign layer1_out[2263] = layer0_out[2958];
    assign layer1_out[2264] = ~layer0_out[3582] | layer0_out[3583];
    assign layer1_out[2265] = ~(layer0_out[1901] & layer0_out[1902]);
    assign layer1_out[2266] = layer0_out[7020];
    assign layer1_out[2267] = layer0_out[7311];
    assign layer1_out[2268] = layer0_out[3615];
    assign layer1_out[2269] = layer0_out[4169] & layer0_out[4170];
    assign layer1_out[2270] = ~layer0_out[1138] | layer0_out[1137];
    assign layer1_out[2271] = ~layer0_out[6930] | layer0_out[6929];
    assign layer1_out[2272] = ~(layer0_out[6490] & layer0_out[6491]);
    assign layer1_out[2273] = ~layer0_out[896] | layer0_out[895];
    assign layer1_out[2274] = layer0_out[1352] & layer0_out[1353];
    assign layer1_out[2275] = ~layer0_out[2002];
    assign layer1_out[2276] = ~layer0_out[5064];
    assign layer1_out[2277] = 1'b1;
    assign layer1_out[2278] = layer0_out[3843];
    assign layer1_out[2279] = ~(layer0_out[2295] & layer0_out[2296]);
    assign layer1_out[2280] = ~layer0_out[2831];
    assign layer1_out[2281] = layer0_out[3924];
    assign layer1_out[2282] = layer0_out[5562] | layer0_out[5563];
    assign layer1_out[2283] = ~layer0_out[7369] | layer0_out[7370];
    assign layer1_out[2284] = ~layer0_out[5039];
    assign layer1_out[2285] = layer0_out[3087];
    assign layer1_out[2286] = layer0_out[3068];
    assign layer1_out[2287] = ~(layer0_out[1281] & layer0_out[1282]);
    assign layer1_out[2288] = ~(layer0_out[1676] ^ layer0_out[1677]);
    assign layer1_out[2289] = 1'b0;
    assign layer1_out[2290] = 1'b1;
    assign layer1_out[2291] = layer0_out[7581] ^ layer0_out[7582];
    assign layer1_out[2292] = ~(layer0_out[7136] & layer0_out[7137]);
    assign layer1_out[2293] = ~(layer0_out[2463] ^ layer0_out[2464]);
    assign layer1_out[2294] = layer0_out[5613];
    assign layer1_out[2295] = layer0_out[2239] & ~layer0_out[2238];
    assign layer1_out[2296] = ~(layer0_out[6498] & layer0_out[6499]);
    assign layer1_out[2297] = layer0_out[7877] & ~layer0_out[7878];
    assign layer1_out[2298] = ~(layer0_out[5496] | layer0_out[5497]);
    assign layer1_out[2299] = layer0_out[6833];
    assign layer1_out[2300] = layer0_out[3859];
    assign layer1_out[2301] = ~(layer0_out[6752] | layer0_out[6753]);
    assign layer1_out[2302] = ~(layer0_out[546] ^ layer0_out[547]);
    assign layer1_out[2303] = layer0_out[3104];
    assign layer1_out[2304] = 1'b1;
    assign layer1_out[2305] = ~layer0_out[6071] | layer0_out[6072];
    assign layer1_out[2306] = ~(layer0_out[6282] | layer0_out[6283]);
    assign layer1_out[2307] = ~layer0_out[7926];
    assign layer1_out[2308] = ~layer0_out[4359] | layer0_out[4360];
    assign layer1_out[2309] = layer0_out[5356] | layer0_out[5357];
    assign layer1_out[2310] = ~layer0_out[872] | layer0_out[873];
    assign layer1_out[2311] = ~layer0_out[424] | layer0_out[423];
    assign layer1_out[2312] = ~layer0_out[7665] | layer0_out[7664];
    assign layer1_out[2313] = layer0_out[53];
    assign layer1_out[2314] = layer0_out[6023];
    assign layer1_out[2315] = ~(layer0_out[3422] ^ layer0_out[3423]);
    assign layer1_out[2316] = layer0_out[3632] | layer0_out[3633];
    assign layer1_out[2317] = ~layer0_out[5564];
    assign layer1_out[2318] = layer0_out[1258];
    assign layer1_out[2319] = ~(layer0_out[5486] | layer0_out[5487]);
    assign layer1_out[2320] = layer0_out[2887] & ~layer0_out[2886];
    assign layer1_out[2321] = layer0_out[4447] & layer0_out[4448];
    assign layer1_out[2322] = ~(layer0_out[6147] & layer0_out[6148]);
    assign layer1_out[2323] = layer0_out[7301];
    assign layer1_out[2324] = layer0_out[635] & layer0_out[636];
    assign layer1_out[2325] = layer0_out[1092];
    assign layer1_out[2326] = layer0_out[4674] | layer0_out[4675];
    assign layer1_out[2327] = ~(layer0_out[6977] | layer0_out[6978]);
    assign layer1_out[2328] = 1'b0;
    assign layer1_out[2329] = ~(layer0_out[2991] ^ layer0_out[2992]);
    assign layer1_out[2330] = layer0_out[4745];
    assign layer1_out[2331] = layer0_out[5125];
    assign layer1_out[2332] = ~(layer0_out[4467] | layer0_out[4468]);
    assign layer1_out[2333] = layer0_out[2313] & layer0_out[2314];
    assign layer1_out[2334] = ~(layer0_out[7156] & layer0_out[7157]);
    assign layer1_out[2335] = ~layer0_out[1024];
    assign layer1_out[2336] = layer0_out[4472] & layer0_out[4473];
    assign layer1_out[2337] = ~layer0_out[1336];
    assign layer1_out[2338] = layer0_out[5570] & ~layer0_out[5571];
    assign layer1_out[2339] = ~layer0_out[1953] | layer0_out[1952];
    assign layer1_out[2340] = layer0_out[357] & layer0_out[358];
    assign layer1_out[2341] = layer0_out[4073] & ~layer0_out[4074];
    assign layer1_out[2342] = ~layer0_out[4343];
    assign layer1_out[2343] = ~(layer0_out[34] | layer0_out[35]);
    assign layer1_out[2344] = ~layer0_out[7874];
    assign layer1_out[2345] = ~layer0_out[3400] | layer0_out[3401];
    assign layer1_out[2346] = layer0_out[1414];
    assign layer1_out[2347] = layer0_out[3248];
    assign layer1_out[2348] = layer0_out[1353] & ~layer0_out[1354];
    assign layer1_out[2349] = layer0_out[1458] & layer0_out[1459];
    assign layer1_out[2350] = layer0_out[4669] ^ layer0_out[4670];
    assign layer1_out[2351] = ~(layer0_out[4290] | layer0_out[4291]);
    assign layer1_out[2352] = ~layer0_out[5290] | layer0_out[5291];
    assign layer1_out[2353] = ~layer0_out[6821];
    assign layer1_out[2354] = layer0_out[7842];
    assign layer1_out[2355] = ~(layer0_out[4613] & layer0_out[4614]);
    assign layer1_out[2356] = layer0_out[787] | layer0_out[788];
    assign layer1_out[2357] = ~(layer0_out[883] | layer0_out[884]);
    assign layer1_out[2358] = ~(layer0_out[5602] & layer0_out[5603]);
    assign layer1_out[2359] = ~layer0_out[5142] | layer0_out[5143];
    assign layer1_out[2360] = 1'b0;
    assign layer1_out[2361] = ~(layer0_out[2704] & layer0_out[2705]);
    assign layer1_out[2362] = ~layer0_out[3764];
    assign layer1_out[2363] = ~(layer0_out[169] & layer0_out[170]);
    assign layer1_out[2364] = layer0_out[1647] ^ layer0_out[1648];
    assign layer1_out[2365] = ~layer0_out[2937] | layer0_out[2936];
    assign layer1_out[2366] = ~layer0_out[3844];
    assign layer1_out[2367] = 1'b0;
    assign layer1_out[2368] = layer0_out[1589] | layer0_out[1590];
    assign layer1_out[2369] = ~layer0_out[684] | layer0_out[685];
    assign layer1_out[2370] = ~layer0_out[2962] | layer0_out[2961];
    assign layer1_out[2371] = 1'b1;
    assign layer1_out[2372] = layer0_out[6522] | layer0_out[6523];
    assign layer1_out[2373] = layer0_out[255] & ~layer0_out[256];
    assign layer1_out[2374] = ~(layer0_out[670] & layer0_out[671]);
    assign layer1_out[2375] = ~(layer0_out[5867] | layer0_out[5868]);
    assign layer1_out[2376] = layer0_out[5217] & ~layer0_out[5218];
    assign layer1_out[2377] = layer0_out[5214];
    assign layer1_out[2378] = layer0_out[4681];
    assign layer1_out[2379] = ~layer0_out[2636] | layer0_out[2637];
    assign layer1_out[2380] = layer0_out[6074];
    assign layer1_out[2381] = layer0_out[1284];
    assign layer1_out[2382] = ~(layer0_out[7071] | layer0_out[7072]);
    assign layer1_out[2383] = layer0_out[1187] | layer0_out[1188];
    assign layer1_out[2384] = ~layer0_out[4499] | layer0_out[4500];
    assign layer1_out[2385] = ~(layer0_out[4050] ^ layer0_out[4051]);
    assign layer1_out[2386] = ~layer0_out[4394] | layer0_out[4393];
    assign layer1_out[2387] = ~layer0_out[3238];
    assign layer1_out[2388] = ~layer0_out[7312];
    assign layer1_out[2389] = ~(layer0_out[3139] & layer0_out[3140]);
    assign layer1_out[2390] = layer0_out[2366] & layer0_out[2367];
    assign layer1_out[2391] = ~layer0_out[6134] | layer0_out[6133];
    assign layer1_out[2392] = ~layer0_out[5579];
    assign layer1_out[2393] = ~layer0_out[972];
    assign layer1_out[2394] = ~layer0_out[4925] | layer0_out[4926];
    assign layer1_out[2395] = layer0_out[3438];
    assign layer1_out[2396] = ~(layer0_out[325] | layer0_out[326]);
    assign layer1_out[2397] = ~layer0_out[1244];
    assign layer1_out[2398] = ~(layer0_out[5739] | layer0_out[5740]);
    assign layer1_out[2399] = ~layer0_out[5373] | layer0_out[5372];
    assign layer1_out[2400] = layer0_out[1645] ^ layer0_out[1646];
    assign layer1_out[2401] = layer0_out[5159] ^ layer0_out[5160];
    assign layer1_out[2402] = layer0_out[5799] ^ layer0_out[5800];
    assign layer1_out[2403] = layer0_out[3473] & ~layer0_out[3472];
    assign layer1_out[2404] = layer0_out[2529] | layer0_out[2530];
    assign layer1_out[2405] = layer0_out[6347] | layer0_out[6348];
    assign layer1_out[2406] = layer0_out[1786] & layer0_out[1787];
    assign layer1_out[2407] = layer0_out[4603] & ~layer0_out[4604];
    assign layer1_out[2408] = layer0_out[2351] & ~layer0_out[2350];
    assign layer1_out[2409] = layer0_out[905] ^ layer0_out[906];
    assign layer1_out[2410] = layer0_out[6939] & layer0_out[6940];
    assign layer1_out[2411] = layer0_out[6905] & layer0_out[6906];
    assign layer1_out[2412] = layer0_out[2147] & layer0_out[2148];
    assign layer1_out[2413] = ~layer0_out[4033];
    assign layer1_out[2414] = ~layer0_out[5194] | layer0_out[5193];
    assign layer1_out[2415] = ~layer0_out[2404];
    assign layer1_out[2416] = 1'b1;
    assign layer1_out[2417] = 1'b1;
    assign layer1_out[2418] = ~layer0_out[4522] | layer0_out[4523];
    assign layer1_out[2419] = layer0_out[2564] ^ layer0_out[2565];
    assign layer1_out[2420] = layer0_out[655] & ~layer0_out[654];
    assign layer1_out[2421] = layer0_out[1946] & ~layer0_out[1945];
    assign layer1_out[2422] = layer0_out[4217] & layer0_out[4218];
    assign layer1_out[2423] = layer0_out[5331];
    assign layer1_out[2424] = ~layer0_out[439] | layer0_out[438];
    assign layer1_out[2425] = ~layer0_out[4666] | layer0_out[4665];
    assign layer1_out[2426] = layer0_out[3828] & layer0_out[3829];
    assign layer1_out[2427] = layer0_out[3362];
    assign layer1_out[2428] = ~layer0_out[6774] | layer0_out[6775];
    assign layer1_out[2429] = layer0_out[7013] | layer0_out[7014];
    assign layer1_out[2430] = layer0_out[459] | layer0_out[460];
    assign layer1_out[2431] = ~layer0_out[7929] | layer0_out[7928];
    assign layer1_out[2432] = ~layer0_out[775] | layer0_out[774];
    assign layer1_out[2433] = layer0_out[2611];
    assign layer1_out[2434] = layer0_out[3349];
    assign layer1_out[2435] = ~layer0_out[4307] | layer0_out[4306];
    assign layer1_out[2436] = ~layer0_out[60];
    assign layer1_out[2437] = 1'b0;
    assign layer1_out[2438] = layer0_out[4042] | layer0_out[4043];
    assign layer1_out[2439] = 1'b0;
    assign layer1_out[2440] = layer0_out[1240];
    assign layer1_out[2441] = layer0_out[5165] & layer0_out[5166];
    assign layer1_out[2442] = ~(layer0_out[5342] & layer0_out[5343]);
    assign layer1_out[2443] = layer0_out[1340];
    assign layer1_out[2444] = ~(layer0_out[6218] | layer0_out[6219]);
    assign layer1_out[2445] = layer0_out[2174];
    assign layer1_out[2446] = layer0_out[822] & ~layer0_out[823];
    assign layer1_out[2447] = ~layer0_out[7866];
    assign layer1_out[2448] = layer0_out[380];
    assign layer1_out[2449] = ~(layer0_out[4960] & layer0_out[4961]);
    assign layer1_out[2450] = ~layer0_out[3333] | layer0_out[3332];
    assign layer1_out[2451] = ~layer0_out[6076] | layer0_out[6077];
    assign layer1_out[2452] = ~layer0_out[370];
    assign layer1_out[2453] = ~layer0_out[7611] | layer0_out[7610];
    assign layer1_out[2454] = ~(layer0_out[4814] & layer0_out[4815]);
    assign layer1_out[2455] = layer0_out[7753];
    assign layer1_out[2456] = ~layer0_out[1082] | layer0_out[1081];
    assign layer1_out[2457] = layer0_out[2315];
    assign layer1_out[2458] = ~layer0_out[720];
    assign layer1_out[2459] = layer0_out[5010];
    assign layer1_out[2460] = layer0_out[4089] & ~layer0_out[4090];
    assign layer1_out[2461] = ~(layer0_out[6959] & layer0_out[6960]);
    assign layer1_out[2462] = ~layer0_out[5003] | layer0_out[5002];
    assign layer1_out[2463] = ~layer0_out[6430] | layer0_out[6429];
    assign layer1_out[2464] = ~(layer0_out[5235] & layer0_out[5236]);
    assign layer1_out[2465] = layer0_out[3669] & ~layer0_out[3668];
    assign layer1_out[2466] = layer0_out[2384] & layer0_out[2385];
    assign layer1_out[2467] = layer0_out[7286] & ~layer0_out[7287];
    assign layer1_out[2468] = ~layer0_out[4782];
    assign layer1_out[2469] = layer0_out[1178];
    assign layer1_out[2470] = ~layer0_out[553] | layer0_out[554];
    assign layer1_out[2471] = ~layer0_out[7200] | layer0_out[7201];
    assign layer1_out[2472] = ~(layer0_out[4663] ^ layer0_out[4664]);
    assign layer1_out[2473] = ~layer0_out[6275] | layer0_out[6274];
    assign layer1_out[2474] = ~layer0_out[323];
    assign layer1_out[2475] = ~(layer0_out[2877] ^ layer0_out[2878]);
    assign layer1_out[2476] = ~layer0_out[5088];
    assign layer1_out[2477] = ~layer0_out[3009];
    assign layer1_out[2478] = layer0_out[1201] & layer0_out[1202];
    assign layer1_out[2479] = ~layer0_out[6875];
    assign layer1_out[2480] = layer0_out[2062] & layer0_out[2063];
    assign layer1_out[2481] = ~layer0_out[2264] | layer0_out[2263];
    assign layer1_out[2482] = layer0_out[360] ^ layer0_out[361];
    assign layer1_out[2483] = layer0_out[792] & layer0_out[793];
    assign layer1_out[2484] = ~(layer0_out[7332] | layer0_out[7333]);
    assign layer1_out[2485] = ~layer0_out[1199];
    assign layer1_out[2486] = layer0_out[2526];
    assign layer1_out[2487] = layer0_out[3565] | layer0_out[3566];
    assign layer1_out[2488] = layer0_out[7267];
    assign layer1_out[2489] = layer0_out[4269];
    assign layer1_out[2490] = ~layer0_out[1564];
    assign layer1_out[2491] = layer0_out[6255] & ~layer0_out[6256];
    assign layer1_out[2492] = ~layer0_out[1860];
    assign layer1_out[2493] = layer0_out[5917] & ~layer0_out[5918];
    assign layer1_out[2494] = ~(layer0_out[3137] | layer0_out[3138]);
    assign layer1_out[2495] = ~(layer0_out[7347] | layer0_out[7348]);
    assign layer1_out[2496] = ~layer0_out[2626] | layer0_out[2627];
    assign layer1_out[2497] = 1'b1;
    assign layer1_out[2498] = ~layer0_out[7990];
    assign layer1_out[2499] = ~(layer0_out[2746] & layer0_out[2747]);
    assign layer1_out[2500] = ~(layer0_out[7058] | layer0_out[7059]);
    assign layer1_out[2501] = layer0_out[2501];
    assign layer1_out[2502] = layer0_out[43];
    assign layer1_out[2503] = layer0_out[440] & layer0_out[441];
    assign layer1_out[2504] = ~layer0_out[5037] | layer0_out[5038];
    assign layer1_out[2505] = ~layer0_out[4164];
    assign layer1_out[2506] = layer0_out[6913] | layer0_out[6914];
    assign layer1_out[2507] = layer0_out[6766] & layer0_out[6767];
    assign layer1_out[2508] = layer0_out[420] | layer0_out[421];
    assign layer1_out[2509] = ~layer0_out[2258] | layer0_out[2257];
    assign layer1_out[2510] = layer0_out[3979] & ~layer0_out[3980];
    assign layer1_out[2511] = layer0_out[3771];
    assign layer1_out[2512] = layer0_out[6061];
    assign layer1_out[2513] = layer0_out[5126];
    assign layer1_out[2514] = layer0_out[941];
    assign layer1_out[2515] = ~layer0_out[228] | layer0_out[227];
    assign layer1_out[2516] = layer0_out[4518] & ~layer0_out[4517];
    assign layer1_out[2517] = ~(layer0_out[2375] | layer0_out[2376]);
    assign layer1_out[2518] = ~layer0_out[3728];
    assign layer1_out[2519] = layer0_out[7480];
    assign layer1_out[2520] = layer0_out[1717];
    assign layer1_out[2521] = layer0_out[3835] | layer0_out[3836];
    assign layer1_out[2522] = layer0_out[7986] & layer0_out[7987];
    assign layer1_out[2523] = layer0_out[7623] | layer0_out[7624];
    assign layer1_out[2524] = layer0_out[3462];
    assign layer1_out[2525] = layer0_out[70];
    assign layer1_out[2526] = ~layer0_out[1057] | layer0_out[1058];
    assign layer1_out[2527] = ~layer0_out[6212] | layer0_out[6213];
    assign layer1_out[2528] = layer0_out[1091];
    assign layer1_out[2529] = ~layer0_out[6063];
    assign layer1_out[2530] = ~(layer0_out[44] & layer0_out[45]);
    assign layer1_out[2531] = layer0_out[2562] & ~layer0_out[2561];
    assign layer1_out[2532] = ~layer0_out[1948];
    assign layer1_out[2533] = ~layer0_out[2494] | layer0_out[2495];
    assign layer1_out[2534] = ~layer0_out[6363] | layer0_out[6362];
    assign layer1_out[2535] = layer0_out[6418];
    assign layer1_out[2536] = layer0_out[7451];
    assign layer1_out[2537] = layer0_out[3750] | layer0_out[3751];
    assign layer1_out[2538] = ~(layer0_out[753] | layer0_out[754]);
    assign layer1_out[2539] = ~(layer0_out[2073] ^ layer0_out[2074]);
    assign layer1_out[2540] = layer0_out[1234];
    assign layer1_out[2541] = layer0_out[1656];
    assign layer1_out[2542] = ~layer0_out[7647];
    assign layer1_out[2543] = layer0_out[6774];
    assign layer1_out[2544] = ~(layer0_out[2689] | layer0_out[2690]);
    assign layer1_out[2545] = ~layer0_out[7492];
    assign layer1_out[2546] = ~(layer0_out[6288] & layer0_out[6289]);
    assign layer1_out[2547] = ~layer0_out[5894];
    assign layer1_out[2548] = ~(layer0_out[4686] ^ layer0_out[4687]);
    assign layer1_out[2549] = ~layer0_out[797] | layer0_out[796];
    assign layer1_out[2550] = layer0_out[1943] & ~layer0_out[1942];
    assign layer1_out[2551] = ~(layer0_out[4716] & layer0_out[4717]);
    assign layer1_out[2552] = ~(layer0_out[5941] | layer0_out[5942]);
    assign layer1_out[2553] = layer0_out[4292] & ~layer0_out[4293];
    assign layer1_out[2554] = layer0_out[5585] | layer0_out[5586];
    assign layer1_out[2555] = ~layer0_out[1271];
    assign layer1_out[2556] = layer0_out[810] & ~layer0_out[811];
    assign layer1_out[2557] = layer0_out[597];
    assign layer1_out[2558] = ~(layer0_out[7238] | layer0_out[7239]);
    assign layer1_out[2559] = layer0_out[2344] & ~layer0_out[2345];
    assign layer1_out[2560] = layer0_out[1029];
    assign layer1_out[2561] = ~(layer0_out[5956] & layer0_out[5957]);
    assign layer1_out[2562] = ~layer0_out[5197];
    assign layer1_out[2563] = ~layer0_out[2641] | layer0_out[2640];
    assign layer1_out[2564] = ~(layer0_out[5643] | layer0_out[5644]);
    assign layer1_out[2565] = 1'b0;
    assign layer1_out[2566] = layer0_out[7954] & ~layer0_out[7953];
    assign layer1_out[2567] = ~layer0_out[7319] | layer0_out[7320];
    assign layer1_out[2568] = ~(layer0_out[1625] | layer0_out[1626]);
    assign layer1_out[2569] = ~layer0_out[898];
    assign layer1_out[2570] = ~(layer0_out[4843] ^ layer0_out[4844]);
    assign layer1_out[2571] = layer0_out[2089] & ~layer0_out[2088];
    assign layer1_out[2572] = layer0_out[7341] ^ layer0_out[7342];
    assign layer1_out[2573] = layer0_out[1019] & layer0_out[1020];
    assign layer1_out[2574] = ~(layer0_out[2119] | layer0_out[2120]);
    assign layer1_out[2575] = ~layer0_out[3692];
    assign layer1_out[2576] = ~layer0_out[3773] | layer0_out[3774];
    assign layer1_out[2577] = ~layer0_out[5251];
    assign layer1_out[2578] = 1'b1;
    assign layer1_out[2579] = layer0_out[4697] ^ layer0_out[4698];
    assign layer1_out[2580] = layer0_out[5769];
    assign layer1_out[2581] = layer0_out[3890];
    assign layer1_out[2582] = layer0_out[7000];
    assign layer1_out[2583] = layer0_out[5566];
    assign layer1_out[2584] = ~(layer0_out[2596] & layer0_out[2597]);
    assign layer1_out[2585] = ~(layer0_out[3214] ^ layer0_out[3215]);
    assign layer1_out[2586] = 1'b0;
    assign layer1_out[2587] = ~layer0_out[3697];
    assign layer1_out[2588] = ~layer0_out[4063];
    assign layer1_out[2589] = layer0_out[2821];
    assign layer1_out[2590] = ~(layer0_out[6299] ^ layer0_out[6300]);
    assign layer1_out[2591] = ~layer0_out[1868];
    assign layer1_out[2592] = ~layer0_out[6455];
    assign layer1_out[2593] = ~(layer0_out[3592] | layer0_out[3593]);
    assign layer1_out[2594] = 1'b0;
    assign layer1_out[2595] = layer0_out[4622];
    assign layer1_out[2596] = layer0_out[7133] | layer0_out[7134];
    assign layer1_out[2597] = layer0_out[2421];
    assign layer1_out[2598] = 1'b0;
    assign layer1_out[2599] = ~(layer0_out[505] ^ layer0_out[506]);
    assign layer1_out[2600] = ~layer0_out[587];
    assign layer1_out[2601] = layer0_out[7569] & ~layer0_out[7570];
    assign layer1_out[2602] = 1'b1;
    assign layer1_out[2603] = ~layer0_out[1627] | layer0_out[1626];
    assign layer1_out[2604] = layer0_out[7018] & ~layer0_out[7017];
    assign layer1_out[2605] = layer0_out[6765] & layer0_out[6766];
    assign layer1_out[2606] = ~(layer0_out[7942] & layer0_out[7943]);
    assign layer1_out[2607] = layer0_out[1723];
    assign layer1_out[2608] = layer0_out[2096];
    assign layer1_out[2609] = ~layer0_out[2659];
    assign layer1_out[2610] = layer0_out[7711] ^ layer0_out[7712];
    assign layer1_out[2611] = layer0_out[5181] & ~layer0_out[5182];
    assign layer1_out[2612] = layer0_out[6705] & ~layer0_out[6706];
    assign layer1_out[2613] = layer0_out[2937] & ~layer0_out[2938];
    assign layer1_out[2614] = layer0_out[3498] & ~layer0_out[3497];
    assign layer1_out[2615] = layer0_out[2692] & ~layer0_out[2693];
    assign layer1_out[2616] = ~layer0_out[1495] | layer0_out[1494];
    assign layer1_out[2617] = ~layer0_out[4365] | layer0_out[4364];
    assign layer1_out[2618] = ~layer0_out[1172] | layer0_out[1171];
    assign layer1_out[2619] = layer0_out[585] & ~layer0_out[584];
    assign layer1_out[2620] = ~layer0_out[6034];
    assign layer1_out[2621] = ~layer0_out[83] | layer0_out[82];
    assign layer1_out[2622] = ~(layer0_out[6925] ^ layer0_out[6926]);
    assign layer1_out[2623] = ~(layer0_out[2700] & layer0_out[2701]);
    assign layer1_out[2624] = ~layer0_out[1742] | layer0_out[1741];
    assign layer1_out[2625] = layer0_out[6279] | layer0_out[6280];
    assign layer1_out[2626] = ~layer0_out[6643] | layer0_out[6644];
    assign layer1_out[2627] = ~(layer0_out[7103] & layer0_out[7104]);
    assign layer1_out[2628] = ~(layer0_out[6427] | layer0_out[6428]);
    assign layer1_out[2629] = layer0_out[6757] & ~layer0_out[6756];
    assign layer1_out[2630] = ~layer0_out[692];
    assign layer1_out[2631] = layer0_out[6494] | layer0_out[6495];
    assign layer1_out[2632] = layer0_out[5534];
    assign layer1_out[2633] = ~layer0_out[2973] | layer0_out[2974];
    assign layer1_out[2634] = ~layer0_out[3973] | layer0_out[3972];
    assign layer1_out[2635] = ~layer0_out[5533] | layer0_out[5534];
    assign layer1_out[2636] = ~layer0_out[4654] | layer0_out[4653];
    assign layer1_out[2637] = ~(layer0_out[4506] | layer0_out[4507]);
    assign layer1_out[2638] = 1'b1;
    assign layer1_out[2639] = 1'b1;
    assign layer1_out[2640] = layer0_out[4132] & ~layer0_out[4133];
    assign layer1_out[2641] = layer0_out[2278];
    assign layer1_out[2642] = ~layer0_out[1297];
    assign layer1_out[2643] = layer0_out[2910] & ~layer0_out[2909];
    assign layer1_out[2644] = ~(layer0_out[545] & layer0_out[546]);
    assign layer1_out[2645] = ~(layer0_out[7149] ^ layer0_out[7150]);
    assign layer1_out[2646] = ~layer0_out[3539];
    assign layer1_out[2647] = layer0_out[56];
    assign layer1_out[2648] = ~layer0_out[2652] | layer0_out[2651];
    assign layer1_out[2649] = ~layer0_out[2432];
    assign layer1_out[2650] = ~layer0_out[3354];
    assign layer1_out[2651] = ~layer0_out[2816] | layer0_out[2817];
    assign layer1_out[2652] = layer0_out[6906];
    assign layer1_out[2653] = layer0_out[3838] & ~layer0_out[3837];
    assign layer1_out[2654] = layer0_out[7558];
    assign layer1_out[2655] = layer0_out[4181] & ~layer0_out[4180];
    assign layer1_out[2656] = ~layer0_out[6743];
    assign layer1_out[2657] = layer0_out[4558];
    assign layer1_out[2658] = layer0_out[947];
    assign layer1_out[2659] = layer0_out[7779] & ~layer0_out[7780];
    assign layer1_out[2660] = ~(layer0_out[1400] | layer0_out[1401]);
    assign layer1_out[2661] = ~(layer0_out[2361] ^ layer0_out[2362]);
    assign layer1_out[2662] = ~layer0_out[828] | layer0_out[829];
    assign layer1_out[2663] = ~(layer0_out[2776] | layer0_out[2777]);
    assign layer1_out[2664] = layer0_out[5391];
    assign layer1_out[2665] = layer0_out[5641] | layer0_out[5642];
    assign layer1_out[2666] = ~(layer0_out[4005] | layer0_out[4006]);
    assign layer1_out[2667] = layer0_out[5592];
    assign layer1_out[2668] = layer0_out[2385];
    assign layer1_out[2669] = layer0_out[7578] | layer0_out[7579];
    assign layer1_out[2670] = layer0_out[7625];
    assign layer1_out[2671] = ~(layer0_out[3685] ^ layer0_out[3686]);
    assign layer1_out[2672] = layer0_out[6984];
    assign layer1_out[2673] = layer0_out[935] ^ layer0_out[936];
    assign layer1_out[2674] = ~layer0_out[730];
    assign layer1_out[2675] = ~layer0_out[4583] | layer0_out[4582];
    assign layer1_out[2676] = ~(layer0_out[0] | layer0_out[2]);
    assign layer1_out[2677] = ~(layer0_out[7315] | layer0_out[7316]);
    assign layer1_out[2678] = 1'b1;
    assign layer1_out[2679] = layer0_out[168];
    assign layer1_out[2680] = layer0_out[4516] ^ layer0_out[4517];
    assign layer1_out[2681] = ~layer0_out[5254] | layer0_out[5255];
    assign layer1_out[2682] = ~(layer0_out[3691] | layer0_out[3692]);
    assign layer1_out[2683] = layer0_out[5423] & ~layer0_out[5424];
    assign layer1_out[2684] = layer0_out[4260];
    assign layer1_out[2685] = layer0_out[7562] & ~layer0_out[7563];
    assign layer1_out[2686] = ~layer0_out[4044] | layer0_out[4045];
    assign layer1_out[2687] = layer0_out[2765] & ~layer0_out[2766];
    assign layer1_out[2688] = layer0_out[403];
    assign layer1_out[2689] = layer0_out[2857] & ~layer0_out[2858];
    assign layer1_out[2690] = layer0_out[1880] & ~layer0_out[1881];
    assign layer1_out[2691] = layer0_out[4158] & ~layer0_out[4159];
    assign layer1_out[2692] = 1'b1;
    assign layer1_out[2693] = ~layer0_out[7930] | layer0_out[7929];
    assign layer1_out[2694] = layer0_out[1073];
    assign layer1_out[2695] = layer0_out[6153] | layer0_out[6154];
    assign layer1_out[2696] = layer0_out[6805];
    assign layer1_out[2697] = layer0_out[3193] ^ layer0_out[3194];
    assign layer1_out[2698] = ~layer0_out[4677];
    assign layer1_out[2699] = ~layer0_out[6505];
    assign layer1_out[2700] = layer0_out[6604];
    assign layer1_out[2701] = layer0_out[668] & ~layer0_out[667];
    assign layer1_out[2702] = ~(layer0_out[1611] ^ layer0_out[1612]);
    assign layer1_out[2703] = layer0_out[4925] & ~layer0_out[4924];
    assign layer1_out[2704] = layer0_out[1175];
    assign layer1_out[2705] = layer0_out[1683] & ~layer0_out[1682];
    assign layer1_out[2706] = ~layer0_out[4558] | layer0_out[4557];
    assign layer1_out[2707] = ~(layer0_out[1222] | layer0_out[1223]);
    assign layer1_out[2708] = ~layer0_out[6276] | layer0_out[6277];
    assign layer1_out[2709] = ~layer0_out[1010] | layer0_out[1009];
    assign layer1_out[2710] = 1'b0;
    assign layer1_out[2711] = 1'b1;
    assign layer1_out[2712] = ~(layer0_out[5730] ^ layer0_out[5731]);
    assign layer1_out[2713] = layer0_out[3500] & ~layer0_out[3501];
    assign layer1_out[2714] = ~layer0_out[959];
    assign layer1_out[2715] = ~(layer0_out[7293] & layer0_out[7294]);
    assign layer1_out[2716] = ~layer0_out[4861];
    assign layer1_out[2717] = ~(layer0_out[98] | layer0_out[99]);
    assign layer1_out[2718] = layer0_out[6748];
    assign layer1_out[2719] = ~layer0_out[714];
    assign layer1_out[2720] = ~(layer0_out[6311] & layer0_out[6312]);
    assign layer1_out[2721] = ~layer0_out[5624] | layer0_out[5625];
    assign layer1_out[2722] = ~(layer0_out[7004] & layer0_out[7005]);
    assign layer1_out[2723] = ~layer0_out[3782] | layer0_out[3781];
    assign layer1_out[2724] = layer0_out[2840] ^ layer0_out[2841];
    assign layer1_out[2725] = layer0_out[5734];
    assign layer1_out[2726] = layer0_out[6529];
    assign layer1_out[2727] = 1'b0;
    assign layer1_out[2728] = ~(layer0_out[5067] | layer0_out[5068]);
    assign layer1_out[2729] = layer0_out[6024];
    assign layer1_out[2730] = layer0_out[7062] & layer0_out[7063];
    assign layer1_out[2731] = layer0_out[7911] | layer0_out[7912];
    assign layer1_out[2732] = ~layer0_out[6459];
    assign layer1_out[2733] = ~(layer0_out[610] & layer0_out[611]);
    assign layer1_out[2734] = ~layer0_out[196];
    assign layer1_out[2735] = layer0_out[3420];
    assign layer1_out[2736] = layer0_out[2679] & ~layer0_out[2678];
    assign layer1_out[2737] = layer0_out[2531] & ~layer0_out[2532];
    assign layer1_out[2738] = layer0_out[2724] & ~layer0_out[2723];
    assign layer1_out[2739] = layer0_out[1731] & layer0_out[1732];
    assign layer1_out[2740] = 1'b0;
    assign layer1_out[2741] = ~(layer0_out[7447] & layer0_out[7448]);
    assign layer1_out[2742] = layer0_out[3498];
    assign layer1_out[2743] = layer0_out[830] & layer0_out[831];
    assign layer1_out[2744] = ~(layer0_out[1515] | layer0_out[1516]);
    assign layer1_out[2745] = ~layer0_out[7874] | layer0_out[7875];
    assign layer1_out[2746] = layer0_out[408] & layer0_out[409];
    assign layer1_out[2747] = ~layer0_out[1635];
    assign layer1_out[2748] = layer0_out[3633] | layer0_out[3634];
    assign layer1_out[2749] = ~layer0_out[2074] | layer0_out[2075];
    assign layer1_out[2750] = ~(layer0_out[7092] | layer0_out[7093]);
    assign layer1_out[2751] = layer0_out[7967];
    assign layer1_out[2752] = layer0_out[4883] | layer0_out[4884];
    assign layer1_out[2753] = layer0_out[1960] | layer0_out[1961];
    assign layer1_out[2754] = ~layer0_out[3602] | layer0_out[3601];
    assign layer1_out[2755] = layer0_out[6264];
    assign layer1_out[2756] = ~(layer0_out[806] & layer0_out[807]);
    assign layer1_out[2757] = ~layer0_out[288] | layer0_out[289];
    assign layer1_out[2758] = ~layer0_out[2375];
    assign layer1_out[2759] = layer0_out[5488] & ~layer0_out[5487];
    assign layer1_out[2760] = ~layer0_out[5189];
    assign layer1_out[2761] = layer0_out[2890] | layer0_out[2891];
    assign layer1_out[2762] = layer0_out[2500] ^ layer0_out[2501];
    assign layer1_out[2763] = ~(layer0_out[3496] | layer0_out[3497]);
    assign layer1_out[2764] = ~(layer0_out[3504] | layer0_out[3505]);
    assign layer1_out[2765] = 1'b0;
    assign layer1_out[2766] = layer0_out[2169];
    assign layer1_out[2767] = layer0_out[3030];
    assign layer1_out[2768] = ~layer0_out[6158] | layer0_out[6157];
    assign layer1_out[2769] = layer0_out[2979] & ~layer0_out[2978];
    assign layer1_out[2770] = ~(layer0_out[2082] | layer0_out[2083]);
    assign layer1_out[2771] = ~(layer0_out[1891] & layer0_out[1892]);
    assign layer1_out[2772] = 1'b0;
    assign layer1_out[2773] = ~layer0_out[3333];
    assign layer1_out[2774] = layer0_out[6484] | layer0_out[6485];
    assign layer1_out[2775] = layer0_out[529];
    assign layer1_out[2776] = layer0_out[908];
    assign layer1_out[2777] = layer0_out[1752] & layer0_out[1753];
    assign layer1_out[2778] = ~(layer0_out[4982] & layer0_out[4983]);
    assign layer1_out[2779] = layer0_out[7056];
    assign layer1_out[2780] = ~layer0_out[2343];
    assign layer1_out[2781] = layer0_out[2021] | layer0_out[2022];
    assign layer1_out[2782] = ~(layer0_out[2072] | layer0_out[2073]);
    assign layer1_out[2783] = ~layer0_out[4035];
    assign layer1_out[2784] = layer0_out[4725] | layer0_out[4726];
    assign layer1_out[2785] = ~layer0_out[6073] | layer0_out[6072];
    assign layer1_out[2786] = 1'b1;
    assign layer1_out[2787] = ~layer0_out[878] | layer0_out[879];
    assign layer1_out[2788] = layer0_out[6057] & ~layer0_out[6058];
    assign layer1_out[2789] = ~(layer0_out[5102] & layer0_out[5103]);
    assign layer1_out[2790] = ~layer0_out[3545] | layer0_out[3546];
    assign layer1_out[2791] = layer0_out[7902];
    assign layer1_out[2792] = layer0_out[503] | layer0_out[504];
    assign layer1_out[2793] = ~layer0_out[2913] | layer0_out[2914];
    assign layer1_out[2794] = ~layer0_out[4968] | layer0_out[4967];
    assign layer1_out[2795] = layer0_out[974];
    assign layer1_out[2796] = ~layer0_out[4708];
    assign layer1_out[2797] = layer0_out[2698] | layer0_out[2699];
    assign layer1_out[2798] = layer0_out[6592] | layer0_out[6593];
    assign layer1_out[2799] = ~layer0_out[130];
    assign layer1_out[2800] = ~layer0_out[6704];
    assign layer1_out[2801] = 1'b1;
    assign layer1_out[2802] = layer0_out[3534] & ~layer0_out[3533];
    assign layer1_out[2803] = ~layer0_out[6048] | layer0_out[6049];
    assign layer1_out[2804] = ~layer0_out[223];
    assign layer1_out[2805] = 1'b0;
    assign layer1_out[2806] = layer0_out[5984] & ~layer0_out[5985];
    assign layer1_out[2807] = layer0_out[1457];
    assign layer1_out[2808] = ~(layer0_out[1244] | layer0_out[1245]);
    assign layer1_out[2809] = ~layer0_out[4798];
    assign layer1_out[2810] = layer0_out[2492];
    assign layer1_out[2811] = 1'b0;
    assign layer1_out[2812] = layer0_out[2335] & layer0_out[2336];
    assign layer1_out[2813] = layer0_out[191];
    assign layer1_out[2814] = layer0_out[1836] & layer0_out[1837];
    assign layer1_out[2815] = layer0_out[3221] | layer0_out[3222];
    assign layer1_out[2816] = ~(layer0_out[4659] & layer0_out[4660]);
    assign layer1_out[2817] = layer0_out[7475] | layer0_out[7476];
    assign layer1_out[2818] = layer0_out[5903] | layer0_out[5904];
    assign layer1_out[2819] = ~layer0_out[2296];
    assign layer1_out[2820] = layer0_out[6890];
    assign layer1_out[2821] = ~layer0_out[4381];
    assign layer1_out[2822] = layer0_out[158] ^ layer0_out[159];
    assign layer1_out[2823] = layer0_out[4122];
    assign layer1_out[2824] = ~layer0_out[2931];
    assign layer1_out[2825] = ~layer0_out[5918];
    assign layer1_out[2826] = ~(layer0_out[6292] ^ layer0_out[6293]);
    assign layer1_out[2827] = ~layer0_out[5777];
    assign layer1_out[2828] = ~layer0_out[5675];
    assign layer1_out[2829] = layer0_out[3460] & ~layer0_out[3461];
    assign layer1_out[2830] = layer0_out[3369] & ~layer0_out[3368];
    assign layer1_out[2831] = ~layer0_out[1208] | layer0_out[1209];
    assign layer1_out[2832] = ~(layer0_out[1302] & layer0_out[1303]);
    assign layer1_out[2833] = layer0_out[3339];
    assign layer1_out[2834] = ~layer0_out[3042];
    assign layer1_out[2835] = ~layer0_out[6995];
    assign layer1_out[2836] = ~layer0_out[4537];
    assign layer1_out[2837] = layer0_out[5637];
    assign layer1_out[2838] = layer0_out[6842];
    assign layer1_out[2839] = ~layer0_out[5149] | layer0_out[5150];
    assign layer1_out[2840] = ~(layer0_out[7283] ^ layer0_out[7284]);
    assign layer1_out[2841] = layer0_out[5229] & ~layer0_out[5228];
    assign layer1_out[2842] = layer0_out[3300] & layer0_out[3301];
    assign layer1_out[2843] = layer0_out[7364] ^ layer0_out[7365];
    assign layer1_out[2844] = layer0_out[4453] & ~layer0_out[4454];
    assign layer1_out[2845] = layer0_out[3780] & layer0_out[3781];
    assign layer1_out[2846] = layer0_out[6508] ^ layer0_out[6509];
    assign layer1_out[2847] = layer0_out[1373] ^ layer0_out[1374];
    assign layer1_out[2848] = ~layer0_out[5446] | layer0_out[5445];
    assign layer1_out[2849] = 1'b1;
    assign layer1_out[2850] = layer0_out[1672] & ~layer0_out[1671];
    assign layer1_out[2851] = layer0_out[4294] ^ layer0_out[4295];
    assign layer1_out[2852] = ~layer0_out[6921] | layer0_out[6920];
    assign layer1_out[2853] = layer0_out[3704];
    assign layer1_out[2854] = layer0_out[1375] ^ layer0_out[1376];
    assign layer1_out[2855] = layer0_out[1322] ^ layer0_out[1323];
    assign layer1_out[2856] = ~layer0_out[5326];
    assign layer1_out[2857] = ~layer0_out[3673];
    assign layer1_out[2858] = layer0_out[6821] | layer0_out[6822];
    assign layer1_out[2859] = layer0_out[4786] & ~layer0_out[4787];
    assign layer1_out[2860] = layer0_out[3245];
    assign layer1_out[2861] = ~(layer0_out[3470] ^ layer0_out[3471]);
    assign layer1_out[2862] = ~layer0_out[4350];
    assign layer1_out[2863] = layer0_out[3470] & ~layer0_out[3469];
    assign layer1_out[2864] = ~layer0_out[4429];
    assign layer1_out[2865] = ~(layer0_out[6254] ^ layer0_out[6255]);
    assign layer1_out[2866] = ~layer0_out[737];
    assign layer1_out[2867] = ~(layer0_out[4599] | layer0_out[4600]);
    assign layer1_out[2868] = ~layer0_out[457] | layer0_out[456];
    assign layer1_out[2869] = layer0_out[6598] & ~layer0_out[6599];
    assign layer1_out[2870] = ~layer0_out[5043];
    assign layer1_out[2871] = ~layer0_out[4179];
    assign layer1_out[2872] = layer0_out[7809] & layer0_out[7810];
    assign layer1_out[2873] = ~layer0_out[4910] | layer0_out[4909];
    assign layer1_out[2874] = ~layer0_out[7854];
    assign layer1_out[2875] = ~(layer0_out[4765] | layer0_out[4766]);
    assign layer1_out[2876] = ~layer0_out[4597] | layer0_out[4596];
    assign layer1_out[2877] = layer0_out[7154];
    assign layer1_out[2878] = layer0_out[5568];
    assign layer1_out[2879] = layer0_out[3299] & ~layer0_out[3298];
    assign layer1_out[2880] = layer0_out[7599] ^ layer0_out[7600];
    assign layer1_out[2881] = layer0_out[6687] & ~layer0_out[6688];
    assign layer1_out[2882] = ~(layer0_out[6971] ^ layer0_out[6972]);
    assign layer1_out[2883] = layer0_out[305];
    assign layer1_out[2884] = layer0_out[5515] & ~layer0_out[5514];
    assign layer1_out[2885] = layer0_out[735] | layer0_out[736];
    assign layer1_out[2886] = 1'b1;
    assign layer1_out[2887] = layer0_out[425];
    assign layer1_out[2888] = layer0_out[1992] | layer0_out[1993];
    assign layer1_out[2889] = layer0_out[640] & ~layer0_out[641];
    assign layer1_out[2890] = ~(layer0_out[2568] | layer0_out[2569]);
    assign layer1_out[2891] = layer0_out[1679] & layer0_out[1680];
    assign layer1_out[2892] = layer0_out[4717] & ~layer0_out[4718];
    assign layer1_out[2893] = ~(layer0_out[1739] ^ layer0_out[1740]);
    assign layer1_out[2894] = ~(layer0_out[3156] & layer0_out[3157]);
    assign layer1_out[2895] = ~(layer0_out[777] ^ layer0_out[778]);
    assign layer1_out[2896] = layer0_out[6885] & layer0_out[6886];
    assign layer1_out[2897] = layer0_out[6117] & layer0_out[6118];
    assign layer1_out[2898] = ~layer0_out[4618];
    assign layer1_out[2899] = layer0_out[262] ^ layer0_out[263];
    assign layer1_out[2900] = ~layer0_out[7425] | layer0_out[7424];
    assign layer1_out[2901] = ~layer0_out[1165];
    assign layer1_out[2902] = ~layer0_out[7737] | layer0_out[7736];
    assign layer1_out[2903] = layer0_out[5804] & ~layer0_out[5803];
    assign layer1_out[2904] = ~layer0_out[3915];
    assign layer1_out[2905] = layer0_out[4787];
    assign layer1_out[2906] = ~layer0_out[802] | layer0_out[801];
    assign layer1_out[2907] = ~layer0_out[436] | layer0_out[437];
    assign layer1_out[2908] = ~(layer0_out[1410] & layer0_out[1411]);
    assign layer1_out[2909] = layer0_out[1654];
    assign layer1_out[2910] = layer0_out[7164] ^ layer0_out[7165];
    assign layer1_out[2911] = ~layer0_out[5365] | layer0_out[5366];
    assign layer1_out[2912] = ~layer0_out[6657] | layer0_out[6658];
    assign layer1_out[2913] = ~layer0_out[2] | layer0_out[1];
    assign layer1_out[2914] = layer0_out[2553];
    assign layer1_out[2915] = layer0_out[1990] | layer0_out[1991];
    assign layer1_out[2916] = ~(layer0_out[7705] | layer0_out[7706]);
    assign layer1_out[2917] = layer0_out[6054];
    assign layer1_out[2918] = ~(layer0_out[5328] ^ layer0_out[5329]);
    assign layer1_out[2919] = ~layer0_out[6521];
    assign layer1_out[2920] = ~(layer0_out[5926] & layer0_out[5927]);
    assign layer1_out[2921] = layer0_out[1463];
    assign layer1_out[2922] = ~(layer0_out[2896] & layer0_out[2897]);
    assign layer1_out[2923] = layer0_out[2136] & ~layer0_out[2135];
    assign layer1_out[2924] = layer0_out[7596];
    assign layer1_out[2925] = layer0_out[2547] & ~layer0_out[2546];
    assign layer1_out[2926] = ~(layer0_out[4325] & layer0_out[4326]);
    assign layer1_out[2927] = layer0_out[5122];
    assign layer1_out[2928] = ~layer0_out[7919] | layer0_out[7920];
    assign layer1_out[2929] = layer0_out[4755];
    assign layer1_out[2930] = ~layer0_out[5835];
    assign layer1_out[2931] = layer0_out[4609] & ~layer0_out[4608];
    assign layer1_out[2932] = ~layer0_out[739] | layer0_out[738];
    assign layer1_out[2933] = layer0_out[6084] | layer0_out[6085];
    assign layer1_out[2934] = ~layer0_out[6092];
    assign layer1_out[2935] = layer0_out[2827] & ~layer0_out[2826];
    assign layer1_out[2936] = layer0_out[2648] & ~layer0_out[2647];
    assign layer1_out[2937] = layer0_out[7580] & layer0_out[7581];
    assign layer1_out[2938] = layer0_out[2082];
    assign layer1_out[2939] = layer0_out[1706] | layer0_out[1707];
    assign layer1_out[2940] = ~layer0_out[6032];
    assign layer1_out[2941] = ~(layer0_out[4455] & layer0_out[4456]);
    assign layer1_out[2942] = 1'b0;
    assign layer1_out[2943] = ~layer0_out[3959];
    assign layer1_out[2944] = ~layer0_out[6045];
    assign layer1_out[2945] = 1'b1;
    assign layer1_out[2946] = layer0_out[5881];
    assign layer1_out[2947] = layer0_out[1255] & layer0_out[1256];
    assign layer1_out[2948] = layer0_out[4240];
    assign layer1_out[2949] = ~layer0_out[5585] | layer0_out[5584];
    assign layer1_out[2950] = ~layer0_out[2956];
    assign layer1_out[2951] = layer0_out[613] & layer0_out[614];
    assign layer1_out[2952] = layer0_out[5407] & ~layer0_out[5408];
    assign layer1_out[2953] = ~(layer0_out[1491] & layer0_out[1492]);
    assign layer1_out[2954] = ~layer0_out[7838];
    assign layer1_out[2955] = layer0_out[4301];
    assign layer1_out[2956] = layer0_out[5238] & ~layer0_out[5239];
    assign layer1_out[2957] = layer0_out[5341] & ~layer0_out[5340];
    assign layer1_out[2958] = ~(layer0_out[6478] | layer0_out[6479]);
    assign layer1_out[2959] = layer0_out[350] & ~layer0_out[351];
    assign layer1_out[2960] = layer0_out[1672];
    assign layer1_out[2961] = layer0_out[2959] & ~layer0_out[2960];
    assign layer1_out[2962] = layer0_out[7403];
    assign layer1_out[2963] = ~layer0_out[4951] | layer0_out[4952];
    assign layer1_out[2964] = layer0_out[2650] & ~layer0_out[2649];
    assign layer1_out[2965] = ~layer0_out[1649];
    assign layer1_out[2966] = 1'b1;
    assign layer1_out[2967] = ~layer0_out[5557];
    assign layer1_out[2968] = layer0_out[5384] & layer0_out[5385];
    assign layer1_out[2969] = ~(layer0_out[1637] & layer0_out[1638]);
    assign layer1_out[2970] = ~(layer0_out[1858] | layer0_out[1859]);
    assign layer1_out[2971] = layer0_out[2550] & ~layer0_out[2551];
    assign layer1_out[2972] = ~(layer0_out[3848] | layer0_out[3849]);
    assign layer1_out[2973] = ~(layer0_out[7612] | layer0_out[7613]);
    assign layer1_out[2974] = 1'b1;
    assign layer1_out[2975] = ~layer0_out[3467];
    assign layer1_out[2976] = layer0_out[6649] & layer0_out[6650];
    assign layer1_out[2977] = layer0_out[5419] | layer0_out[5420];
    assign layer1_out[2978] = 1'b1;
    assign layer1_out[2979] = ~(layer0_out[1766] | layer0_out[1767]);
    assign layer1_out[2980] = layer0_out[1023];
    assign layer1_out[2981] = ~(layer0_out[2614] | layer0_out[2615]);
    assign layer1_out[2982] = 1'b0;
    assign layer1_out[2983] = layer0_out[5000] & ~layer0_out[5001];
    assign layer1_out[2984] = layer0_out[147];
    assign layer1_out[2985] = layer0_out[6648] & layer0_out[6649];
    assign layer1_out[2986] = layer0_out[577] & layer0_out[578];
    assign layer1_out[2987] = layer0_out[4993];
    assign layer1_out[2988] = 1'b1;
    assign layer1_out[2989] = ~(layer0_out[5768] ^ layer0_out[5769]);
    assign layer1_out[2990] = 1'b1;
    assign layer1_out[2991] = ~(layer0_out[4394] ^ layer0_out[4395]);
    assign layer1_out[2992] = ~layer0_out[3136];
    assign layer1_out[2993] = layer0_out[6431];
    assign layer1_out[2994] = layer0_out[5438] & ~layer0_out[5439];
    assign layer1_out[2995] = layer0_out[7877];
    assign layer1_out[2996] = ~(layer0_out[6450] | layer0_out[6451]);
    assign layer1_out[2997] = ~(layer0_out[5635] | layer0_out[5636]);
    assign layer1_out[2998] = layer0_out[3275] | layer0_out[3276];
    assign layer1_out[2999] = layer0_out[2091] | layer0_out[2092];
    assign layer1_out[3000] = layer0_out[2133];
    assign layer1_out[3001] = layer0_out[3524] & ~layer0_out[3523];
    assign layer1_out[3002] = layer0_out[378];
    assign layer1_out[3003] = layer0_out[2902] & ~layer0_out[2901];
    assign layer1_out[3004] = ~layer0_out[5999];
    assign layer1_out[3005] = ~layer0_out[6080];
    assign layer1_out[3006] = 1'b1;
    assign layer1_out[3007] = layer0_out[1265];
    assign layer1_out[3008] = ~layer0_out[5515];
    assign layer1_out[3009] = 1'b1;
    assign layer1_out[3010] = layer0_out[5589];
    assign layer1_out[3011] = ~(layer0_out[24] ^ layer0_out[25]);
    assign layer1_out[3012] = layer0_out[2392] | layer0_out[2393];
    assign layer1_out[3013] = layer0_out[3803];
    assign layer1_out[3014] = ~(layer0_out[206] & layer0_out[207]);
    assign layer1_out[3015] = layer0_out[7013] & ~layer0_out[7012];
    assign layer1_out[3016] = layer0_out[990];
    assign layer1_out[3017] = layer0_out[6195] | layer0_out[6196];
    assign layer1_out[3018] = ~(layer0_out[3083] & layer0_out[3084]);
    assign layer1_out[3019] = ~layer0_out[3384];
    assign layer1_out[3020] = ~layer0_out[2831] | layer0_out[2830];
    assign layer1_out[3021] = ~layer0_out[3428] | layer0_out[3429];
    assign layer1_out[3022] = layer0_out[7980] & layer0_out[7981];
    assign layer1_out[3023] = layer0_out[6513];
    assign layer1_out[3024] = layer0_out[7292] & layer0_out[7293];
    assign layer1_out[3025] = ~layer0_out[7041];
    assign layer1_out[3026] = ~(layer0_out[6314] | layer0_out[6315]);
    assign layer1_out[3027] = layer0_out[6371] ^ layer0_out[6372];
    assign layer1_out[3028] = layer0_out[356];
    assign layer1_out[3029] = ~(layer0_out[4678] | layer0_out[4679]);
    assign layer1_out[3030] = layer0_out[4264] & ~layer0_out[4265];
    assign layer1_out[3031] = ~(layer0_out[4605] | layer0_out[4606]);
    assign layer1_out[3032] = ~layer0_out[2712];
    assign layer1_out[3033] = layer0_out[3829] & layer0_out[3830];
    assign layer1_out[3034] = layer0_out[30] & ~layer0_out[31];
    assign layer1_out[3035] = layer0_out[5207] & layer0_out[5208];
    assign layer1_out[3036] = layer0_out[6010] & ~layer0_out[6011];
    assign layer1_out[3037] = ~layer0_out[7078];
    assign layer1_out[3038] = layer0_out[5978] & layer0_out[5979];
    assign layer1_out[3039] = layer0_out[1195] & ~layer0_out[1194];
    assign layer1_out[3040] = layer0_out[3943] & ~layer0_out[3942];
    assign layer1_out[3041] = ~layer0_out[1198];
    assign layer1_out[3042] = ~(layer0_out[1869] & layer0_out[1870]);
    assign layer1_out[3043] = ~layer0_out[3226];
    assign layer1_out[3044] = layer0_out[54];
    assign layer1_out[3045] = 1'b1;
    assign layer1_out[3046] = layer0_out[892];
    assign layer1_out[3047] = layer0_out[423];
    assign layer1_out[3048] = ~(layer0_out[783] & layer0_out[784]);
    assign layer1_out[3049] = layer0_out[5670] & layer0_out[5671];
    assign layer1_out[3050] = layer0_out[1083] | layer0_out[1084];
    assign layer1_out[3051] = ~layer0_out[2759];
    assign layer1_out[3052] = ~layer0_out[4480];
    assign layer1_out[3053] = ~(layer0_out[3761] ^ layer0_out[3762]);
    assign layer1_out[3054] = layer0_out[5872] & ~layer0_out[5873];
    assign layer1_out[3055] = 1'b1;
    assign layer1_out[3056] = ~(layer0_out[4246] & layer0_out[4247]);
    assign layer1_out[3057] = ~layer0_out[6615];
    assign layer1_out[3058] = layer0_out[5104] | layer0_out[5105];
    assign layer1_out[3059] = ~layer0_out[7769] | layer0_out[7768];
    assign layer1_out[3060] = ~layer0_out[967];
    assign layer1_out[3061] = ~(layer0_out[7906] & layer0_out[7907]);
    assign layer1_out[3062] = layer0_out[7146];
    assign layer1_out[3063] = ~layer0_out[5353];
    assign layer1_out[3064] = layer0_out[3403] ^ layer0_out[3404];
    assign layer1_out[3065] = layer0_out[3663];
    assign layer1_out[3066] = layer0_out[526] | layer0_out[527];
    assign layer1_out[3067] = ~layer0_out[1169];
    assign layer1_out[3068] = layer0_out[5796] & ~layer0_out[5797];
    assign layer1_out[3069] = layer0_out[6337] & ~layer0_out[6338];
    assign layer1_out[3070] = layer0_out[390] & ~layer0_out[389];
    assign layer1_out[3071] = ~layer0_out[1534] | layer0_out[1533];
    assign layer1_out[3072] = ~layer0_out[6739];
    assign layer1_out[3073] = 1'b0;
    assign layer1_out[3074] = layer0_out[3091] & ~layer0_out[3090];
    assign layer1_out[3075] = ~(layer0_out[2948] & layer0_out[2949]);
    assign layer1_out[3076] = ~layer0_out[6841];
    assign layer1_out[3077] = ~layer0_out[1883];
    assign layer1_out[3078] = 1'b1;
    assign layer1_out[3079] = 1'b1;
    assign layer1_out[3080] = ~layer0_out[6375];
    assign layer1_out[3081] = ~layer0_out[5173] | layer0_out[5172];
    assign layer1_out[3082] = layer0_out[7151] & layer0_out[7152];
    assign layer1_out[3083] = layer0_out[7497] & layer0_out[7498];
    assign layer1_out[3084] = ~(layer0_out[1791] & layer0_out[1792]);
    assign layer1_out[3085] = ~layer0_out[7674];
    assign layer1_out[3086] = ~layer0_out[516];
    assign layer1_out[3087] = layer0_out[4009] ^ layer0_out[4010];
    assign layer1_out[3088] = layer0_out[1813] & ~layer0_out[1812];
    assign layer1_out[3089] = ~(layer0_out[5986] & layer0_out[5987]);
    assign layer1_out[3090] = 1'b0;
    assign layer1_out[3091] = layer0_out[6818];
    assign layer1_out[3092] = ~layer0_out[3521];
    assign layer1_out[3093] = ~layer0_out[6758] | layer0_out[6759];
    assign layer1_out[3094] = ~layer0_out[4555];
    assign layer1_out[3095] = ~layer0_out[7891] | layer0_out[7892];
    assign layer1_out[3096] = 1'b0;
    assign layer1_out[3097] = layer0_out[1069];
    assign layer1_out[3098] = ~layer0_out[7365];
    assign layer1_out[3099] = ~(layer0_out[1641] ^ layer0_out[1642]);
    assign layer1_out[3100] = layer0_out[4615];
    assign layer1_out[3101] = ~(layer0_out[2897] ^ layer0_out[2898]);
    assign layer1_out[3102] = layer0_out[4845];
    assign layer1_out[3103] = ~layer0_out[4415] | layer0_out[4414];
    assign layer1_out[3104] = ~layer0_out[3195];
    assign layer1_out[3105] = layer0_out[3537];
    assign layer1_out[3106] = ~(layer0_out[3216] | layer0_out[3217]);
    assign layer1_out[3107] = layer0_out[6718];
    assign layer1_out[3108] = layer0_out[3093] ^ layer0_out[3094];
    assign layer1_out[3109] = ~layer0_out[3818];
    assign layer1_out[3110] = ~(layer0_out[7938] | layer0_out[7939]);
    assign layer1_out[3111] = ~(layer0_out[3984] | layer0_out[3985]);
    assign layer1_out[3112] = ~layer0_out[6725];
    assign layer1_out[3113] = layer0_out[1139] & layer0_out[1140];
    assign layer1_out[3114] = ~layer0_out[7791] | layer0_out[7792];
    assign layer1_out[3115] = layer0_out[1084];
    assign layer1_out[3116] = layer0_out[1292] & ~layer0_out[1291];
    assign layer1_out[3117] = ~layer0_out[1801] | layer0_out[1800];
    assign layer1_out[3118] = ~layer0_out[7885];
    assign layer1_out[3119] = layer0_out[4732] | layer0_out[4733];
    assign layer1_out[3120] = ~layer0_out[7873] | layer0_out[7872];
    assign layer1_out[3121] = ~layer0_out[6668];
    assign layer1_out[3122] = ~layer0_out[4973] | layer0_out[4972];
    assign layer1_out[3123] = layer0_out[1841] & ~layer0_out[1842];
    assign layer1_out[3124] = layer0_out[5721] & ~layer0_out[5722];
    assign layer1_out[3125] = ~(layer0_out[952] ^ layer0_out[953]);
    assign layer1_out[3126] = layer0_out[5057] | layer0_out[5058];
    assign layer1_out[3127] = ~(layer0_out[5293] & layer0_out[5294]);
    assign layer1_out[3128] = layer0_out[1312] & ~layer0_out[1311];
    assign layer1_out[3129] = layer0_out[5911];
    assign layer1_out[3130] = ~(layer0_out[7066] & layer0_out[7067]);
    assign layer1_out[3131] = layer0_out[2899] & layer0_out[2900];
    assign layer1_out[3132] = ~(layer0_out[497] & layer0_out[498]);
    assign layer1_out[3133] = ~layer0_out[2545] | layer0_out[2544];
    assign layer1_out[3134] = ~layer0_out[4548] | layer0_out[4547];
    assign layer1_out[3135] = ~layer0_out[4225];
    assign layer1_out[3136] = layer0_out[677];
    assign layer1_out[3137] = layer0_out[1254] & layer0_out[1255];
    assign layer1_out[3138] = layer0_out[4594] & layer0_out[4595];
    assign layer1_out[3139] = ~layer0_out[700];
    assign layer1_out[3140] = layer0_out[4193];
    assign layer1_out[3141] = layer0_out[3536] & layer0_out[3537];
    assign layer1_out[3142] = ~layer0_out[7142] | layer0_out[7143];
    assign layer1_out[3143] = layer0_out[3621] & layer0_out[3622];
    assign layer1_out[3144] = layer0_out[271] & ~layer0_out[270];
    assign layer1_out[3145] = ~layer0_out[1838];
    assign layer1_out[3146] = layer0_out[4038] & layer0_out[4039];
    assign layer1_out[3147] = layer0_out[3379];
    assign layer1_out[3148] = ~layer0_out[3286] | layer0_out[3287];
    assign layer1_out[3149] = layer0_out[6685];
    assign layer1_out[3150] = layer0_out[1776];
    assign layer1_out[3151] = layer0_out[334] & layer0_out[335];
    assign layer1_out[3152] = ~(layer0_out[4615] & layer0_out[4616]);
    assign layer1_out[3153] = layer0_out[2320] ^ layer0_out[2321];
    assign layer1_out[3154] = layer0_out[6100];
    assign layer1_out[3155] = layer0_out[6573] & ~layer0_out[6572];
    assign layer1_out[3156] = layer0_out[6070] & ~layer0_out[6071];
    assign layer1_out[3157] = ~layer0_out[374] | layer0_out[373];
    assign layer1_out[3158] = layer0_out[5201] & ~layer0_out[5202];
    assign layer1_out[3159] = ~(layer0_out[3147] | layer0_out[3148]);
    assign layer1_out[3160] = layer0_out[7225] & ~layer0_out[7226];
    assign layer1_out[3161] = ~layer0_out[4627];
    assign layer1_out[3162] = layer0_out[2667];
    assign layer1_out[3163] = layer0_out[6042] & layer0_out[6043];
    assign layer1_out[3164] = layer0_out[6095] & ~layer0_out[6094];
    assign layer1_out[3165] = ~layer0_out[1833];
    assign layer1_out[3166] = ~layer0_out[3889];
    assign layer1_out[3167] = layer0_out[957];
    assign layer1_out[3168] = ~layer0_out[5373];
    assign layer1_out[3169] = ~layer0_out[7];
    assign layer1_out[3170] = 1'b1;
    assign layer1_out[3171] = ~layer0_out[2226] | layer0_out[2225];
    assign layer1_out[3172] = ~layer0_out[1394];
    assign layer1_out[3173] = ~(layer0_out[7080] | layer0_out[7081]);
    assign layer1_out[3174] = ~layer0_out[4467];
    assign layer1_out[3175] = ~(layer0_out[113] | layer0_out[114]);
    assign layer1_out[3176] = ~(layer0_out[7715] | layer0_out[7716]);
    assign layer1_out[3177] = layer0_out[4378] & layer0_out[4379];
    assign layer1_out[3178] = layer0_out[3241] ^ layer0_out[3242];
    assign layer1_out[3179] = ~layer0_out[6217] | layer0_out[6216];
    assign layer1_out[3180] = ~layer0_out[2141] | layer0_out[2140];
    assign layer1_out[3181] = ~layer0_out[6552];
    assign layer1_out[3182] = layer0_out[6574];
    assign layer1_out[3183] = ~layer0_out[2626] | layer0_out[2625];
    assign layer1_out[3184] = ~(layer0_out[4579] & layer0_out[4580]);
    assign layer1_out[3185] = ~layer0_out[3197] | layer0_out[3196];
    assign layer1_out[3186] = 1'b0;
    assign layer1_out[3187] = layer0_out[7636];
    assign layer1_out[3188] = ~(layer0_out[7916] ^ layer0_out[7917]);
    assign layer1_out[3189] = ~layer0_out[3571];
    assign layer1_out[3190] = layer0_out[6413] & ~layer0_out[6414];
    assign layer1_out[3191] = ~(layer0_out[5706] & layer0_out[5707]);
    assign layer1_out[3192] = layer0_out[4389] & ~layer0_out[4390];
    assign layer1_out[3193] = ~(layer0_out[2810] ^ layer0_out[2811]);
    assign layer1_out[3194] = ~layer0_out[1203];
    assign layer1_out[3195] = ~layer0_out[934] | layer0_out[933];
    assign layer1_out[3196] = layer0_out[2233] & ~layer0_out[2232];
    assign layer1_out[3197] = layer0_out[2648];
    assign layer1_out[3198] = ~layer0_out[5976];
    assign layer1_out[3199] = layer0_out[6403] & layer0_out[6404];
    assign layer1_out[3200] = layer0_out[6416];
    assign layer1_out[3201] = ~(layer0_out[2532] | layer0_out[2533]);
    assign layer1_out[3202] = ~layer0_out[4067];
    assign layer1_out[3203] = layer0_out[5291];
    assign layer1_out[3204] = ~layer0_out[5786] | layer0_out[5787];
    assign layer1_out[3205] = ~layer0_out[2403] | layer0_out[2404];
    assign layer1_out[3206] = layer0_out[6350];
    assign layer1_out[3207] = layer0_out[3153] & layer0_out[3154];
    assign layer1_out[3208] = ~layer0_out[4426];
    assign layer1_out[3209] = layer0_out[7564];
    assign layer1_out[3210] = layer0_out[1527] & ~layer0_out[1526];
    assign layer1_out[3211] = layer0_out[2984] & layer0_out[2985];
    assign layer1_out[3212] = layer0_out[4316] | layer0_out[4317];
    assign layer1_out[3213] = ~(layer0_out[594] & layer0_out[595]);
    assign layer1_out[3214] = ~layer0_out[1140] | layer0_out[1141];
    assign layer1_out[3215] = layer0_out[1370] | layer0_out[1371];
    assign layer1_out[3216] = 1'b1;
    assign layer1_out[3217] = ~layer0_out[1238];
    assign layer1_out[3218] = layer0_out[7544];
    assign layer1_out[3219] = ~(layer0_out[7888] | layer0_out[7889]);
    assign layer1_out[3220] = ~(layer0_out[7670] & layer0_out[7671]);
    assign layer1_out[3221] = layer0_out[6148] ^ layer0_out[6149];
    assign layer1_out[3222] = ~layer0_out[874];
    assign layer1_out[3223] = ~(layer0_out[25] | layer0_out[26]);
    assign layer1_out[3224] = ~(layer0_out[1472] & layer0_out[1473]);
    assign layer1_out[3225] = ~layer0_out[2827] | layer0_out[2828];
    assign layer1_out[3226] = ~layer0_out[2719] | layer0_out[2720];
    assign layer1_out[3227] = layer0_out[6410] & layer0_out[6411];
    assign layer1_out[3228] = ~layer0_out[4710];
    assign layer1_out[3229] = ~layer0_out[6868];
    assign layer1_out[3230] = layer0_out[6806] & layer0_out[6807];
    assign layer1_out[3231] = ~(layer0_out[7514] & layer0_out[7515]);
    assign layer1_out[3232] = ~layer0_out[6510] | layer0_out[6511];
    assign layer1_out[3233] = layer0_out[3751] & ~layer0_out[3752];
    assign layer1_out[3234] = 1'b0;
    assign layer1_out[3235] = layer0_out[3955];
    assign layer1_out[3236] = layer0_out[7005];
    assign layer1_out[3237] = ~layer0_out[2217];
    assign layer1_out[3238] = layer0_out[1599];
    assign layer1_out[3239] = layer0_out[7653] & ~layer0_out[7652];
    assign layer1_out[3240] = 1'b0;
    assign layer1_out[3241] = ~(layer0_out[5649] & layer0_out[5650]);
    assign layer1_out[3242] = ~layer0_out[1157];
    assign layer1_out[3243] = layer0_out[497];
    assign layer1_out[3244] = layer0_out[7322] | layer0_out[7323];
    assign layer1_out[3245] = layer0_out[1079] & layer0_out[1080];
    assign layer1_out[3246] = 1'b1;
    assign layer1_out[3247] = layer0_out[6102];
    assign layer1_out[3248] = layer0_out[6875] & ~layer0_out[6874];
    assign layer1_out[3249] = ~(layer0_out[6193] | layer0_out[6194]);
    assign layer1_out[3250] = ~(layer0_out[7626] | layer0_out[7627]);
    assign layer1_out[3251] = layer0_out[2950];
    assign layer1_out[3252] = ~(layer0_out[5671] | layer0_out[5672]);
    assign layer1_out[3253] = ~layer0_out[822];
    assign layer1_out[3254] = layer0_out[1577] | layer0_out[1578];
    assign layer1_out[3255] = layer0_out[1712] & layer0_out[1713];
    assign layer1_out[3256] = ~(layer0_out[3846] & layer0_out[3847]);
    assign layer1_out[3257] = ~(layer0_out[3824] | layer0_out[3825]);
    assign layer1_out[3258] = layer0_out[5049] | layer0_out[5050];
    assign layer1_out[3259] = ~layer0_out[7392];
    assign layer1_out[3260] = layer0_out[1224];
    assign layer1_out[3261] = ~(layer0_out[7455] | layer0_out[7456]);
    assign layer1_out[3262] = layer0_out[5066];
    assign layer1_out[3263] = ~layer0_out[3466];
    assign layer1_out[3264] = ~(layer0_out[1309] | layer0_out[1310]);
    assign layer1_out[3265] = layer0_out[5548];
    assign layer1_out[3266] = ~layer0_out[6713];
    assign layer1_out[3267] = ~(layer0_out[1663] ^ layer0_out[1664]);
    assign layer1_out[3268] = ~(layer0_out[7229] & layer0_out[7230]);
    assign layer1_out[3269] = layer0_out[4507];
    assign layer1_out[3270] = ~layer0_out[953];
    assign layer1_out[3271] = ~layer0_out[7121];
    assign layer1_out[3272] = 1'b1;
    assign layer1_out[3273] = layer0_out[3981] & ~layer0_out[3982];
    assign layer1_out[3274] = ~(layer0_out[4728] & layer0_out[4729]);
    assign layer1_out[3275] = layer0_out[4574] | layer0_out[4575];
    assign layer1_out[3276] = layer0_out[1547];
    assign layer1_out[3277] = layer0_out[572] & layer0_out[573];
    assign layer1_out[3278] = layer0_out[4262] | layer0_out[4263];
    assign layer1_out[3279] = layer0_out[4542] & ~layer0_out[4541];
    assign layer1_out[3280] = ~(layer0_out[5969] | layer0_out[5970]);
    assign layer1_out[3281] = ~layer0_out[6444];
    assign layer1_out[3282] = layer0_out[6604] & ~layer0_out[6605];
    assign layer1_out[3283] = 1'b0;
    assign layer1_out[3284] = layer0_out[719] ^ layer0_out[720];
    assign layer1_out[3285] = layer0_out[4332];
    assign layer1_out[3286] = ~layer0_out[2164];
    assign layer1_out[3287] = ~(layer0_out[4449] & layer0_out[4450]);
    assign layer1_out[3288] = ~layer0_out[1721];
    assign layer1_out[3289] = ~layer0_out[7420];
    assign layer1_out[3290] = layer0_out[4287];
    assign layer1_out[3291] = ~layer0_out[4866];
    assign layer1_out[3292] = layer0_out[3482];
    assign layer1_out[3293] = layer0_out[295] | layer0_out[296];
    assign layer1_out[3294] = layer0_out[5176] & ~layer0_out[5175];
    assign layer1_out[3295] = ~(layer0_out[254] & layer0_out[255]);
    assign layer1_out[3296] = ~layer0_out[2126];
    assign layer1_out[3297] = ~(layer0_out[2409] | layer0_out[2410]);
    assign layer1_out[3298] = ~(layer0_out[2528] | layer0_out[2529]);
    assign layer1_out[3299] = layer0_out[4312] ^ layer0_out[4313];
    assign layer1_out[3300] = layer0_out[1034];
    assign layer1_out[3301] = ~(layer0_out[1217] & layer0_out[1218]);
    assign layer1_out[3302] = ~layer0_out[717];
    assign layer1_out[3303] = ~(layer0_out[4045] & layer0_out[4046]);
    assign layer1_out[3304] = ~(layer0_out[4929] | layer0_out[4930]);
    assign layer1_out[3305] = layer0_out[4598];
    assign layer1_out[3306] = 1'b1;
    assign layer1_out[3307] = 1'b1;
    assign layer1_out[3308] = ~layer0_out[5038];
    assign layer1_out[3309] = layer0_out[7554];
    assign layer1_out[3310] = ~layer0_out[1301] | layer0_out[1300];
    assign layer1_out[3311] = layer0_out[2573] ^ layer0_out[2574];
    assign layer1_out[3312] = ~layer0_out[5276];
    assign layer1_out[3313] = layer0_out[4155] & ~layer0_out[4156];
    assign layer1_out[3314] = layer0_out[2733] & ~layer0_out[2732];
    assign layer1_out[3315] = layer0_out[3837];
    assign layer1_out[3316] = ~layer0_out[6859] | layer0_out[6860];
    assign layer1_out[3317] = layer0_out[3911] & ~layer0_out[3910];
    assign layer1_out[3318] = layer0_out[740] | layer0_out[741];
    assign layer1_out[3319] = layer0_out[2734];
    assign layer1_out[3320] = ~layer0_out[1402];
    assign layer1_out[3321] = layer0_out[1476];
    assign layer1_out[3322] = layer0_out[2644];
    assign layer1_out[3323] = layer0_out[2398] | layer0_out[2399];
    assign layer1_out[3324] = ~(layer0_out[2695] & layer0_out[2696]);
    assign layer1_out[3325] = layer0_out[5680];
    assign layer1_out[3326] = layer0_out[5927];
    assign layer1_out[3327] = ~(layer0_out[5820] & layer0_out[5821]);
    assign layer1_out[3328] = ~layer0_out[429];
    assign layer1_out[3329] = layer0_out[5253] & ~layer0_out[5252];
    assign layer1_out[3330] = ~layer0_out[913];
    assign layer1_out[3331] = layer0_out[415] & ~layer0_out[414];
    assign layer1_out[3332] = layer0_out[5659];
    assign layer1_out[3333] = layer0_out[951] & layer0_out[952];
    assign layer1_out[3334] = layer0_out[7370] | layer0_out[7371];
    assign layer1_out[3335] = ~layer0_out[4832] | layer0_out[4833];
    assign layer1_out[3336] = layer0_out[3857] & ~layer0_out[3856];
    assign layer1_out[3337] = 1'b0;
    assign layer1_out[3338] = layer0_out[2292];
    assign layer1_out[3339] = layer0_out[7077];
    assign layer1_out[3340] = ~(layer0_out[5826] & layer0_out[5827]);
    assign layer1_out[3341] = layer0_out[7231];
    assign layer1_out[3342] = layer0_out[5117] ^ layer0_out[5118];
    assign layer1_out[3343] = ~(layer0_out[4323] & layer0_out[4324]);
    assign layer1_out[3344] = ~layer0_out[7866] | layer0_out[7867];
    assign layer1_out[3345] = layer0_out[4137] | layer0_out[4138];
    assign layer1_out[3346] = ~layer0_out[7532];
    assign layer1_out[3347] = ~layer0_out[1338];
    assign layer1_out[3348] = ~layer0_out[6922] | layer0_out[6921];
    assign layer1_out[3349] = ~layer0_out[6712] | layer0_out[6713];
    assign layer1_out[3350] = layer0_out[7685] | layer0_out[7686];
    assign layer1_out[3351] = layer0_out[2844] & layer0_out[2845];
    assign layer1_out[3352] = ~layer0_out[5074] | layer0_out[5073];
    assign layer1_out[3353] = layer0_out[7749];
    assign layer1_out[3354] = layer0_out[1037] & layer0_out[1038];
    assign layer1_out[3355] = layer0_out[5239] & layer0_out[5240];
    assign layer1_out[3356] = ~layer0_out[2941];
    assign layer1_out[3357] = ~layer0_out[1875];
    assign layer1_out[3358] = ~(layer0_out[3036] ^ layer0_out[3037]);
    assign layer1_out[3359] = layer0_out[6631];
    assign layer1_out[3360] = layer0_out[935];
    assign layer1_out[3361] = layer0_out[3463];
    assign layer1_out[3362] = layer0_out[7246];
    assign layer1_out[3363] = ~(layer0_out[5052] | layer0_out[5053]);
    assign layer1_out[3364] = layer0_out[889] & layer0_out[890];
    assign layer1_out[3365] = 1'b0;
    assign layer1_out[3366] = layer0_out[6600] ^ layer0_out[6601];
    assign layer1_out[3367] = layer0_out[1256] & ~layer0_out[1257];
    assign layer1_out[3368] = layer0_out[3525] | layer0_out[3526];
    assign layer1_out[3369] = ~layer0_out[3809];
    assign layer1_out[3370] = ~layer0_out[7598];
    assign layer1_out[3371] = layer0_out[1960];
    assign layer1_out[3372] = ~layer0_out[3072] | layer0_out[3071];
    assign layer1_out[3373] = ~(layer0_out[6415] | layer0_out[6416]);
    assign layer1_out[3374] = layer0_out[7252];
    assign layer1_out[3375] = 1'b1;
    assign layer1_out[3376] = ~layer0_out[970] | layer0_out[969];
    assign layer1_out[3377] = ~(layer0_out[114] | layer0_out[115]);
    assign layer1_out[3378] = ~layer0_out[5299];
    assign layer1_out[3379] = ~layer0_out[180];
    assign layer1_out[3380] = layer0_out[1715] & layer0_out[1716];
    assign layer1_out[3381] = ~(layer0_out[6447] & layer0_out[6448]);
    assign layer1_out[3382] = layer0_out[6154] | layer0_out[6155];
    assign layer1_out[3383] = layer0_out[3429] & ~layer0_out[3430];
    assign layer1_out[3384] = layer0_out[2939] | layer0_out[2940];
    assign layer1_out[3385] = 1'b0;
    assign layer1_out[3386] = ~(layer0_out[6295] | layer0_out[6296]);
    assign layer1_out[3387] = layer0_out[950] & ~layer0_out[949];
    assign layer1_out[3388] = layer0_out[3000] | layer0_out[3001];
    assign layer1_out[3389] = layer0_out[1684] & ~layer0_out[1683];
    assign layer1_out[3390] = layer0_out[221] & ~layer0_out[220];
    assign layer1_out[3391] = layer0_out[5316];
    assign layer1_out[3392] = layer0_out[3897] & layer0_out[3898];
    assign layer1_out[3393] = ~layer0_out[7767] | layer0_out[7766];
    assign layer1_out[3394] = layer0_out[4983];
    assign layer1_out[3395] = layer0_out[5446] & ~layer0_out[5447];
    assign layer1_out[3396] = ~layer0_out[1847] | layer0_out[1848];
    assign layer1_out[3397] = layer0_out[7188] | layer0_out[7189];
    assign layer1_out[3398] = layer0_out[1734];
    assign layer1_out[3399] = ~layer0_out[5839] | layer0_out[5838];
    assign layer1_out[3400] = 1'b1;
    assign layer1_out[3401] = ~layer0_out[3267] | layer0_out[3266];
    assign layer1_out[3402] = ~layer0_out[1535];
    assign layer1_out[3403] = ~layer0_out[5275];
    assign layer1_out[3404] = layer0_out[2446] | layer0_out[2447];
    assign layer1_out[3405] = ~layer0_out[7221];
    assign layer1_out[3406] = ~layer0_out[4971];
    assign layer1_out[3407] = layer0_out[926];
    assign layer1_out[3408] = ~layer0_out[4636];
    assign layer1_out[3409] = layer0_out[6233];
    assign layer1_out[3410] = layer0_out[1444] & layer0_out[1445];
    assign layer1_out[3411] = ~(layer0_out[2964] | layer0_out[2965]);
    assign layer1_out[3412] = layer0_out[5845];
    assign layer1_out[3413] = ~(layer0_out[7007] & layer0_out[7008]);
    assign layer1_out[3414] = layer0_out[3912] & ~layer0_out[3913];
    assign layer1_out[3415] = 1'b1;
    assign layer1_out[3416] = ~layer0_out[6115] | layer0_out[6114];
    assign layer1_out[3417] = ~(layer0_out[3908] ^ layer0_out[3909]);
    assign layer1_out[3418] = ~(layer0_out[5729] ^ layer0_out[5730]);
    assign layer1_out[3419] = ~layer0_out[3555];
    assign layer1_out[3420] = ~layer0_out[4676] | layer0_out[4677];
    assign layer1_out[3421] = layer0_out[129] & layer0_out[130];
    assign layer1_out[3422] = ~layer0_out[3092] | layer0_out[3091];
    assign layer1_out[3423] = ~layer0_out[4021] | layer0_out[4020];
    assign layer1_out[3424] = ~layer0_out[4579] | layer0_out[4578];
    assign layer1_out[3425] = ~layer0_out[2895] | layer0_out[2896];
    assign layer1_out[3426] = ~layer0_out[856];
    assign layer1_out[3427] = layer0_out[6737] & ~layer0_out[6736];
    assign layer1_out[3428] = layer0_out[7546] & ~layer0_out[7545];
    assign layer1_out[3429] = 1'b1;
    assign layer1_out[3430] = ~(layer0_out[6612] & layer0_out[6613]);
    assign layer1_out[3431] = ~layer0_out[2933] | layer0_out[2934];
    assign layer1_out[3432] = ~(layer0_out[3468] & layer0_out[3469]);
    assign layer1_out[3433] = layer0_out[5426] ^ layer0_out[5427];
    assign layer1_out[3434] = layer0_out[7975] ^ layer0_out[7976];
    assign layer1_out[3435] = layer0_out[326] & ~layer0_out[327];
    assign layer1_out[3436] = ~(layer0_out[615] ^ layer0_out[616]);
    assign layer1_out[3437] = ~layer0_out[6676] | layer0_out[6677];
    assign layer1_out[3438] = layer0_out[3407] & layer0_out[3408];
    assign layer1_out[3439] = ~(layer0_out[1778] & layer0_out[1779]);
    assign layer1_out[3440] = layer0_out[4147] & ~layer0_out[4146];
    assign layer1_out[3441] = layer0_out[956];
    assign layer1_out[3442] = layer0_out[7048];
    assign layer1_out[3443] = ~layer0_out[7090] | layer0_out[7091];
    assign layer1_out[3444] = layer0_out[1719];
    assign layer1_out[3445] = 1'b1;
    assign layer1_out[3446] = ~layer0_out[861];
    assign layer1_out[3447] = ~layer0_out[5257] | layer0_out[5258];
    assign layer1_out[3448] = layer0_out[1884] | layer0_out[1885];
    assign layer1_out[3449] = layer0_out[6291];
    assign layer1_out[3450] = ~(layer0_out[2347] | layer0_out[2348]);
    assign layer1_out[3451] = ~(layer0_out[2891] & layer0_out[2892]);
    assign layer1_out[3452] = layer0_out[3575];
    assign layer1_out[3453] = ~(layer0_out[5137] ^ layer0_out[5138]);
    assign layer1_out[3454] = layer0_out[3584];
    assign layer1_out[3455] = layer0_out[7997];
    assign layer1_out[3456] = 1'b0;
    assign layer1_out[3457] = ~(layer0_out[2716] & layer0_out[2717]);
    assign layer1_out[3458] = layer0_out[4824] | layer0_out[4825];
    assign layer1_out[3459] = layer0_out[4600] & ~layer0_out[4601];
    assign layer1_out[3460] = layer0_out[6828];
    assign layer1_out[3461] = ~layer0_out[6339];
    assign layer1_out[3462] = ~(layer0_out[643] ^ layer0_out[644]);
    assign layer1_out[3463] = layer0_out[3353] | layer0_out[3354];
    assign layer1_out[3464] = 1'b0;
    assign layer1_out[3465] = ~layer0_out[5670];
    assign layer1_out[3466] = layer0_out[6823] & ~layer0_out[6822];
    assign layer1_out[3467] = ~layer0_out[3251] | layer0_out[3250];
    assign layer1_out[3468] = layer0_out[443] & ~layer0_out[444];
    assign layer1_out[3469] = layer0_out[1139] & ~layer0_out[1138];
    assign layer1_out[3470] = layer0_out[6749];
    assign layer1_out[3471] = layer0_out[5300] | layer0_out[5301];
    assign layer1_out[3472] = ~layer0_out[1050] | layer0_out[1049];
    assign layer1_out[3473] = ~layer0_out[3210];
    assign layer1_out[3474] = ~layer0_out[2987];
    assign layer1_out[3475] = layer0_out[1030] | layer0_out[1031];
    assign layer1_out[3476] = layer0_out[2019] & ~layer0_out[2020];
    assign layer1_out[3477] = layer0_out[3613];
    assign layer1_out[3478] = layer0_out[4504] & layer0_out[4505];
    assign layer1_out[3479] = layer0_out[7272] | layer0_out[7273];
    assign layer1_out[3480] = ~(layer0_out[6691] | layer0_out[6692]);
    assign layer1_out[3481] = layer0_out[2215];
    assign layer1_out[3482] = layer0_out[5893];
    assign layer1_out[3483] = ~layer0_out[7980];
    assign layer1_out[3484] = ~layer0_out[5622] | layer0_out[5621];
    assign layer1_out[3485] = layer0_out[5361] & layer0_out[5362];
    assign layer1_out[3486] = 1'b1;
    assign layer1_out[3487] = layer0_out[2317] & ~layer0_out[2316];
    assign layer1_out[3488] = layer0_out[354];
    assign layer1_out[3489] = ~layer0_out[1939];
    assign layer1_out[3490] = ~layer0_out[4109];
    assign layer1_out[3491] = layer0_out[3753];
    assign layer1_out[3492] = 1'b0;
    assign layer1_out[3493] = layer0_out[6814] & ~layer0_out[6813];
    assign layer1_out[3494] = ~layer0_out[662];
    assign layer1_out[3495] = layer0_out[6022] & ~layer0_out[6021];
    assign layer1_out[3496] = layer0_out[1771] ^ layer0_out[1772];
    assign layer1_out[3497] = ~layer0_out[825];
    assign layer1_out[3498] = layer0_out[1623];
    assign layer1_out[3499] = ~(layer0_out[7216] | layer0_out[7217]);
    assign layer1_out[3500] = layer0_out[7663];
    assign layer1_out[3501] = ~(layer0_out[1426] | layer0_out[1427]);
    assign layer1_out[3502] = layer0_out[5651];
    assign layer1_out[3503] = ~layer0_out[1072] | layer0_out[1071];
    assign layer1_out[3504] = ~(layer0_out[4448] | layer0_out[4449]);
    assign layer1_out[3505] = ~layer0_out[6321];
    assign layer1_out[3506] = layer0_out[7708] & layer0_out[7709];
    assign layer1_out[3507] = 1'b1;
    assign layer1_out[3508] = layer0_out[2682];
    assign layer1_out[3509] = ~layer0_out[6371];
    assign layer1_out[3510] = ~layer0_out[2027] | layer0_out[2026];
    assign layer1_out[3511] = ~(layer0_out[1799] ^ layer0_out[1800]);
    assign layer1_out[3512] = 1'b1;
    assign layer1_out[3513] = ~layer0_out[4802] | layer0_out[4803];
    assign layer1_out[3514] = ~(layer0_out[1898] | layer0_out[1899]);
    assign layer1_out[3515] = ~layer0_out[6923] | layer0_out[6922];
    assign layer1_out[3516] = ~layer0_out[3308] | layer0_out[3309];
    assign layer1_out[3517] = layer0_out[2659];
    assign layer1_out[3518] = layer0_out[5518] & ~layer0_out[5519];
    assign layer1_out[3519] = layer0_out[2974];
    assign layer1_out[3520] = layer0_out[574];
    assign layer1_out[3521] = ~layer0_out[412] | layer0_out[413];
    assign layer1_out[3522] = ~layer0_out[5185] | layer0_out[5186];
    assign layer1_out[3523] = ~layer0_out[7088] | layer0_out[7087];
    assign layer1_out[3524] = 1'b0;
    assign layer1_out[3525] = ~(layer0_out[7318] | layer0_out[7319]);
    assign layer1_out[3526] = ~layer0_out[3817] | layer0_out[3816];
    assign layer1_out[3527] = ~layer0_out[1158];
    assign layer1_out[3528] = ~(layer0_out[6442] | layer0_out[6443]);
    assign layer1_out[3529] = layer0_out[2982] & layer0_out[2983];
    assign layer1_out[3530] = layer0_out[6863];
    assign layer1_out[3531] = ~(layer0_out[3722] | layer0_out[3723]);
    assign layer1_out[3532] = ~(layer0_out[3593] & layer0_out[3594]);
    assign layer1_out[3533] = layer0_out[4551];
    assign layer1_out[3534] = layer0_out[3045] & layer0_out[3046];
    assign layer1_out[3535] = ~layer0_out[5852] | layer0_out[5851];
    assign layer1_out[3536] = 1'b1;
    assign layer1_out[3537] = 1'b1;
    assign layer1_out[3538] = ~(layer0_out[184] | layer0_out[185]);
    assign layer1_out[3539] = layer0_out[6646] & ~layer0_out[6647];
    assign layer1_out[3540] = ~(layer0_out[5985] | layer0_out[5986]);
    assign layer1_out[3541] = ~layer0_out[1877] | layer0_out[1876];
    assign layer1_out[3542] = layer0_out[820] & layer0_out[821];
    assign layer1_out[3543] = layer0_out[3111];
    assign layer1_out[3544] = 1'b0;
    assign layer1_out[3545] = layer0_out[5055];
    assign layer1_out[3546] = ~(layer0_out[355] ^ layer0_out[356]);
    assign layer1_out[3547] = 1'b0;
    assign layer1_out[3548] = layer0_out[4964];
    assign layer1_out[3549] = layer0_out[1069] | layer0_out[1070];
    assign layer1_out[3550] = layer0_out[6001];
    assign layer1_out[3551] = layer0_out[6665] ^ layer0_out[6666];
    assign layer1_out[3552] = ~layer0_out[6186];
    assign layer1_out[3553] = ~layer0_out[5025];
    assign layer1_out[3554] = layer0_out[786] & ~layer0_out[787];
    assign layer1_out[3555] = ~(layer0_out[3433] & layer0_out[3434]);
    assign layer1_out[3556] = ~(layer0_out[1326] ^ layer0_out[1327]);
    assign layer1_out[3557] = layer0_out[239];
    assign layer1_out[3558] = ~(layer0_out[5601] | layer0_out[5602]);
    assign layer1_out[3559] = ~layer0_out[5447] | layer0_out[5448];
    assign layer1_out[3560] = layer0_out[662] ^ layer0_out[663];
    assign layer1_out[3561] = layer0_out[1976];
    assign layer1_out[3562] = layer0_out[6699] & layer0_out[6700];
    assign layer1_out[3563] = layer0_out[4837] & ~layer0_out[4836];
    assign layer1_out[3564] = ~(layer0_out[6709] & layer0_out[6710]);
    assign layer1_out[3565] = layer0_out[7169];
    assign layer1_out[3566] = layer0_out[6219] & ~layer0_out[6220];
    assign layer1_out[3567] = ~layer0_out[1541] | layer0_out[1540];
    assign layer1_out[3568] = layer0_out[3115] ^ layer0_out[3116];
    assign layer1_out[3569] = layer0_out[6978] | layer0_out[6979];
    assign layer1_out[3570] = layer0_out[6470] & ~layer0_out[6471];
    assign layer1_out[3571] = layer0_out[6589] | layer0_out[6590];
    assign layer1_out[3572] = ~layer0_out[4491];
    assign layer1_out[3573] = ~layer0_out[7048];
    assign layer1_out[3574] = ~layer0_out[5989];
    assign layer1_out[3575] = layer0_out[5237] & ~layer0_out[5236];
    assign layer1_out[3576] = layer0_out[1640];
    assign layer1_out[3577] = layer0_out[4954] | layer0_out[4955];
    assign layer1_out[3578] = ~(layer0_out[2990] | layer0_out[2991]);
    assign layer1_out[3579] = ~layer0_out[5758];
    assign layer1_out[3580] = 1'b0;
    assign layer1_out[3581] = ~layer0_out[7542];
    assign layer1_out[3582] = ~layer0_out[6079];
    assign layer1_out[3583] = ~layer0_out[5385];
    assign layer1_out[3584] = ~(layer0_out[6846] | layer0_out[6847]);
    assign layer1_out[3585] = layer0_out[629] & layer0_out[630];
    assign layer1_out[3586] = ~layer0_out[7389] | layer0_out[7390];
    assign layer1_out[3587] = ~(layer0_out[3475] & layer0_out[3476]);
    assign layer1_out[3588] = ~layer0_out[5286];
    assign layer1_out[3589] = layer0_out[2202] | layer0_out[2203];
    assign layer1_out[3590] = layer0_out[795] & ~layer0_out[796];
    assign layer1_out[3591] = ~layer0_out[7566];
    assign layer1_out[3592] = layer0_out[6755];
    assign layer1_out[3593] = layer0_out[1957];
    assign layer1_out[3594] = ~layer0_out[7818] | layer0_out[7817];
    assign layer1_out[3595] = layer0_out[1906] & layer0_out[1907];
    assign layer1_out[3596] = layer0_out[4195] ^ layer0_out[4196];
    assign layer1_out[3597] = ~(layer0_out[6155] & layer0_out[6156]);
    assign layer1_out[3598] = ~layer0_out[3458];
    assign layer1_out[3599] = ~(layer0_out[7276] ^ layer0_out[7277]);
    assign layer1_out[3600] = layer0_out[6620] & ~layer0_out[6619];
    assign layer1_out[3601] = layer0_out[6504];
    assign layer1_out[3602] = ~layer0_out[7655] | layer0_out[7654];
    assign layer1_out[3603] = ~layer0_out[660];
    assign layer1_out[3604] = ~layer0_out[1999] | layer0_out[2000];
    assign layer1_out[3605] = layer0_out[7690] & ~layer0_out[7689];
    assign layer1_out[3606] = layer0_out[6955] | layer0_out[6956];
    assign layer1_out[3607] = ~layer0_out[2541];
    assign layer1_out[3608] = layer0_out[4085] & ~layer0_out[4084];
    assign layer1_out[3609] = ~(layer0_out[46] ^ layer0_out[47]);
    assign layer1_out[3610] = ~layer0_out[1677] | layer0_out[1678];
    assign layer1_out[3611] = ~layer0_out[1375] | layer0_out[1374];
    assign layer1_out[3612] = ~layer0_out[2774] | layer0_out[2773];
    assign layer1_out[3613] = layer0_out[4509] & ~layer0_out[4508];
    assign layer1_out[3614] = layer0_out[1144] & ~layer0_out[1143];
    assign layer1_out[3615] = ~layer0_out[3945];
    assign layer1_out[3616] = layer0_out[7984] & layer0_out[7985];
    assign layer1_out[3617] = layer0_out[1533];
    assign layer1_out[3618] = ~layer0_out[6545];
    assign layer1_out[3619] = ~layer0_out[5983] | layer0_out[5984];
    assign layer1_out[3620] = layer0_out[7316] & layer0_out[7317];
    assign layer1_out[3621] = ~layer0_out[7698] | layer0_out[7699];
    assign layer1_out[3622] = 1'b0;
    assign layer1_out[3623] = ~layer0_out[2917] | layer0_out[2916];
    assign layer1_out[3624] = ~layer0_out[2967] | layer0_out[2966];
    assign layer1_out[3625] = layer0_out[5763] & layer0_out[5764];
    assign layer1_out[3626] = layer0_out[3795];
    assign layer1_out[3627] = layer0_out[2811];
    assign layer1_out[3628] = layer0_out[6087] & layer0_out[6088];
    assign layer1_out[3629] = ~(layer0_out[249] | layer0_out[250]);
    assign layer1_out[3630] = ~(layer0_out[2499] & layer0_out[2500]);
    assign layer1_out[3631] = layer0_out[1027] ^ layer0_out[1028];
    assign layer1_out[3632] = ~layer0_out[2364] | layer0_out[2365];
    assign layer1_out[3633] = layer0_out[7860] | layer0_out[7861];
    assign layer1_out[3634] = layer0_out[6184] ^ layer0_out[6185];
    assign layer1_out[3635] = layer0_out[7050] & ~layer0_out[7051];
    assign layer1_out[3636] = ~layer0_out[1983];
    assign layer1_out[3637] = layer0_out[6103] | layer0_out[6104];
    assign layer1_out[3638] = ~(layer0_out[3776] | layer0_out[3777]);
    assign layer1_out[3639] = layer0_out[3612] & layer0_out[3613];
    assign layer1_out[3640] = layer0_out[7594] & layer0_out[7595];
    assign layer1_out[3641] = layer0_out[2993];
    assign layer1_out[3642] = layer0_out[5431] ^ layer0_out[5432];
    assign layer1_out[3643] = ~(layer0_out[2587] & layer0_out[2588]);
    assign layer1_out[3644] = ~layer0_out[6929] | layer0_out[6928];
    assign layer1_out[3645] = ~layer0_out[565];
    assign layer1_out[3646] = layer0_out[6239] & ~layer0_out[6238];
    assign layer1_out[3647] = ~layer0_out[3473];
    assign layer1_out[3648] = layer0_out[446] | layer0_out[447];
    assign layer1_out[3649] = ~layer0_out[5384];
    assign layer1_out[3650] = layer0_out[3296];
    assign layer1_out[3651] = ~layer0_out[5305];
    assign layer1_out[3652] = layer0_out[5165];
    assign layer1_out[3653] = layer0_out[204] & ~layer0_out[203];
    assign layer1_out[3654] = layer0_out[967] | layer0_out[968];
    assign layer1_out[3655] = ~layer0_out[6135] | layer0_out[6134];
    assign layer1_out[3656] = layer0_out[7513] & layer0_out[7514];
    assign layer1_out[3657] = layer0_out[1851];
    assign layer1_out[3658] = layer0_out[6268] | layer0_out[6269];
    assign layer1_out[3659] = layer0_out[4238];
    assign layer1_out[3660] = layer0_out[4739] & ~layer0_out[4740];
    assign layer1_out[3661] = layer0_out[3080] | layer0_out[3081];
    assign layer1_out[3662] = layer0_out[3963] & ~layer0_out[3962];
    assign layer1_out[3663] = layer0_out[7703] & layer0_out[7704];
    assign layer1_out[3664] = layer0_out[4054] & ~layer0_out[4055];
    assign layer1_out[3665] = ~(layer0_out[1384] ^ layer0_out[1385]);
    assign layer1_out[3666] = 1'b0;
    assign layer1_out[3667] = layer0_out[1280] & ~layer0_out[1279];
    assign layer1_out[3668] = 1'b0;
    assign layer1_out[3669] = ~(layer0_out[1840] | layer0_out[1841]);
    assign layer1_out[3670] = layer0_out[4369];
    assign layer1_out[3671] = layer0_out[5085] | layer0_out[5086];
    assign layer1_out[3672] = ~(layer0_out[2210] & layer0_out[2211]);
    assign layer1_out[3673] = ~layer0_out[7985] | layer0_out[7986];
    assign layer1_out[3674] = layer0_out[7747] & ~layer0_out[7746];
    assign layer1_out[3675] = ~(layer0_out[754] ^ layer0_out[755]);
    assign layer1_out[3676] = layer0_out[893] & layer0_out[894];
    assign layer1_out[3677] = layer0_out[5378];
    assign layer1_out[3678] = ~layer0_out[4947];
    assign layer1_out[3679] = layer0_out[3453] & ~layer0_out[3452];
    assign layer1_out[3680] = ~layer0_out[3733];
    assign layer1_out[3681] = layer0_out[1119] & layer0_out[1120];
    assign layer1_out[3682] = layer0_out[5222];
    assign layer1_out[3683] = ~(layer0_out[5792] & layer0_out[5793]);
    assign layer1_out[3684] = ~layer0_out[979];
    assign layer1_out[3685] = ~layer0_out[1413];
    assign layer1_out[3686] = ~layer0_out[2111] | layer0_out[2112];
    assign layer1_out[3687] = ~layer0_out[364] | layer0_out[365];
    assign layer1_out[3688] = layer0_out[2279] & layer0_out[2280];
    assign layer1_out[3689] = layer0_out[7896] ^ layer0_out[7897];
    assign layer1_out[3690] = layer0_out[7754];
    assign layer1_out[3691] = layer0_out[6497] ^ layer0_out[6498];
    assign layer1_out[3692] = ~layer0_out[5470] | layer0_out[5471];
    assign layer1_out[3693] = layer0_out[3845] ^ layer0_out[3846];
    assign layer1_out[3694] = layer0_out[4968];
    assign layer1_out[3695] = layer0_out[544] & layer0_out[545];
    assign layer1_out[3696] = ~(layer0_out[5652] & layer0_out[5653]);
    assign layer1_out[3697] = ~layer0_out[2781];
    assign layer1_out[3698] = layer0_out[986] & layer0_out[987];
    assign layer1_out[3699] = ~(layer0_out[3387] | layer0_out[3388]);
    assign layer1_out[3700] = ~layer0_out[2472];
    assign layer1_out[3701] = ~(layer0_out[1651] | layer0_out[1652]);
    assign layer1_out[3702] = layer0_out[3278] | layer0_out[3279];
    assign layer1_out[3703] = ~layer0_out[4102] | layer0_out[4101];
    assign layer1_out[3704] = ~layer0_out[7703] | layer0_out[7702];
    assign layer1_out[3705] = ~(layer0_out[6496] | layer0_out[6497]);
    assign layer1_out[3706] = 1'b1;
    assign layer1_out[3707] = layer0_out[4032] | layer0_out[4033];
    assign layer1_out[3708] = ~layer0_out[3005];
    assign layer1_out[3709] = ~layer0_out[1156];
    assign layer1_out[3710] = ~(layer0_out[5887] ^ layer0_out[5888]);
    assign layer1_out[3711] = 1'b0;
    assign layer1_out[3712] = ~layer0_out[7714];
    assign layer1_out[3713] = layer0_out[3244];
    assign layer1_out[3714] = layer0_out[6205] ^ layer0_out[6206];
    assign layer1_out[3715] = ~layer0_out[603] | layer0_out[602];
    assign layer1_out[3716] = 1'b0;
    assign layer1_out[3717] = ~layer0_out[3505];
    assign layer1_out[3718] = 1'b0;
    assign layer1_out[3719] = layer0_out[1333];
    assign layer1_out[3720] = layer0_out[4647] & ~layer0_out[4646];
    assign layer1_out[3721] = layer0_out[6912] & ~layer0_out[6911];
    assign layer1_out[3722] = layer0_out[1271];
    assign layer1_out[3723] = ~layer0_out[3983] | layer0_out[3982];
    assign layer1_out[3724] = ~layer0_out[7434];
    assign layer1_out[3725] = 1'b0;
    assign layer1_out[3726] = layer0_out[2100] & ~layer0_out[2099];
    assign layer1_out[3727] = layer0_out[3370] & ~layer0_out[3371];
    assign layer1_out[3728] = 1'b0;
    assign layer1_out[3729] = ~layer0_out[6943];
    assign layer1_out[3730] = layer0_out[919] & ~layer0_out[920];
    assign layer1_out[3731] = ~layer0_out[678];
    assign layer1_out[3732] = layer0_out[5814] & layer0_out[5815];
    assign layer1_out[3733] = layer0_out[5061] & ~layer0_out[5062];
    assign layer1_out[3734] = layer0_out[1159] & ~layer0_out[1158];
    assign layer1_out[3735] = ~layer0_out[6751] | layer0_out[6752];
    assign layer1_out[3736] = ~(layer0_out[3040] & layer0_out[3041]);
    assign layer1_out[3737] = layer0_out[7587];
    assign layer1_out[3738] = ~layer0_out[387] | layer0_out[388];
    assign layer1_out[3739] = layer0_out[4549] | layer0_out[4550];
    assign layer1_out[3740] = 1'b0;
    assign layer1_out[3741] = layer0_out[3786];
    assign layer1_out[3742] = 1'b1;
    assign layer1_out[3743] = 1'b1;
    assign layer1_out[3744] = 1'b0;
    assign layer1_out[3745] = layer0_out[4330] & ~layer0_out[4329];
    assign layer1_out[3746] = layer0_out[5797];
    assign layer1_out[3747] = layer0_out[2146] & layer0_out[2147];
    assign layer1_out[3748] = layer0_out[2006];
    assign layer1_out[3749] = ~layer0_out[2823] | layer0_out[2822];
    assign layer1_out[3750] = ~layer0_out[7161];
    assign layer1_out[3751] = ~layer0_out[142] | layer0_out[143];
    assign layer1_out[3752] = 1'b0;
    assign layer1_out[3753] = layer0_out[5060] & ~layer0_out[5061];
    assign layer1_out[3754] = layer0_out[1471] & ~layer0_out[1470];
    assign layer1_out[3755] = layer0_out[4933] ^ layer0_out[4934];
    assign layer1_out[3756] = 1'b0;
    assign layer1_out[3757] = ~(layer0_out[3053] | layer0_out[3054]);
    assign layer1_out[3758] = layer0_out[4880] | layer0_out[4881];
    assign layer1_out[3759] = ~layer0_out[5463] | layer0_out[5464];
    assign layer1_out[3760] = ~layer0_out[4021];
    assign layer1_out[3761] = ~layer0_out[5990];
    assign layer1_out[3762] = ~(layer0_out[6323] ^ layer0_out[6324]);
    assign layer1_out[3763] = ~layer0_out[2056];
    assign layer1_out[3764] = layer0_out[289] & layer0_out[290];
    assign layer1_out[3765] = ~layer0_out[3496];
    assign layer1_out[3766] = ~layer0_out[7864] | layer0_out[7863];
    assign layer1_out[3767] = layer0_out[5731] | layer0_out[5732];
    assign layer1_out[3768] = layer0_out[5170] & ~layer0_out[5169];
    assign layer1_out[3769] = layer0_out[3694] | layer0_out[3695];
    assign layer1_out[3770] = layer0_out[347] & ~layer0_out[348];
    assign layer1_out[3771] = layer0_out[2521] ^ layer0_out[2522];
    assign layer1_out[3772] = layer0_out[3916];
    assign layer1_out[3773] = ~layer0_out[874];
    assign layer1_out[3774] = layer0_out[1829] & ~layer0_out[1828];
    assign layer1_out[3775] = layer0_out[6886] ^ layer0_out[6887];
    assign layer1_out[3776] = ~layer0_out[5246];
    assign layer1_out[3777] = 1'b1;
    assign layer1_out[3778] = ~layer0_out[3657];
    assign layer1_out[3779] = layer0_out[7264];
    assign layer1_out[3780] = ~(layer0_out[7203] | layer0_out[7204]);
    assign layer1_out[3781] = ~layer0_out[4371];
    assign layer1_out[3782] = layer0_out[5131] | layer0_out[5132];
    assign layer1_out[3783] = ~(layer0_out[600] ^ layer0_out[601]);
    assign layer1_out[3784] = layer0_out[2045] ^ layer0_out[2046];
    assign layer1_out[3785] = ~(layer0_out[4816] | layer0_out[4817]);
    assign layer1_out[3786] = ~layer0_out[4471] | layer0_out[4470];
    assign layer1_out[3787] = ~(layer0_out[5806] & layer0_out[5807]);
    assign layer1_out[3788] = layer0_out[537];
    assign layer1_out[3789] = ~layer0_out[5207] | layer0_out[5206];
    assign layer1_out[3790] = layer0_out[6170] & ~layer0_out[6169];
    assign layer1_out[3791] = layer0_out[4161];
    assign layer1_out[3792] = ~(layer0_out[6851] ^ layer0_out[6852]);
    assign layer1_out[3793] = ~layer0_out[1572] | layer0_out[1571];
    assign layer1_out[3794] = 1'b0;
    assign layer1_out[3795] = ~layer0_out[7393] | layer0_out[7392];
    assign layer1_out[3796] = ~layer0_out[7813] | layer0_out[7812];
    assign layer1_out[3797] = layer0_out[2159] | layer0_out[2160];
    assign layer1_out[3798] = ~layer0_out[1425];
    assign layer1_out[3799] = ~(layer0_out[750] & layer0_out[751]);
    assign layer1_out[3800] = ~(layer0_out[4263] & layer0_out[4264]);
    assign layer1_out[3801] = ~layer0_out[3696];
    assign layer1_out[3802] = ~layer0_out[2418];
    assign layer1_out[3803] = ~(layer0_out[7500] | layer0_out[7501]);
    assign layer1_out[3804] = layer0_out[6056];
    assign layer1_out[3805] = 1'b1;
    assign layer1_out[3806] = ~(layer0_out[2023] | layer0_out[2024]);
    assign layer1_out[3807] = ~layer0_out[6901];
    assign layer1_out[3808] = layer0_out[358];
    assign layer1_out[3809] = layer0_out[3894];
    assign layer1_out[3810] = ~(layer0_out[6838] | layer0_out[6839]);
    assign layer1_out[3811] = ~(layer0_out[7887] | layer0_out[7888]);
    assign layer1_out[3812] = 1'b1;
    assign layer1_out[3813] = layer0_out[5492] & ~layer0_out[5493];
    assign layer1_out[3814] = layer0_out[7386] & ~layer0_out[7385];
    assign layer1_out[3815] = layer0_out[1006];
    assign layer1_out[3816] = ~layer0_out[5273];
    assign layer1_out[3817] = ~layer0_out[4605] | layer0_out[4604];
    assign layer1_out[3818] = ~layer0_out[5683] | layer0_out[5684];
    assign layer1_out[3819] = layer0_out[5973];
    assign layer1_out[3820] = ~layer0_out[4893] | layer0_out[4894];
    assign layer1_out[3821] = ~layer0_out[1930];
    assign layer1_out[3822] = ~layer0_out[1534] | layer0_out[1535];
    assign layer1_out[3823] = layer0_out[4831] & ~layer0_out[4830];
    assign layer1_out[3824] = layer0_out[2266] | layer0_out[2267];
    assign layer1_out[3825] = 1'b1;
    assign layer1_out[3826] = ~layer0_out[1653];
    assign layer1_out[3827] = ~(layer0_out[4569] | layer0_out[4570]);
    assign layer1_out[3828] = layer0_out[4500] & layer0_out[4501];
    assign layer1_out[3829] = ~layer0_out[1827];
    assign layer1_out[3830] = ~layer0_out[2312];
    assign layer1_out[3831] = ~layer0_out[7718];
    assign layer1_out[3832] = ~layer0_out[6344] | layer0_out[6345];
    assign layer1_out[3833] = ~layer0_out[1050] | layer0_out[1051];
    assign layer1_out[3834] = layer0_out[501] & layer0_out[502];
    assign layer1_out[3835] = ~(layer0_out[2980] ^ layer0_out[2981]);
    assign layer1_out[3836] = layer0_out[3408] & ~layer0_out[3409];
    assign layer1_out[3837] = ~layer0_out[4268];
    assign layer1_out[3838] = layer0_out[612] ^ layer0_out[613];
    assign layer1_out[3839] = layer0_out[4142] & ~layer0_out[4141];
    assign layer1_out[3840] = ~(layer0_out[7608] | layer0_out[7609]);
    assign layer1_out[3841] = layer0_out[3440] | layer0_out[3441];
    assign layer1_out[3842] = ~(layer0_out[5220] | layer0_out[5221]);
    assign layer1_out[3843] = ~layer0_out[2238];
    assign layer1_out[3844] = ~layer0_out[6983] | layer0_out[6982];
    assign layer1_out[3845] = layer0_out[3293] & ~layer0_out[3292];
    assign layer1_out[3846] = ~layer0_out[865];
    assign layer1_out[3847] = ~layer0_out[6825];
    assign layer1_out[3848] = ~layer0_out[440] | layer0_out[439];
    assign layer1_out[3849] = layer0_out[7991] & ~layer0_out[7990];
    assign layer1_out[3850] = 1'b1;
    assign layer1_out[3851] = layer0_out[1486];
    assign layer1_out[3852] = layer0_out[509];
    assign layer1_out[3853] = 1'b0;
    assign layer1_out[3854] = layer0_out[5499];
    assign layer1_out[3855] = ~(layer0_out[672] ^ layer0_out[673]);
    assign layer1_out[3856] = ~layer0_out[6116] | layer0_out[6115];
    assign layer1_out[3857] = layer0_out[6365] | layer0_out[6366];
    assign layer1_out[3858] = 1'b0;
    assign layer1_out[3859] = layer0_out[2003] & layer0_out[2004];
    assign layer1_out[3860] = ~layer0_out[7743] | layer0_out[7744];
    assign layer1_out[3861] = ~layer0_out[1974] | layer0_out[1973];
    assign layer1_out[3862] = 1'b1;
    assign layer1_out[3863] = ~(layer0_out[4987] & layer0_out[4988]);
    assign layer1_out[3864] = layer0_out[7577] & ~layer0_out[7578];
    assign layer1_out[3865] = ~(layer0_out[7845] & layer0_out[7846]);
    assign layer1_out[3866] = ~layer0_out[5677];
    assign layer1_out[3867] = layer0_out[3862] & ~layer0_out[3861];
    assign layer1_out[3868] = ~(layer0_out[7859] | layer0_out[7860]);
    assign layer1_out[3869] = ~layer0_out[7262] | layer0_out[7261];
    assign layer1_out[3870] = ~layer0_out[5910] | layer0_out[5911];
    assign layer1_out[3871] = ~layer0_out[6708] | layer0_out[6707];
    assign layer1_out[3872] = layer0_out[5203] & ~layer0_out[5204];
    assign layer1_out[3873] = ~(layer0_out[3740] & layer0_out[3741]);
    assign layer1_out[3874] = layer0_out[219] & layer0_out[220];
    assign layer1_out[3875] = layer0_out[7494];
    assign layer1_out[3876] = layer0_out[157] | layer0_out[158];
    assign layer1_out[3877] = 1'b1;
    assign layer1_out[3878] = ~(layer0_out[6422] ^ layer0_out[6423]);
    assign layer1_out[3879] = ~layer0_out[1242] | layer0_out[1241];
    assign layer1_out[3880] = ~(layer0_out[5432] | layer0_out[5433]);
    assign layer1_out[3881] = ~layer0_out[7323];
    assign layer1_out[3882] = ~layer0_out[7687] | layer0_out[7686];
    assign layer1_out[3883] = ~(layer0_out[4921] | layer0_out[4922]);
    assign layer1_out[3884] = layer0_out[4134];
    assign layer1_out[3885] = layer0_out[6761] & ~layer0_out[6760];
    assign layer1_out[3886] = layer0_out[4571] & layer0_out[4572];
    assign layer1_out[3887] = layer0_out[2606] & ~layer0_out[2605];
    assign layer1_out[3888] = layer0_out[1614] & ~layer0_out[1613];
    assign layer1_out[3889] = layer0_out[6009] ^ layer0_out[6010];
    assign layer1_out[3890] = ~(layer0_out[7458] ^ layer0_out[7459]);
    assign layer1_out[3891] = layer0_out[4689] | layer0_out[4690];
    assign layer1_out[3892] = layer0_out[4205] | layer0_out[4206];
    assign layer1_out[3893] = layer0_out[6836] ^ layer0_out[6837];
    assign layer1_out[3894] = layer0_out[5458] | layer0_out[5459];
    assign layer1_out[3895] = ~layer0_out[594];
    assign layer1_out[3896] = ~layer0_out[6562] | layer0_out[6561];
    assign layer1_out[3897] = layer0_out[2054] & ~layer0_out[2055];
    assign layer1_out[3898] = ~layer0_out[6551];
    assign layer1_out[3899] = ~layer0_out[4473];
    assign layer1_out[3900] = layer0_out[20] & ~layer0_out[19];
    assign layer1_out[3901] = layer0_out[341];
    assign layer1_out[3902] = layer0_out[1773] & ~layer0_out[1772];
    assign layer1_out[3903] = layer0_out[1420] & ~layer0_out[1419];
    assign layer1_out[3904] = ~layer0_out[7417] | layer0_out[7418];
    assign layer1_out[3905] = layer0_out[2507] & ~layer0_out[2506];
    assign layer1_out[3906] = ~(layer0_out[4656] ^ layer0_out[4657]);
    assign layer1_out[3907] = ~layer0_out[4842] | layer0_out[4841];
    assign layer1_out[3908] = ~layer0_out[3931] | layer0_out[3930];
    assign layer1_out[3909] = layer0_out[1369] & ~layer0_out[1368];
    assign layer1_out[3910] = layer0_out[7871];
    assign layer1_out[3911] = ~layer0_out[2290];
    assign layer1_out[3912] = layer0_out[5162];
    assign layer1_out[3913] = layer0_out[4281];
    assign layer1_out[3914] = ~(layer0_out[5174] & layer0_out[5175]);
    assign layer1_out[3915] = ~layer0_out[6977] | layer0_out[6976];
    assign layer1_out[3916] = ~layer0_out[2919];
    assign layer1_out[3917] = ~(layer0_out[6015] ^ layer0_out[6016]);
    assign layer1_out[3918] = layer0_out[4055] & ~layer0_out[4056];
    assign layer1_out[3919] = ~(layer0_out[7697] ^ layer0_out[7698]);
    assign layer1_out[3920] = ~(layer0_out[1126] | layer0_out[1127]);
    assign layer1_out[3921] = layer0_out[3727];
    assign layer1_out[3922] = layer0_out[6953] & ~layer0_out[6952];
    assign layer1_out[3923] = layer0_out[5198];
    assign layer1_out[3924] = layer0_out[5841] & layer0_out[5842];
    assign layer1_out[3925] = ~(layer0_out[512] & layer0_out[513]);
    assign layer1_out[3926] = layer0_out[3619] & ~layer0_out[3620];
    assign layer1_out[3927] = layer0_out[7077];
    assign layer1_out[3928] = ~(layer0_out[6812] & layer0_out[6813]);
    assign layer1_out[3929] = ~layer0_out[5934] | layer0_out[5935];
    assign layer1_out[3930] = layer0_out[7962] ^ layer0_out[7963];
    assign layer1_out[3931] = layer0_out[6319] & layer0_out[6320];
    assign layer1_out[3932] = ~layer0_out[1780];
    assign layer1_out[3933] = layer0_out[6501] ^ layer0_out[6502];
    assign layer1_out[3934] = layer0_out[3565];
    assign layer1_out[3935] = layer0_out[7477];
    assign layer1_out[3936] = ~layer0_out[604];
    assign layer1_out[3937] = layer0_out[6202] & ~layer0_out[6201];
    assign layer1_out[3938] = layer0_out[3069] | layer0_out[3070];
    assign layer1_out[3939] = layer0_out[7210] & layer0_out[7211];
    assign layer1_out[3940] = layer0_out[5028];
    assign layer1_out[3941] = layer0_out[1665];
    assign layer1_out[3942] = 1'b0;
    assign layer1_out[3943] = ~layer0_out[4142] | layer0_out[4143];
    assign layer1_out[3944] = ~(layer0_out[4223] | layer0_out[4224]);
    assign layer1_out[3945] = ~(layer0_out[4535] & layer0_out[4536]);
    assign layer1_out[3946] = ~layer0_out[5452];
    assign layer1_out[3947] = layer0_out[3346] & ~layer0_out[3345];
    assign layer1_out[3948] = layer0_out[6533];
    assign layer1_out[3949] = layer0_out[1991] & layer0_out[1992];
    assign layer1_out[3950] = layer0_out[4501];
    assign layer1_out[3951] = layer0_out[5095];
    assign layer1_out[3952] = layer0_out[1633] & ~layer0_out[1634];
    assign layer1_out[3953] = ~layer0_out[3985] | layer0_out[3986];
    assign layer1_out[3954] = ~(layer0_out[7921] | layer0_out[7922]);
    assign layer1_out[3955] = ~(layer0_out[7337] & layer0_out[7338]);
    assign layer1_out[3956] = ~layer0_out[860] | layer0_out[861];
    assign layer1_out[3957] = ~(layer0_out[6741] & layer0_out[6742]);
    assign layer1_out[3958] = 1'b1;
    assign layer1_out[3959] = layer0_out[5544];
    assign layer1_out[3960] = ~layer0_out[6669];
    assign layer1_out[3961] = layer0_out[3294] & layer0_out[3295];
    assign layer1_out[3962] = ~(layer0_out[5579] ^ layer0_out[5580]);
    assign layer1_out[3963] = layer0_out[4694] | layer0_out[4695];
    assign layer1_out[3964] = ~(layer0_out[7638] | layer0_out[7639]);
    assign layer1_out[3965] = layer0_out[5889];
    assign layer1_out[3966] = layer0_out[6041];
    assign layer1_out[3967] = 1'b1;
    assign layer1_out[3968] = ~layer0_out[589];
    assign layer1_out[3969] = ~layer0_out[4147];
    assign layer1_out[3970] = ~layer0_out[3919];
    assign layer1_out[3971] = ~layer0_out[6328];
    assign layer1_out[3972] = ~layer0_out[7815] | layer0_out[7816];
    assign layer1_out[3973] = ~layer0_out[7300] | layer0_out[7299];
    assign layer1_out[3974] = layer0_out[3827];
    assign layer1_out[3975] = ~layer0_out[1591];
    assign layer1_out[3976] = ~layer0_out[6861] | layer0_out[6860];
    assign layer1_out[3977] = ~layer0_out[2341] | layer0_out[2340];
    assign layer1_out[3978] = layer0_out[5371];
    assign layer1_out[3979] = layer0_out[6518] & ~layer0_out[6517];
    assign layer1_out[3980] = layer0_out[7528];
    assign layer1_out[3981] = ~layer0_out[5853];
    assign layer1_out[3982] = 1'b0;
    assign layer1_out[3983] = ~layer0_out[4594] | layer0_out[4593];
    assign layer1_out[3984] = layer0_out[348];
    assign layer1_out[3985] = layer0_out[3995] & ~layer0_out[3996];
    assign layer1_out[3986] = layer0_out[838] & ~layer0_out[837];
    assign layer1_out[3987] = 1'b1;
    assign layer1_out[3988] = ~(layer0_out[3070] ^ layer0_out[3071]);
    assign layer1_out[3989] = ~layer0_out[3718] | layer0_out[3717];
    assign layer1_out[3990] = layer0_out[6248] | layer0_out[6249];
    assign layer1_out[3991] = ~layer0_out[443] | layer0_out[442];
    assign layer1_out[3992] = layer0_out[7969] & layer0_out[7970];
    assign layer1_out[3993] = layer0_out[3426];
    assign layer1_out[3994] = ~layer0_out[7722] | layer0_out[7721];
    assign layer1_out[3995] = layer0_out[202] & ~layer0_out[201];
    assign layer1_out[3996] = layer0_out[7144];
    assign layer1_out[3997] = ~layer0_out[728];
    assign layer1_out[3998] = ~layer0_out[1226];
    assign layer1_out[3999] = layer0_out[3176] & layer0_out[3177];
    assign layer1_out[4000] = layer0_out[3146];
    assign layer1_out[4001] = layer0_out[6357];
    assign layer1_out[4002] = ~(layer0_out[1658] & layer0_out[1659]);
    assign layer1_out[4003] = layer0_out[7090] & ~layer0_out[7089];
    assign layer1_out[4004] = layer0_out[5501] & ~layer0_out[5502];
    assign layer1_out[4005] = ~(layer0_out[3167] & layer0_out[3168]);
    assign layer1_out[4006] = ~layer0_out[3289];
    assign layer1_out[4007] = ~layer0_out[3207] | layer0_out[3206];
    assign layer1_out[4008] = layer0_out[2735] & ~layer0_out[2736];
    assign layer1_out[4009] = ~layer0_out[5605];
    assign layer1_out[4010] = layer0_out[2383] | layer0_out[2384];
    assign layer1_out[4011] = layer0_out[1114] & layer0_out[1115];
    assign layer1_out[4012] = ~layer0_out[5541];
    assign layer1_out[4013] = layer0_out[3499] & ~layer0_out[3500];
    assign layer1_out[4014] = layer0_out[2371];
    assign layer1_out[4015] = ~layer0_out[268];
    assign layer1_out[4016] = 1'b1;
    assign layer1_out[4017] = ~layer0_out[1233];
    assign layer1_out[4018] = layer0_out[479];
    assign layer1_out[4019] = ~(layer0_out[3708] | layer0_out[3709]);
    assign layer1_out[4020] = ~layer0_out[3517] | layer0_out[3518];
    assign layer1_out[4021] = ~layer0_out[3879] | layer0_out[3880];
    assign layer1_out[4022] = layer0_out[2114] ^ layer0_out[2115];
    assign layer1_out[4023] = layer0_out[5445];
    assign layer1_out[4024] = layer0_out[3269];
    assign layer1_out[4025] = layer0_out[205] & ~layer0_out[204];
    assign layer1_out[4026] = ~layer0_out[6111];
    assign layer1_out[4027] = ~(layer0_out[6680] ^ layer0_out[6681]);
    assign layer1_out[4028] = layer0_out[5894] & layer0_out[5895];
    assign layer1_out[4029] = ~layer0_out[2814];
    assign layer1_out[4030] = ~(layer0_out[3885] & layer0_out[3886]);
    assign layer1_out[4031] = layer0_out[1162] & ~layer0_out[1161];
    assign layer1_out[4032] = ~layer0_out[2221];
    assign layer1_out[4033] = ~layer0_out[2985] | layer0_out[2986];
    assign layer1_out[4034] = layer0_out[4457];
    assign layer1_out[4035] = ~(layer0_out[6387] & layer0_out[6388]);
    assign layer1_out[4036] = layer0_out[7502] & ~layer0_out[7501];
    assign layer1_out[4037] = ~layer0_out[1087];
    assign layer1_out[4038] = ~layer0_out[1748];
    assign layer1_out[4039] = layer0_out[7591] & ~layer0_out[7592];
    assign layer1_out[4040] = ~(layer0_out[2043] | layer0_out[2044]);
    assign layer1_out[4041] = layer0_out[951];
    assign layer1_out[4042] = layer0_out[5966];
    assign layer1_out[4043] = layer0_out[2220] & ~layer0_out[2219];
    assign layer1_out[4044] = ~(layer0_out[3741] ^ layer0_out[3742]);
    assign layer1_out[4045] = ~(layer0_out[308] | layer0_out[309]);
    assign layer1_out[4046] = layer0_out[1570];
    assign layer1_out[4047] = layer0_out[4085] & ~layer0_out[4086];
    assign layer1_out[4048] = ~layer0_out[2933] | layer0_out[2932];
    assign layer1_out[4049] = layer0_out[426] | layer0_out[427];
    assign layer1_out[4050] = layer0_out[3640] & layer0_out[3641];
    assign layer1_out[4051] = ~layer0_out[7073] | layer0_out[7074];
    assign layer1_out[4052] = ~(layer0_out[5101] | layer0_out[5102]);
    assign layer1_out[4053] = ~layer0_out[6912] | layer0_out[6913];
    assign layer1_out[4054] = layer0_out[694];
    assign layer1_out[4055] = layer0_out[2855] & ~layer0_out[2854];
    assign layer1_out[4056] = ~layer0_out[4334];
    assign layer1_out[4057] = ~(layer0_out[391] | layer0_out[392]);
    assign layer1_out[4058] = layer0_out[7723] & ~layer0_out[7722];
    assign layer1_out[4059] = ~(layer0_out[5163] | layer0_out[5164]);
    assign layer1_out[4060] = ~(layer0_out[2633] | layer0_out[2634]);
    assign layer1_out[4061] = layer0_out[155] ^ layer0_out[156];
    assign layer1_out[4062] = layer0_out[3251] | layer0_out[3252];
    assign layer1_out[4063] = ~layer0_out[2254] | layer0_out[2253];
    assign layer1_out[4064] = ~(layer0_out[5041] & layer0_out[5042]);
    assign layer1_out[4065] = layer0_out[2601];
    assign layer1_out[4066] = ~layer0_out[5285] | layer0_out[5284];
    assign layer1_out[4067] = ~layer0_out[7298] | layer0_out[7297];
    assign layer1_out[4068] = ~(layer0_out[7284] & layer0_out[7285]);
    assign layer1_out[4069] = layer0_out[7345] & ~layer0_out[7346];
    assign layer1_out[4070] = layer0_out[5063] & ~layer0_out[5062];
    assign layer1_out[4071] = ~layer0_out[4986] | layer0_out[4985];
    assign layer1_out[4072] = layer0_out[1128];
    assign layer1_out[4073] = ~layer0_out[3477];
    assign layer1_out[4074] = layer0_out[5832];
    assign layer1_out[4075] = ~(layer0_out[5498] ^ layer0_out[5499]);
    assign layer1_out[4076] = ~layer0_out[503];
    assign layer1_out[4077] = layer0_out[4293] & layer0_out[4294];
    assign layer1_out[4078] = layer0_out[318] | layer0_out[319];
    assign layer1_out[4079] = ~layer0_out[5805];
    assign layer1_out[4080] = ~(layer0_out[7275] ^ layer0_out[7276]);
    assign layer1_out[4081] = ~(layer0_out[7383] ^ layer0_out[7384]);
    assign layer1_out[4082] = ~layer0_out[5592];
    assign layer1_out[4083] = ~layer0_out[5191] | layer0_out[5190];
    assign layer1_out[4084] = ~(layer0_out[4094] ^ layer0_out[4095]);
    assign layer1_out[4085] = ~layer0_out[7949];
    assign layer1_out[4086] = layer0_out[5782] & ~layer0_out[5781];
    assign layer1_out[4087] = ~layer0_out[6729] | layer0_out[6728];
    assign layer1_out[4088] = layer0_out[4357] & ~layer0_out[4356];
    assign layer1_out[4089] = ~layer0_out[5553];
    assign layer1_out[4090] = layer0_out[4885] & ~layer0_out[4884];
    assign layer1_out[4091] = layer0_out[1236] | layer0_out[1237];
    assign layer1_out[4092] = ~layer0_out[2031];
    assign layer1_out[4093] = layer0_out[2208];
    assign layer1_out[4094] = ~(layer0_out[2422] ^ layer0_out[2423]);
    assign layer1_out[4095] = layer0_out[3831];
    assign layer1_out[4096] = layer0_out[1546];
    assign layer1_out[4097] = layer0_out[1528];
    assign layer1_out[4098] = ~layer0_out[7696];
    assign layer1_out[4099] = ~layer0_out[6224] | layer0_out[6225];
    assign layer1_out[4100] = ~layer0_out[3665] | layer0_out[3666];
    assign layer1_out[4101] = ~(layer0_out[7613] ^ layer0_out[7614]);
    assign layer1_out[4102] = layer0_out[323];
    assign layer1_out[4103] = 1'b1;
    assign layer1_out[4104] = layer0_out[2411];
    assign layer1_out[4105] = layer0_out[2665] & ~layer0_out[2666];
    assign layer1_out[4106] = layer0_out[3706];
    assign layer1_out[4107] = ~(layer0_out[4324] & layer0_out[4325]);
    assign layer1_out[4108] = layer0_out[257] & ~layer0_out[256];
    assign layer1_out[4109] = ~layer0_out[6653];
    assign layer1_out[4110] = 1'b1;
    assign layer1_out[4111] = ~layer0_out[7827] | layer0_out[7828];
    assign layer1_out[4112] = layer0_out[5352];
    assign layer1_out[4113] = layer0_out[5641];
    assign layer1_out[4114] = layer0_out[281] | layer0_out[282];
    assign layer1_out[4115] = layer0_out[675] & ~layer0_out[674];
    assign layer1_out[4116] = layer0_out[3789];
    assign layer1_out[4117] = layer0_out[1242] & layer0_out[1243];
    assign layer1_out[4118] = ~layer0_out[5559];
    assign layer1_out[4119] = layer0_out[7826];
    assign layer1_out[4120] = ~(layer0_out[630] | layer0_out[631]);
    assign layer1_out[4121] = ~layer0_out[7138];
    assign layer1_out[4122] = ~layer0_out[7162] | layer0_out[7163];
    assign layer1_out[4123] = layer0_out[4564];
    assign layer1_out[4124] = layer0_out[5184];
    assign layer1_out[4125] = ~layer0_out[3507];
    assign layer1_out[4126] = ~(layer0_out[3766] ^ layer0_out[3767]);
    assign layer1_out[4127] = layer0_out[3018];
    assign layer1_out[4128] = ~layer0_out[5349];
    assign layer1_out[4129] = layer0_out[6660] & layer0_out[6661];
    assign layer1_out[4130] = layer0_out[129];
    assign layer1_out[4131] = ~layer0_out[3883];
    assign layer1_out[4132] = ~layer0_out[5756] | layer0_out[5757];
    assign layer1_out[4133] = layer0_out[2162] & ~layer0_out[2163];
    assign layer1_out[4134] = layer0_out[5437];
    assign layer1_out[4135] = layer0_out[401] & layer0_out[402];
    assign layer1_out[4136] = layer0_out[7653] & layer0_out[7654];
    assign layer1_out[4137] = 1'b0;
    assign layer1_out[4138] = ~(layer0_out[1051] | layer0_out[1052]);
    assign layer1_out[4139] = ~layer0_out[2024];
    assign layer1_out[4140] = ~(layer0_out[286] | layer0_out[287]);
    assign layer1_out[4141] = ~layer0_out[329];
    assign layer1_out[4142] = layer0_out[2562] & layer0_out[2563];
    assign layer1_out[4143] = ~layer0_out[5823];
    assign layer1_out[4144] = layer0_out[2250];
    assign layer1_out[4145] = ~(layer0_out[5425] | layer0_out[5426]);
    assign layer1_out[4146] = ~layer0_out[4333];
    assign layer1_out[4147] = layer0_out[4285];
    assign layer1_out[4148] = ~layer0_out[1131];
    assign layer1_out[4149] = layer0_out[3998] & layer0_out[3999];
    assign layer1_out[4150] = layer0_out[2570] & ~layer0_out[2571];
    assign layer1_out[4151] = layer0_out[557] & layer0_out[558];
    assign layer1_out[4152] = ~(layer0_out[7871] & layer0_out[7872]);
    assign layer1_out[4153] = layer0_out[5013];
    assign layer1_out[4154] = ~layer0_out[3102];
    assign layer1_out[4155] = layer0_out[4274] & layer0_out[4275];
    assign layer1_out[4156] = ~layer0_out[405];
    assign layer1_out[4157] = layer0_out[819] | layer0_out[820];
    assign layer1_out[4158] = layer0_out[3697] & ~layer0_out[3698];
    assign layer1_out[4159] = layer0_out[37];
    assign layer1_out[4160] = layer0_out[7621] ^ layer0_out[7622];
    assign layer1_out[4161] = layer0_out[1478] & ~layer0_out[1477];
    assign layer1_out[4162] = layer0_out[3131];
    assign layer1_out[4163] = ~(layer0_out[3554] & layer0_out[3555]);
    assign layer1_out[4164] = ~layer0_out[4699] | layer0_out[4698];
    assign layer1_out[4165] = ~(layer0_out[3112] | layer0_out[3113]);
    assign layer1_out[4166] = layer0_out[4518];
    assign layer1_out[4167] = layer0_out[3648] & layer0_out[3649];
    assign layer1_out[4168] = 1'b0;
    assign layer1_out[4169] = layer0_out[3064];
    assign layer1_out[4170] = ~(layer0_out[1072] & layer0_out[1073]);
    assign layer1_out[4171] = ~layer0_out[6242] | layer0_out[6243];
    assign layer1_out[4172] = layer0_out[760] & ~layer0_out[761];
    assign layer1_out[4173] = ~layer0_out[1843] | layer0_out[1842];
    assign layer1_out[4174] = layer0_out[3337] & layer0_out[3338];
    assign layer1_out[4175] = ~(layer0_out[7498] | layer0_out[7499]);
    assign layer1_out[4176] = ~layer0_out[3267] | layer0_out[3268];
    assign layer1_out[4177] = ~layer0_out[2769];
    assign layer1_out[4178] = ~layer0_out[2863];
    assign layer1_out[4179] = ~layer0_out[13] | layer0_out[14];
    assign layer1_out[4180] = ~layer0_out[7104] | layer0_out[7105];
    assign layer1_out[4181] = layer0_out[5473];
    assign layer1_out[4182] = 1'b0;
    assign layer1_out[4183] = layer0_out[946] & ~layer0_out[945];
    assign layer1_out[4184] = ~layer0_out[171];
    assign layer1_out[4185] = ~layer0_out[3867];
    assign layer1_out[4186] = ~layer0_out[1806];
    assign layer1_out[4187] = ~layer0_out[7031];
    assign layer1_out[4188] = ~layer0_out[3045] | layer0_out[3044];
    assign layer1_out[4189] = ~layer0_out[5589] | layer0_out[5590];
    assign layer1_out[4190] = layer0_out[1146] & ~layer0_out[1145];
    assign layer1_out[4191] = 1'b0;
    assign layer1_out[4192] = layer0_out[7785];
    assign layer1_out[4193] = ~(layer0_out[3870] ^ layer0_out[3871]);
    assign layer1_out[4194] = layer0_out[1421] & ~layer0_out[1420];
    assign layer1_out[4195] = layer0_out[454];
    assign layer1_out[4196] = ~layer0_out[2714];
    assign layer1_out[4197] = ~layer0_out[6332];
    assign layer1_out[4198] = layer0_out[790] & layer0_out[791];
    assign layer1_out[4199] = ~(layer0_out[3977] ^ layer0_out[3978]);
    assign layer1_out[4200] = layer0_out[3634] | layer0_out[3635];
    assign layer1_out[4201] = layer0_out[6192];
    assign layer1_out[4202] = ~layer0_out[3393];
    assign layer1_out[4203] = ~(layer0_out[1963] | layer0_out[1964]);
    assign layer1_out[4204] = ~(layer0_out[634] & layer0_out[635]);
    assign layer1_out[4205] = ~(layer0_out[7359] | layer0_out[7360]);
    assign layer1_out[4206] = layer0_out[7043] ^ layer0_out[7044];
    assign layer1_out[4207] = layer0_out[3392] | layer0_out[3393];
    assign layer1_out[4208] = ~layer0_out[4927] | layer0_out[4928];
    assign layer1_out[4209] = layer0_out[7913] & ~layer0_out[7912];
    assign layer1_out[4210] = ~layer0_out[284];
    assign layer1_out[4211] = layer0_out[6556];
    assign layer1_out[4212] = ~(layer0_out[7550] | layer0_out[7551]);
    assign layer1_out[4213] = layer0_out[4704];
    assign layer1_out[4214] = layer0_out[1702] ^ layer0_out[1703];
    assign layer1_out[4215] = ~layer0_out[2050];
    assign layer1_out[4216] = ~layer0_out[7489] | layer0_out[7490];
    assign layer1_out[4217] = layer0_out[5735] | layer0_out[5736];
    assign layer1_out[4218] = ~layer0_out[7634] | layer0_out[7635];
    assign layer1_out[4219] = layer0_out[6834] | layer0_out[6835];
    assign layer1_out[4220] = ~(layer0_out[6768] ^ layer0_out[6769]);
    assign layer1_out[4221] = 1'b1;
    assign layer1_out[4222] = layer0_out[7739] & layer0_out[7740];
    assign layer1_out[4223] = ~(layer0_out[1005] | layer0_out[1006]);
    assign layer1_out[4224] = ~layer0_out[134] | layer0_out[133];
    assign layer1_out[4225] = layer0_out[3668];
    assign layer1_out[4226] = layer0_out[5957] & ~layer0_out[5958];
    assign layer1_out[4227] = ~(layer0_out[3917] | layer0_out[3918]);
    assign layer1_out[4228] = layer0_out[7135];
    assign layer1_out[4229] = ~layer0_out[1276] | layer0_out[1277];
    assign layer1_out[4230] = layer0_out[6493];
    assign layer1_out[4231] = ~layer0_out[1603] | layer0_out[1604];
    assign layer1_out[4232] = layer0_out[7897] & layer0_out[7898];
    assign layer1_out[4233] = ~layer0_out[1517];
    assign layer1_out[4234] = layer0_out[3678] | layer0_out[3679];
    assign layer1_out[4235] = ~layer0_out[5058] | layer0_out[5059];
    assign layer1_out[4236] = layer0_out[5312] & layer0_out[5313];
    assign layer1_out[4237] = ~layer0_out[3574];
    assign layer1_out[4238] = 1'b1;
    assign layer1_out[4239] = layer0_out[3624];
    assign layer1_out[4240] = layer0_out[2283] & layer0_out[2284];
    assign layer1_out[4241] = ~layer0_out[5103] | layer0_out[5104];
    assign layer1_out[4242] = layer0_out[7187];
    assign layer1_out[4243] = layer0_out[48];
    assign layer1_out[4244] = ~layer0_out[1417] | layer0_out[1418];
    assign layer1_out[4245] = layer0_out[183] ^ layer0_out[184];
    assign layer1_out[4246] = ~layer0_out[7439];
    assign layer1_out[4247] = layer0_out[2623];
    assign layer1_out[4248] = ~layer0_out[2444] | layer0_out[2445];
    assign layer1_out[4249] = ~layer0_out[1961] | layer0_out[1962];
    assign layer1_out[4250] = ~(layer0_out[788] | layer0_out[789]);
    assign layer1_out[4251] = ~layer0_out[144] | layer0_out[145];
    assign layer1_out[4252] = ~(layer0_out[2740] | layer0_out[2741]);
    assign layer1_out[4253] = layer0_out[198] & ~layer0_out[197];
    assign layer1_out[4254] = layer0_out[6252] | layer0_out[6253];
    assign layer1_out[4255] = layer0_out[3542];
    assign layer1_out[4256] = 1'b1;
    assign layer1_out[4257] = layer0_out[7344] & layer0_out[7345];
    assign layer1_out[4258] = layer0_out[1058] ^ layer0_out[1059];
    assign layer1_out[4259] = ~(layer0_out[2849] & layer0_out[2850]);
    assign layer1_out[4260] = layer0_out[3287];
    assign layer1_out[4261] = ~(layer0_out[4811] & layer0_out[4812]);
    assign layer1_out[4262] = ~layer0_out[5253];
    assign layer1_out[4263] = layer0_out[5335] | layer0_out[5336];
    assign layer1_out[4264] = ~(layer0_out[7081] & layer0_out[7082]);
    assign layer1_out[4265] = layer0_out[3673] & ~layer0_out[3672];
    assign layer1_out[4266] = 1'b1;
    assign layer1_out[4267] = layer0_out[2537] | layer0_out[2538];
    assign layer1_out[4268] = layer0_out[543] | layer0_out[544];
    assign layer1_out[4269] = layer0_out[381] | layer0_out[382];
    assign layer1_out[4270] = ~layer0_out[7606];
    assign layer1_out[4271] = ~layer0_out[6327];
    assign layer1_out[4272] = layer0_out[5434] & layer0_out[5435];
    assign layer1_out[4273] = layer0_out[5336];
    assign layer1_out[4274] = layer0_out[7761];
    assign layer1_out[4275] = layer0_out[7050] & ~layer0_out[7049];
    assign layer1_out[4276] = ~layer0_out[2294] | layer0_out[2295];
    assign layer1_out[4277] = ~layer0_out[5145];
    assign layer1_out[4278] = ~layer0_out[5224];
    assign layer1_out[4279] = 1'b1;
    assign layer1_out[4280] = 1'b1;
    assign layer1_out[4281] = layer0_out[4461];
    assign layer1_out[4282] = layer0_out[2976] ^ layer0_out[2977];
    assign layer1_out[4283] = layer0_out[6844] | layer0_out[6845];
    assign layer1_out[4284] = ~layer0_out[3303];
    assign layer1_out[4285] = layer0_out[4939];
    assign layer1_out[4286] = ~(layer0_out[6359] & layer0_out[6360]);
    assign layer1_out[4287] = layer0_out[6567];
    assign layer1_out[4288] = layer0_out[1844] & ~layer0_out[1845];
    assign layer1_out[4289] = layer0_out[7227];
    assign layer1_out[4290] = ~layer0_out[709] | layer0_out[710];
    assign layer1_out[4291] = ~layer0_out[2196] | layer0_out[2195];
    assign layer1_out[4292] = ~layer0_out[3127] | layer0_out[3128];
    assign layer1_out[4293] = layer0_out[4658] | layer0_out[4659];
    assign layer1_out[4294] = layer0_out[2914];
    assign layer1_out[4295] = ~(layer0_out[4373] ^ layer0_out[4374]);
    assign layer1_out[4296] = ~layer0_out[4353] | layer0_out[4354];
    assign layer1_out[4297] = ~(layer0_out[6119] | layer0_out[6120]);
    assign layer1_out[4298] = layer0_out[4153];
    assign layer1_out[4299] = layer0_out[5824];
    assign layer1_out[4300] = layer0_out[3327];
    assign layer1_out[4301] = layer0_out[3217];
    assign layer1_out[4302] = layer0_out[5420] & ~layer0_out[5421];
    assign layer1_out[4303] = layer0_out[2221] | layer0_out[2222];
    assign layer1_out[4304] = ~layer0_out[1918];
    assign layer1_out[4305] = layer0_out[110];
    assign layer1_out[4306] = ~layer0_out[5843];
    assign layer1_out[4307] = ~layer0_out[1579];
    assign layer1_out[4308] = ~(layer0_out[5891] & layer0_out[5892]);
    assign layer1_out[4309] = ~layer0_out[4626] | layer0_out[4625];
    assign layer1_out[4310] = ~(layer0_out[6355] | layer0_out[6356]);
    assign layer1_out[4311] = layer0_out[2803];
    assign layer1_out[4312] = layer0_out[781] & ~layer0_out[782];
    assign layer1_out[4313] = ~(layer0_out[843] & layer0_out[844]);
    assign layer1_out[4314] = layer0_out[4327] & ~layer0_out[4326];
    assign layer1_out[4315] = ~layer0_out[5287] | layer0_out[5286];
    assign layer1_out[4316] = ~layer0_out[7426] | layer0_out[7427];
    assign layer1_out[4317] = ~layer0_out[7674];
    assign layer1_out[4318] = layer0_out[6445] & ~layer0_out[6444];
    assign layer1_out[4319] = layer0_out[7477];
    assign layer1_out[4320] = ~layer0_out[1625] | layer0_out[1624];
    assign layer1_out[4321] = ~layer0_out[5463] | layer0_out[5462];
    assign layer1_out[4322] = ~layer0_out[3730] | layer0_out[3731];
    assign layer1_out[4323] = ~(layer0_out[1529] & layer0_out[1530]);
    assign layer1_out[4324] = layer0_out[5491];
    assign layer1_out[4325] = layer0_out[3445] | layer0_out[3446];
    assign layer1_out[4326] = layer0_out[6979];
    assign layer1_out[4327] = layer0_out[7884] ^ layer0_out[7885];
    assign layer1_out[4328] = layer0_out[2124] ^ layer0_out[2125];
    assign layer1_out[4329] = layer0_out[3649] ^ layer0_out[3650];
    assign layer1_out[4330] = layer0_out[6108] | layer0_out[6109];
    assign layer1_out[4331] = layer0_out[6171];
    assign layer1_out[4332] = ~(layer0_out[6721] | layer0_out[6722]);
    assign layer1_out[4333] = ~layer0_out[1734] | layer0_out[1733];
    assign layer1_out[4334] = layer0_out[2010];
    assign layer1_out[4335] = ~layer0_out[6915];
    assign layer1_out[4336] = ~(layer0_out[5507] ^ layer0_out[5508]);
    assign layer1_out[4337] = ~(layer0_out[912] ^ layer0_out[913]);
    assign layer1_out[4338] = ~layer0_out[3895];
    assign layer1_out[4339] = layer0_out[7510] & ~layer0_out[7511];
    assign layer1_out[4340] = ~layer0_out[5464];
    assign layer1_out[4341] = ~(layer0_out[1067] | layer0_out[1068]);
    assign layer1_out[4342] = layer0_out[478];
    assign layer1_out[4343] = 1'b0;
    assign layer1_out[4344] = layer0_out[2229] ^ layer0_out[2230];
    assign layer1_out[4345] = layer0_out[3361];
    assign layer1_out[4346] = ~(layer0_out[2724] | layer0_out[2725]);
    assign layer1_out[4347] = ~layer0_out[2619];
    assign layer1_out[4348] = ~(layer0_out[6361] & layer0_out[6362]);
    assign layer1_out[4349] = layer0_out[3557] & ~layer0_out[3556];
    assign layer1_out[4350] = layer0_out[6739] | layer0_out[6740];
    assign layer1_out[4351] = layer0_out[1491];
    assign layer1_out[4352] = ~layer0_out[7661];
    assign layer1_out[4353] = ~layer0_out[559] | layer0_out[558];
    assign layer1_out[4354] = layer0_out[2618];
    assign layer1_out[4355] = layer0_out[6363] & layer0_out[6364];
    assign layer1_out[4356] = ~layer0_out[5618] | layer0_out[5617];
    assign layer1_out[4357] = layer0_out[3757];
    assign layer1_out[4358] = ~layer0_out[3364];
    assign layer1_out[4359] = ~layer0_out[524] | layer0_out[525];
    assign layer1_out[4360] = ~layer0_out[7449] | layer0_out[7448];
    assign layer1_out[4361] = layer0_out[900];
    assign layer1_out[4362] = ~(layer0_out[4366] | layer0_out[4367]);
    assign layer1_out[4363] = ~layer0_out[6489] | layer0_out[6490];
    assign layer1_out[4364] = ~layer0_out[7906] | layer0_out[7905];
    assign layer1_out[4365] = layer0_out[399] & ~layer0_out[400];
    assign layer1_out[4366] = ~(layer0_out[5770] & layer0_out[5771]);
    assign layer1_out[4367] = layer0_out[7713] & ~layer0_out[7712];
    assign layer1_out[4368] = ~layer0_out[2776];
    assign layer1_out[4369] = layer0_out[275] & ~layer0_out[274];
    assign layer1_out[4370] = ~(layer0_out[1319] & layer0_out[1320]);
    assign layer1_out[4371] = ~(layer0_out[1095] & layer0_out[1096]);
    assign layer1_out[4372] = ~layer0_out[6395] | layer0_out[6396];
    assign layer1_out[4373] = ~layer0_out[2806] | layer0_out[2807];
    assign layer1_out[4374] = 1'b0;
    assign layer1_out[4375] = ~layer0_out[1347] | layer0_out[1346];
    assign layer1_out[4376] = layer0_out[6515] & ~layer0_out[6514];
    assign layer1_out[4377] = layer0_out[1637];
    assign layer1_out[4378] = ~layer0_out[2363];
    assign layer1_out[4379] = layer0_out[6265] ^ layer0_out[6266];
    assign layer1_out[4380] = 1'b1;
    assign layer1_out[4381] = layer0_out[2441] & layer0_out[2442];
    assign layer1_out[4382] = ~layer0_out[3178];
    assign layer1_out[4383] = layer0_out[7124] & ~layer0_out[7125];
    assign layer1_out[4384] = layer0_out[7158] ^ layer0_out[7159];
    assign layer1_out[4385] = layer0_out[7334] & ~layer0_out[7333];
    assign layer1_out[4386] = ~layer0_out[7744] | layer0_out[7745];
    assign layer1_out[4387] = layer0_out[5144] & ~layer0_out[5143];
    assign layer1_out[4388] = layer0_out[4818];
    assign layer1_out[4389] = layer0_out[1403] & layer0_out[1404];
    assign layer1_out[4390] = layer0_out[3587] | layer0_out[3588];
    assign layer1_out[4391] = layer0_out[887] ^ layer0_out[888];
    assign layer1_out[4392] = 1'b1;
    assign layer1_out[4393] = ~layer0_out[2177];
    assign layer1_out[4394] = layer0_out[4266] & ~layer0_out[4265];
    assign layer1_out[4395] = ~(layer0_out[4511] & layer0_out[4512]);
    assign layer1_out[4396] = ~layer0_out[7606] | layer0_out[7607];
    assign layer1_out[4397] = ~(layer0_out[5358] | layer0_out[5359]);
    assign layer1_out[4398] = ~layer0_out[6723] | layer0_out[6724];
    assign layer1_out[4399] = layer0_out[5645];
    assign layer1_out[4400] = ~(layer0_out[3310] & layer0_out[3311]);
    assign layer1_out[4401] = 1'b0;
    assign layer1_out[4402] = layer0_out[211] | layer0_out[212];
    assign layer1_out[4403] = layer0_out[6934] & ~layer0_out[6933];
    assign layer1_out[4404] = layer0_out[344] | layer0_out[345];
    assign layer1_out[4405] = ~(layer0_out[2944] & layer0_out[2945]);
    assign layer1_out[4406] = 1'b1;
    assign layer1_out[4407] = layer0_out[3352] | layer0_out[3353];
    assign layer1_out[4408] = layer0_out[6537] & layer0_out[6538];
    assign layer1_out[4409] = ~layer0_out[2264];
    assign layer1_out[4410] = ~(layer0_out[4525] ^ layer0_out[4526]);
    assign layer1_out[4411] = ~layer0_out[2842] | layer0_out[2843];
    assign layer1_out[4412] = ~(layer0_out[1285] & layer0_out[1286]);
    assign layer1_out[4413] = layer0_out[6560] & ~layer0_out[6559];
    assign layer1_out[4414] = 1'b1;
    assign layer1_out[4415] = ~layer0_out[5049];
    assign layer1_out[4416] = layer0_out[4062];
    assign layer1_out[4417] = ~(layer0_out[6396] & layer0_out[6397]);
    assign layer1_out[4418] = 1'b1;
    assign layer1_out[4419] = layer0_out[4812] & layer0_out[4813];
    assign layer1_out[4420] = ~layer0_out[3999];
    assign layer1_out[4421] = layer0_out[3863] & ~layer0_out[3864];
    assign layer1_out[4422] = layer0_out[5155];
    assign layer1_out[4423] = layer0_out[7587];
    assign layer1_out[4424] = ~(layer0_out[1047] ^ layer0_out[1048]);
    assign layer1_out[4425] = layer0_out[6576];
    assign layer1_out[4426] = layer0_out[704];
    assign layer1_out[4427] = layer0_out[3729] & ~layer0_out[3730];
    assign layer1_out[4428] = layer0_out[7459] | layer0_out[7460];
    assign layer1_out[4429] = layer0_out[7714] | layer0_out[7715];
    assign layer1_out[4430] = layer0_out[1055];
    assign layer1_out[4431] = ~layer0_out[7571];
    assign layer1_out[4432] = layer0_out[3376];
    assign layer1_out[4433] = layer0_out[451] | layer0_out[452];
    assign layer1_out[4434] = ~layer0_out[6596];
    assign layer1_out[4435] = layer0_out[2832] & ~layer0_out[2833];
    assign layer1_out[4436] = ~(layer0_out[371] & layer0_out[372]);
    assign layer1_out[4437] = layer0_out[3033];
    assign layer1_out[4438] = 1'b0;
    assign layer1_out[4439] = ~layer0_out[6305];
    assign layer1_out[4440] = layer0_out[1883];
    assign layer1_out[4441] = 1'b0;
    assign layer1_out[4442] = layer0_out[5924] | layer0_out[5925];
    assign layer1_out[4443] = ~layer0_out[4864] | layer0_out[4863];
    assign layer1_out[4444] = ~layer0_out[2853];
    assign layer1_out[4445] = ~(layer0_out[4850] | layer0_out[4851]);
    assign layer1_out[4446] = layer0_out[5115];
    assign layer1_out[4447] = 1'b0;
    assign layer1_out[4448] = ~layer0_out[3191];
    assign layer1_out[4449] = 1'b1;
    assign layer1_out[4450] = 1'b0;
    assign layer1_out[4451] = layer0_out[6336] & ~layer0_out[6337];
    assign layer1_out[4452] = layer0_out[6746];
    assign layer1_out[4453] = ~(layer0_out[3242] & layer0_out[3243]);
    assign layer1_out[4454] = ~layer0_out[2558] | layer0_out[2557];
    assign layer1_out[4455] = ~layer0_out[572];
    assign layer1_out[4456] = ~layer0_out[1213];
    assign layer1_out[4457] = layer0_out[2145] & layer0_out[2146];
    assign layer1_out[4458] = ~layer0_out[6380];
    assign layer1_out[4459] = layer0_out[7112] | layer0_out[7113];
    assign layer1_out[4460] = ~layer0_out[259] | layer0_out[260];
    assign layer1_out[4461] = ~layer0_out[5795] | layer0_out[5794];
    assign layer1_out[4462] = layer0_out[3737];
    assign layer1_out[4463] = 1'b0;
    assign layer1_out[4464] = 1'b1;
    assign layer1_out[4465] = ~(layer0_out[6206] & layer0_out[6207]);
    assign layer1_out[4466] = ~layer0_out[2517];
    assign layer1_out[4467] = ~(layer0_out[2654] ^ layer0_out[2655]);
    assign layer1_out[4468] = ~(layer0_out[598] | layer0_out[599]);
    assign layer1_out[4469] = layer0_out[4514] ^ layer0_out[4515];
    assign layer1_out[4470] = layer0_out[5977];
    assign layer1_out[4471] = layer0_out[4268] ^ layer0_out[4269];
    assign layer1_out[4472] = ~layer0_out[2339] | layer0_out[2340];
    assign layer1_out[4473] = layer0_out[6910] & ~layer0_out[6909];
    assign layer1_out[4474] = ~layer0_out[6633] | layer0_out[6634];
    assign layer1_out[4475] = layer0_out[4891];
    assign layer1_out[4476] = layer0_out[65] & layer0_out[66];
    assign layer1_out[4477] = ~(layer0_out[807] | layer0_out[808]);
    assign layer1_out[4478] = ~layer0_out[3343] | layer0_out[3344];
    assign layer1_out[4479] = ~layer0_out[3052] | layer0_out[3053];
    assign layer1_out[4480] = ~layer0_out[1189];
    assign layer1_out[4481] = ~layer0_out[2677];
    assign layer1_out[4482] = ~(layer0_out[6981] | layer0_out[6982]);
    assign layer1_out[4483] = layer0_out[3543];
    assign layer1_out[4484] = ~layer0_out[6853] | layer0_out[6852];
    assign layer1_out[4485] = layer0_out[3073];
    assign layer1_out[4486] = ~(layer0_out[6132] ^ layer0_out[6133]);
    assign layer1_out[4487] = layer0_out[4628] ^ layer0_out[4629];
    assign layer1_out[4488] = layer0_out[4086] | layer0_out[4087];
    assign layer1_out[4489] = ~layer0_out[3367] | layer0_out[3366];
    assign layer1_out[4490] = ~layer0_out[3264];
    assign layer1_out[4491] = layer0_out[7127] & ~layer0_out[7126];
    assign layer1_out[4492] = layer0_out[6527] & layer0_out[6528];
    assign layer1_out[4493] = ~layer0_out[1606] | layer0_out[1605];
    assign layer1_out[4494] = ~(layer0_out[2460] & layer0_out[2461]);
    assign layer1_out[4495] = ~layer0_out[3065] | layer0_out[3066];
    assign layer1_out[4496] = layer0_out[3163] ^ layer0_out[3164];
    assign layer1_out[4497] = ~layer0_out[3984];
    assign layer1_out[4498] = ~layer0_out[7114];
    assign layer1_out[4499] = layer0_out[2799];
    assign layer1_out[4500] = ~layer0_out[479] | layer0_out[480];
    assign layer1_out[4501] = ~layer0_out[1644];
    assign layer1_out[4502] = ~(layer0_out[3227] & layer0_out[3228]);
    assign layer1_out[4503] = layer0_out[1496] & ~layer0_out[1497];
    assign layer1_out[4504] = ~layer0_out[7969] | layer0_out[7968];
    assign layer1_out[4505] = layer0_out[3580];
    assign layer1_out[4506] = ~(layer0_out[1986] & layer0_out[1987]);
    assign layer1_out[4507] = ~(layer0_out[3283] & layer0_out[3284]);
    assign layer1_out[4508] = ~layer0_out[1686];
    assign layer1_out[4509] = layer0_out[2767] ^ layer0_out[2768];
    assign layer1_out[4510] = layer0_out[620] & layer0_out[621];
    assign layer1_out[4511] = ~(layer0_out[3160] & layer0_out[3161]);
    assign layer1_out[4512] = ~layer0_out[5561] | layer0_out[5560];
    assign layer1_out[4513] = layer0_out[5970] & ~layer0_out[5971];
    assign layer1_out[4514] = ~layer0_out[2736];
    assign layer1_out[4515] = ~(layer0_out[975] & layer0_out[976]);
    assign layer1_out[4516] = layer0_out[1808];
    assign layer1_out[4517] = layer0_out[227];
    assign layer1_out[4518] = layer0_out[5863] & ~layer0_out[5862];
    assign layer1_out[4519] = ~(layer0_out[2709] | layer0_out[2710]);
    assign layer1_out[4520] = ~layer0_out[6486];
    assign layer1_out[4521] = ~layer0_out[2258];
    assign layer1_out[4522] = ~(layer0_out[2875] | layer0_out[2876]);
    assign layer1_out[4523] = layer0_out[3822] & ~layer0_out[3823];
    assign layer1_out[4524] = layer0_out[7596];
    assign layer1_out[4525] = ~layer0_out[7428];
    assign layer1_out[4526] = ~layer0_out[6375];
    assign layer1_out[4527] = layer0_out[3699];
    assign layer1_out[4528] = ~(layer0_out[3264] ^ layer0_out[3265]);
    assign layer1_out[4529] = ~layer0_out[7718] | layer0_out[7719];
    assign layer1_out[4530] = layer0_out[5750] | layer0_out[5751];
    assign layer1_out[4531] = ~layer0_out[5460];
    assign layer1_out[4532] = 1'b1;
    assign layer1_out[4533] = layer0_out[5869];
    assign layer1_out[4534] = ~layer0_out[6285] | layer0_out[6284];
    assign layer1_out[4535] = ~(layer0_out[5992] & layer0_out[5993]);
    assign layer1_out[4536] = ~(layer0_out[5607] | layer0_out[5608]);
    assign layer1_out[4537] = ~layer0_out[5607];
    assign layer1_out[4538] = ~(layer0_out[1268] & layer0_out[1269]);
    assign layer1_out[4539] = ~(layer0_out[3551] | layer0_out[3552]);
    assign layer1_out[4540] = layer0_out[3974] | layer0_out[3975];
    assign layer1_out[4541] = layer0_out[362] | layer0_out[363];
    assign layer1_out[4542] = ~layer0_out[4937];
    assign layer1_out[4543] = ~layer0_out[4222];
    assign layer1_out[4544] = ~(layer0_out[7409] ^ layer0_out[7410]);
    assign layer1_out[4545] = layer0_out[1905] & ~layer0_out[1904];
    assign layer1_out[4546] = layer0_out[7039];
    assign layer1_out[4547] = ~layer0_out[246] | layer0_out[247];
    assign layer1_out[4548] = ~(layer0_out[6266] & layer0_out[6267]);
    assign layer1_out[4549] = ~layer0_out[6434] | layer0_out[6435];
    assign layer1_out[4550] = layer0_out[7520] & ~layer0_out[7521];
    assign layer1_out[4551] = layer0_out[1341] & layer0_out[1342];
    assign layer1_out[4552] = 1'b0;
    assign layer1_out[4553] = ~(layer0_out[3180] | layer0_out[3181]);
    assign layer1_out[4554] = ~layer0_out[3330];
    assign layer1_out[4555] = layer0_out[6584] & ~layer0_out[6585];
    assign layer1_out[4556] = layer0_out[243];
    assign layer1_out[4557] = layer0_out[1274];
    assign layer1_out[4558] = ~layer0_out[6711] | layer0_out[6710];
    assign layer1_out[4559] = layer0_out[6178];
    assign layer1_out[4560] = layer0_out[7972] & layer0_out[7973];
    assign layer1_out[4561] = layer0_out[218] | layer0_out[219];
    assign layer1_out[4562] = layer0_out[1378];
    assign layer1_out[4563] = ~(layer0_out[7511] & layer0_out[7512]);
    assign layer1_out[4564] = layer0_out[549] & layer0_out[550];
    assign layer1_out[4565] = layer0_out[1487];
    assign layer1_out[4566] = ~(layer0_out[1314] & layer0_out[1315]);
    assign layer1_out[4567] = layer0_out[4931] & ~layer0_out[4932];
    assign layer1_out[4568] = 1'b1;
    assign layer1_out[4569] = ~(layer0_out[4648] & layer0_out[4649]);
    assign layer1_out[4570] = layer0_out[5311] & layer0_out[5312];
    assign layer1_out[4571] = layer0_out[2364] & ~layer0_out[2363];
    assign layer1_out[4572] = layer0_out[3512] | layer0_out[3513];
    assign layer1_out[4573] = layer0_out[2514] & ~layer0_out[2515];
    assign layer1_out[4574] = 1'b1;
    assign layer1_out[4575] = ~layer0_out[2282];
    assign layer1_out[4576] = layer0_out[1268];
    assign layer1_out[4577] = layer0_out[4899];
    assign layer1_out[4578] = layer0_out[418] & ~layer0_out[417];
    assign layer1_out[4579] = layer0_out[4629];
    assign layer1_out[4580] = layer0_out[3625] | layer0_out[3626];
    assign layer1_out[4581] = layer0_out[1576] | layer0_out[1577];
    assign layer1_out[4582] = layer0_out[2916] & ~layer0_out[2915];
    assign layer1_out[4583] = 1'b0;
    assign layer1_out[4584] = layer0_out[141] & layer0_out[142];
    assign layer1_out[4585] = layer0_out[7060];
    assign layer1_out[4586] = ~layer0_out[7452];
    assign layer1_out[4587] = layer0_out[7102] | layer0_out[7103];
    assign layer1_out[4588] = ~(layer0_out[4534] & layer0_out[4535]);
    assign layer1_out[4589] = ~layer0_out[6768];
    assign layer1_out[4590] = ~layer0_out[1355] | layer0_out[1356];
    assign layer1_out[4591] = layer0_out[2105] & layer0_out[2106];
    assign layer1_out[4592] = ~(layer0_out[5995] & layer0_out[5996]);
    assign layer1_out[4593] = layer0_out[6232] & ~layer0_out[6231];
    assign layer1_out[4594] = layer0_out[5653];
    assign layer1_out[4595] = layer0_out[4320];
    assign layer1_out[4596] = ~layer0_out[652] | layer0_out[651];
    assign layer1_out[4597] = layer0_out[2797] & ~layer0_out[2796];
    assign layer1_out[4598] = layer0_out[2183] | layer0_out[2184];
    assign layer1_out[4599] = layer0_out[7700];
    assign layer1_out[4600] = 1'b1;
    assign layer1_out[4601] = layer0_out[2370] & ~layer0_out[2369];
    assign layer1_out[4602] = ~layer0_out[7773] | layer0_out[7774];
    assign layer1_out[4603] = ~(layer0_out[6123] & layer0_out[6124]);
    assign layer1_out[4604] = ~layer0_out[5690] | layer0_out[5689];
    assign layer1_out[4605] = ~(layer0_out[2155] & layer0_out[2156]);
    assign layer1_out[4606] = layer0_out[3480];
    assign layer1_out[4607] = ~layer0_out[3750] | layer0_out[3749];
    assign layer1_out[4608] = layer0_out[5654] & layer0_out[5655];
    assign layer1_out[4609] = ~layer0_out[1915];
    assign layer1_out[4610] = layer0_out[7393] & ~layer0_out[7394];
    assign layer1_out[4611] = ~layer0_out[5428] | layer0_out[5429];
    assign layer1_out[4612] = layer0_out[333] | layer0_out[334];
    assign layer1_out[4613] = layer0_out[6376] & ~layer0_out[6377];
    assign layer1_out[4614] = ~layer0_out[4644];
    assign layer1_out[4615] = ~layer0_out[4383] | layer0_out[4384];
    assign layer1_out[4616] = ~layer0_out[3438];
    assign layer1_out[4617] = ~layer0_out[2001];
    assign layer1_out[4618] = layer0_out[7822] & ~layer0_out[7821];
    assign layer1_out[4619] = layer0_out[897] | layer0_out[898];
    assign layer1_out[4620] = ~(layer0_out[4198] ^ layer0_out[4199]);
    assign layer1_out[4621] = ~layer0_out[3929];
    assign layer1_out[4622] = ~layer0_out[3373];
    assign layer1_out[4623] = layer0_out[1227] & layer0_out[1228];
    assign layer1_out[4624] = ~(layer0_out[2774] | layer0_out[2775]);
    assign layer1_out[4625] = ~(layer0_out[4082] | layer0_out[4083]);
    assign layer1_out[4626] = ~(layer0_out[7925] | layer0_out[7926]);
    assign layer1_out[4627] = ~layer0_out[112] | layer0_out[111];
    assign layer1_out[4628] = ~layer0_out[5598] | layer0_out[5597];
    assign layer1_out[4629] = layer0_out[4584];
    assign layer1_out[4630] = ~(layer0_out[7211] | layer0_out[7212]);
    assign layer1_out[4631] = layer0_out[5248] & layer0_out[5249];
    assign layer1_out[4632] = 1'b1;
    assign layer1_out[4633] = layer0_out[1463] & ~layer0_out[1462];
    assign layer1_out[4634] = ~layer0_out[6999] | layer0_out[6998];
    assign layer1_out[4635] = layer0_out[7326];
    assign layer1_out[4636] = 1'b1;
    assign layer1_out[4637] = ~layer0_out[3313];
    assign layer1_out[4638] = layer0_out[51] | layer0_out[52];
    assign layer1_out[4639] = ~(layer0_out[5240] | layer0_out[5241]);
    assign layer1_out[4640] = layer0_out[1370];
    assign layer1_out[4641] = ~layer0_out[5739];
    assign layer1_out[4642] = layer0_out[2795] & ~layer0_out[2796];
    assign layer1_out[4643] = ~layer0_out[1740];
    assign layer1_out[4644] = 1'b0;
    assign layer1_out[4645] = ~layer0_out[4184] | layer0_out[4185];
    assign layer1_out[4646] = ~(layer0_out[80] & layer0_out[81]);
    assign layer1_out[4647] = ~(layer0_out[4687] ^ layer0_out[4688]);
    assign layer1_out[4648] = ~layer0_out[611] | layer0_out[612];
    assign layer1_out[4649] = ~layer0_out[6988];
    assign layer1_out[4650] = ~layer0_out[3927] | layer0_out[3928];
    assign layer1_out[4651] = layer0_out[5327];
    assign layer1_out[4652] = ~layer0_out[3721];
    assign layer1_out[4653] = ~layer0_out[7942];
    assign layer1_out[4654] = ~(layer0_out[74] & layer0_out[75]);
    assign layer1_out[4655] = layer0_out[309] & ~layer0_out[310];
    assign layer1_out[4656] = layer0_out[539] | layer0_out[540];
    assign layer1_out[4657] = ~(layer0_out[148] | layer0_out[149]);
    assign layer1_out[4658] = layer0_out[4801];
    assign layer1_out[4659] = ~(layer0_out[7733] | layer0_out[7734]);
    assign layer1_out[4660] = ~(layer0_out[2731] & layer0_out[2732]);
    assign layer1_out[4661] = layer0_out[1880];
    assign layer1_out[4662] = ~layer0_out[2097];
    assign layer1_out[4663] = ~(layer0_out[4733] ^ layer0_out[4734]);
    assign layer1_out[4664] = ~layer0_out[2157];
    assign layer1_out[4665] = layer0_out[6296] | layer0_out[6297];
    assign layer1_out[4666] = ~layer0_out[4969];
    assign layer1_out[4667] = layer0_out[3920] & ~layer0_out[3921];
    assign layer1_out[4668] = ~(layer0_out[7794] & layer0_out[7795]);
    assign layer1_out[4669] = ~(layer0_out[5659] | layer0_out[5660]);
    assign layer1_out[4670] = ~(layer0_out[3542] | layer0_out[3543]);
    assign layer1_out[4671] = ~(layer0_out[3804] | layer0_out[3805]);
    assign layer1_out[4672] = ~layer0_out[2098];
    assign layer1_out[4673] = layer0_out[6963];
    assign layer1_out[4674] = ~layer0_out[7494];
    assign layer1_out[4675] = layer0_out[7597] & ~layer0_out[7598];
    assign layer1_out[4676] = ~(layer0_out[832] & layer0_out[833]);
    assign layer1_out[4677] = ~(layer0_out[1363] | layer0_out[1364]);
    assign layer1_out[4678] = layer0_out[1606] ^ layer0_out[1607];
    assign layer1_out[4679] = ~layer0_out[3759] | layer0_out[3760];
    assign layer1_out[4680] = layer0_out[3922];
    assign layer1_out[4681] = layer0_out[2257];
    assign layer1_out[4682] = layer0_out[2857] & ~layer0_out[2856];
    assign layer1_out[4683] = layer0_out[4001];
    assign layer1_out[4684] = ~(layer0_out[1787] | layer0_out[1788]);
    assign layer1_out[4685] = layer0_out[1026];
    assign layer1_out[4686] = layer0_out[91] ^ layer0_out[92];
    assign layer1_out[4687] = ~layer0_out[772];
    assign layer1_out[4688] = layer0_out[6895] ^ layer0_out[6896];
    assign layer1_out[4689] = layer0_out[4989] & ~layer0_out[4990];
    assign layer1_out[4690] = ~layer0_out[4932];
    assign layer1_out[4691] = ~layer0_out[3185];
    assign layer1_out[4692] = ~layer0_out[1220] | layer0_out[1221];
    assign layer1_out[4693] = 1'b0;
    assign layer1_out[4694] = layer0_out[2612] & ~layer0_out[2613];
    assign layer1_out[4695] = layer0_out[1924];
    assign layer1_out[4696] = ~(layer0_out[3155] | layer0_out[3156]);
    assign layer1_out[4697] = layer0_out[1816] & layer0_out[1817];
    assign layer1_out[4698] = ~(layer0_out[3954] | layer0_out[3955]);
    assign layer1_out[4699] = 1'b1;
    assign layer1_out[4700] = ~(layer0_out[7197] | layer0_out[7198]);
    assign layer1_out[4701] = ~layer0_out[3787];
    assign layer1_out[4702] = layer0_out[5714] & layer0_out[5715];
    assign layer1_out[4703] = 1'b1;
    assign layer1_out[4704] = layer0_out[1521] & layer0_out[1522];
    assign layer1_out[4705] = ~layer0_out[1520] | layer0_out[1519];
    assign layer1_out[4706] = layer0_out[3501] & layer0_out[3502];
    assign layer1_out[4707] = layer0_out[2743];
    assign layer1_out[4708] = ~(layer0_out[1907] & layer0_out[1908]);
    assign layer1_out[4709] = ~layer0_out[4313];
    assign layer1_out[4710] = layer0_out[5133] & ~layer0_out[5134];
    assign layer1_out[4711] = ~layer0_out[4697];
    assign layer1_out[4712] = layer0_out[7207];
    assign layer1_out[4713] = ~layer0_out[3561];
    assign layer1_out[4714] = layer0_out[416] & ~layer0_out[415];
    assign layer1_out[4715] = ~layer0_out[4505];
    assign layer1_out[4716] = ~layer0_out[1855];
    assign layer1_out[4717] = layer0_out[5212] & ~layer0_out[5213];
    assign layer1_out[4718] = ~layer0_out[4976];
    assign layer1_out[4719] = layer0_out[1622] ^ layer0_out[1623];
    assign layer1_out[4720] = layer0_out[4989];
    assign layer1_out[4721] = ~layer0_out[2739];
    assign layer1_out[4722] = layer0_out[6614];
    assign layer1_out[4723] = layer0_out[4120] & layer0_out[4121];
    assign layer1_out[4724] = layer0_out[916];
    assign layer1_out[4725] = layer0_out[685];
    assign layer1_out[4726] = layer0_out[1378] & ~layer0_out[1377];
    assign layer1_out[4727] = ~layer0_out[4896] | layer0_out[4897];
    assign layer1_out[4728] = ~layer0_out[528];
    assign layer1_out[4729] = layer0_out[2755] & ~layer0_out[2756];
    assign layer1_out[4730] = layer0_out[4601] ^ layer0_out[4602];
    assign layer1_out[4731] = layer0_out[6651];
    assign layer1_out[4732] = ~layer0_out[2099];
    assign layer1_out[4733] = 1'b0;
    assign layer1_out[4734] = ~(layer0_out[5531] ^ layer0_out[5532]);
    assign layer1_out[4735] = ~layer0_out[4783] | layer0_out[4784];
    assign layer1_out[4736] = ~layer0_out[1169];
    assign layer1_out[4737] = ~layer0_out[7802];
    assign layer1_out[4738] = ~layer0_out[7006];
    assign layer1_out[4739] = layer0_out[1661] & ~layer0_out[1662];
    assign layer1_out[4740] = ~layer0_out[2269] | layer0_out[2268];
    assign layer1_out[4741] = layer0_out[5493] & ~layer0_out[5494];
    assign layer1_out[4742] = ~layer0_out[6168] | layer0_out[6169];
    assign layer1_out[4743] = layer0_out[4485] | layer0_out[4486];
    assign layer1_out[4744] = layer0_out[5760] | layer0_out[5761];
    assign layer1_out[4745] = layer0_out[266] & ~layer0_out[265];
    assign layer1_out[4746] = ~(layer0_out[5110] & layer0_out[5111]);
    assign layer1_out[4747] = layer0_out[6840];
    assign layer1_out[4748] = layer0_out[2670];
    assign layer1_out[4749] = layer0_out[2172] | layer0_out[2173];
    assign layer1_out[4750] = ~(layer0_out[173] ^ layer0_out[174]);
    assign layer1_out[4751] = ~layer0_out[3669];
    assign layer1_out[4752] = layer0_out[1785] | layer0_out[1786];
    assign layer1_out[4753] = ~(layer0_out[6373] ^ layer0_out[6374]);
    assign layer1_out[4754] = layer0_out[4716];
    assign layer1_out[4755] = ~layer0_out[2585] | layer0_out[2584];
    assign layer1_out[4756] = ~layer0_out[6273] | layer0_out[6274];
    assign layer1_out[4757] = layer0_out[2204];
    assign layer1_out[4758] = ~layer0_out[1947];
    assign layer1_out[4759] = layer0_out[132];
    assign layer1_out[4760] = layer0_out[4819];
    assign layer1_out[4761] = layer0_out[187] & ~layer0_out[186];
    assign layer1_out[4762] = ~(layer0_out[1392] & layer0_out[1393]);
    assign layer1_out[4763] = layer0_out[5874] | layer0_out[5875];
    assign layer1_out[4764] = layer0_out[3519];
    assign layer1_out[4765] = ~(layer0_out[2226] & layer0_out[2227]);
    assign layer1_out[4766] = layer0_out[6335];
    assign layer1_out[4767] = layer0_out[2684];
    assign layer1_out[4768] = layer0_out[3317] & ~layer0_out[3318];
    assign layer1_out[4769] = layer0_out[7571] | layer0_out[7572];
    assign layer1_out[4770] = layer0_out[5700] | layer0_out[5701];
    assign layer1_out[4771] = layer0_out[2239] ^ layer0_out[2240];
    assign layer1_out[4772] = layer0_out[4776];
    assign layer1_out[4773] = ~layer0_out[4958];
    assign layer1_out[4774] = ~layer0_out[1017];
    assign layer1_out[4775] = ~layer0_out[5959] | layer0_out[5960];
    assign layer1_out[4776] = layer0_out[5261];
    assign layer1_out[4777] = ~layer0_out[7857] | layer0_out[7856];
    assign layer1_out[4778] = layer0_out[1389] & ~layer0_out[1390];
    assign layer1_out[4779] = layer0_out[1458];
    assign layer1_out[4780] = layer0_out[2119] & ~layer0_out[2118];
    assign layer1_out[4781] = layer0_out[3480] & layer0_out[3481];
    assign layer1_out[4782] = ~layer0_out[2650] | layer0_out[2651];
    assign layer1_out[4783] = layer0_out[467] & ~layer0_out[466];
    assign layer1_out[4784] = ~layer0_out[461];
    assign layer1_out[4785] = layer0_out[2934];
    assign layer1_out[4786] = ~layer0_out[6500];
    assign layer1_out[4787] = layer0_out[5661] & ~layer0_out[5660];
    assign layer1_out[4788] = 1'b0;
    assign layer1_out[4789] = ~layer0_out[4208];
    assign layer1_out[4790] = layer0_out[5610] & ~layer0_out[5611];
    assign layer1_out[4791] = ~layer0_out[4719];
    assign layer1_out[4792] = layer0_out[5341];
    assign layer1_out[4793] = ~layer0_out[3731];
    assign layer1_out[4794] = layer0_out[2652];
    assign layer1_out[4795] = layer0_out[7011] & ~layer0_out[7012];
    assign layer1_out[4796] = layer0_out[4149] & ~layer0_out[4150];
    assign layer1_out[4797] = ~layer0_out[7351];
    assign layer1_out[4798] = ~layer0_out[6994];
    assign layer1_out[4799] = 1'b1;
    assign layer1_out[4800] = layer0_out[869] | layer0_out[870];
    assign layer1_out[4801] = ~layer0_out[3929];
    assign layer1_out[4802] = layer0_out[5441] & layer0_out[5442];
    assign layer1_out[4803] = ~layer0_out[1826];
    assign layer1_out[4804] = layer0_out[1279];
    assign layer1_out[4805] = layer0_out[7687];
    assign layer1_out[4806] = ~layer0_out[5298] | layer0_out[5297];
    assign layer1_out[4807] = layer0_out[6331] & ~layer0_out[6330];
    assign layer1_out[4808] = ~layer0_out[653];
    assign layer1_out[4809] = ~layer0_out[3449];
    assign layer1_out[4810] = layer0_out[141];
    assign layer1_out[4811] = layer0_out[7983];
    assign layer1_out[4812] = layer0_out[7408] | layer0_out[7409];
    assign layer1_out[4813] = layer0_out[2552];
    assign layer1_out[4814] = ~(layer0_out[7579] ^ layer0_out[7580]);
    assign layer1_out[4815] = layer0_out[3850] | layer0_out[3851];
    assign layer1_out[4816] = 1'b1;
    assign layer1_out[4817] = layer0_out[1988];
    assign layer1_out[4818] = ~layer0_out[6996];
    assign layer1_out[4819] = layer0_out[4538] & ~layer0_out[4539];
    assign layer1_out[4820] = ~(layer0_out[1545] | layer0_out[1546]);
    assign layer1_out[4821] = ~layer0_out[4315] | layer0_out[4314];
    assign layer1_out[4822] = ~layer0_out[2780] | layer0_out[2781];
    assign layer1_out[4823] = layer0_out[3990];
    assign layer1_out[4824] = ~layer0_out[5656] | layer0_out[5655];
    assign layer1_out[4825] = layer0_out[296] & ~layer0_out[297];
    assign layer1_out[4826] = ~(layer0_out[2928] | layer0_out[2929]);
    assign layer1_out[4827] = layer0_out[2892] & ~layer0_out[2893];
    assign layer1_out[4828] = layer0_out[5479] | layer0_out[5480];
    assign layer1_out[4829] = layer0_out[848] & ~layer0_out[849];
    assign layer1_out[4830] = ~(layer0_out[6302] & layer0_out[6303]);
    assign layer1_out[4831] = layer0_out[7880] ^ layer0_out[7881];
    assign layer1_out[4832] = layer0_out[5167];
    assign layer1_out[4833] = layer0_out[3436] & ~layer0_out[3435];
    assign layer1_out[4834] = layer0_out[435] | layer0_out[436];
    assign layer1_out[4835] = ~layer0_out[4790];
    assign layer1_out[4836] = ~(layer0_out[6467] & layer0_out[6468]);
    assign layer1_out[4837] = ~(layer0_out[7824] ^ layer0_out[7825]);
    assign layer1_out[4838] = layer0_out[7829] & layer0_out[7830];
    assign layer1_out[4839] = ~layer0_out[3875] | layer0_out[3874];
    assign layer1_out[4840] = layer0_out[523];
    assign layer1_out[4841] = ~layer0_out[2640];
    assign layer1_out[4842] = layer0_out[3596];
    assign layer1_out[4843] = ~layer0_out[7382] | layer0_out[7381];
    assign layer1_out[4844] = 1'b0;
    assign layer1_out[4845] = ~(layer0_out[5072] & layer0_out[5073]);
    assign layer1_out[4846] = ~layer0_out[325] | layer0_out[324];
    assign layer1_out[4847] = 1'b0;
    assign layer1_out[4848] = layer0_out[7676] | layer0_out[7677];
    assign layer1_out[4849] = ~(layer0_out[2218] | layer0_out[2219]);
    assign layer1_out[4850] = ~layer0_out[4486];
    assign layer1_out[4851] = ~(layer0_out[5435] & layer0_out[5436]);
    assign layer1_out[4852] = layer0_out[5390];
    assign layer1_out[4853] = ~layer0_out[2834];
    assign layer1_out[4854] = ~(layer0_out[5611] | layer0_out[5612]);
    assign layer1_out[4855] = ~layer0_out[5053] | layer0_out[5054];
    assign layer1_out[4856] = layer0_out[406];
    assign layer1_out[4857] = ~layer0_out[1995] | layer0_out[1994];
    assign layer1_out[4858] = layer0_out[2760] & layer0_out[2761];
    assign layer1_out[4859] = 1'b0;
    assign layer1_out[4860] = ~(layer0_out[2609] | layer0_out[2610]);
    assign layer1_out[4861] = layer0_out[1651] & ~layer0_out[1650];
    assign layer1_out[4862] = layer0_out[7699] ^ layer0_out[7700];
    assign layer1_out[4863] = 1'b1;
    assign layer1_out[4864] = ~layer0_out[7415];
    assign layer1_out[4865] = layer0_out[1115];
    assign layer1_out[4866] = ~layer0_out[4280];
    assign layer1_out[4867] = ~(layer0_out[3638] ^ layer0_out[3639]);
    assign layer1_out[4868] = 1'b1;
    assign layer1_out[4869] = ~(layer0_out[5294] & layer0_out[5295]);
    assign layer1_out[4870] = ~layer0_out[6925] | layer0_out[6924];
    assign layer1_out[4871] = ~layer0_out[2465];
    assign layer1_out[4872] = ~layer0_out[7434];
    assign layer1_out[4873] = layer0_out[5932] | layer0_out[5933];
    assign layer1_out[4874] = layer0_out[367] & ~layer0_out[368];
    assign layer1_out[4875] = 1'b1;
    assign layer1_out[4876] = layer0_out[7401] & ~layer0_out[7402];
    assign layer1_out[4877] = ~layer0_out[6058] | layer0_out[6059];
    assign layer1_out[4878] = layer0_out[2391] & ~layer0_out[2390];
    assign layer1_out[4879] = layer0_out[5922] ^ layer0_out[5923];
    assign layer1_out[4880] = ~(layer0_out[2309] | layer0_out[2310]);
    assign layer1_out[4881] = ~(layer0_out[5209] & layer0_out[5210]);
    assign layer1_out[4882] = ~layer0_out[1076];
    assign layer1_out[4883] = layer0_out[731] ^ layer0_out[732];
    assign layer1_out[4884] = 1'b0;
    assign layer1_out[4885] = 1'b1;
    assign layer1_out[4886] = ~layer0_out[2596];
    assign layer1_out[4887] = layer0_out[2720] & ~layer0_out[2721];
    assign layer1_out[4888] = ~layer0_out[7266] | layer0_out[7265];
    assign layer1_out[4889] = layer0_out[3942];
    assign layer1_out[4890] = ~layer0_out[3215];
    assign layer1_out[4891] = layer0_out[5293];
    assign layer1_out[4892] = 1'b1;
    assign layer1_out[4893] = 1'b1;
    assign layer1_out[4894] = layer0_out[3059];
    assign layer1_out[4895] = layer0_out[6582];
    assign layer1_out[4896] = 1'b0;
    assign layer1_out[4897] = ~layer0_out[3026];
    assign layer1_out[4898] = layer0_out[4027];
    assign layer1_out[4899] = layer0_out[4911];
    assign layer1_out[4900] = 1'b0;
    assign layer1_out[4901] = layer0_out[1262] & layer0_out[1263];
    assign layer1_out[4902] = layer0_out[6282] & ~layer0_out[6281];
    assign layer1_out[4903] = ~(layer0_out[6937] | layer0_out[6938]);
    assign layer1_out[4904] = ~layer0_out[1147] | layer0_out[1148];
    assign layer1_out[4905] = ~layer0_out[4405];
    assign layer1_out[4906] = ~layer0_out[5913] | layer0_out[5912];
    assign layer1_out[4907] = layer0_out[3664] & layer0_out[3665];
    assign layer1_out[4908] = layer0_out[4057] | layer0_out[4058];
    assign layer1_out[4909] = ~layer0_out[944];
    assign layer1_out[4910] = layer0_out[6181] & ~layer0_out[6182];
    assign layer1_out[4911] = layer0_out[6787];
    assign layer1_out[4912] = ~layer0_out[588] | layer0_out[589];
    assign layer1_out[4913] = ~layer0_out[1332] | layer0_out[1331];
    assign layer1_out[4914] = ~(layer0_out[7667] ^ layer0_out[7668]);
    assign layer1_out[4915] = ~layer0_out[4152];
    assign layer1_out[4916] = ~(layer0_out[4013] | layer0_out[4014]);
    assign layer1_out[4917] = layer0_out[3423];
    assign layer1_out[4918] = 1'b1;
    assign layer1_out[4919] = layer0_out[3341];
    assign layer1_out[4920] = ~(layer0_out[6673] | layer0_out[6674]);
    assign layer1_out[4921] = ~layer0_out[7641];
    assign layer1_out[4922] = ~(layer0_out[3081] | layer0_out[3082]);
    assign layer1_out[4923] = layer0_out[4230] & ~layer0_out[4229];
    assign layer1_out[4924] = ~(layer0_out[7171] ^ layer0_out[7172]);
    assign layer1_out[4925] = layer0_out[2911];
    assign layer1_out[4926] = layer0_out[6686] & ~layer0_out[6685];
    assign layer1_out[4927] = ~(layer0_out[2434] & layer0_out[2435]);
    assign layer1_out[4928] = layer0_out[7182];
    assign layer1_out[4929] = ~layer0_out[5468];
    assign layer1_out[4930] = layer0_out[7358] & layer0_out[7359];
    assign layer1_out[4931] = ~(layer0_out[3122] & layer0_out[3123]);
    assign layer1_out[4932] = ~(layer0_out[7198] & layer0_out[7199]);
    assign layer1_out[4933] = layer0_out[2406];
    assign layer1_out[4934] = ~layer0_out[1857] | layer0_out[1858];
    assign layer1_out[4935] = ~layer0_out[1764] | layer0_out[1765];
    assign layer1_out[4936] = layer0_out[1983] ^ layer0_out[1984];
    assign layer1_out[4937] = ~layer0_out[3079] | layer0_out[3080];
    assign layer1_out[4938] = layer0_out[5490];
    assign layer1_out[4939] = ~layer0_out[7506] | layer0_out[7505];
    assign layer1_out[4940] = ~(layer0_out[7546] & layer0_out[7547]);
    assign layer1_out[4941] = layer0_out[6344] & ~layer0_out[6343];
    assign layer1_out[4942] = ~layer0_out[4748] | layer0_out[4747];
    assign layer1_out[4943] = ~(layer0_out[124] | layer0_out[125]);
    assign layer1_out[4944] = layer0_out[3682] & ~layer0_out[3681];
    assign layer1_out[4945] = layer0_out[3149] & layer0_out[3150];
    assign layer1_out[4946] = layer0_out[555];
    assign layer1_out[4947] = ~layer0_out[6081] | layer0_out[6082];
    assign layer1_out[4948] = ~(layer0_out[7184] & layer0_out[7185]);
    assign layer1_out[4949] = layer0_out[226] & ~layer0_out[225];
    assign layer1_out[4950] = 1'b0;
    assign layer1_out[4951] = ~(layer0_out[6068] & layer0_out[6069]);
    assign layer1_out[4952] = ~layer0_out[5608];
    assign layer1_out[4953] = ~layer0_out[5831];
    assign layer1_out[4954] = ~(layer0_out[921] & layer0_out[922]);
    assign layer1_out[4955] = layer0_out[384] & ~layer0_out[385];
    assign layer1_out[4956] = layer0_out[4305];
    assign layer1_out[4957] = ~layer0_out[4714];
    assign layer1_out[4958] = layer0_out[2800];
    assign layer1_out[4959] = 1'b0;
    assign layer1_out[4960] = layer0_out[2016] & ~layer0_out[2017];
    assign layer1_out[4961] = 1'b0;
    assign layer1_out[4962] = layer0_out[4419];
    assign layer1_out[4963] = layer0_out[1434] & layer0_out[1435];
    assign layer1_out[4964] = layer0_out[5766] & layer0_out[5767];
    assign layer1_out[4965] = layer0_out[647] & ~layer0_out[646];
    assign layer1_out[4966] = ~layer0_out[6183] | layer0_out[6182];
    assign layer1_out[4967] = layer0_out[2289] & ~layer0_out[2288];
    assign layer1_out[4968] = 1'b1;
    assign layer1_out[4969] = ~(layer0_out[5899] & layer0_out[5900]);
    assign layer1_out[4970] = ~layer0_out[6651] | layer0_out[6652];
    assign layer1_out[4971] = layer0_out[1295] ^ layer0_out[1296];
    assign layer1_out[4972] = 1'b0;
    assign layer1_out[4973] = ~(layer0_out[1185] & layer0_out[1186]);
    assign layer1_out[4974] = ~(layer0_out[5782] & layer0_out[5783]);
    assign layer1_out[4975] = ~layer0_out[2962] | layer0_out[2963];
    assign layer1_out[4976] = layer0_out[6894];
    assign layer1_out[4977] = ~layer0_out[1504] | layer0_out[1505];
    assign layer1_out[4978] = layer0_out[346];
    assign layer1_out[4979] = ~layer0_out[2844];
    assign layer1_out[4980] = ~layer0_out[3628];
    assign layer1_out[4981] = layer0_out[2818];
    assign layer1_out[4982] = ~layer0_out[6093] | layer0_out[6094];
    assign layer1_out[4983] = layer0_out[2330] | layer0_out[2331];
    assign layer1_out[4984] = ~(layer0_out[1895] ^ layer0_out[1896]);
    assign layer1_out[4985] = layer0_out[4588];
    assign layer1_out[4986] = layer0_out[4672] & ~layer0_out[4673];
    assign layer1_out[4987] = ~(layer0_out[1289] | layer0_out[1290]);
    assign layer1_out[4988] = layer0_out[2405] & layer0_out[2406];
    assign layer1_out[4989] = ~layer0_out[7194];
    assign layer1_out[4990] = ~(layer0_out[5595] & layer0_out[5596]);
    assign layer1_out[4991] = layer0_out[242] & ~layer0_out[241];
    assign layer1_out[4992] = ~(layer0_out[1674] & layer0_out[1675]);
    assign layer1_out[4993] = ~(layer0_out[5657] & layer0_out[5658]);
    assign layer1_out[4994] = ~layer0_out[2674];
    assign layer1_out[4995] = ~layer0_out[1768];
    assign layer1_out[4996] = layer0_out[2149] & ~layer0_out[2148];
    assign layer1_out[4997] = layer0_out[5020];
    assign layer1_out[4998] = ~layer0_out[5127] | layer0_out[5128];
    assign layer1_out[4999] = layer0_out[3200] & layer0_out[3201];
    assign layer1_out[5000] = ~(layer0_out[1794] | layer0_out[1795]);
    assign layer1_out[5001] = 1'b1;
    assign layer1_out[5002] = ~layer0_out[4913];
    assign layer1_out[5003] = ~layer0_out[7168] | layer0_out[7167];
    assign layer1_out[5004] = layer0_out[4211] & ~layer0_out[4210];
    assign layer1_out[5005] = layer0_out[6000];
    assign layer1_out[5006] = layer0_out[7593] & layer0_out[7594];
    assign layer1_out[5007] = 1'b1;
    assign layer1_out[5008] = layer0_out[6940] & ~layer0_out[6941];
    assign layer1_out[5009] = layer0_out[4018] & ~layer0_out[4017];
    assign layer1_out[5010] = layer0_out[1930] & layer0_out[1931];
    assign layer1_out[5011] = ~layer0_out[4271];
    assign layer1_out[5012] = ~(layer0_out[413] & layer0_out[414]);
    assign layer1_out[5013] = layer0_out[3467];
    assign layer1_out[5014] = layer0_out[7628] ^ layer0_out[7629];
    assign layer1_out[5015] = layer0_out[4277] & ~layer0_out[4278];
    assign layer1_out[5016] = ~(layer0_out[7127] ^ layer0_out[7128]);
    assign layer1_out[5017] = ~(layer0_out[1502] & layer0_out[1503]);
    assign layer1_out[5018] = ~(layer0_out[5320] & layer0_out[5321]);
    assign layer1_out[5019] = ~layer0_out[4475];
    assign layer1_out[5020] = 1'b1;
    assign layer1_out[5021] = ~layer0_out[553] | layer0_out[552];
    assign layer1_out[5022] = layer0_out[6152];
    assign layer1_out[5023] = ~layer0_out[3852];
    assign layer1_out[5024] = ~(layer0_out[4859] ^ layer0_out[4860]);
    assign layer1_out[5025] = ~layer0_out[5324];
    assign layer1_out[5026] = 1'b0;
    assign layer1_out[5027] = ~layer0_out[6721] | layer0_out[6720];
    assign layer1_out[5028] = layer0_out[883] & ~layer0_out[882];
    assign layer1_out[5029] = layer0_out[6254];
    assign layer1_out[5030] = layer0_out[7243] ^ layer0_out[7244];
    assign layer1_out[5031] = layer0_out[7692] & ~layer0_out[7691];
    assign layer1_out[5032] = layer0_out[463] & ~layer0_out[464];
    assign layer1_out[5033] = ~layer0_out[4074];
    assign layer1_out[5034] = ~layer0_out[1660];
    assign layer1_out[5035] = ~layer0_out[5335];
    assign layer1_out[5036] = 1'b1;
    assign layer1_out[5037] = 1'b0;
    assign layer1_out[5038] = layer0_out[3207] & layer0_out[3208];
    assign layer1_out[5039] = layer0_out[5742];
    assign layer1_out[5040] = layer0_out[3019] & layer0_out[3020];
    assign layer1_out[5041] = ~(layer0_out[6495] | layer0_out[6496]);
    assign layer1_out[5042] = ~(layer0_out[5538] | layer0_out[5539]);
    assign layer1_out[5043] = ~layer0_out[5975] | layer0_out[5976];
    assign layer1_out[5044] = layer0_out[1632];
    assign layer1_out[5045] = ~layer0_out[1736];
    assign layer1_out[5046] = ~(layer0_out[7836] ^ layer0_out[7837]);
    assign layer1_out[5047] = ~layer0_out[3841] | layer0_out[3842];
    assign layer1_out[5048] = ~(layer0_out[315] & layer0_out[316]);
    assign layer1_out[5049] = layer0_out[6635];
    assign layer1_out[5050] = ~(layer0_out[6624] ^ layer0_out[6625]);
    assign layer1_out[5051] = ~layer0_out[5946];
    assign layer1_out[5052] = ~layer0_out[4190];
    assign layer1_out[5053] = layer0_out[6210] & ~layer0_out[6209];
    assign layer1_out[5054] = layer0_out[26] | layer0_out[27];
    assign layer1_out[5055] = ~layer0_out[2278];
    assign layer1_out[5056] = layer0_out[2319] | layer0_out[2320];
    assign layer1_out[5057] = ~layer0_out[748];
    assign layer1_out[5058] = ~layer0_out[2901];
    assign layer1_out[5059] = layer0_out[6676];
    assign layer1_out[5060] = ~(layer0_out[2771] | layer0_out[2772]);
    assign layer1_out[5061] = ~(layer0_out[3329] & layer0_out[3330]);
    assign layer1_out[5062] = ~layer0_out[4315] | layer0_out[4316];
    assign layer1_out[5063] = layer0_out[4617] & layer0_out[4618];
    assign layer1_out[5064] = layer0_out[1937];
    assign layer1_out[5065] = ~layer0_out[4417] | layer0_out[4418];
    assign layer1_out[5066] = ~layer0_out[2358];
    assign layer1_out[5067] = layer0_out[6358] ^ layer0_out[6359];
    assign layer1_out[5068] = ~layer0_out[4475];
    assign layer1_out[5069] = ~layer0_out[4570];
    assign layer1_out[5070] = ~layer0_out[7884] | layer0_out[7883];
    assign layer1_out[5071] = layer0_out[6790] ^ layer0_out[6791];
    assign layer1_out[5072] = 1'b1;
    assign layer1_out[5073] = 1'b0;
    assign layer1_out[5074] = layer0_out[2506];
    assign layer1_out[5075] = ~layer0_out[5720] | layer0_out[5719];
    assign layer1_out[5076] = ~layer0_out[2116];
    assign layer1_out[5077] = ~(layer0_out[5075] & layer0_out[5076]);
    assign layer1_out[5078] = layer0_out[7274] & ~layer0_out[7275];
    assign layer1_out[5079] = layer0_out[7368] & ~layer0_out[7369];
    assign layer1_out[5080] = ~layer0_out[5828] | layer0_out[5827];
    assign layer1_out[5081] = ~layer0_out[2917];
    assign layer1_out[5082] = ~layer0_out[2284];
    assign layer1_out[5083] = layer0_out[1751] & ~layer0_out[1750];
    assign layer1_out[5084] = ~layer0_out[4022] | layer0_out[4023];
    assign layer1_out[5085] = layer0_out[1176] | layer0_out[1177];
    assign layer1_out[5086] = layer0_out[710] & layer0_out[711];
    assign layer1_out[5087] = ~(layer0_out[7656] ^ layer0_out[7657]);
    assign layer1_out[5088] = layer0_out[41];
    assign layer1_out[5089] = layer0_out[2421] & ~layer0_out[2422];
    assign layer1_out[5090] = ~(layer0_out[2151] | layer0_out[2152]);
    assign layer1_out[5091] = layer0_out[1824] & layer0_out[1825];
    assign layer1_out[5092] = layer0_out[3839];
    assign layer1_out[5093] = ~(layer0_out[1294] & layer0_out[1295]);
    assign layer1_out[5094] = ~layer0_out[5141];
    assign layer1_out[5095] = ~layer0_out[6323];
    assign layer1_out[5096] = layer0_out[5132];
    assign layer1_out[5097] = layer0_out[1709] & ~layer0_out[1710];
    assign layer1_out[5098] = layer0_out[1032] & ~layer0_out[1031];
    assign layer1_out[5099] = 1'b1;
    assign layer1_out[5100] = ~layer0_out[3013];
    assign layer1_out[5101] = 1'b1;
    assign layer1_out[5102] = ~layer0_out[6146];
    assign layer1_out[5103] = layer0_out[6797] & layer0_out[6798];
    assign layer1_out[5104] = ~layer0_out[2599];
    assign layer1_out[5105] = layer0_out[7483];
    assign layer1_out[5106] = layer0_out[6264] | layer0_out[6265];
    assign layer1_out[5107] = ~(layer0_out[4412] ^ layer0_out[4413]);
    assign layer1_out[5108] = 1'b1;
    assign layer1_out[5109] = ~layer0_out[1872];
    assign layer1_out[5110] = layer0_out[1020];
    assign layer1_out[5111] = layer0_out[5777] & layer0_out[5778];
    assign layer1_out[5112] = layer0_out[6482] | layer0_out[6483];
    assign layer1_out[5113] = 1'b0;
    assign layer1_out[5114] = ~(layer0_out[3290] & layer0_out[3291]);
    assign layer1_out[5115] = ~layer0_out[5966];
    assign layer1_out[5116] = 1'b1;
    assign layer1_out[5117] = layer0_out[4627] & ~layer0_out[4628];
    assign layer1_out[5118] = ~layer0_out[4754];
    assign layer1_out[5119] = layer0_out[369] ^ layer0_out[370];
    assign layer1_out[5120] = ~layer0_out[2835];
    assign layer1_out[5121] = layer0_out[1845];
    assign layer1_out[5122] = ~layer0_out[5076] | layer0_out[5077];
    assign layer1_out[5123] = layer0_out[3568] & ~layer0_out[3567];
    assign layer1_out[5124] = layer0_out[2290] | layer0_out[2291];
    assign layer1_out[5125] = ~layer0_out[2514] | layer0_out[2513];
    assign layer1_out[5126] = layer0_out[6731] & ~layer0_out[6730];
    assign layer1_out[5127] = layer0_out[770] & ~layer0_out[769];
    assign layer1_out[5128] = layer0_out[7823];
    assign layer1_out[5129] = layer0_out[16];
    assign layer1_out[5130] = layer0_out[4560] & layer0_out[4561];
    assign layer1_out[5131] = layer0_out[4820] | layer0_out[4821];
    assign layer1_out[5132] = ~layer0_out[3166];
    assign layer1_out[5133] = layer0_out[7022] | layer0_out[7023];
    assign layer1_out[5134] = layer0_out[3760] & layer0_out[3761];
    assign layer1_out[5135] = ~layer0_out[617];
    assign layer1_out[5136] = ~layer0_out[7949];
    assign layer1_out[5137] = ~layer0_out[6983];
    assign layer1_out[5138] = 1'b0;
    assign layer1_out[5139] = ~layer0_out[6346];
    assign layer1_out[5140] = ~layer0_out[3551] | layer0_out[3550];
    assign layer1_out[5141] = layer0_out[7530] & layer0_out[7531];
    assign layer1_out[5142] = layer0_out[6781] & ~layer0_out[6780];
    assign layer1_out[5143] = ~(layer0_out[1461] | layer0_out[1462]);
    assign layer1_out[5144] = layer0_out[4695] | layer0_out[4696];
    assign layer1_out[5145] = layer0_out[7782] & ~layer0_out[7783];
    assign layer1_out[5146] = layer0_out[7844] & ~layer0_out[7845];
    assign layer1_out[5147] = layer0_out[1823] | layer0_out[1824];
    assign layer1_out[5148] = ~(layer0_out[1941] | layer0_out[1942]);
    assign layer1_out[5149] = ~layer0_out[5941] | layer0_out[5940];
    assign layer1_out[5150] = ~layer0_out[6078];
    assign layer1_out[5151] = layer0_out[4608] & ~layer0_out[4607];
    assign layer1_out[5152] = 1'b0;
    assign layer1_out[5153] = ~(layer0_out[3675] | layer0_out[3676]);
    assign layer1_out[5154] = ~layer0_out[2409];
    assign layer1_out[5155] = layer0_out[1523] & layer0_out[1524];
    assign layer1_out[5156] = 1'b0;
    assign layer1_out[5157] = ~layer0_out[7735];
    assign layer1_out[5158] = layer0_out[5829] & ~layer0_out[5830];
    assign layer1_out[5159] = layer0_out[7670] & ~layer0_out[7669];
    assign layer1_out[5160] = ~(layer0_out[5289] & layer0_out[5290]);
    assign layer1_out[5161] = layer0_out[3800] & ~layer0_out[3799];
    assign layer1_out[5162] = ~layer0_out[799];
    assign layer1_out[5163] = layer0_out[2579];
    assign layer1_out[5164] = layer0_out[3819] & ~layer0_out[3818];
    assign layer1_out[5165] = layer0_out[7250] | layer0_out[7251];
    assign layer1_out[5166] = layer0_out[3643];
    assign layer1_out[5167] = ~layer0_out[884] | layer0_out[885];
    assign layer1_out[5168] = ~layer0_out[6075];
    assign layer1_out[5169] = ~layer0_out[1556];
    assign layer1_out[5170] = layer0_out[2172] & ~layer0_out[2171];
    assign layer1_out[5171] = 1'b0;
    assign layer1_out[5172] = layer0_out[989] & ~layer0_out[988];
    assign layer1_out[5173] = layer0_out[4023] & ~layer0_out[4024];
    assign layer1_out[5174] = layer0_out[1846] ^ layer0_out[1847];
    assign layer1_out[5175] = layer0_out[4065];
    assign layer1_out[5176] = layer0_out[3523] & ~layer0_out[3522];
    assign layer1_out[5177] = ~(layer0_out[5953] | layer0_out[5954]);
    assign layer1_out[5178] = layer0_out[7524] & layer0_out[7525];
    assign layer1_out[5179] = layer0_out[3757];
    assign layer1_out[5180] = layer0_out[2478] & layer0_out[2479];
    assign layer1_out[5181] = 1'b1;
    assign layer1_out[5182] = 1'b0;
    assign layer1_out[5183] = ~layer0_out[4953];
    assign layer1_out[5184] = ~(layer0_out[2957] | layer0_out[2958]);
    assign layer1_out[5185] = ~(layer0_out[5711] | layer0_out[5712]);
    assign layer1_out[5186] = ~layer0_out[5718];
    assign layer1_out[5187] = layer0_out[3302] ^ layer0_out[3303];
    assign layer1_out[5188] = layer0_out[2078] | layer0_out[2079];
    assign layer1_out[5189] = layer0_out[7751] & ~layer0_out[7750];
    assign layer1_out[5190] = ~layer0_out[4311];
    assign layer1_out[5191] = layer0_out[7195] ^ layer0_out[7196];
    assign layer1_out[5192] = layer0_out[6863] ^ layer0_out[6864];
    assign layer1_out[5193] = 1'b0;
    assign layer1_out[5194] = layer0_out[1813] & ~layer0_out[1814];
    assign layer1_out[5195] = layer0_out[4773] & ~layer0_out[4772];
    assign layer1_out[5196] = 1'b1;
    assign layer1_out[5197] = ~layer0_out[7646];
    assign layer1_out[5198] = layer0_out[2525];
    assign layer1_out[5199] = layer0_out[7630] & ~layer0_out[7631];
    assign layer1_out[5200] = layer0_out[4684] & ~layer0_out[4683];
    assign layer1_out[5201] = ~layer0_out[3068];
    assign layer1_out[5202] = layer0_out[1802] & layer0_out[1803];
    assign layer1_out[5203] = ~layer0_out[5949] | layer0_out[5950];
    assign layer1_out[5204] = ~layer0_out[7502];
    assign layer1_out[5205] = layer0_out[961] & ~layer0_out[960];
    assign layer1_out[5206] = ~(layer0_out[756] ^ layer0_out[757]);
    assign layer1_out[5207] = ~layer0_out[5309];
    assign layer1_out[5208] = layer0_out[2286] & layer0_out[2287];
    assign layer1_out[5209] = ~layer0_out[5613];
    assign layer1_out[5210] = layer0_out[932];
    assign layer1_out[5211] = ~layer0_out[767];
    assign layer1_out[5212] = ~layer0_out[4584];
    assign layer1_out[5213] = layer0_out[5] & ~layer0_out[4];
    assign layer1_out[5214] = ~(layer0_out[1743] & layer0_out[1744]);
    assign layer1_out[5215] = ~layer0_out[3170] | layer0_out[3169];
    assign layer1_out[5216] = layer0_out[762] & ~layer0_out[763];
    assign layer1_out[5217] = ~(layer0_out[7788] & layer0_out[7789]);
    assign layer1_out[5218] = layer0_out[7192];
    assign layer1_out[5219] = ~layer0_out[5228];
    assign layer1_out[5220] = layer0_out[3099] & ~layer0_out[3100];
    assign layer1_out[5221] = layer0_out[7313] & layer0_out[7314];
    assign layer1_out[5222] = ~layer0_out[4724];
    assign layer1_out[5223] = layer0_out[5908] & layer0_out[5909];
    assign layer1_out[5224] = layer0_out[5017] & ~layer0_out[5016];
    assign layer1_out[5225] = ~layer0_out[458];
    assign layer1_out[5226] = layer0_out[3483] & layer0_out[3484];
    assign layer1_out[5227] = 1'b1;
    assign layer1_out[5228] = ~layer0_out[2249] | layer0_out[2250];
    assign layer1_out[5229] = layer0_out[258] | layer0_out[259];
    assign layer1_out[5230] = ~layer0_out[2414];
    assign layer1_out[5231] = layer0_out[4177] & ~layer0_out[4178];
    assign layer1_out[5232] = layer0_out[6128] | layer0_out[6129];
    assign layer1_out[5233] = layer0_out[3636] | layer0_out[3637];
    assign layer1_out[5234] = ~layer0_out[4094] | layer0_out[4093];
    assign layer1_out[5235] = ~layer0_out[1872];
    assign layer1_out[5236] = ~layer0_out[2591];
    assign layer1_out[5237] = layer0_out[2081] & ~layer0_out[2080];
    assign layer1_out[5238] = layer0_out[5748] & ~layer0_out[5747];
    assign layer1_out[5239] = layer0_out[1758];
    assign layer1_out[5240] = ~layer0_out[6140] | layer0_out[6139];
    assign layer1_out[5241] = ~(layer0_out[2772] | layer0_out[2773]);
    assign layer1_out[5242] = ~layer0_out[6236];
    assign layer1_out[5243] = ~layer0_out[965] | layer0_out[966];
    assign layer1_out[5244] = layer0_out[294] | layer0_out[295];
    assign layer1_out[5245] = ~(layer0_out[1619] | layer0_out[1620]);
    assign layer1_out[5246] = layer0_out[306] & layer0_out[307];
    assign layer1_out[5247] = ~layer0_out[3146] | layer0_out[3147];
    assign layer1_out[5248] = layer0_out[2158];
    assign layer1_out[5249] = layer0_out[1738];
    assign layer1_out[5250] = ~layer0_out[5709] | layer0_out[5708];
    assign layer1_out[5251] = layer0_out[4838];
    assign layer1_out[5252] = layer0_out[6664] & ~layer0_out[6663];
    assign layer1_out[5253] = layer0_out[3717];
    assign layer1_out[5254] = layer0_out[3677] & layer0_out[3678];
    assign layer1_out[5255] = ~layer0_out[6674];
    assign layer1_out[5256] = ~layer0_out[850];
    assign layer1_out[5257] = layer0_out[2758] & ~layer0_out[2757];
    assign layer1_out[5258] = layer0_out[689] | layer0_out[690];
    assign layer1_out[5259] = ~layer0_out[6397];
    assign layer1_out[5260] = layer0_out[1630] | layer0_out[1631];
    assign layer1_out[5261] = layer0_out[3860] & ~layer0_out[3861];
    assign layer1_out[5262] = layer0_out[6180] ^ layer0_out[6181];
    assign layer1_out[5263] = ~layer0_out[7180];
    assign layer1_out[5264] = ~layer0_out[96] | layer0_out[95];
    assign layer1_out[5265] = ~layer0_out[6007] | layer0_out[6006];
    assign layer1_out[5266] = 1'b0;
    assign layer1_out[5267] = ~(layer0_out[1299] | layer0_out[1300]);
    assign layer1_out[5268] = ~(layer0_out[2425] & layer0_out[2426]);
    assign layer1_out[5269] = 1'b1;
    assign layer1_out[5270] = layer0_out[2209];
    assign layer1_out[5271] = ~(layer0_out[2013] | layer0_out[2014]);
    assign layer1_out[5272] = ~layer0_out[7298] | layer0_out[7299];
    assign layer1_out[5273] = layer0_out[3852] | layer0_out[3853];
    assign layer1_out[5274] = ~layer0_out[56];
    assign layer1_out[5275] = ~layer0_out[4843];
    assign layer1_out[5276] = ~(layer0_out[3560] & layer0_out[3561]);
    assign layer1_out[5277] = ~layer0_out[1262] | layer0_out[1261];
    assign layer1_out[5278] = ~(layer0_out[1944] & layer0_out[1945]);
    assign layer1_out[5279] = 1'b0;
    assign layer1_out[5280] = 1'b1;
    assign layer1_out[5281] = layer0_out[4058] & ~layer0_out[4059];
    assign layer1_out[5282] = layer0_out[4622];
    assign layer1_out[5283] = ~layer0_out[4785];
    assign layer1_out[5284] = layer0_out[1934];
    assign layer1_out[5285] = ~layer0_out[5092] | layer0_out[5093];
    assign layer1_out[5286] = ~layer0_out[48];
    assign layer1_out[5287] = ~(layer0_out[3938] | layer0_out[3939]);
    assign layer1_out[5288] = ~layer0_out[7019];
    assign layer1_out[5289] = ~layer0_out[6392];
    assign layer1_out[5290] = layer0_out[5605] & ~layer0_out[5604];
    assign layer1_out[5291] = ~layer0_out[7256];
    assign layer1_out[5292] = ~layer0_out[5708] | layer0_out[5707];
    assign layer1_out[5293] = ~layer0_out[4871];
    assign layer1_out[5294] = layer0_out[3442];
    assign layer1_out[5295] = ~layer0_out[713] | layer0_out[714];
    assign layer1_out[5296] = layer0_out[5027] & ~layer0_out[5026];
    assign layer1_out[5297] = layer0_out[7249] & layer0_out[7250];
    assign layer1_out[5298] = ~(layer0_out[7453] | layer0_out[7454]);
    assign layer1_out[5299] = layer0_out[7506] | layer0_out[7507];
    assign layer1_out[5300] = ~layer0_out[5575] | layer0_out[5576];
    assign layer1_out[5301] = layer0_out[5248] & ~layer0_out[5247];
    assign layer1_out[5302] = layer0_out[7789];
    assign layer1_out[5303] = ~layer0_out[926] | layer0_out[927];
    assign layer1_out[5304] = layer0_out[7950] & layer0_out[7951];
    assign layer1_out[5305] = ~(layer0_out[7083] & layer0_out[7084]);
    assign layer1_out[5306] = layer0_out[2460];
    assign layer1_out[5307] = 1'b0;
    assign layer1_out[5308] = layer0_out[4204];
    assign layer1_out[5309] = layer0_out[1569] & ~layer0_out[1570];
    assign layer1_out[5310] = ~layer0_out[6294] | layer0_out[6295];
    assign layer1_out[5311] = 1'b1;
    assign layer1_out[5312] = ~layer0_out[7260];
    assign layer1_out[5313] = ~(layer0_out[4007] ^ layer0_out[4008]);
    assign layer1_out[5314] = ~layer0_out[3605] | layer0_out[3606];
    assign layer1_out[5315] = ~(layer0_out[3030] | layer0_out[3031]);
    assign layer1_out[5316] = ~layer0_out[36] | layer0_out[37];
    assign layer1_out[5317] = layer0_out[5513];
    assign layer1_out[5318] = layer0_out[3006] & ~layer0_out[3005];
    assign layer1_out[5319] = layer0_out[2673] & ~layer0_out[2674];
    assign layer1_out[5320] = layer0_out[7025];
    assign layer1_out[5321] = layer0_out[3690] & layer0_out[3691];
    assign layer1_out[5322] = ~layer0_out[2921];
    assign layer1_out[5323] = layer0_out[7122];
    assign layer1_out[5324] = ~(layer0_out[4815] ^ layer0_out[4816]);
    assign layer1_out[5325] = layer0_out[7900] | layer0_out[7901];
    assign layer1_out[5326] = ~(layer0_out[1548] & layer0_out[1549]);
    assign layer1_out[5327] = ~(layer0_out[5537] | layer0_out[5538]);
    assign layer1_out[5328] = ~layer0_out[4010];
    assign layer1_out[5329] = ~(layer0_out[4451] & layer0_out[4452]);
    assign layer1_out[5330] = ~(layer0_out[7239] & layer0_out[7240]);
    assign layer1_out[5331] = layer0_out[6881] & layer0_out[6882];
    assign layer1_out[5332] = layer0_out[3769] & ~layer0_out[3768];
    assign layer1_out[5333] = ~(layer0_out[6888] | layer0_out[6889]);
    assign layer1_out[5334] = 1'b0;
    assign layer1_out[5335] = ~layer0_out[4346] | layer0_out[4345];
    assign layer1_out[5336] = layer0_out[7481];
    assign layer1_out[5337] = ~layer0_out[2368] | layer0_out[2367];
    assign layer1_out[5338] = layer0_out[6203];
    assign layer1_out[5339] = layer0_out[5476];
    assign layer1_out[5340] = ~(layer0_out[457] | layer0_out[458]);
    assign layer1_out[5341] = layer0_out[2935];
    assign layer1_out[5342] = layer0_out[6726] & layer0_out[6727];
    assign layer1_out[5343] = ~(layer0_out[5556] ^ layer0_out[5557]);
    assign layer1_out[5344] = ~layer0_out[4854];
    assign layer1_out[5345] = ~(layer0_out[3107] & layer0_out[3108]);
    assign layer1_out[5346] = layer0_out[1466] ^ layer0_out[1467];
    assign layer1_out[5347] = ~layer0_out[6858] | layer0_out[6857];
    assign layer1_out[5348] = ~(layer0_out[6597] | layer0_out[6598]);
    assign layer1_out[5349] = ~layer0_out[4025];
    assign layer1_out[5350] = ~layer0_out[7292] | layer0_out[7291];
    assign layer1_out[5351] = 1'b1;
    assign layer1_out[5352] = layer0_out[566] & ~layer0_out[567];
    assign layer1_out[5353] = ~layer0_out[6635];
    assign layer1_out[5354] = ~(layer0_out[5454] & layer0_out[5455]);
    assign layer1_out[5355] = layer0_out[1701] | layer0_out[1702];
    assign layer1_out[5356] = ~layer0_out[6451] | layer0_out[6452];
    assign layer1_out[5357] = layer0_out[839];
    assign layer1_out[5358] = layer0_out[2880];
    assign layer1_out[5359] = layer0_out[2977];
    assign layer1_out[5360] = ~(layer0_out[7168] & layer0_out[7169]);
    assign layer1_out[5361] = ~layer0_out[6107];
    assign layer1_out[5362] = layer0_out[1859];
    assign layer1_out[5363] = 1'b0;
    assign layer1_out[5364] = ~layer0_out[1948];
    assign layer1_out[5365] = layer0_out[6970];
    assign layer1_out[5366] = ~(layer0_out[2267] | layer0_out[2268]);
    assign layer1_out[5367] = ~layer0_out[968];
    assign layer1_out[5368] = layer0_out[7977] & ~layer0_out[7976];
    assign layer1_out[5369] = layer0_out[2783] & ~layer0_out[2782];
    assign layer1_out[5370] = layer0_out[4081] | layer0_out[4082];
    assign layer1_out[5371] = layer0_out[6690];
    assign layer1_out[5372] = layer0_out[1927] | layer0_out[1928];
    assign layer1_out[5373] = layer0_out[3968] | layer0_out[3969];
    assign layer1_out[5374] = layer0_out[1448];
    assign layer1_out[5375] = ~(layer0_out[4731] & layer0_out[4732]);
    assign layer1_out[5376] = layer0_out[7399] | layer0_out[7400];
    assign layer1_out[5377] = 1'b0;
    assign layer1_out[5378] = layer0_out[4209];
    assign layer1_out[5379] = ~(layer0_out[6251] ^ layer0_out[6252]);
    assign layer1_out[5380] = layer0_out[1123];
    assign layer1_out[5381] = ~(layer0_out[657] & layer0_out[658]);
    assign layer1_out[5382] = layer0_out[2018] & ~layer0_out[2019];
    assign layer1_out[5383] = ~layer0_out[4242];
    assign layer1_out[5384] = layer0_out[6326] & ~layer0_out[6325];
    assign layer1_out[5385] = layer0_out[3017];
    assign layer1_out[5386] = 1'b0;
    assign layer1_out[5387] = ~layer0_out[4435] | layer0_out[4434];
    assign layer1_out[5388] = ~layer0_out[1145] | layer0_out[1144];
    assign layer1_out[5389] = layer0_out[5639] & ~layer0_out[5640];
    assign layer1_out[5390] = layer0_out[4088];
    assign layer1_out[5391] = ~(layer0_out[310] ^ layer0_out[311]);
    assign layer1_out[5392] = ~(layer0_out[330] ^ layer0_out[331]);
    assign layer1_out[5393] = ~(layer0_out[4633] | layer0_out[4634]);
    assign layer1_out[5394] = layer0_out[4917] | layer0_out[4918];
    assign layer1_out[5395] = layer0_out[1903] & ~layer0_out[1902];
    assign layer1_out[5396] = layer0_out[6765];
    assign layer1_out[5397] = layer0_out[2390];
    assign layer1_out[5398] = layer0_out[4156];
    assign layer1_out[5399] = 1'b0;
    assign layer1_out[5400] = ~layer0_out[6391];
    assign layer1_out[5401] = ~(layer0_out[3170] | layer0_out[3171]);
    assign layer1_out[5402] = ~layer0_out[2084] | layer0_out[2085];
    assign layer1_out[5403] = layer0_out[626] | layer0_out[627];
    assign layer1_out[5404] = layer0_out[1357] ^ layer0_out[1358];
    assign layer1_out[5405] = 1'b0;
    assign layer1_out[5406] = layer0_out[7708];
    assign layer1_out[5407] = layer0_out[4375];
    assign layer1_out[5408] = ~(layer0_out[1406] | layer0_out[1407]);
    assign layer1_out[5409] = ~layer0_out[6474];
    assign layer1_out[5410] = ~layer0_out[5685] | layer0_out[5684];
    assign layer1_out[5411] = layer0_out[4706] & layer0_out[4707];
    assign layer1_out[5412] = 1'b0;
    assign layer1_out[5413] = layer0_out[4856] | layer0_out[4857];
    assign layer1_out[5414] = ~layer0_out[6271];
    assign layer1_out[5415] = ~layer0_out[2523];
    assign layer1_out[5416] = layer0_out[4382] & ~layer0_out[4383];
    assign layer1_out[5417] = ~(layer0_out[1832] ^ layer0_out[1833]);
    assign layer1_out[5418] = layer0_out[2048] & ~layer0_out[2047];
    assign layer1_out[5419] = ~(layer0_out[2401] & layer0_out[2402]);
    assign layer1_out[5420] = layer0_out[352];
    assign layer1_out[5421] = layer0_out[6419];
    assign layer1_out[5422] = ~layer0_out[6468];
    assign layer1_out[5423] = layer0_out[6667] ^ layer0_out[6668];
    assign layer1_out[5424] = layer0_out[3023] & layer0_out[3024];
    assign layer1_out[5425] = ~layer0_out[974] | layer0_out[975];
    assign layer1_out[5426] = layer0_out[4891];
    assign layer1_out[5427] = layer0_out[3774] | layer0_out[3775];
    assign layer1_out[5428] = layer0_out[3085] & layer0_out[3086];
    assign layer1_out[5429] = ~layer0_out[3029] | layer0_out[3028];
    assign layer1_out[5430] = 1'b0;
    assign layer1_out[5431] = ~layer0_out[7180];
    assign layer1_out[5432] = ~(layer0_out[1979] | layer0_out[1980]);
    assign layer1_out[5433] = ~layer0_out[7895];
    assign layer1_out[5434] = ~layer0_out[1168];
    assign layer1_out[5435] = 1'b0;
    assign layer1_out[5436] = 1'b0;
    assign layer1_out[5437] = ~layer0_out[6081];
    assign layer1_out[5438] = ~layer0_out[237];
    assign layer1_out[5439] = 1'b0;
    assign layer1_out[5440] = layer0_out[4868] & layer0_out[4869];
    assign layer1_out[5441] = ~layer0_out[5376] | layer0_out[5375];
    assign layer1_out[5442] = layer0_out[5656] | layer0_out[5657];
    assign layer1_out[5443] = layer0_out[570] ^ layer0_out[571];
    assign layer1_out[5444] = layer0_out[7974];
    assign layer1_out[5445] = layer0_out[610];
    assign layer1_out[5446] = ~(layer0_out[6783] ^ layer0_out[6784]);
    assign layer1_out[5447] = ~layer0_out[6587] | layer0_out[6586];
    assign layer1_out[5448] = ~(layer0_out[4851] | layer0_out[4852]);
    assign layer1_out[5449] = layer0_out[4220] & ~layer0_out[4221];
    assign layer1_out[5450] = ~layer0_out[6684] | layer0_out[6683];
    assign layer1_out[5451] = layer0_out[561];
    assign layer1_out[5452] = ~layer0_out[153];
    assign layer1_out[5453] = layer0_out[3158];
    assign layer1_out[5454] = ~(layer0_out[803] | layer0_out[804]);
    assign layer1_out[5455] = 1'b1;
    assign layer1_out[5456] = layer0_out[2691] & layer0_out[2692];
    assign layer1_out[5457] = layer0_out[534];
    assign layer1_out[5458] = layer0_out[657];
    assign layer1_out[5459] = layer0_out[5774] ^ layer0_out[5775];
    assign layer1_out[5460] = layer0_out[7861] & ~layer0_out[7862];
    assign layer1_out[5461] = ~layer0_out[2474];
    assign layer1_out[5462] = ~(layer0_out[5405] ^ layer0_out[5406]);
    assign layer1_out[5463] = layer0_out[4886] & ~layer0_out[4885];
    assign layer1_out[5464] = layer0_out[7999] & ~layer0_out[7998];
    assign layer1_out[5465] = ~(layer0_out[4566] ^ layer0_out[4567]);
    assign layer1_out[5466] = ~layer0_out[3361];
    assign layer1_out[5467] = layer0_out[2496];
    assign layer1_out[5468] = layer0_out[6557] & layer0_out[6558];
    assign layer1_out[5469] = layer0_out[4172] | layer0_out[4173];
    assign layer1_out[5470] = layer0_out[1349] | layer0_out[1350];
    assign layer1_out[5471] = ~layer0_out[3971];
    assign layer1_out[5472] = layer0_out[233] & ~layer0_out[234];
    assign layer1_out[5473] = layer0_out[3224] & ~layer0_out[3225];
    assign layer1_out[5474] = ~layer0_out[7755];
    assign layer1_out[5475] = ~layer0_out[359];
    assign layer1_out[5476] = layer0_out[7851];
    assign layer1_out[5477] = ~layer0_out[7361] | layer0_out[7360];
    assign layer1_out[5478] = ~(layer0_out[5886] | layer0_out[5887]);
    assign layer1_out[5479] = ~layer0_out[7110];
    assign layer1_out[5480] = layer0_out[4736] | layer0_out[4737];
    assign layer1_out[5481] = ~(layer0_out[3401] | layer0_out[3402]);
    assign layer1_out[5482] = layer0_out[4515];
    assign layer1_out[5483] = ~layer0_out[319];
    assign layer1_out[5484] = ~layer0_out[930] | layer0_out[931];
    assign layer1_out[5485] = layer0_out[5686] & layer0_out[5687];
    assign layer1_out[5486] = layer0_out[4233];
    assign layer1_out[5487] = ~layer0_out[1647] | layer0_out[1646];
    assign layer1_out[5488] = ~layer0_out[1583] | layer0_out[1584];
    assign layer1_out[5489] = layer0_out[1320];
    assign layer1_out[5490] = layer0_out[7424] & ~layer0_out[7423];
    assign layer1_out[5491] = ~layer0_out[6917] | layer0_out[6918];
    assign layer1_out[5492] = ~layer0_out[5477] | layer0_out[5478];
    assign layer1_out[5493] = 1'b1;
    assign layer1_out[5494] = layer0_out[6240];
    assign layer1_out[5495] = layer0_out[6640] | layer0_out[6641];
    assign layer1_out[5496] = ~(layer0_out[4014] | layer0_out[4015]);
    assign layer1_out[5497] = ~layer0_out[2741] | layer0_out[2742];
    assign layer1_out[5498] = layer0_out[7804] ^ layer0_out[7805];
    assign layer1_out[5499] = ~(layer0_out[7960] | layer0_out[7961]);
    assign layer1_out[5500] = ~layer0_out[3988] | layer0_out[3989];
    assign layer1_out[5501] = ~layer0_out[3323] | layer0_out[3324];
    assign layer1_out[5502] = layer0_out[741] | layer0_out[742];
    assign layer1_out[5503] = 1'b0;
    assign layer1_out[5504] = layer0_out[3431];
    assign layer1_out[5505] = layer0_out[1867] | layer0_out[1868];
    assign layer1_out[5506] = layer0_out[2941];
    assign layer1_out[5507] = layer0_out[1968] & ~layer0_out[1969];
    assign layer1_out[5508] = ~layer0_out[6411];
    assign layer1_out[5509] = ~layer0_out[3305];
    assign layer1_out[5510] = 1'b1;
    assign layer1_out[5511] = ~(layer0_out[1356] & layer0_out[1357]);
    assign layer1_out[5512] = ~(layer0_out[5942] & layer0_out[5943]);
    assign layer1_out[5513] = layer0_out[5871];
    assign layer1_out[5514] = 1'b1;
    assign layer1_out[5515] = ~layer0_out[4889] | layer0_out[4888];
    assign layer1_out[5516] = ~layer0_out[1161] | layer0_out[1160];
    assign layer1_out[5517] = layer0_out[6388] ^ layer0_out[6389];
    assign layer1_out[5518] = ~layer0_out[1193] | layer0_out[1192];
    assign layer1_out[5519] = ~(layer0_out[2164] & layer0_out[2165]);
    assign layer1_out[5520] = 1'b1;
    assign layer1_out[5521] = layer0_out[1181];
    assign layer1_out[5522] = ~(layer0_out[1916] ^ layer0_out[1917]);
    assign layer1_out[5523] = layer0_out[3623] | layer0_out[3624];
    assign layer1_out[5524] = ~(layer0_out[1405] & layer0_out[1406]);
    assign layer1_out[5525] = 1'b1;
    assign layer1_out[5526] = 1'b0;
    assign layer1_out[5527] = ~(layer0_out[5510] & layer0_out[5511]);
    assign layer1_out[5528] = ~(layer0_out[929] ^ layer0_out[930]);
    assign layer1_out[5529] = layer0_out[6936] & ~layer0_out[6937];
    assign layer1_out[5530] = layer0_out[4684] & ~layer0_out[4685];
    assign layer1_out[5531] = ~layer0_out[4878];
    assign layer1_out[5532] = 1'b1;
    assign layer1_out[5533] = ~(layer0_out[4778] | layer0_out[4779]);
    assign layer1_out[5534] = ~(layer0_out[1621] | layer0_out[1622]);
    assign layer1_out[5535] = layer0_out[5454];
    assign layer1_out[5536] = layer0_out[1893] & layer0_out[1894];
    assign layer1_out[5537] = ~layer0_out[3268] | layer0_out[3269];
    assign layer1_out[5538] = layer0_out[7947] & ~layer0_out[7946];
    assign layer1_out[5539] = layer0_out[3299] | layer0_out[3300];
    assign layer1_out[5540] = ~(layer0_out[6402] & layer0_out[6403]);
    assign layer1_out[5541] = ~layer0_out[474];
    assign layer1_out[5542] = layer0_out[6830] & ~layer0_out[6831];
    assign layer1_out[5543] = ~layer0_out[3535] | layer0_out[3536];
    assign layer1_out[5544] = ~layer0_out[7038] | layer0_out[7037];
    assign layer1_out[5545] = layer0_out[3284] & layer0_out[3285];
    assign layer1_out[5546] = ~(layer0_out[6716] & layer0_out[6717]);
    assign layer1_out[5547] = ~layer0_out[5788];
    assign layer1_out[5548] = layer0_out[2971];
    assign layer1_out[5549] = ~(layer0_out[222] & layer0_out[223]);
    assign layer1_out[5550] = layer0_out[6364] & layer0_out[6365];
    assign layer1_out[5551] = layer0_out[5734];
    assign layer1_out[5552] = layer0_out[5949] & ~layer0_out[5948];
    assign layer1_out[5553] = layer0_out[2247];
    assign layer1_out[5554] = ~layer0_out[3584];
    assign layer1_out[5555] = 1'b0;
    assign layer1_out[5556] = 1'b1;
    assign layer1_out[5557] = layer0_out[3569];
    assign layer1_out[5558] = ~(layer0_out[5369] | layer0_out[5370]);
    assign layer1_out[5559] = layer0_out[5915] | layer0_out[5916];
    assign layer1_out[5560] = ~layer0_out[1748];
    assign layer1_out[5561] = ~layer0_out[4945];
    assign layer1_out[5562] = ~layer0_out[1465] | layer0_out[1466];
    assign layer1_out[5563] = ~layer0_out[1314] | layer0_out[1313];
    assign layer1_out[5564] = ~layer0_out[520] | layer0_out[521];
    assign layer1_out[5565] = ~layer0_out[2861] | layer0_out[2860];
    assign layer1_out[5566] = ~layer0_out[1561] | layer0_out[1560];
    assign layer1_out[5567] = ~layer0_out[3986] | layer0_out[3987];
    assign layer1_out[5568] = ~layer0_out[3159];
    assign layer1_out[5569] = layer0_out[4185];
    assign layer1_out[5570] = layer0_out[6773];
    assign layer1_out[5571] = ~layer0_out[579] | layer0_out[578];
    assign layer1_out[5572] = layer0_out[7855] & ~layer0_out[7854];
    assign layer1_out[5573] = layer0_out[4970] & ~layer0_out[4971];
    assign layer1_out[5574] = ~(layer0_out[6882] & layer0_out[6883]);
    assign layer1_out[5575] = layer0_out[7354] & ~layer0_out[7353];
    assign layer1_out[5576] = layer0_out[4322] & ~layer0_out[4321];
    assign layer1_out[5577] = layer0_out[7635] & ~layer0_out[7636];
    assign layer1_out[5578] = layer0_out[3096];
    assign layer1_out[5579] = ~layer0_out[7513];
    assign layer1_out[5580] = ~layer0_out[3119];
    assign layer1_out[5581] = ~layer0_out[3775];
    assign layer1_out[5582] = layer0_out[6400] & ~layer0_out[6399];
    assign layer1_out[5583] = layer0_out[5946];
    assign layer1_out[5584] = ~(layer0_out[4309] | layer0_out[4310]);
    assign layer1_out[5585] = ~layer0_out[2473] | layer0_out[2472];
    assign layer1_out[5586] = 1'b1;
    assign layer1_out[5587] = 1'b1;
    assign layer1_out[5588] = layer0_out[3712] | layer0_out[3713];
    assign layer1_out[5589] = ~(layer0_out[4642] | layer0_out[4643]);
    assign layer1_out[5590] = ~layer0_out[2549] | layer0_out[2548];
    assign layer1_out[5591] = layer0_out[4288] ^ layer0_out[4289];
    assign layer1_out[5592] = layer0_out[5070] & ~layer0_out[5071];
    assign layer1_out[5593] = ~layer0_out[2922];
    assign layer1_out[5594] = ~(layer0_out[3315] & layer0_out[3316]);
    assign layer1_out[5595] = layer0_out[705] | layer0_out[706];
    assign layer1_out[5596] = layer0_out[928] & layer0_out[929];
    assign layer1_out[5597] = layer0_out[5715] | layer0_out[5716];
    assign layer1_out[5598] = ~(layer0_out[6421] | layer0_out[6422]);
    assign layer1_out[5599] = ~(layer0_out[6160] & layer0_out[6161]);
    assign layer1_out[5600] = ~layer0_out[278] | layer0_out[279];
    assign layer1_out[5601] = ~(layer0_out[6502] ^ layer0_out[6503]);
    assign layer1_out[5602] = layer0_out[2444];
    assign layer1_out[5603] = ~layer0_out[3823] | layer0_out[3824];
    assign layer1_out[5604] = ~layer0_out[6662];
    assign layer1_out[5605] = ~layer0_out[6871];
    assign layer1_out[5606] = ~(layer0_out[342] | layer0_out[343]);
    assign layer1_out[5607] = ~layer0_out[4667] | layer0_out[4668];
    assign layer1_out[5608] = layer0_out[3319];
    assign layer1_out[5609] = layer0_out[3488] & ~layer0_out[3489];
    assign layer1_out[5610] = ~layer0_out[2002];
    assign layer1_out[5611] = ~layer0_out[5029] | layer0_out[5028];
    assign layer1_out[5612] = layer0_out[4780] ^ layer0_out[4781];
    assign layer1_out[5613] = layer0_out[4035] & ~layer0_out[4034];
    assign layer1_out[5614] = layer0_out[3203] & ~layer0_out[3204];
    assign layer1_out[5615] = layer0_out[2251];
    assign layer1_out[5616] = ~layer0_out[1629];
    assign layer1_out[5617] = ~layer0_out[1065] | layer0_out[1066];
    assign layer1_out[5618] = ~layer0_out[5406] | layer0_out[5407];
    assign layer1_out[5619] = ~layer0_out[272];
    assign layer1_out[5620] = layer0_out[3052];
    assign layer1_out[5621] = ~(layer0_out[4121] & layer0_out[4122]);
    assign layer1_out[5622] = ~layer0_out[2085] | layer0_out[2086];
    assign layer1_out[5623] = layer0_out[932] & ~layer0_out[933];
    assign layer1_out[5624] = ~layer0_out[4794];
    assign layer1_out[5625] = layer0_out[664] & ~layer0_out[663];
    assign layer1_out[5626] = ~(layer0_out[4436] & layer0_out[4437]);
    assign layer1_out[5627] = ~(layer0_out[3581] ^ layer0_out[3582]);
    assign layer1_out[5628] = layer0_out[7847] & ~layer0_out[7848];
    assign layer1_out[5629] = layer0_out[6973] | layer0_out[6974];
    assign layer1_out[5630] = layer0_out[7792] & ~layer0_out[7793];
    assign layer1_out[5631] = ~layer0_out[6259] | layer0_out[6260];
    assign layer1_out[5632] = 1'b0;
    assign layer1_out[5633] = ~layer0_out[7395] | layer0_out[7396];
    assign layer1_out[5634] = layer0_out[7137] ^ layer0_out[7138];
    assign layer1_out[5635] = layer0_out[521] & ~layer0_out[522];
    assign layer1_out[5636] = layer0_out[6168];
    assign layer1_out[5637] = layer0_out[3117];
    assign layer1_out[5638] = ~layer0_out[5214] | layer0_out[5215];
    assign layer1_out[5639] = ~layer0_out[5698];
    assign layer1_out[5640] = layer0_out[4711] & layer0_out[4712];
    assign layer1_out[5641] = 1'b0;
    assign layer1_out[5642] = 1'b0;
    assign layer1_out[5643] = 1'b0;
    assign layer1_out[5644] = layer0_out[1014];
    assign layer1_out[5645] = layer0_out[4132];
    assign layer1_out[5646] = 1'b1;
    assign layer1_out[5647] = layer0_out[1725] | layer0_out[1726];
    assign layer1_out[5648] = ~layer0_out[5497];
    assign layer1_out[5649] = ~(layer0_out[4487] ^ layer0_out[4488]);
    assign layer1_out[5650] = ~layer0_out[3655];
    assign layer1_out[5651] = ~layer0_out[1980] | layer0_out[1981];
    assign layer1_out[5652] = layer0_out[2867];
    assign layer1_out[5653] = layer0_out[1888] | layer0_out[1889];
    assign layer1_out[5654] = ~layer0_out[6481];
    assign layer1_out[5655] = ~layer0_out[576];
    assign layer1_out[5656] = layer0_out[7822] & layer0_out[7823];
    assign layer1_out[5657] = ~(layer0_out[5852] ^ layer0_out[5853]);
    assign layer1_out[5658] = layer0_out[5139] | layer0_out[5140];
    assign layer1_out[5659] = ~layer0_out[7178] | layer0_out[7179];
    assign layer1_out[5660] = ~(layer0_out[5461] & layer0_out[5462]);
    assign layer1_out[5661] = ~(layer0_out[1124] & layer0_out[1125]);
    assign layer1_out[5662] = ~layer0_out[2426];
    assign layer1_out[5663] = ~layer0_out[2102];
    assign layer1_out[5664] = ~layer0_out[2544] | layer0_out[2543];
    assign layer1_out[5665] = layer0_out[1815] ^ layer0_out[1816];
    assign layer1_out[5666] = ~layer0_out[7573];
    assign layer1_out[5667] = ~(layer0_out[2252] & layer0_out[2253]);
    assign layer1_out[5668] = layer0_out[5471] & layer0_out[5472];
    assign layer1_out[5669] = ~layer0_out[299] | layer0_out[300];
    assign layer1_out[5670] = 1'b0;
    assign layer1_out[5671] = layer0_out[6851] & ~layer0_out[6850];
    assign layer1_out[5672] = ~layer0_out[316];
    assign layer1_out[5673] = layer0_out[7114] & ~layer0_out[7115];
    assign layer1_out[5674] = ~layer0_out[6167];
    assign layer1_out[5675] = layer0_out[1344] & ~layer0_out[1343];
    assign layer1_out[5676] = layer0_out[5004] ^ layer0_out[5005];
    assign layer1_out[5677] = layer0_out[3459] | layer0_out[3460];
    assign layer1_out[5678] = layer0_out[2261] & ~layer0_out[2262];
    assign layer1_out[5679] = layer0_out[2644] & ~layer0_out[2643];
    assign layer1_out[5680] = layer0_out[565];
    assign layer1_out[5681] = ~(layer0_out[5242] & layer0_out[5243]);
    assign layer1_out[5682] = 1'b0;
    assign layer1_out[5683] = ~layer0_out[2750] | layer0_out[2751];
    assign layer1_out[5684] = ~layer0_out[44];
    assign layer1_out[5685] = layer0_out[7329] | layer0_out[7330];
    assign layer1_out[5686] = layer0_out[5080] & ~layer0_out[5081];
    assign layer1_out[5687] = ~(layer0_out[7775] | layer0_out[7776]);
    assign layer1_out[5688] = layer0_out[3340] & ~layer0_out[3341];
    assign layer1_out[5689] = ~(layer0_out[1531] & layer0_out[1532]);
    assign layer1_out[5690] = layer0_out[862] & ~layer0_out[863];
    assign layer1_out[5691] = layer0_out[3288] & ~layer0_out[3289];
    assign layer1_out[5692] = layer0_out[3585] & ~layer0_out[3586];
    assign layer1_out[5693] = layer0_out[7331];
    assign layer1_out[5694] = layer0_out[2477] | layer0_out[2478];
    assign layer1_out[5695] = ~layer0_out[3098] | layer0_out[3099];
    assign layer1_out[5696] = ~layer0_out[5056];
    assign layer1_out[5697] = ~layer0_out[5681] | layer0_out[5682];
    assign layer1_out[5698] = layer0_out[6450] & ~layer0_out[6449];
    assign layer1_out[5699] = ~(layer0_out[5879] ^ layer0_out[5880]);
    assign layer1_out[5700] = ~(layer0_out[7478] | layer0_out[7479]);
    assign layer1_out[5701] = layer0_out[1572] | layer0_out[1573];
    assign layer1_out[5702] = layer0_out[536] | layer0_out[537];
    assign layer1_out[5703] = layer0_out[3277] ^ layer0_out[3278];
    assign layer1_out[5704] = ~layer0_out[4767];
    assign layer1_out[5705] = ~layer0_out[5665];
    assign layer1_out[5706] = ~layer0_out[7064] | layer0_out[7063];
    assign layer1_out[5707] = layer0_out[844] & layer0_out[845];
    assign layer1_out[5708] = layer0_out[3871];
    assign layer1_out[5709] = layer0_out[2470];
    assign layer1_out[5710] = ~layer0_out[4164];
    assign layer1_out[5711] = layer0_out[6200];
    assign layer1_out[5712] = ~layer0_out[3511];
    assign layer1_out[5713] = ~(layer0_out[5485] & layer0_out[5486]);
    assign layer1_out[5714] = layer0_out[4941] & layer0_out[4942];
    assign layer1_out[5715] = layer0_out[6197];
    assign layer1_out[5716] = ~layer0_out[2792];
    assign layer1_out[5717] = layer0_out[2542] & ~layer0_out[2541];
    assign layer1_out[5718] = ~layer0_out[4527] | layer0_out[4528];
    assign layer1_out[5719] = layer0_out[7325] & ~layer0_out[7324];
    assign layer1_out[5720] = layer0_out[2436];
    assign layer1_out[5721] = layer0_out[4661];
    assign layer1_out[5722] = ~(layer0_out[7246] & layer0_out[7247]);
    assign layer1_out[5723] = ~layer0_out[1175];
    assign layer1_out[5724] = 1'b1;
    assign layer1_out[5725] = layer0_out[7129] | layer0_out[7130];
    assign layer1_out[5726] = layer0_out[4292] & ~layer0_out[4291];
    assign layer1_out[5727] = ~layer0_out[3783] | layer0_out[3782];
    assign layer1_out[5728] = ~layer0_out[5451];
    assign layer1_out[5729] = layer0_out[5369];
    assign layer1_out[5730] = layer0_out[3454] ^ layer0_out[3455];
    assign layer1_out[5731] = layer0_out[1599] | layer0_out[1600];
    assign layer1_out[5732] = layer0_out[6931];
    assign layer1_out[5733] = layer0_out[5100] & ~layer0_out[5101];
    assign layer1_out[5734] = layer0_out[3462] & ~layer0_out[3463];
    assign layer1_out[5735] = ~layer0_out[3233];
    assign layer1_out[5736] = layer0_out[4552];
    assign layer1_out[5737] = layer0_out[7795];
    assign layer1_out[5738] = layer0_out[1103] | layer0_out[1104];
    assign layer1_out[5739] = layer0_out[2999] & ~layer0_out[2998];
    assign layer1_out[5740] = ~layer0_out[1039];
    assign layer1_out[5741] = layer0_out[3991] & ~layer0_out[3992];
    assign layer1_out[5742] = layer0_out[5628];
    assign layer1_out[5743] = layer0_out[3367];
    assign layer1_out[5744] = layer0_out[1044];
    assign layer1_out[5745] = layer0_out[1828];
    assign layer1_out[5746] = layer0_out[6932] & ~layer0_out[6933];
    assign layer1_out[5747] = layer0_out[6693] & ~layer0_out[6692];
    assign layer1_out[5748] = layer0_out[4107];
    assign layer1_out[5749] = 1'b1;
    assign layer1_out[5750] = layer0_out[7085] ^ layer0_out[7086];
    assign layer1_out[5751] = ~layer0_out[211];
    assign layer1_out[5752] = 1'b1;
    assign layer1_out[5753] = layer0_out[5523];
    assign layer1_out[5754] = layer0_out[2427] & layer0_out[2428];
    assign layer1_out[5755] = layer0_out[7199];
    assign layer1_out[5756] = 1'b0;
    assign layer1_out[5757] = ~layer0_out[5484];
    assign layer1_out[5758] = ~layer0_out[1094];
    assign layer1_out[5759] = ~layer0_out[477] | layer0_out[476];
    assign layer1_out[5760] = layer0_out[4520] | layer0_out[4521];
    assign layer1_out[5761] = layer0_out[7372];
    assign layer1_out[5762] = layer0_out[5916];
    assign layer1_out[5763] = ~(layer0_out[7961] ^ layer0_out[7962]);
    assign layer1_out[5764] = ~layer0_out[7241];
    assign layer1_out[5765] = layer0_out[6688] & layer0_out[6689];
    assign layer1_out[5766] = layer0_out[3658] ^ layer0_out[3659];
    assign layer1_out[5767] = ~layer0_out[7782];
    assign layer1_out[5768] = ~layer0_out[1395];
    assign layer1_out[5769] = layer0_out[1214];
    assign layer1_out[5770] = layer0_out[5724] & ~layer0_out[5723];
    assign layer1_out[5771] = ~layer0_out[3563];
    assign layer1_out[5772] = layer0_out[1433] & ~layer0_out[1432];
    assign layer1_out[5773] = ~layer0_out[6608] | layer0_out[6607];
    assign layer1_out[5774] = layer0_out[4168] & ~layer0_out[4169];
    assign layer1_out[5775] = layer0_out[7680] & layer0_out[7681];
    assign layer1_out[5776] = layer0_out[5033] | layer0_out[5034];
    assign layer1_out[5777] = ~layer0_out[5046] | layer0_out[5047];
    assign layer1_out[5778] = layer0_out[5909] | layer0_out[5910];
    assign layer1_out[5779] = ~layer0_out[3589] | layer0_out[3590];
    assign layer1_out[5780] = ~(layer0_out[5837] | layer0_out[5838]);
    assign layer1_out[5781] = layer0_out[2837] & ~layer0_out[2838];
    assign layer1_out[5782] = layer0_out[3103] & ~layer0_out[3104];
    assign layer1_out[5783] = ~(layer0_out[7271] | layer0_out[7272]);
    assign layer1_out[5784] = layer0_out[7052] & layer0_out[7053];
    assign layer1_out[5785] = ~layer0_out[3893] | layer0_out[3892];
    assign layer1_out[5786] = layer0_out[4946] & ~layer0_out[4947];
    assign layer1_out[5787] = ~(layer0_out[1542] | layer0_out[1543]);
    assign layer1_out[5788] = ~layer0_out[399] | layer0_out[398];
    assign layer1_out[5789] = layer0_out[4705] & ~layer0_out[4706];
    assign layer1_out[5790] = ~layer0_out[4919] | layer0_out[4920];
    assign layer1_out[5791] = ~(layer0_out[1479] & layer0_out[1480]);
    assign layer1_out[5792] = layer0_out[4858] & ~layer0_out[4859];
    assign layer1_out[5793] = ~layer0_out[1718];
    assign layer1_out[5794] = layer0_out[7065] ^ layer0_out[7066];
    assign layer1_out[5795] = ~layer0_out[39] | layer0_out[40];
    assign layer1_out[5796] = ~(layer0_out[3456] | layer0_out[3457]);
    assign layer1_out[5797] = ~layer0_out[3745] | layer0_out[3744];
    assign layer1_out[5798] = 1'b1;
    assign layer1_out[5799] = ~layer0_out[3404] | layer0_out[3405];
    assign layer1_out[5800] = 1'b1;
    assign layer1_out[5801] = layer0_out[2997] | layer0_out[2998];
    assign layer1_out[5802] = ~layer0_out[680];
    assign layer1_out[5803] = ~(layer0_out[1338] & layer0_out[1339]);
    assign layer1_out[5804] = layer0_out[6957];
    assign layer1_out[5805] = ~layer0_out[3208] | layer0_out[3209];
    assign layer1_out[5806] = layer0_out[6288];
    assign layer1_out[5807] = layer0_out[4436];
    assign layer1_out[5808] = 1'b1;
    assign layer1_out[5809] = ~layer0_out[3176] | layer0_out[3175];
    assign layer1_out[5810] = ~layer0_out[1925] | layer0_out[1926];
    assign layer1_out[5811] = layer0_out[5374] ^ layer0_out[5375];
    assign layer1_out[5812] = ~(layer0_out[3027] ^ layer0_out[3028]);
    assign layer1_out[5813] = 1'b0;
    assign layer1_out[5814] = ~(layer0_out[6366] & layer0_out[6367]);
    assign layer1_out[5815] = ~layer0_out[2433];
    assign layer1_out[5816] = layer0_out[1003] | layer0_out[1004];
    assign layer1_out[5817] = ~layer0_out[7777];
    assign layer1_out[5818] = ~layer0_out[2828];
    assign layer1_out[5819] = ~(layer0_out[7045] & layer0_out[7046]);
    assign layer1_out[5820] = ~layer0_out[187];
    assign layer1_out[5821] = ~(layer0_out[5745] ^ layer0_out[5746]);
    assign layer1_out[5822] = layer0_out[3988] & ~layer0_out[3987];
    assign layer1_out[5823] = ~(layer0_out[2298] & layer0_out[2299]);
    assign layer1_out[5824] = layer0_out[1148] | layer0_out[1149];
    assign layer1_out[5825] = layer0_out[7097] & layer0_out[7098];
    assign layer1_out[5826] = ~layer0_out[3396];
    assign layer1_out[5827] = layer0_out[6834];
    assign layer1_out[5828] = ~(layer0_out[6304] & layer0_out[6305]);
    assign layer1_out[5829] = layer0_out[2580] | layer0_out[2581];
    assign layer1_out[5830] = ~layer0_out[7430];
    assign layer1_out[5831] = 1'b0;
    assign layer1_out[5832] = layer0_out[6053];
    assign layer1_out[5833] = ~(layer0_out[5468] ^ layer0_out[5469]);
    assign layer1_out[5834] = ~layer0_out[5204] | layer0_out[5205];
    assign layer1_out[5835] = ~(layer0_out[5875] | layer0_out[5876]);
    assign layer1_out[5836] = ~layer0_out[4577];
    assign layer1_out[5837] = ~layer0_out[6454] | layer0_out[6453];
    assign layer1_out[5838] = layer0_out[1459] & layer0_out[1460];
    assign layer1_out[5839] = 1'b0;
    assign layer1_out[5840] = layer0_out[2709];
    assign layer1_out[5841] = layer0_out[3528];
    assign layer1_out[5842] = ~layer0_out[2668];
    assign layer1_out[5843] = ~layer0_out[6630];
    assign layer1_out[5844] = layer0_out[6901];
    assign layer1_out[5845] = layer0_out[6389] | layer0_out[6390];
    assign layer1_out[5846] = ~layer0_out[5937] | layer0_out[5936];
    assign layer1_out[5847] = layer0_out[2483];
    assign layer1_out[5848] = ~(layer0_out[5779] ^ layer0_out[5780]);
    assign layer1_out[5849] = layer0_out[6195] & ~layer0_out[6194];
    assign layer1_out[5850] = ~layer0_out[6353] | layer0_out[6354];
    assign layer1_out[5851] = layer0_out[6270];
    assign layer1_out[5852] = 1'b1;
    assign layer1_out[5853] = layer0_out[470] & ~layer0_out[471];
    assign layer1_out[5854] = layer0_out[850] | layer0_out[851];
    assign layer1_out[5855] = layer0_out[1098];
    assign layer1_out[5856] = layer0_out[4438];
    assign layer1_out[5857] = layer0_out[6579] & ~layer0_out[6578];
    assign layer1_out[5858] = ~layer0_out[3513];
    assign layer1_out[5859] = layer0_out[5080];
    assign layer1_out[5860] = layer0_out[7442];
    assign layer1_out[5861] = layer0_out[7993];
    assign layer1_out[5862] = layer0_out[387];
    assign layer1_out[5863] = ~layer0_out[5519] | layer0_out[5520];
    assign layer1_out[5864] = layer0_out[5413];
    assign layer1_out[5865] = layer0_out[3158] & ~layer0_out[3157];
    assign layer1_out[5866] = ~(layer0_out[3864] ^ layer0_out[3865]);
    assign layer1_out[5867] = layer0_out[4331] ^ layer0_out[4332];
    assign layer1_out[5868] = layer0_out[3219] & ~layer0_out[3218];
    assign layer1_out[5869] = layer0_out[7849] & ~layer0_out[7848];
    assign layer1_out[5870] = ~layer0_out[811] | layer0_out[812];
    assign layer1_out[5871] = layer0_out[3054];
    assign layer1_out[5872] = ~(layer0_out[653] | layer0_out[654]);
    assign layer1_out[5873] = 1'b0;
    assign layer1_out[5874] = ~layer0_out[7955] | layer0_out[7956];
    assign layer1_out[5875] = ~layer0_out[2142];
    assign layer1_out[5876] = ~layer0_out[4095];
    assign layer1_out[5877] = ~layer0_out[58] | layer0_out[57];
    assign layer1_out[5878] = ~layer0_out[7954];
    assign layer1_out[5879] = ~layer0_out[3061];
    assign layer1_out[5880] = layer0_out[915] & ~layer0_out[914];
    assign layer1_out[5881] = ~(layer0_out[4866] | layer0_out[4867]);
    assign layer1_out[5882] = 1'b0;
    assign layer1_out[5883] = ~layer0_out[7932] | layer0_out[7931];
    assign layer1_out[5884] = layer0_out[3796];
    assign layer1_out[5885] = ~layer0_out[5922];
    assign layer1_out[5886] = ~(layer0_out[5282] & layer0_out[5283]);
    assign layer1_out[5887] = ~layer0_out[4037];
    assign layer1_out[5888] = ~layer0_out[4721];
    assign layer1_out[5889] = layer0_out[4441];
    assign layer1_out[5890] = layer0_out[6548];
    assign layer1_out[5891] = layer0_out[6221] & ~layer0_out[6220];
    assign layer1_out[5892] = layer0_out[7026];
    assign layer1_out[5893] = ~layer0_out[6592] | layer0_out[6591];
    assign layer1_out[5894] = ~layer0_out[5931];
    assign layer1_out[5895] = ~layer0_out[3963];
    assign layer1_out[5896] = layer0_out[601];
    assign layer1_out[5897] = layer0_out[4479] | layer0_out[4480];
    assign layer1_out[5898] = ~(layer0_out[580] & layer0_out[581]);
    assign layer1_out[5899] = layer0_out[282] & layer0_out[283];
    assign layer1_out[5900] = ~layer0_out[6819];
    assign layer1_out[5901] = layer0_out[4182] | layer0_out[4183];
    assign layer1_out[5902] = layer0_out[6410];
    assign layer1_out[5903] = layer0_out[4477] & ~layer0_out[4478];
    assign layer1_out[5904] = layer0_out[7685];
    assign layer1_out[5905] = ~layer0_out[744] | layer0_out[745];
    assign layer1_out[5906] = layer0_out[1479] & ~layer0_out[1478];
    assign layer1_out[5907] = layer0_out[5542] | layer0_out[5543];
    assign layer1_out[5908] = ~layer0_out[3426] | layer0_out[3427];
    assign layer1_out[5909] = ~layer0_out[3901];
    assign layer1_out[5910] = ~layer0_out[2584];
    assign layer1_out[5911] = layer0_out[2512];
    assign layer1_out[5912] = layer0_out[1482];
    assign layer1_out[5913] = ~(layer0_out[6217] & layer0_out[6218]);
    assign layer1_out[5914] = layer0_out[2451] ^ layer0_out[2452];
    assign layer1_out[5915] = 1'b0;
    assign layer1_out[5916] = ~layer0_out[911];
    assign layer1_out[5917] = ~layer0_out[4753] | layer0_out[4752];
    assign layer1_out[5918] = layer0_out[6065];
    assign layer1_out[5919] = ~layer0_out[7446];
    assign layer1_out[5920] = ~layer0_out[1324] | layer0_out[1323];
    assign layer1_out[5921] = ~layer0_out[1035] | layer0_out[1036];
    assign layer1_out[5922] = ~layer0_out[6259] | layer0_out[6258];
    assign layer1_out[5923] = layer0_out[4714] & ~layer0_out[4713];
    assign layer1_out[5924] = layer0_out[7091];
    assign layer1_out[5925] = 1'b0;
    assign layer1_out[5926] = layer0_out[5798];
    assign layer1_out[5927] = layer0_out[108] ^ layer0_out[109];
    assign layer1_out[5928] = ~layer0_out[2837];
    assign layer1_out[5929] = ~(layer0_out[481] | layer0_out[482]);
    assign layer1_out[5930] = layer0_out[3679] & layer0_out[3680];
    assign layer1_out[5931] = ~(layer0_out[5244] | layer0_out[5245]);
    assign layer1_out[5932] = ~layer0_out[2457] | layer0_out[2456];
    assign layer1_out[5933] = layer0_out[4092];
    assign layer1_out[5934] = ~layer0_out[5323];
    assign layer1_out[5935] = ~layer0_out[4581] | layer0_out[4580];
    assign layer1_out[5936] = layer0_out[354];
    assign layer1_out[5937] = layer0_out[2662];
    assign layer1_out[5938] = ~layer0_out[7659];
    assign layer1_out[5939] = layer0_out[3604] & ~layer0_out[3605];
    assign layer1_out[5940] = layer0_out[3509];
    assign layer1_out[5941] = ~layer0_out[7520] | layer0_out[7519];
    assign layer1_out[5942] = ~layer0_out[4414];
    assign layer1_out[5943] = layer0_out[488] & layer0_out[489];
    assign layer1_out[5944] = ~(layer0_out[959] | layer0_out[960]);
    assign layer1_out[5945] = ~(layer0_out[2848] | layer0_out[2849]);
    assign layer1_out[5946] = ~(layer0_out[3652] & layer0_out[3653]);
    assign layer1_out[5947] = ~(layer0_out[1184] | layer0_out[1185]);
    assign layer1_out[5948] = layer0_out[7053] ^ layer0_out[7054];
    assign layer1_out[5949] = layer0_out[6543] & layer0_out[6544];
    assign layer1_out[5950] = ~(layer0_out[7386] & layer0_out[7387]);
    assign layer1_out[5951] = ~(layer0_out[4135] ^ layer0_out[4136]);
    assign layer1_out[5952] = layer0_out[3339];
    assign layer1_out[5953] = ~(layer0_out[5018] | layer0_out[5019]);
    assign layer1_out[5954] = ~(layer0_out[2885] & layer0_out[2886]);
    assign layer1_out[5955] = ~(layer0_out[3630] & layer0_out[3631]);
    assign layer1_out[5956] = layer0_out[6908];
    assign layer1_out[5957] = ~(layer0_out[3416] & layer0_out[3417]);
    assign layer1_out[5958] = ~layer0_out[722];
    assign layer1_out[5959] = ~layer0_out[6005];
    assign layer1_out[5960] = ~(layer0_out[5344] ^ layer0_out[5345]);
    assign layer1_out[5961] = ~layer0_out[7748];
    assign layer1_out[5962] = 1'b0;
    assign layer1_out[5963] = 1'b0;
    assign layer1_out[5964] = layer0_out[2414];
    assign layer1_out[5965] = ~(layer0_out[1627] & layer0_out[1628]);
    assign layer1_out[5966] = layer0_out[5858] & layer0_out[5859];
    assign layer1_out[5967] = ~layer0_out[1398] | layer0_out[1399];
    assign layer1_out[5968] = layer0_out[2714];
    assign layer1_out[5969] = ~layer0_out[7131];
    assign layer1_out[5970] = ~(layer0_out[2190] & layer0_out[2191]);
    assign layer1_out[5971] = ~layer0_out[7819];
    assign layer1_out[5972] = layer0_out[445] | layer0_out[446];
    assign layer1_out[5973] = layer0_out[4337] | layer0_out[4338];
    assign layer1_out[5974] = ~layer0_out[2594] | layer0_out[2595];
    assign layer1_out[5975] = ~layer0_out[5457] | layer0_out[5458];
    assign layer1_out[5976] = layer0_out[7551] ^ layer0_out[7552];
    assign layer1_out[5977] = ~(layer0_out[4437] ^ layer0_out[4438]);
    assign layer1_out[5978] = ~layer0_out[1849] | layer0_out[1850];
    assign layer1_out[5979] = layer0_out[3210];
    assign layer1_out[5980] = ~layer0_out[2744];
    assign layer1_out[5981] = ~layer0_out[2682] | layer0_out[2683];
    assign layer1_out[5982] = ~(layer0_out[9] | layer0_out[10]);
    assign layer1_out[5983] = layer0_out[5332] | layer0_out[5333];
    assign layer1_out[5984] = ~layer0_out[7148] | layer0_out[7147];
    assign layer1_out[5985] = ~(layer0_out[3514] ^ layer0_out[3515]);
    assign layer1_out[5986] = ~(layer0_out[7832] & layer0_out[7833]);
    assign layer1_out[5987] = ~layer0_out[2632];
    assign layer1_out[5988] = ~layer0_out[3936];
    assign layer1_out[5989] = layer0_out[5440] & ~layer0_out[5439];
    assign layer1_out[5990] = layer0_out[6706] | layer0_out[6707];
    assign layer1_out[5991] = ~layer0_out[59];
    assign layer1_out[5992] = layer0_out[6959];
    assign layer1_out[5993] = layer0_out[2968] ^ layer0_out[2969];
    assign layer1_out[5994] = 1'b1;
    assign layer1_out[5995] = ~(layer0_out[2388] | layer0_out[2389]);
    assign layer1_out[5996] = ~layer0_out[1447] | layer0_out[1446];
    assign layer1_out[5997] = ~(layer0_out[7486] ^ layer0_out[7487]);
    assign layer1_out[5998] = 1'b1;
    assign layer1_out[5999] = ~layer0_out[2167];
    assign layer1_out[6000] = layer0_out[7252] & layer0_out[7253];
    assign layer1_out[6001] = ~layer0_out[2703];
    assign layer1_out[6002] = ~(layer0_out[7108] & layer0_out[7109]);
    assign layer1_out[6003] = ~(layer0_out[2275] & layer0_out[2276]);
    assign layer1_out[6004] = layer0_out[7609];
    assign layer1_out[6005] = layer0_out[5504] | layer0_out[5505];
    assign layer1_out[6006] = ~(layer0_out[7799] | layer0_out[7800]);
    assign layer1_out[6007] = layer0_out[791];
    assign layer1_out[6008] = layer0_out[462] | layer0_out[463];
    assign layer1_out[6009] = ~(layer0_out[7805] ^ layer0_out[7806]);
    assign layer1_out[6010] = ~layer0_out[5052] | layer0_out[5051];
    assign layer1_out[6011] = ~layer0_out[7474] | layer0_out[7475];
    assign layer1_out[6012] = ~layer0_out[905];
    assign layer1_out[6013] = layer0_out[6378];
    assign layer1_out[6014] = ~(layer0_out[3748] ^ layer0_out[3749]);
    assign layer1_out[6015] = layer0_out[5442] & ~layer0_out[5443];
    assign layer1_out[6016] = 1'b0;
    assign layer1_out[6017] = layer0_out[2402] & ~layer0_out[2403];
    assign layer1_out[6018] = 1'b1;
    assign layer1_out[6019] = layer0_out[4298] & ~layer0_out[4299];
    assign layer1_out[6020] = ~layer0_out[7548];
    assign layer1_out[6021] = layer0_out[6056];
    assign layer1_out[6022] = layer0_out[4701];
    assign layer1_out[6023] = layer0_out[2481];
    assign layer1_out[6024] = layer0_out[1111] | layer0_out[1112];
    assign layer1_out[6025] = layer0_out[2751] & ~layer0_out[2752];
    assign layer1_out[6026] = layer0_out[4126] & ~layer0_out[4125];
    assign layer1_out[6027] = ~layer0_out[5324] | layer0_out[5323];
    assign layer1_out[6028] = ~layer0_out[836];
    assign layer1_out[6029] = layer0_out[4175] ^ layer0_out[4176];
    assign layer1_out[6030] = 1'b0;
    assign layer1_out[6031] = layer0_out[6457] & layer0_out[6458];
    assign layer1_out[6032] = layer0_out[7297];
    assign layer1_out[6033] = ~(layer0_out[1328] & layer0_out[1329]);
    assign layer1_out[6034] = ~layer0_out[5209] | layer0_out[5208];
    assign layer1_out[6035] = layer0_out[3562];
    assign layer1_out[6036] = 1'b1;
    assign layer1_out[6037] = ~layer0_out[840];
    assign layer1_out[6038] = ~layer0_out[7283];
    assign layer1_out[6039] = layer0_out[1771] & ~layer0_out[1770];
    assign layer1_out[6040] = ~layer0_out[6691];
    assign layer1_out[6041] = ~(layer0_out[6439] & layer0_out[6440]);
    assign layer1_out[6042] = layer0_out[6856];
    assign layer1_out[6043] = layer0_out[4317] ^ layer0_out[4318];
    assign layer1_out[6044] = layer0_out[1557] ^ layer0_out[1558];
    assign layer1_out[6045] = layer0_out[7273];
    assign layer1_out[6046] = layer0_out[1431] ^ layer0_out[1432];
    assign layer1_out[6047] = ~layer0_out[2469] | layer0_out[2470];
    assign layer1_out[6048] = ~layer0_out[1125];
    assign layer1_out[6049] = 1'b0;
    assign layer1_out[6050] = layer0_out[1580];
    assign layer1_out[6051] = layer0_out[106] & layer0_out[107];
    assign layer1_out[6052] = ~(layer0_out[3007] & layer0_out[3008]);
    assign layer1_out[6053] = layer0_out[383] & layer0_out[384];
    assign layer1_out[6054] = layer0_out[4804] & ~layer0_out[4805];
    assign layer1_out[6055] = layer0_out[6142] & ~layer0_out[6143];
    assign layer1_out[6056] = 1'b1;
    assign layer1_out[6057] = layer0_out[7245] & ~layer0_out[7244];
    assign layer1_out[6058] = ~layer0_out[5351] | layer0_out[5350];
    assign layer1_out[6059] = layer0_out[7241];
    assign layer1_out[6060] = ~layer0_out[212];
    assign layer1_out[6061] = ~(layer0_out[2044] & layer0_out[2045]);
    assign layer1_out[6062] = ~layer0_out[3101];
    assign layer1_out[6063] = layer0_out[5645];
    assign layer1_out[6064] = layer0_out[4723];
    assign layer1_out[6065] = layer0_out[5580] | layer0_out[5581];
    assign layer1_out[6066] = layer0_out[1654];
    assign layer1_out[6067] = layer0_out[5455];
    assign layer1_out[6068] = layer0_out[6459];
    assign layer1_out[6069] = ~layer0_out[3509];
    assign layer1_out[6070] = ~layer0_out[6246] | layer0_out[6245];
    assign layer1_out[6071] = layer0_out[6672] ^ layer0_out[6673];
    assign layer1_out[6072] = ~(layer0_out[6795] & layer0_out[6796]);
    assign layer1_out[6073] = layer0_out[1021];
    assign layer1_out[6074] = 1'b0;
    assign layer1_out[6075] = layer0_out[4831] & layer0_out[4832];
    assign layer1_out[6076] = layer0_out[6818];
    assign layer1_out[6077] = layer0_out[3039] & ~layer0_out[3040];
    assign layer1_out[6078] = layer0_out[1539];
    assign layer1_out[6079] = ~layer0_out[2095];
    assign layer1_out[6080] = ~layer0_out[2764];
    assign layer1_out[6081] = layer0_out[6491] & ~layer0_out[6492];
    assign layer1_out[6082] = layer0_out[2573];
    assign layer1_out[6083] = layer0_out[5833] ^ layer0_out[5834];
    assign layer1_out[6084] = ~layer0_out[4129] | layer0_out[4130];
    assign layer1_out[6085] = layer0_out[780] & layer0_out[781];
    assign layer1_out[6086] = layer0_out[1632] ^ layer0_out[1633];
    assign layer1_out[6087] = layer0_out[3990] ^ layer0_out[3991];
    assign layer1_out[6088] = layer0_out[3544] & ~layer0_out[3545];
    assign layer1_out[6089] = ~layer0_out[1730] | layer0_out[1729];
    assign layer1_out[6090] = ~layer0_out[949] | layer0_out[948];
    assign layer1_out[6091] = ~layer0_out[1425] | layer0_out[1426];
    assign layer1_out[6092] = layer0_out[5299] | layer0_out[5300];
    assign layer1_out[6093] = layer0_out[2735];
    assign layer1_out[6094] = layer0_out[2465];
    assign layer1_out[6095] = ~layer0_out[6172] | layer0_out[6171];
    assign layer1_out[6096] = layer0_out[230] | layer0_out[231];
    assign layer1_out[6097] = ~layer0_out[2549] | layer0_out[2550];
    assign layer1_out[6098] = ~(layer0_out[349] | layer0_out[350]);
    assign layer1_out[6099] = layer0_out[6646] & ~layer0_out[6645];
    assign layer1_out[6100] = layer0_out[3758] | layer0_out[3759];
    assign layer1_out[6101] = ~layer0_out[4403];
    assign layer1_out[6102] = layer0_out[4855] | layer0_out[4856];
    assign layer1_out[6103] = ~layer0_out[6424];
    assign layer1_out[6104] = ~layer0_out[6464];
    assign layer1_out[6105] = ~layer0_out[2269];
    assign layer1_out[6106] = 1'b0;
    assign layer1_out[6107] = 1'b1;
    assign layer1_out[6108] = ~layer0_out[3789];
    assign layer1_out[6109] = ~layer0_out[5929] | layer0_out[5928];
    assign layer1_out[6110] = layer0_out[1304] ^ layer0_out[1305];
    assign layer1_out[6111] = layer0_out[291];
    assign layer1_out[6112] = ~(layer0_out[4068] & layer0_out[4069]);
    assign layer1_out[6113] = layer0_out[1969];
    assign layer1_out[6114] = ~layer0_out[7310] | layer0_out[7309];
    assign layer1_out[6115] = ~(layer0_out[1275] & layer0_out[1276]);
    assign layer1_out[6116] = ~(layer0_out[1776] ^ layer0_out[1777]);
    assign layer1_out[6117] = ~(layer0_out[4027] | layer0_out[4028]);
    assign layer1_out[6118] = layer0_out[2598];
    assign layer1_out[6119] = ~(layer0_out[4260] & layer0_out[4261]);
    assign layer1_out[6120] = ~layer0_out[3811];
    assign layer1_out[6121] = ~layer0_out[7362] | layer0_out[7361];
    assign layer1_out[6122] = 1'b0;
    assign layer1_out[6123] = ~(layer0_out[2381] | layer0_out[2382]);
    assign layer1_out[6124] = ~(layer0_out[2325] ^ layer0_out[2326]);
    assign layer1_out[6125] = ~(layer0_out[2627] ^ layer0_out[2628]);
    assign layer1_out[6126] = layer0_out[7174] | layer0_out[7175];
    assign layer1_out[6127] = layer0_out[3444] ^ layer0_out[3445];
    assign layer1_out[6128] = layer0_out[5517];
    assign layer1_out[6129] = ~layer0_out[3724];
    assign layer1_out[6130] = layer0_out[3965] & layer0_out[3966];
    assign layer1_out[6131] = layer0_out[4803] & ~layer0_out[4804];
    assign layer1_out[6132] = ~layer0_out[4886];
    assign layer1_out[6133] = ~layer0_out[22] | layer0_out[23];
    assign layer1_out[6134] = ~layer0_out[2707];
    assign layer1_out[6135] = layer0_out[7464] ^ layer0_out[7465];
    assign layer1_out[6136] = ~layer0_out[1866] | layer0_out[1865];
    assign layer1_out[6137] = ~(layer0_out[4920] & layer0_out[4921]);
    assign layer1_out[6138] = layer0_out[6511] | layer0_out[6512];
    assign layer1_out[6139] = ~layer0_out[5158];
    assign layer1_out[6140] = ~layer0_out[6893] | layer0_out[6892];
    assign layer1_out[6141] = ~layer0_out[3533] | layer0_out[3532];
    assign layer1_out[6142] = ~layer0_out[2771];
    assign layer1_out[6143] = ~(layer0_out[3038] | layer0_out[3039]);
    assign layer1_out[6144] = layer0_out[1848];
    assign layer1_out[6145] = ~(layer0_out[1364] ^ layer0_out[1365]);
    assign layer1_out[6146] = layer0_out[2835] & layer0_out[2836];
    assign layer1_out[6147] = layer0_out[7549] | layer0_out[7550];
    assign layer1_out[6148] = ~layer0_out[6306] | layer0_out[6307];
    assign layer1_out[6149] = layer0_out[275] & ~layer0_out[276];
    assign layer1_out[6150] = layer0_out[5705];
    assign layer1_out[6151] = ~(layer0_out[5873] | layer0_out[5874]);
    assign layer1_out[6152] = layer0_out[4140];
    assign layer1_out[6153] = layer0_out[7112];
    assign layer1_out[6154] = layer0_out[4346] ^ layer0_out[4347];
    assign layer1_out[6155] = ~layer0_out[3043] | layer0_out[3044];
    assign layer1_out[6156] = 1'b1;
    assign layer1_out[6157] = layer0_out[4762] & ~layer0_out[4761];
    assign layer1_out[6158] = layer0_out[7055] ^ layer0_out[7056];
    assign layer1_out[6159] = ~(layer0_out[5950] | layer0_out[5951]);
    assign layer1_out[6160] = ~(layer0_out[4025] | layer0_out[4026]);
    assign layer1_out[6161] = layer0_out[2379] & ~layer0_out[2380];
    assign layer1_out[6162] = layer0_out[9];
    assign layer1_out[6163] = layer0_out[2509];
    assign layer1_out[6164] = ~layer0_out[6151];
    assign layer1_out[6165] = ~(layer0_out[5338] ^ layer0_out[5339]);
    assign layer1_out[6166] = ~layer0_out[1062];
    assign layer1_out[6167] = ~layer0_out[4064] | layer0_out[4063];
    assign layer1_out[6168] = ~layer0_out[1222] | layer0_out[1221];
    assign layer1_out[6169] = layer0_out[41] | layer0_out[42];
    assign layer1_out[6170] = ~layer0_out[1727];
    assign layer1_out[6171] = layer0_out[509];
    assign layer1_out[6172] = ~layer0_out[2446] | layer0_out[2445];
    assign layer1_out[6173] = layer0_out[733] & ~layer0_out[734];
    assign layer1_out[6174] = ~layer0_out[2028];
    assign layer1_out[6175] = ~layer0_out[3093] | layer0_out[3092];
    assign layer1_out[6176] = ~layer0_out[7499];
    assign layer1_out[6177] = layer0_out[4724] & ~layer0_out[4725];
    assign layer1_out[6178] = ~layer0_out[3764] | layer0_out[3763];
    assign layer1_out[6179] = ~layer0_out[5930] | layer0_out[5931];
    assign layer1_out[6180] = layer0_out[599] ^ layer0_out[600];
    assign layer1_out[6181] = layer0_out[2061];
    assign layer1_out[6182] = ~layer0_out[7373];
    assign layer1_out[6183] = ~(layer0_out[5661] & layer0_out[5662]);
    assign layer1_out[6184] = layer0_out[5250];
    assign layer1_out[6185] = layer0_out[7603] & ~layer0_out[7602];
    assign layer1_out[6186] = layer0_out[2987] | layer0_out[2988];
    assign layer1_out[6187] = 1'b0;
    assign layer1_out[6188] = ~(layer0_out[752] ^ layer0_out[753]);
    assign layer1_out[6189] = layer0_out[3314];
    assign layer1_out[6190] = ~layer0_out[7992] | layer0_out[7991];
    assign layer1_out[6191] = layer0_out[63];
    assign layer1_out[6192] = ~layer0_out[5182];
    assign layer1_out[6193] = ~layer0_out[1596];
    assign layer1_out[6194] = 1'b1;
    assign layer1_out[6195] = layer0_out[2307];
    assign layer1_out[6196] = ~layer0_out[4084];
    assign layer1_out[6197] = layer0_out[1012] & layer0_out[1013];
    assign layer1_out[6198] = layer0_out[3374] & ~layer0_out[3375];
    assign layer1_out[6199] = ~layer0_out[5249];
    assign layer1_out[6200] = layer0_out[105] & layer0_out[106];
    assign layer1_out[6201] = ~layer0_out[6927];
    assign layer1_out[6202] = layer0_out[1684] ^ layer0_out[1685];
    assign layer1_out[6203] = ~layer0_out[4348] | layer0_out[4349];
    assign layer1_out[6204] = layer0_out[1573];
    assign layer1_out[6205] = 1'b0;
    assign layer1_out[6206] = ~(layer0_out[1077] ^ layer0_out[1078]);
    assign layer1_out[6207] = ~layer0_out[2393];
    assign layer1_out[6208] = ~layer0_out[7944];
    assign layer1_out[6209] = ~(layer0_out[5522] & layer0_out[5523]);
    assign layer1_out[6210] = ~layer0_out[2438];
    assign layer1_out[6211] = ~layer0_out[4075] | layer0_out[4076];
    assign layer1_out[6212] = layer0_out[1886];
    assign layer1_out[6213] = ~layer0_out[3612];
    assign layer1_out[6214] = layer0_out[3390];
    assign layer1_out[6215] = ~layer0_out[4442] | layer0_out[4443];
    assign layer1_out[6216] = ~(layer0_out[3725] ^ layer0_out[3726]);
    assign layer1_out[6217] = ~(layer0_out[229] | layer0_out[230]);
    assign layer1_out[6218] = layer0_out[6910] & layer0_out[6911];
    assign layer1_out[6219] = layer0_out[4246] & ~layer0_out[4245];
    assign layer1_out[6220] = layer0_out[4251] & ~layer0_out[4250];
    assign layer1_out[6221] = ~(layer0_out[4680] | layer0_out[4681]);
    assign layer1_out[6222] = layer0_out[1984] & layer0_out[1985];
    assign layer1_out[6223] = 1'b1;
    assign layer1_out[6224] = layer0_out[216] & ~layer0_out[217];
    assign layer1_out[6225] = layer0_out[6622] & layer0_out[6623];
    assign layer1_out[6226] = 1'b1;
    assign layer1_out[6227] = ~(layer0_out[5722] ^ layer0_out[5723]);
    assign layer1_out[6228] = ~layer0_out[4952] | layer0_out[4953];
    assign layer1_out[6229] = layer0_out[894];
    assign layer1_out[6230] = layer0_out[6825] | layer0_out[6826];
    assign layer1_out[6231] = layer0_out[400];
    assign layer1_out[6232] = layer0_out[7892] & layer0_out[7893];
    assign layer1_out[6233] = layer0_out[6590];
    assign layer1_out[6234] = layer0_out[7079];
    assign layer1_out[6235] = layer0_out[6563] & layer0_out[6564];
    assign layer1_out[6236] = layer0_out[1196] | layer0_out[1197];
    assign layer1_out[6237] = ~layer0_out[6473] | layer0_out[6474];
    assign layer1_out[6238] = ~(layer0_out[2492] & layer0_out[2493]);
    assign layer1_out[6239] = layer0_out[1817] ^ layer0_out[1818];
    assign layer1_out[6240] = ~(layer0_out[6190] | layer0_out[6191]);
    assign layer1_out[6241] = layer0_out[3174] ^ layer0_out[3175];
    assign layer1_out[6242] = ~(layer0_out[1467] | layer0_out[1468]);
    assign layer1_out[6243] = ~(layer0_out[6213] | layer0_out[6214]);
    assign layer1_out[6244] = layer0_out[7720] & ~layer0_out[7719];
    assign layer1_out[6245] = layer0_out[2186];
    assign layer1_out[6246] = ~(layer0_out[2324] & layer0_out[2325]);
    assign layer1_out[6247] = ~(layer0_out[5403] | layer0_out[5404]);
    assign layer1_out[6248] = layer0_out[841];
    assign layer1_out[6249] = 1'b1;
    assign layer1_out[6250] = ~(layer0_out[2065] & layer0_out[2066]);
    assign layer1_out[6251] = ~(layer0_out[5823] ^ layer0_out[5824]);
    assign layer1_out[6252] = ~layer0_out[4137] | layer0_out[4136];
    assign layer1_out[6253] = ~layer0_out[5991] | layer0_out[5992];
    assign layer1_out[6254] = layer0_out[4029];
    assign layer1_out[6255] = ~layer0_out[1194] | layer0_out[1193];
    assign layer1_out[6256] = layer0_out[2372] & ~layer0_out[2373];
    assign layer1_out[6257] = ~(layer0_out[5476] & layer0_out[5477]);
    assign layer1_out[6258] = ~layer0_out[1530];
    assign layer1_out[6259] = layer0_out[1484] | layer0_out[1485];
    assign layer1_out[6260] = ~(layer0_out[5982] | layer0_out[5983]);
    assign layer1_out[6261] = ~layer0_out[7073] | layer0_out[7072];
    assign layer1_out[6262] = layer0_out[4009];
    assign layer1_out[6263] = layer0_out[179] & ~layer0_out[180];
    assign layer1_out[6264] = ~layer0_out[3629];
    assign layer1_out[6265] = ~layer0_out[2994] | layer0_out[2993];
    assign layer1_out[6266] = ~layer0_out[7829];
    assign layer1_out[6267] = ~(layer0_out[5166] & layer0_out[5167]);
    assign layer1_out[6268] = layer0_out[5784];
    assign layer1_out[6269] = ~(layer0_out[2166] | layer0_out[2167]);
    assign layer1_out[6270] = layer0_out[2117];
    assign layer1_out[6271] = ~(layer0_out[5633] & layer0_out[5634]);
    assign layer1_out[6272] = ~layer0_out[2077];
    assign layer1_out[6273] = ~(layer0_out[7907] & layer0_out[7908]);
    assign layer1_out[6274] = ~(layer0_out[2467] & layer0_out[2468]);
    assign layer1_out[6275] = ~(layer0_out[885] | layer0_out[886]);
    assign layer1_out[6276] = layer0_out[1316];
    assign layer1_out[6277] = ~layer0_out[3283] | layer0_out[3282];
    assign layer1_out[6278] = layer0_out[5566] & layer0_out[5567];
    assign layer1_out[6279] = ~(layer0_out[2825] & layer0_out[2826]);
    assign layer1_out[6280] = 1'b0;
    assign layer1_out[6281] = 1'b1;
    assign layer1_out[6282] = layer0_out[5116] & layer0_out[5117];
    assign layer1_out[6283] = ~layer0_out[771];
    assign layer1_out[6284] = ~layer0_out[2411] | layer0_out[2412];
    assign layer1_out[6285] = ~layer0_out[4171] | layer0_out[4172];
    assign layer1_out[6286] = layer0_out[6241] | layer0_out[6242];
    assign layer1_out[6287] = ~layer0_out[5516] | layer0_out[5517];
    assign layer1_out[6288] = layer0_out[7526] & layer0_out[7527];
    assign layer1_out[6289] = ~layer0_out[997];
    assign layer1_out[6290] = layer0_out[6316] | layer0_out[6317];
    assign layer1_out[6291] = layer0_out[2726] ^ layer0_out[2727];
    assign layer1_out[6292] = layer0_out[843] & ~layer0_out[842];
    assign layer1_out[6293] = ~(layer0_out[3940] & layer0_out[3941]);
    assign layer1_out[6294] = ~layer0_out[4763];
    assign layer1_out[6295] = layer0_out[2272] & ~layer0_out[2273];
    assign layer1_out[6296] = ~layer0_out[3511];
    assign layer1_out[6297] = ~(layer0_out[6677] ^ layer0_out[6678]);
    assign layer1_out[6298] = layer0_out[1568] & ~layer0_out[1567];
    assign layer1_out[6299] = layer0_out[4744];
    assign layer1_out[6300] = layer0_out[2454] & layer0_out[2455];
    assign layer1_out[6301] = ~layer0_out[5107];
    assign layer1_out[6302] = ~layer0_out[3876];
    assign layer1_out[6303] = ~layer0_out[5008] | layer0_out[5007];
    assign layer1_out[6304] = ~(layer0_out[3896] | layer0_out[3897]);
    assign layer1_out[6305] = layer0_out[6796];
    assign layer1_out[6306] = ~layer0_out[5111];
    assign layer1_out[6307] = ~layer0_out[1151] | layer0_out[1150];
    assign layer1_out[6308] = layer0_out[2386] & layer0_out[2387];
    assign layer1_out[6309] = layer0_out[3271] & ~layer0_out[3270];
    assign layer1_out[6310] = layer0_out[5423];
    assign layer1_out[6311] = ~(layer0_out[687] | layer0_out[688]);
    assign layer1_out[6312] = layer0_out[1118] & ~layer0_out[1119];
    assign layer1_out[6313] = layer0_out[2235] & layer0_out[2236];
    assign layer1_out[6314] = layer0_out[65] & ~layer0_out[64];
    assign layer1_out[6315] = ~(layer0_out[6384] & layer0_out[6385]);
    assign layer1_out[6316] = layer0_out[6545] | layer0_out[6546];
    assign layer1_out[6317] = layer0_out[4730];
    assign layer1_out[6318] = ~(layer0_out[2851] | layer0_out[2852]);
    assign layer1_out[6319] = ~layer0_out[4731];
    assign layer1_out[6320] = ~layer0_out[7903] | layer0_out[7904];
    assign layer1_out[6321] = layer0_out[3252] & ~layer0_out[3253];
    assign layer1_out[6322] = layer0_out[3479];
    assign layer1_out[6323] = layer0_out[4582];
    assign layer1_out[6324] = layer0_out[7995] & ~layer0_out[7996];
    assign layer1_out[6325] = ~layer0_out[2301];
    assign layer1_out[6326] = layer0_out[2068];
    assign layer1_out[6327] = layer0_out[3344];
    assign layer1_out[6328] = ~layer0_out[6848] | layer0_out[6847];
    assign layer1_out[6329] = ~layer0_out[5979];
    assign layer1_out[6330] = ~(layer0_out[1498] & layer0_out[1499]);
    assign layer1_out[6331] = 1'b1;
    assign layer1_out[6332] = layer0_out[1415] & ~layer0_out[1414];
    assign layer1_out[6333] = ~(layer0_out[6369] | layer0_out[6370]);
    assign layer1_out[6334] = layer0_out[2593];
    assign layer1_out[6335] = layer0_out[532];
    assign layer1_out[6336] = layer0_out[5395];
    assign layer1_out[6337] = layer0_out[2527] & layer0_out[2528];
    assign layer1_out[6338] = layer0_out[6153] & ~layer0_out[6152];
    assign layer1_out[6339] = ~layer0_out[4363];
    assign layer1_out[6340] = ~(layer0_out[5113] ^ layer0_out[5114]);
    assign layer1_out[6341] = layer0_out[6038];
    assign layer1_out[6342] = ~layer0_out[6041] | layer0_out[6042];
    assign layer1_out[6343] = ~layer0_out[4154];
    assign layer1_out[6344] = ~layer0_out[137] | layer0_out[136];
    assign layer1_out[6345] = layer0_out[2599] & ~layer0_out[2600];
    assign layer1_out[6346] = layer0_out[2670] | layer0_out[2671];
    assign layer1_out[6347] = ~(layer0_out[5141] | layer0_out[5142]);
    assign layer1_out[6348] = layer0_out[4497];
    assign layer1_out[6349] = layer0_out[6652] ^ layer0_out[6653];
    assign layer1_out[6350] = layer0_out[4358] | layer0_out[4359];
    assign layer1_out[6351] = ~layer0_out[6872] | layer0_out[6873];
    assign layer1_out[6352] = ~layer0_out[5072];
    assign layer1_out[6353] = ~(layer0_out[1280] & layer0_out[1281]);
    assign layer1_out[6354] = layer0_out[3947] & layer0_out[3948];
    assign layer1_out[6355] = layer0_out[292] & layer0_out[293];
    assign layer1_out[6356] = ~layer0_out[4139] | layer0_out[4138];
    assign layer1_out[6357] = layer0_out[7432] | layer0_out[7433];
    assign layer1_out[6358] = ~layer0_out[5362] | layer0_out[5363];
    assign layer1_out[6359] = ~layer0_out[6718] | layer0_out[6717];
    assign layer1_out[6360] = 1'b1;
    assign layer1_out[6361] = layer0_out[6062];
    assign layer1_out[6362] = 1'b0;
    assign layer1_out[6363] = layer0_out[4432] & ~layer0_out[4431];
    assign layer1_out[6364] = layer0_out[4357] | layer0_out[4358];
    assign layer1_out[6365] = ~layer0_out[6446];
    assign layer1_out[6366] = layer0_out[3939] & layer0_out[3940];
    assign layer1_out[6367] = 1'b1;
    assign layer1_out[6368] = layer0_out[116] & ~layer0_out[117];
    assign layer1_out[6369] = ~layer0_out[5313] | layer0_out[5314];
    assign layer1_out[6370] = ~layer0_out[1101];
    assign layer1_out[6371] = layer0_out[4906] & ~layer0_out[4905];
    assign layer1_out[6372] = ~(layer0_out[6331] ^ layer0_out[6332]);
    assign layer1_out[6373] = layer0_out[4544] & ~layer0_out[4545];
    assign layer1_out[6374] = ~layer0_out[5610];
    assign layer1_out[6375] = ~layer0_out[3164];
    assign layer1_out[6376] = 1'b1;
    assign layer1_out[6377] = layer0_out[3840] & ~layer0_out[3841];
    assign layer1_out[6378] = layer0_out[2538] | layer0_out[2539];
    assign layer1_out[6379] = ~(layer0_out[217] | layer0_out[218]);
    assign layer1_out[6380] = layer0_out[4611];
    assign layer1_out[6381] = ~layer0_out[7540] | layer0_out[7539];
    assign layer1_out[6382] = layer0_out[4926] & layer0_out[4927];
    assign layer1_out[6383] = ~(layer0_out[2869] | layer0_out[2870]);
    assign layer1_out[6384] = ~layer0_out[1153] | layer0_out[1154];
    assign layer1_out[6385] = ~(layer0_out[5749] & layer0_out[5750]);
    assign layer1_out[6386] = ~(layer0_out[4837] & layer0_out[4838]);
    assign layer1_out[6387] = ~(layer0_out[3701] | layer0_out[3702]);
    assign layer1_out[6388] = layer0_out[3142] & layer0_out[3143];
    assign layer1_out[6389] = ~(layer0_out[6247] & layer0_out[6248]);
    assign layer1_out[6390] = layer0_out[3671] & layer0_out[3672];
    assign layer1_out[6391] = ~layer0_out[682] | layer0_out[683];
    assign layer1_out[6392] = layer0_out[2723] & ~layer0_out[2722];
    assign layer1_out[6393] = ~layer0_out[1469] | layer0_out[1470];
    assign layer1_out[6394] = ~layer0_out[1507] | layer0_out[1506];
    assign layer1_out[6395] = ~layer0_out[4073];
    assign layer1_out[6396] = ~layer0_out[2847] | layer0_out[2848];
    assign layer1_out[6397] = layer0_out[2457];
    assign layer1_out[6398] = ~layer0_out[5590];
    assign layer1_out[6399] = ~layer0_out[4490];
    assign layer1_out[6400] = 1'b0;
    assign layer1_out[6401] = ~layer0_out[5603];
    assign layer1_out[6402] = ~(layer0_out[5527] | layer0_out[5528]);
    assign layer1_out[6403] = ~layer0_out[7146];
    assign layer1_out[6404] = layer0_out[5573] & ~layer0_out[5574];
    assign layer1_out[6405] = layer0_out[1416] & layer0_out[1417];
    assign layer1_out[6406] = layer0_out[4144] & ~layer0_out[4143];
    assign layer1_out[6407] = ~layer0_out[7431] | layer0_out[7432];
    assign layer1_out[6408] = layer0_out[2292];
    assign layer1_out[6409] = layer0_out[1045] & layer0_out[1046];
    assign layer1_out[6410] = layer0_out[5051];
    assign layer1_out[6411] = layer0_out[5929] & ~layer0_out[5930];
    assign layer1_out[6412] = layer0_out[269] & layer0_out[270];
    assign layer1_out[6413] = 1'b0;
    assign layer1_out[6414] = ~(layer0_out[2884] | layer0_out[2885]);
    assign layer1_out[6415] = ~layer0_out[2638];
    assign layer1_out[6416] = layer0_out[7875] ^ layer0_out[7876];
    assign layer1_out[6417] = layer0_out[59];
    assign layer1_out[6418] = ~(layer0_out[4623] & layer0_out[4624]);
    assign layer1_out[6419] = ~layer0_out[6836];
    assign layer1_out[6420] = ~layer0_out[4152] | layer0_out[4151];
    assign layer1_out[6421] = layer0_out[1852];
    assign layer1_out[6422] = ~layer0_out[5279] | layer0_out[5278];
    assign layer1_out[6423] = ~layer0_out[5919];
    assign layer1_out[6424] = ~(layer0_out[63] | layer0_out[64]);
    assign layer1_out[6425] = layer0_out[2276] & layer0_out[2277];
    assign layer1_out[6426] = layer0_out[776] & ~layer0_out[777];
    assign layer1_out[6427] = layer0_out[6531];
    assign layer1_out[6428] = layer0_out[4591];
    assign layer1_out[6429] = ~layer0_out[2233];
    assign layer1_out[6430] = ~layer0_out[254] | layer0_out[253];
    assign layer1_out[6431] = layer0_out[5847] | layer0_out[5848];
    assign layer1_out[6432] = ~layer0_out[3874];
    assign layer1_out[6433] = layer0_out[542];
    assign layer1_out[6434] = layer0_out[4935] & ~layer0_out[4936];
    assign layer1_out[6435] = layer0_out[1475];
    assign layer1_out[6436] = layer0_out[3324] & layer0_out[3325];
    assign layer1_out[6437] = 1'b1;
    assign layer1_out[6438] = layer0_out[3259];
    assign layer1_out[6439] = ~(layer0_out[7002] & layer0_out[7003]);
    assign layer1_out[6440] = layer0_out[2634] & ~layer0_out[2635];
    assign layer1_out[6441] = layer0_out[548] & ~layer0_out[549];
    assign layer1_out[6442] = ~layer0_out[6433] | layer0_out[6432];
    assign layer1_out[6443] = layer0_out[5402] ^ layer0_out[5403];
    assign layer1_out[6444] = ~(layer0_out[6658] | layer0_out[6659]);
    assign layer1_out[6445] = layer0_out[1108] ^ layer0_out[1109];
    assign layer1_out[6446] = layer0_out[6554];
    assign layer1_out[6447] = layer0_out[5727];
    assign layer1_out[6448] = ~layer0_out[5964] | layer0_out[5965];
    assign layer1_out[6449] = layer0_out[1412] & ~layer0_out[1411];
    assign layer1_out[6450] = ~(layer0_out[4874] & layer0_out[4875]);
    assign layer1_out[6451] = ~(layer0_out[6641] | layer0_out[6642]);
    assign layer1_out[6452] = ~layer0_out[6783] | layer0_out[6782];
    assign layer1_out[6453] = 1'b1;
    assign layer1_out[6454] = ~layer0_out[4273];
    assign layer1_out[6455] = ~layer0_out[3872] | layer0_out[3873];
    assign layer1_out[6456] = layer0_out[2038] & ~layer0_out[2039];
    assign layer1_out[6457] = layer0_out[2282] & layer0_out[2283];
    assign layer1_out[6458] = layer0_out[474];
    assign layer1_out[6459] = layer0_out[6158] | layer0_out[6159];
    assign layer1_out[6460] = ~layer0_out[5803] | layer0_out[5802];
    assign layer1_out[6461] = ~layer0_out[395];
    assign layer1_out[6462] = ~(layer0_out[7724] | layer0_out[7725]);
    assign layer1_out[6463] = ~layer0_out[1784];
    assign layer1_out[6464] = ~layer0_out[1696] | layer0_out[1697];
    assign layer1_out[6465] = ~layer0_out[7939] | layer0_out[7940];
    assign layer1_out[6466] = ~layer0_out[7769] | layer0_out[7770];
    assign layer1_out[6467] = ~layer0_out[703];
    assign layer1_out[6468] = layer0_out[3801];
    assign layer1_out[6469] = ~(layer0_out[21] ^ layer0_out[22]);
    assign layer1_out[6470] = ~(layer0_out[2586] | layer0_out[2587]);
    assign layer1_out[6471] = ~layer0_out[3960];
    assign layer1_out[6472] = layer0_out[6309] & layer0_out[6310];
    assign layer1_out[6473] = ~layer0_out[5542] | layer0_out[5541];
    assign layer1_out[6474] = layer0_out[2631] ^ layer0_out[2632];
    assign layer1_out[6475] = layer0_out[151];
    assign layer1_out[6476] = ~(layer0_out[7641] | layer0_out[7642]);
    assign layer1_out[6477] = layer0_out[3108];
    assign layer1_out[6478] = ~layer0_out[4848];
    assign layer1_out[6479] = layer0_out[6408];
    assign layer1_out[6480] = layer0_out[6858] | layer0_out[6859];
    assign layer1_out[6481] = layer0_out[3106] ^ layer0_out[3107];
    assign layer1_out[6482] = layer0_out[6036];
    assign layer1_out[6483] = layer0_out[4071];
    assign layer1_out[6484] = layer0_out[5851];
    assign layer1_out[6485] = ~layer0_out[5975];
    assign layer1_out[6486] = ~layer0_out[5000];
    assign layer1_out[6487] = ~layer0_out[3654];
    assign layer1_out[6488] = ~layer0_out[4288];
    assign layer1_out[6489] = layer0_out[6454] | layer0_out[6455];
    assign layer1_out[6490] = layer0_out[3446] & layer0_out[3447];
    assign layer1_out[6491] = layer0_out[7567] & layer0_out[7568];
    assign layer1_out[6492] = ~(layer0_out[7213] & layer0_out[7214]);
    assign layer1_out[6493] = layer0_out[1499] & layer0_out[1500];
    assign layer1_out[6494] = ~layer0_out[5009];
    assign layer1_out[6495] = layer0_out[5457] & ~layer0_out[5456];
    assign layer1_out[6496] = layer0_out[2996];
    assign layer1_out[6497] = layer0_out[327] | layer0_out[328];
    assign layer1_out[6498] = layer0_out[7052];
    assign layer1_out[6499] = ~layer0_out[7933];
    assign layer1_out[6500] = layer0_out[1036] ^ layer0_out[1037];
    assign layer1_out[6501] = ~layer0_out[1041];
    assign layer1_out[6502] = ~layer0_out[7152];
    assign layer1_out[6503] = layer0_out[7304];
    assign layer1_out[6504] = layer0_out[1931] ^ layer0_out[1932];
    assign layer1_out[6505] = layer0_out[7095] & layer0_out[7096];
    assign layer1_out[6506] = layer0_out[429] | layer0_out[430];
    assign layer1_out[6507] = ~layer0_out[2783] | layer0_out[2784];
    assign layer1_out[6508] = layer0_out[280];
    assign layer1_out[6509] = layer0_out[3420] ^ layer0_out[3421];
    assign layer1_out[6510] = ~(layer0_out[7150] & layer0_out[7151]);
    assign layer1_out[6511] = ~layer0_out[7948];
    assign layer1_out[6512] = layer0_out[3608];
    assign layer1_out[6513] = layer0_out[3722] & ~layer0_out[3721];
    assign layer1_out[6514] = layer0_out[5848] & ~layer0_out[5849];
    assign layer1_out[6515] = layer0_out[4797] & layer0_out[4798];
    assign layer1_out[6516] = ~(layer0_out[2577] ^ layer0_out[2578]);
    assign layer1_out[6517] = layer0_out[7575] & ~layer0_out[7574];
    assign layer1_out[6518] = layer0_out[7737];
    assign layer1_out[6519] = layer0_out[5593];
    assign layer1_out[6520] = layer0_out[6013];
    assign layer1_out[6521] = layer0_out[7094];
    assign layer1_out[6522] = ~layer0_out[6367];
    assign layer1_out[6523] = ~(layer0_out[4127] | layer0_out[4128]);
    assign layer1_out[6524] = layer0_out[628] & ~layer0_out[627];
    assign layer1_out[6525] = ~(layer0_out[6211] ^ layer0_out[6212]);
    assign layer1_out[6526] = ~layer0_out[6309];
    assign layer1_out[6527] = ~layer0_out[1208];
    assign layer1_out[6528] = ~(layer0_out[1981] | layer0_out[1982]);
    assign layer1_out[6529] = 1'b1;
    assign layer1_out[6530] = ~layer0_out[2345] | layer0_out[2346];
    assign layer1_out[6531] = layer0_out[5444] & ~layer0_out[5443];
    assign layer1_out[6532] = layer0_out[2545] & layer0_out[2546];
    assign layer1_out[6533] = layer0_out[2143] & layer0_out[2144];
    assign layer1_out[6534] = ~(layer0_out[4320] & layer0_out[4321]);
    assign layer1_out[6535] = layer0_out[4433] | layer0_out[4434];
    assign layer1_out[6536] = layer0_out[525] | layer0_out[526];
    assign layer1_out[6537] = layer0_out[5409];
    assign layer1_out[6538] = ~layer0_out[6216];
    assign layer1_out[6539] = layer0_out[7387];
    assign layer1_out[6540] = ~layer0_out[2012] | layer0_out[2013];
    assign layer1_out[6541] = ~layer0_out[6380] | layer0_out[6381];
    assign layer1_out[6542] = ~(layer0_out[623] & layer0_out[624]);
    assign layer1_out[6543] = 1'b1;
    assign layer1_out[6544] = ~layer0_out[6954];
    assign layer1_out[6545] = ~layer0_out[4366];
    assign layer1_out[6546] = ~layer0_out[2790];
    assign layer1_out[6547] = ~layer0_out[3455];
    assign layer1_out[6548] = ~layer0_out[2127];
    assign layer1_out[6549] = layer0_out[1153] & ~layer0_out[1152];
    assign layer1_out[6550] = 1'b1;
    assign layer1_out[6551] = layer0_out[3444] & ~layer0_out[3443];
    assign layer1_out[6552] = layer0_out[5415] & ~layer0_out[5416];
    assign layer1_out[6553] = layer0_out[5774];
    assign layer1_out[6554] = layer0_out[3609] & layer0_out[3610];
    assign layer1_out[6555] = layer0_out[1951] | layer0_out[1952];
    assign layer1_out[6556] = layer0_out[7249] & ~layer0_out[7248];
    assign layer1_out[6557] = ~layer0_out[5813];
    assign layer1_out[6558] = ~layer0_out[1240] | layer0_out[1241];
    assign layer1_out[6559] = ~(layer0_out[3869] ^ layer0_out[3870]);
    assign layer1_out[6560] = layer0_out[5785] ^ layer0_out[5786];
    assign layer1_out[6561] = layer0_out[6540];
    assign layer1_out[6562] = layer0_out[99] | layer0_out[100];
    assign layer1_out[6563] = layer0_out[4620] & layer0_out[4621];
    assign layer1_out[6564] = layer0_out[2966];
    assign layer1_out[6565] = layer0_out[3676];
    assign layer1_out[6566] = ~layer0_out[5674];
    assign layer1_out[6567] = ~layer0_out[7101];
    assign layer1_out[6568] = ~layer0_out[4385];
    assign layer1_out[6569] = ~(layer0_out[3618] | layer0_out[3619]);
    assign layer1_out[6570] = layer0_out[5843] & ~layer0_out[5844];
    assign layer1_out[6571] = layer0_out[1551];
    assign layer1_out[6572] = 1'b0;
    assign layer1_out[6573] = layer0_out[27];
    assign layer1_out[6574] = layer0_out[3128];
    assign layer1_out[6575] = ~(layer0_out[729] & layer0_out[730]);
    assign layer1_out[6576] = ~layer0_out[464];
    assign layer1_out[6577] = layer0_out[3913] ^ layer0_out[3914];
    assign layer1_out[6578] = layer0_out[5958] ^ layer0_out[5959];
    assign layer1_out[6579] = 1'b0;
    assign layer1_out[6580] = layer0_out[6116] ^ layer0_out[6117];
    assign layer1_out[6581] = ~(layer0_out[2489] | layer0_out[2490]);
    assign layer1_out[6582] = layer0_out[336] & layer0_out[337];
    assign layer1_out[6583] = ~layer0_out[5575];
    assign layer1_out[6584] = layer0_out[2149] & layer0_out[2150];
    assign layer1_out[6585] = ~layer0_out[5440] | layer0_out[5441];
    assign layer1_out[6586] = layer0_out[3307] & ~layer0_out[3306];
    assign layer1_out[6587] = ~layer0_out[4982];
    assign layer1_out[6588] = layer0_out[1553] | layer0_out[1554];
    assign layer1_out[6589] = ~layer0_out[1896] | layer0_out[1897];
    assign layer1_out[6590] = layer0_out[5382];
    assign layer1_out[6591] = layer0_out[6609];
    assign layer1_out[6592] = layer0_out[1430] | layer0_out[1431];
    assign layer1_out[6593] = layer0_out[3946] & ~layer0_out[3947];
    assign layer1_out[6594] = layer0_out[910];
    assign layer1_out[6595] = layer0_out[5187] & ~layer0_out[5188];
    assign layer1_out[6596] = layer0_out[7071];
    assign layer1_out[6597] = ~layer0_out[6655] | layer0_out[6656];
    assign layer1_out[6598] = layer0_out[7444] & ~layer0_out[7443];
    assign layer1_out[6599] = ~layer0_out[963] | layer0_out[964];
    assign layer1_out[6600] = layer0_out[189];
    assign layer1_out[6601] = layer0_out[303];
    assign layer1_out[6602] = ~layer0_out[291] | layer0_out[290];
    assign layer1_out[6603] = 1'b0;
    assign layer1_out[6604] = ~layer0_out[7472] | layer0_out[7471];
    assign layer1_out[6605] = ~layer0_out[7850] | layer0_out[7849];
    assign layer1_out[6606] = layer0_out[5260];
    assign layer1_out[6607] = ~layer0_out[5279];
    assign layer1_out[6608] = ~(layer0_out[6202] ^ layer0_out[6203]);
    assign layer1_out[6609] = layer0_out[5690];
    assign layer1_out[6610] = ~layer0_out[4103];
    assign layer1_out[6611] = ~layer0_out[5488] | layer0_out[5489];
    assign layer1_out[6612] = layer0_out[3906] ^ layer0_out[3907];
    assign layer1_out[6613] = 1'b1;
    assign layer1_out[6614] = layer0_out[2128] & ~layer0_out[2127];
    assign layer1_out[6615] = layer0_out[7730] & layer0_out[7731];
    assign layer1_out[6616] = layer0_out[6118] & layer0_out[6119];
    assign layer1_out[6617] = layer0_out[815] | layer0_out[816];
    assign layer1_out[6618] = ~layer0_out[3884];
    assign layer1_out[6619] = layer0_out[7659] ^ layer0_out[7660];
    assign layer1_out[6620] = layer0_out[4411] & ~layer0_out[4410];
    assign layer1_out[6621] = ~layer0_out[4519];
    assign layer1_out[6622] = ~(layer0_out[3211] & layer0_out[3212]);
    assign layer1_out[6623] = ~layer0_out[7353] | layer0_out[7352];
    assign layer1_out[6624] = 1'b1;
    assign layer1_out[6625] = ~layer0_out[6275] | layer0_out[6276];
    assign layer1_out[6626] = ~layer0_out[3881];
    assign layer1_out[6627] = ~layer0_out[4118];
    assign layer1_out[6628] = layer0_out[5093];
    assign layer1_out[6629] = layer0_out[1697];
    assign layer1_out[6630] = layer0_out[2493] ^ layer0_out[2494];
    assign layer1_out[6631] = layer0_out[5395];
    assign layer1_out[6632] = ~(layer0_out[4230] & layer0_out[4231]);
    assign layer1_out[6633] = 1'b0;
    assign layer1_out[6634] = layer0_out[888] | layer0_out[889];
    assign layer1_out[6635] = ~layer0_out[4995] | layer0_out[4996];
    assign layer1_out[6636] = ~(layer0_out[581] | layer0_out[582]);
    assign layer1_out[6637] = ~layer0_out[7729];
    assign layer1_out[6638] = layer0_out[4749];
    assign layer1_out[6639] = ~(layer0_out[6946] & layer0_out[6947]);
    assign layer1_out[6640] = layer0_out[2490];
    assign layer1_out[6641] = ~layer0_out[3491];
    assign layer1_out[6642] = 1'b0;
    assign layer1_out[6643] = ~(layer0_out[215] & layer0_out[216]);
    assign layer1_out[6644] = ~layer0_out[6261];
    assign layer1_out[6645] = layer0_out[7732];
    assign layer1_out[6646] = layer0_out[6300];
    assign layer1_out[6647] = ~layer0_out[3309];
    assign layer1_out[6648] = layer0_out[2067];
    assign layer1_out[6649] = ~layer0_out[6803] | layer0_out[6804];
    assign layer1_out[6650] = ~(layer0_out[4914] ^ layer0_out[4915]);
    assign layer1_out[6651] = layer0_out[96] & layer0_out[97];
    assign layer1_out[6652] = ~(layer0_out[3772] & layer0_out[3773]);
    assign layer1_out[6653] = ~layer0_out[2248];
    assign layer1_out[6654] = ~layer0_out[4741];
    assign layer1_out[6655] = ~layer0_out[5360] | layer0_out[5361];
    assign layer1_out[6656] = layer0_out[804];
    assign layer1_out[6657] = layer0_out[6784] & ~layer0_out[6785];
    assign layer1_out[6658] = ~layer0_out[1217];
    assign layer1_out[6659] = layer0_out[7416] & ~layer0_out[7417];
    assign layer1_out[6660] = ~layer0_out[4835] | layer0_out[4834];
    assign layer1_out[6661] = layer0_out[1873] & ~layer0_out[1874];
    assign layer1_out[6662] = layer0_out[5371];
    assign layer1_out[6663] = layer0_out[985] & ~layer0_out[984];
    assign layer1_out[6664] = ~layer0_out[1911];
    assign layer1_out[6665] = layer0_out[3502];
    assign layer1_out[6666] = ~layer0_out[7761] | layer0_out[7760];
    assign layer1_out[6667] = ~layer0_out[2193];
    assign layer1_out[6668] = layer0_out[4675] & layer0_out[4676];
    assign layer1_out[6669] = ~layer0_out[3078];
    assign layer1_out[6670] = layer0_out[5219];
    assign layer1_out[6671] = ~(layer0_out[4465] & layer0_out[4466]);
    assign layer1_out[6672] = ~layer0_out[672] | layer0_out[671];
    assign layer1_out[6673] = ~layer0_out[7124];
    assign layer1_out[6674] = layer0_out[2356] & ~layer0_out[2355];
    assign layer1_out[6675] = layer0_out[3257] | layer0_out[3258];
    assign layer1_out[6676] = 1'b1;
    assign layer1_out[6677] = ~layer0_out[1173];
    assign layer1_out[6678] = layer0_out[2788] & layer0_out[2789];
    assign layer1_out[6679] = layer0_out[6681];
    assign layer1_out[6680] = layer0_out[5705];
    assign layer1_out[6681] = 1'b0;
    assign layer1_out[6682] = ~layer0_out[2430];
    assign layer1_out[6683] = layer0_out[2120] | layer0_out[2121];
    assign layer1_out[6684] = layer0_out[4363] | layer0_out[4364];
    assign layer1_out[6685] = 1'b1;
    assign layer1_out[6686] = layer0_out[213];
    assign layer1_out[6687] = layer0_out[854] | layer0_out[855];
    assign layer1_out[6688] = layer0_out[3645];
    assign layer1_out[6689] = layer0_out[5431] & ~layer0_out[5430];
    assign layer1_out[6690] = layer0_out[758] & ~layer0_out[759];
    assign layer1_out[6691] = ~layer0_out[1575];
    assign layer1_out[6692] = layer0_out[1768];
    assign layer1_out[6693] = layer0_out[6899] & layer0_out[6900];
    assign layer1_out[6694] = layer0_out[964];
    assign layer1_out[6695] = 1'b0;
    assign layer1_out[6696] = ~layer0_out[4123];
    assign layer1_out[6697] = layer0_out[4227] & ~layer0_out[4226];
    assign layer1_out[6698] = layer0_out[3383];
    assign layer1_out[6699] = ~layer0_out[4490] | layer0_out[4491];
    assign layer1_out[6700] = ~layer0_out[5156];
    assign layer1_out[6701] = ~layer0_out[1488] | layer0_out[1487];
    assign layer1_out[6702] = layer0_out[7661];
    assign layer1_out[6703] = ~layer0_out[6552];
    assign layer1_out[6704] = ~layer0_out[1951];
    assign layer1_out[6705] = layer0_out[4254] | layer0_out[4255];
    assign layer1_out[6706] = layer0_out[3082] & layer0_out[3083];
    assign layer1_out[6707] = ~layer0_out[472];
    assign layer1_out[6708] = layer0_out[5160] & ~layer0_out[5161];
    assign layer1_out[6709] = ~layer0_out[7325];
    assign layer1_out[6710] = ~(layer0_out[3915] | layer0_out[3916]);
    assign layer1_out[6711] = layer0_out[6988] & ~layer0_out[6989];
    assign layer1_out[6712] = layer0_out[6310] ^ layer0_out[6311];
    assign layer1_out[6713] = ~layer0_out[1045] | layer0_out[1044];
    assign layer1_out[6714] = ~layer0_out[5903] | layer0_out[5902];
    assign layer1_out[6715] = layer0_out[7740] | layer0_out[7741];
    assign layer1_out[6716] = layer0_out[1925];
    assign layer1_out[6717] = layer0_out[6791] & layer0_out[6792];
    assign layer1_out[6718] = layer0_out[338];
    assign layer1_out[6719] = ~layer0_out[6742];
    assign layer1_out[6720] = ~(layer0_out[1670] | layer0_out[1671]);
    assign layer1_out[6721] = layer0_out[6106] | layer0_out[6107];
    assign layer1_out[6722] = ~layer0_out[6945] | layer0_out[6946];
    assign layer1_out[6723] = ~layer0_out[6352] | layer0_out[6351];
    assign layer1_out[6724] = layer0_out[7620];
    assign layer1_out[6725] = ~layer0_out[248] | layer0_out[247];
    assign layer1_out[6726] = ~layer0_out[6664] | layer0_out[6665];
    assign layer1_out[6727] = layer0_out[7632] | layer0_out[7633];
    assign layer1_out[6728] = layer0_out[6671] ^ layer0_out[6672];
    assign layer1_out[6729] = 1'b0;
    assign layer1_out[6730] = layer0_out[4243];
    assign layer1_out[6731] = ~(layer0_out[6088] & layer0_out[6089]);
    assign layer1_out[6732] = layer0_out[6469];
    assign layer1_out[6733] = ~layer0_out[697] | layer0_out[696];
    assign layer1_out[6734] = layer0_out[4655] ^ layer0_out[4656];
    assign layer1_out[6735] = layer0_out[4956];
    assign layer1_out[6736] = layer0_out[1261];
    assign layer1_out[6737] = layer0_out[4860] & layer0_out[4861];
    assign layer1_out[6738] = layer0_out[6823] | layer0_out[6824];
    assign layer1_out[6739] = layer0_out[5939] & layer0_out[5940];
    assign layer1_out[6740] = 1'b1;
    assign layer1_out[6741] = ~layer0_out[5405] | layer0_out[5404];
    assign layer1_out[6742] = ~(layer0_out[2872] ^ layer0_out[2873]);
    assign layer1_out[6743] = ~layer0_out[5526];
    assign layer1_out[6744] = 1'b1;
    assign layer1_out[6745] = 1'b1;
    assign layer1_out[6746] = layer0_out[6916] | layer0_out[6917];
    assign layer1_out[6747] = layer0_out[4178];
    assign layer1_out[6748] = ~layer0_out[5347] | layer0_out[5348];
    assign layer1_out[6749] = ~layer0_out[6759] | layer0_out[6760];
    assign layer1_out[6750] = layer0_out[2092];
    assign layer1_out[6751] = layer0_out[1536] & ~layer0_out[1537];
    assign layer1_out[6752] = layer0_out[6722] | layer0_out[6723];
    assign layer1_out[6753] = ~layer0_out[4915] | layer0_out[4916];
    assign layer1_out[6754] = ~layer0_out[2008] | layer0_out[2009];
    assign layer1_out[6755] = layer0_out[7806] & ~layer0_out[7807];
    assign layer1_out[6756] = ~(layer0_out[1074] & layer0_out[1075]);
    assign layer1_out[6757] = ~layer0_out[2542] | layer0_out[2543];
    assign layer1_out[6758] = layer0_out[4794] & ~layer0_out[4795];
    assign layer1_out[6759] = ~layer0_out[4261] | layer0_out[4262];
    assign layer1_out[6760] = ~layer0_out[3297];
    assign layer1_out[6761] = 1'b1;
    assign layer1_out[6762] = layer0_out[3770] | layer0_out[3771];
    assign layer1_out[6763] = ~layer0_out[2725];
    assign layer1_out[6764] = layer0_out[4114] & layer0_out[4115];
    assign layer1_out[6765] = layer0_out[2243] ^ layer0_out[2244];
    assign layer1_out[6766] = layer0_out[4906];
    assign layer1_out[6767] = 1'b1;
    assign layer1_out[6768] = ~layer0_out[7838];
    assign layer1_out[6769] = ~layer0_out[2665];
    assign layer1_out[6770] = ~(layer0_out[2424] & layer0_out[2425]);
    assign layer1_out[6771] = layer0_out[4991] & ~layer0_out[4992];
    assign layer1_out[6772] = ~layer0_out[5968] | layer0_out[5967];
    assign layer1_out[6773] = ~(layer0_out[5775] ^ layer0_out[5776]);
    assign layer1_out[6774] = ~layer0_out[2554];
    assign layer1_out[6775] = layer0_out[4400] & ~layer0_out[4401];
    assign layer1_out[6776] = ~layer0_out[7934];
    assign layer1_out[6777] = layer0_out[3682] & layer0_out[3683];
    assign layer1_out[6778] = ~layer0_out[2999];
    assign layer1_out[6779] = layer0_out[3600];
    assign layer1_out[6780] = layer0_out[4183] & layer0_out[4184];
    assign layer1_out[6781] = ~layer0_out[1033] | layer0_out[1032];
    assign layer1_out[6782] = layer0_out[1190] & ~layer0_out[1191];
    assign layer1_out[6783] = ~(layer0_out[6002] ^ layer0_out[6003]);
    assign layer1_out[6784] = layer0_out[1205];
    assign layer1_out[6785] = layer0_out[6472];
    assign layer1_out[6786] = ~(layer0_out[7516] ^ layer0_out[7517]);
    assign layer1_out[6787] = layer0_out[3179] | layer0_out[3180];
    assign layer1_out[6788] = ~(layer0_out[533] | layer0_out[534]);
    assign layer1_out[6789] = 1'b0;
    assign layer1_out[6790] = layer0_out[5412];
    assign layer1_out[6791] = ~(layer0_out[3199] | layer0_out[3200]);
    assign layer1_out[6792] = layer0_out[7549];
    assign layer1_out[6793] = layer0_out[5318];
    assign layer1_out[6794] = layer0_out[7978];
    assign layer1_out[6795] = ~(layer0_out[6702] ^ layer0_out[6703]);
    assign layer1_out[6796] = 1'b1;
    assign layer1_out[6797] = ~(layer0_out[317] & layer0_out[318]);
    assign layer1_out[6798] = ~(layer0_out[5367] ^ layer0_out[5368]);
    assign layer1_out[6799] = ~layer0_out[5345];
    assign layer1_out[6800] = 1'b0;
    assign layer1_out[6801] = layer0_out[3248];
    assign layer1_out[6802] = ~layer0_out[1778];
    assign layer1_out[6803] = ~layer0_out[7257];
    assign layer1_out[6804] = layer0_out[7128] | layer0_out[7129];
    assign layer1_out[6805] = ~layer0_out[2695] | layer0_out[2694];
    assign layer1_out[6806] = ~layer0_out[3926] | layer0_out[3925];
    assign layer1_out[6807] = ~layer0_out[193] | layer0_out[194];
    assign layer1_out[6808] = ~layer0_out[2080] | layer0_out[2079];
    assign layer1_out[6809] = layer0_out[3129] & ~layer0_out[3130];
    assign layer1_out[6810] = 1'b1;
    assign layer1_out[6811] = layer0_out[6846] & ~layer0_out[6845];
    assign layer1_out[6812] = ~(layer0_out[1000] ^ layer0_out[1001]);
    assign layer1_out[6813] = ~layer0_out[2332];
    assign layer1_out[6814] = ~layer0_out[5865];
    assign layer1_out[6815] = layer0_out[3235] & ~layer0_out[3236];
    assign layer1_out[6816] = ~layer0_out[7034] | layer0_out[7035];
    assign layer1_out[6817] = layer0_out[5191] & ~layer0_out[5192];
    assign layer1_out[6818] = layer0_out[694];
    assign layer1_out[6819] = ~layer0_out[1994] | layer0_out[1993];
    assign layer1_out[6820] = ~layer0_out[4882] | layer0_out[4881];
    assign layer1_out[6821] = ~(layer0_out[5550] & layer0_out[5551]);
    assign layer1_out[6822] = layer0_out[4379] & layer0_out[4380];
    assign layer1_out[6823] = ~(layer0_out[2187] & layer0_out[2188]);
    assign layer1_out[6824] = layer0_out[4496] ^ layer0_out[4497];
    assign layer1_out[6825] = ~layer0_out[229];
    assign layer1_out[6826] = layer0_out[5614];
    assign layer1_out[6827] = layer0_out[4426] & ~layer0_out[4425];
    assign layer1_out[6828] = layer0_out[7329];
    assign layer1_out[6829] = ~layer0_out[6705] | layer0_out[6704];
    assign layer1_out[6830] = ~layer0_out[6141] | layer0_out[6140];
    assign layer1_out[6831] = layer0_out[2617] & ~layer0_out[2616];
    assign layer1_out[6832] = layer0_out[6785] & layer0_out[6786];
    assign layer1_out[6833] = ~(layer0_out[5021] | layer0_out[5022]);
    assign layer1_out[6834] = layer0_out[1155];
    assign layer1_out[6835] = layer0_out[3734] & ~layer0_out[3735];
    assign layer1_out[6836] = ~layer0_out[294];
    assign layer1_out[6837] = layer0_out[1797] & layer0_out[1798];
    assign layer1_out[6838] = layer0_out[4206] & ~layer0_out[4207];
    assign layer1_out[6839] = layer0_out[518];
    assign layer1_out[6840] = ~layer0_out[5726];
    assign layer1_out[6841] = ~layer0_out[2656];
    assign layer1_out[6842] = layer0_out[5744] ^ layer0_out[5745];
    assign layer1_out[6843] = layer0_out[7672];
    assign layer1_out[6844] = layer0_out[4266] | layer0_out[4267];
    assign layer1_out[6845] = layer0_out[2802] ^ layer0_out[2803];
    assign layer1_out[6846] = ~layer0_out[3784];
    assign layer1_out[6847] = ~(layer0_out[7496] & layer0_out[7497]);
    assign layer1_out[6848] = ~(layer0_out[5321] & layer0_out[5322]);
    assign layer1_out[6849] = ~(layer0_out[1178] ^ layer0_out[1179]);
    assign layer1_out[6850] = layer0_out[366];
    assign layer1_out[6851] = ~layer0_out[2851];
    assign layer1_out[6852] = layer0_out[3944];
    assign layer1_out[6853] = layer0_out[5685] | layer0_out[5686];
    assign layer1_out[6854] = layer0_out[5288] | layer0_out[5289];
    assign layer1_out[6855] = layer0_out[4828];
    assign layer1_out[6856] = layer0_out[818] & ~layer0_out[817];
    assign layer1_out[6857] = layer0_out[1408];
    assign layer1_out[6858] = ~(layer0_out[6548] & layer0_out[6549]);
    assign layer1_out[6859] = layer0_out[7776] & layer0_out[7777];
    assign layer1_out[6860] = 1'b1;
    assign layer1_out[6861] = layer0_out[5264] & ~layer0_out[5265];
    assign layer1_out[6862] = ~(layer0_out[5741] & layer0_out[5742]);
    assign layer1_out[6863] = layer0_out[1835] | layer0_out[1836];
    assign layer1_out[6864] = 1'b0;
    assign layer1_out[6865] = layer0_out[5128] | layer0_out[5129];
    assign layer1_out[6866] = ~(layer0_out[191] & layer0_out[192]);
    assign layer1_out[6867] = layer0_out[985] & ~layer0_out[986];
    assign layer1_out[6868] = layer0_out[2433] & layer0_out[2434];
    assign layer1_out[6869] = layer0_out[3737] & ~layer0_out[3738];
    assign layer1_out[6870] = ~layer0_out[4852];
    assign layer1_out[6871] = ~layer0_out[5529] | layer0_out[5530];
    assign layer1_out[6872] = ~layer0_out[4923];
    assign layer1_out[6873] = layer0_out[287] & ~layer0_out[288];
    assign layer1_out[6874] = ~layer0_out[146];
    assign layer1_out[6875] = ~layer0_out[391] | layer0_out[390];
    assign layer1_out[6876] = ~layer0_out[136];
    assign layer1_out[6877] = layer0_out[1252] & ~layer0_out[1251];
    assign layer1_out[6878] = ~(layer0_out[1080] ^ layer0_out[1081]);
    assign layer1_out[6879] = layer0_out[5460];
    assign layer1_out[6880] = layer0_out[962] ^ layer0_out[963];
    assign layer1_out[6881] = layer0_out[5728] & layer0_out[5729];
    assign layer1_out[6882] = ~layer0_out[3149] | layer0_out[3148];
    assign layer1_out[6883] = layer0_out[1195] ^ layer0_out[1196];
    assign layer1_out[6884] = layer0_out[3803];
    assign layer1_out[6885] = ~layer0_out[1714];
    assign layer1_out[6886] = ~(layer0_out[3529] | layer0_out[3530]);
    assign layer1_out[6887] = layer0_out[2904] | layer0_out[2905];
    assign layer1_out[6888] = layer0_out[4602] & layer0_out[4603];
    assign layer1_out[6889] = layer0_out[2260] & layer0_out[2261];
    assign layer1_out[6890] = ~layer0_out[1149];
    assign layer1_out[6891] = ~(layer0_out[999] | layer0_out[1000]);
    assign layer1_out[6892] = layer0_out[928];
    assign layer1_out[6893] = ~layer0_out[7008] | layer0_out[7009];
    assign layer1_out[6894] = ~layer0_out[4693];
    assign layer1_out[6895] = ~layer0_out[1065] | layer0_out[1064];
    assign layer1_out[6896] = ~(layer0_out[1724] ^ layer0_out[1725]);
    assign layer1_out[6897] = ~layer0_out[7033];
    assign layer1_out[6898] = layer0_out[6533] & layer0_out[6534];
    assign layer1_out[6899] = ~layer0_out[4318];
    assign layer1_out[6900] = layer0_out[4791] & ~layer0_out[4790];
    assign layer1_out[6901] = layer0_out[1301] ^ layer0_out[1302];
    assign layer1_out[6902] = layer0_out[4998] | layer0_out[4999];
    assign layer1_out[6903] = ~(layer0_out[4355] ^ layer0_out[4356]);
    assign layer1_out[6904] = ~(layer0_out[5576] & layer0_out[5577]);
    assign layer1_out[6905] = ~layer0_out[3532] | layer0_out[3531];
    assign layer1_out[6906] = ~(layer0_out[7437] | layer0_out[7438]);
    assign layer1_out[6907] = ~layer0_out[2590];
    assign layer1_out[6908] = ~(layer0_out[2873] & layer0_out[2874]);
    assign layer1_out[6909] = ~layer0_out[3746];
    assign layer1_out[6910] = 1'b1;
    assign layer1_out[6911] = layer0_out[4648];
    assign layer1_out[6912] = layer0_out[4561] & ~layer0_out[4562];
    assign layer1_out[6913] = layer0_out[3978];
    assign layer1_out[6914] = layer0_out[120];
    assign layer1_out[6915] = layer0_out[119] & ~layer0_out[118];
    assign layer1_out[6916] = layer0_out[703] & ~layer0_out[702];
    assign layer1_out[6917] = ~layer0_out[6340];
    assign layer1_out[6918] = layer0_out[2382];
    assign layer1_out[6919] = ~layer0_out[6902] | layer0_out[6903];
    assign layer1_out[6920] = ~(layer0_out[2761] | layer0_out[2762]);
    assign layer1_out[6921] = ~(layer0_out[6516] & layer0_out[6517]);
    assign layer1_out[6922] = ~(layer0_out[4386] & layer0_out[4387]);
    assign layer1_out[6923] = layer0_out[3687];
    assign layer1_out[6924] = ~layer0_out[2956] | layer0_out[2955];
    assign layer1_out[6925] = layer0_out[4342];
    assign layer1_out[6926] = ~(layer0_out[7068] ^ layer0_out[7069]);
    assign layer1_out[6927] = ~(layer0_out[957] & layer0_out[958]);
    assign layer1_out[6928] = ~layer0_out[1726];
    assign layer1_out[6929] = ~layer0_out[7542];
    assign layer1_out[6930] = ~(layer0_out[3566] | layer0_out[3567]);
    assign layer1_out[6931] = layer0_out[3596];
    assign layer1_out[6932] = ~(layer0_out[4673] ^ layer0_out[4674]);
    assign layer1_out[6933] = layer0_out[7450];
    assign layer1_out[6934] = ~layer0_out[2809] | layer0_out[2810];
    assign layer1_out[6935] = ~layer0_out[1711];
    assign layer1_out[6936] = layer0_out[6221] ^ layer0_out[6222];
    assign layer1_out[6937] = 1'b0;
    assign layer1_out[6938] = ~(layer0_out[2923] | layer0_out[2924]);
    assign layer1_out[6939] = layer0_out[4958] & ~layer0_out[4957];
    assign layer1_out[6940] = ~layer0_out[5756] | layer0_out[5755];
    assign layer1_out[6941] = ~(layer0_out[5233] ^ layer0_out[5234]);
    assign layer1_out[6942] = layer0_out[6286] & layer0_out[6287];
    assign layer1_out[6943] = layer0_out[1509];
    assign layer1_out[6944] = ~(layer0_out[5844] | layer0_out[5845]);
    assign layer1_out[6945] = ~(layer0_out[411] | layer0_out[412]);
    assign layer1_out[6946] = ~layer0_out[2786] | layer0_out[2785];
    assign layer1_out[6947] = 1'b1;
    assign layer1_out[6948] = ~layer0_out[5630];
    assign layer1_out[6949] = layer0_out[4399] ^ layer0_out[4400];
    assign layer1_out[6950] = ~layer0_out[5622] | layer0_out[5623];
    assign layer1_out[6951] = layer0_out[5863] & layer0_out[5864];
    assign layer1_out[6952] = ~layer0_out[2793];
    assign layer1_out[6953] = ~layer0_out[5428] | layer0_out[5427];
    assign layer1_out[6954] = ~layer0_out[2906] | layer0_out[2905];
    assign layer1_out[6955] = layer0_out[4654];
    assign layer1_out[6956] = 1'b0;
    assign layer1_out[6957] = layer0_out[4606] ^ layer0_out[4607];
    assign layer1_out[6958] = layer0_out[3820] & ~layer0_out[3821];
    assign layer1_out[6959] = ~(layer0_out[5273] | layer0_out[5274]);
    assign layer1_out[6960] = layer0_out[5366] & ~layer0_out[5367];
    assign layer1_out[6961] = layer0_out[4769] & ~layer0_out[4768];
    assign layer1_out[6962] = ~layer0_out[3912] | layer0_out[3911];
    assign layer1_out[6963] = 1'b1;
    assign layer1_out[6964] = layer0_out[5469] ^ layer0_out[5470];
    assign layer1_out[6965] = 1'b1;
    assign layer1_out[6966] = layer0_out[4276] | layer0_out[4277];
    assign layer1_out[6967] = ~(layer0_out[1429] ^ layer0_out[1430]);
    assign layer1_out[6968] = ~(layer0_out[4349] & layer0_out[4350]);
    assign layer1_out[6969] = layer0_out[876];
    assign layer1_out[6970] = layer0_out[419] & ~layer0_out[420];
    assign layer1_out[6971] = ~layer0_out[2222];
    assign layer1_out[6972] = layer0_out[1518];
    assign layer1_out[6973] = layer0_out[6196];
    assign layer1_out[6974] = layer0_out[2863];
    assign layer1_out[6975] = ~layer0_out[7923];
    assign layer1_out[6976] = ~(layer0_out[7988] | layer0_out[7989]);
    assign layer1_out[6977] = ~layer0_out[2188] | layer0_out[2189];
    assign layer1_out[6978] = ~layer0_out[260] | layer0_out[261];
    assign layer1_out[6979] = ~layer0_out[1696];
    assign layer1_out[6980] = layer0_out[7820] & ~layer0_out[7819];
    assign layer1_out[6981] = ~layer0_out[3134];
    assign layer1_out[6982] = ~layer0_out[5330] | layer0_out[5329];
    assign layer1_out[6983] = layer0_out[3492];
    assign layer1_out[6984] = layer0_out[6800] ^ layer0_out[6801];
    assign layer1_out[6985] = layer0_out[7656] & ~layer0_out[7655];
    assign layer1_out[6986] = layer0_out[7254] & layer0_out[7255];
    assign layer1_out[6987] = ~layer0_out[1956];
    assign layer1_out[6988] = layer0_out[5020] | layer0_out[5021];
    assign layer1_out[6989] = layer0_out[6406] & ~layer0_out[6405];
    assign layer1_out[6990] = layer0_out[5821] | layer0_out[5822];
    assign layer1_out[6991] = ~layer0_out[4098];
    assign layer1_out[6992] = layer0_out[7662] ^ layer0_out[7663];
    assign layer1_out[6993] = ~layer0_out[1390] | layer0_out[1391];
    assign layer1_out[6994] = ~layer0_out[7058];
    assign layer1_out[6995] = layer0_out[208] & ~layer0_out[207];
    assign layer1_out[6996] = ~layer0_out[3924];
    assign layer1_out[6997] = layer0_out[817];
    assign layer1_out[6998] = ~layer0_out[206];
    assign layer1_out[6999] = ~(layer0_out[3262] & layer0_out[3263]);
    assign layer1_out[7000] = ~(layer0_out[4369] | layer0_out[4370]);
    assign layer1_out[7001] = ~layer0_out[4202];
    assign layer1_out[7002] = layer0_out[4249];
    assign layer1_out[7003] = layer0_out[2297] & layer0_out[2298];
    assign layer1_out[7004] = layer0_out[3255];
    assign layer1_out[7005] = layer0_out[6756] & ~layer0_out[6755];
    assign layer1_out[7006] = ~(layer0_out[1287] | layer0_out[1288]);
    assign layer1_out[7007] = ~(layer0_out[14] & layer0_out[15]);
    assign layer1_out[7008] = ~layer0_out[5482];
    assign layer1_out[7009] = layer0_out[3948];
    assign layer1_out[7010] = layer0_out[4348] & ~layer0_out[4347];
    assign layer1_out[7011] = layer0_out[3166] & layer0_out[3167];
    assign layer1_out[7012] = ~layer0_out[3035];
    assign layer1_out[7013] = layer0_out[4053];
    assign layer1_out[7014] = layer0_out[6869];
    assign layer1_out[7015] = ~layer0_out[5900];
    assign layer1_out[7016] = ~layer0_out[2100];
    assign layer1_out[7017] = ~layer0_out[1509] | layer0_out[1510];
    assign layer1_out[7018] = ~layer0_out[5862];
    assign layer1_out[7019] = ~layer0_out[5013] | layer0_out[5014];
    assign layer1_out[7020] = layer0_out[4666] | layer0_out[4667];
    assign layer1_out[7021] = 1'b0;
    assign layer1_out[7022] = layer0_out[513];
    assign layer1_out[7023] = layer0_out[2792];
    assign layer1_out[7024] = layer0_out[2686];
    assign layer1_out[7025] = ~layer0_out[7508] | layer0_out[7509];
    assign layer1_out[7026] = ~layer0_out[4171] | layer0_out[4170];
    assign layer1_out[7027] = layer0_out[2952];
    assign layer1_out[7028] = layer0_out[4079];
    assign layer1_out[7029] = ~layer0_out[1010] | layer0_out[1011];
    assign layer1_out[7030] = ~(layer0_out[2395] & layer0_out[2396]);
    assign layer1_out[7031] = ~layer0_out[2572] | layer0_out[2571];
    assign layer1_out[7032] = ~layer0_out[7265];
    assign layer1_out[7033] = ~(layer0_out[4416] | layer0_out[4417]);
    assign layer1_out[7034] = ~(layer0_out[7706] & layer0_out[7707]);
    assign layer1_out[7035] = layer0_out[5561] & ~layer0_out[5562];
    assign layer1_out[7036] = layer0_out[1083] & ~layer0_out[1082];
    assign layer1_out[7037] = ~layer0_out[5311];
    assign layer1_out[7038] = ~(layer0_out[538] & layer0_out[539]);
    assign layer1_out[7039] = ~layer0_out[2814] | layer0_out[2815];
    assign layer1_out[7040] = ~(layer0_out[3136] ^ layer0_out[3137]);
    assign layer1_out[7041] = ~(layer0_out[1028] | layer0_out[1029]);
    assign layer1_out[7042] = ~(layer0_out[4940] | layer0_out[4941]);
    assign layer1_out[7043] = layer0_out[7028] & ~layer0_out[7029];
    assign layer1_out[7044] = layer0_out[2875];
    assign layer1_out[7045] = layer0_out[2061] ^ layer0_out[2062];
    assign layer1_out[7046] = ~(layer0_out[5153] & layer0_out[5154]);
    assign layer1_out[7047] = ~(layer0_out[7035] | layer0_out[7036]);
    assign layer1_out[7048] = ~layer0_out[7218];
    assign layer1_out[7049] = ~layer0_out[7270] | layer0_out[7269];
    assign layer1_out[7050] = ~(layer0_out[1269] | layer0_out[1270]);
    assign layer1_out[7051] = ~(layer0_out[1085] & layer0_out[1086]);
    assign layer1_out[7052] = ~layer0_out[3661];
    assign layer1_out[7053] = ~layer0_out[1218] | layer0_out[1219];
    assign layer1_out[7054] = ~(layer0_out[4688] | layer0_out[4689]);
    assign layer1_out[7055] = layer0_out[6680];
    assign layer1_out[7056] = ~(layer0_out[4595] | layer0_out[4596]);
    assign layer1_out[7057] = layer0_out[6540] & ~layer0_out[6539];
    assign layer1_out[7058] = ~(layer0_out[6891] ^ layer0_out[6892]);
    assign layer1_out[7059] = layer0_out[7657];
    assign layer1_out[7060] = ~layer0_out[6462] | layer0_out[6463];
    assign layer1_out[7061] = ~layer0_out[5648];
    assign layer1_out[7062] = ~(layer0_out[937] | layer0_out[938]);
    assign layer1_out[7063] = 1'b1;
    assign layer1_out[7064] = 1'b0;
    assign layer1_out[7065] = layer0_out[6581] | layer0_out[6582];
    assign layer1_out[7066] = layer0_out[1839] & ~layer0_out[1840];
    assign layer1_out[7067] = ~layer0_out[6043] | layer0_out[6044];
    assign layer1_out[7068] = ~(layer0_out[3932] | layer0_out[3933]);
    assign layer1_out[7069] = ~(layer0_out[1811] ^ layer0_out[1812]);
    assign layer1_out[7070] = ~(layer0_out[4338] | layer0_out[4339]);
    assign layer1_out[7071] = ~layer0_out[4276] | layer0_out[4275];
    assign layer1_out[7072] = 1'b0;
    assign layer1_out[7073] = ~layer0_out[4502];
    assign layer1_out[7074] = ~layer0_out[3974];
    assign layer1_out[7075] = layer0_out[507] & ~layer0_out[506];
    assign layer1_out[7076] = ~(layer0_out[5572] & layer0_out[5573]);
    assign layer1_out[7077] = 1'b0;
    assign layer1_out[7078] = ~layer0_out[313] | layer0_out[314];
    assign layer1_out[7079] = layer0_out[1938] & layer0_out[1939];
    assign layer1_out[7080] = layer0_out[6146] & ~layer0_out[6147];
    assign layer1_out[7081] = ~layer0_out[2534] | layer0_out[2533];
    assign layer1_out[7082] = layer0_out[7617] & ~layer0_out[7618];
    assign layer1_out[7083] = layer0_out[1179] & ~layer0_out[1180];
    assign layer1_out[7084] = layer0_out[4296] | layer0_out[4297];
    assign layer1_out[7085] = ~layer0_out[4651];
    assign layer1_out[7086] = layer0_out[123] & layer0_out[124];
    assign layer1_out[7087] = ~layer0_out[33];
    assign layer1_out[7088] = ~layer0_out[3187] | layer0_out[3188];
    assign layer1_out[7089] = ~(layer0_out[2954] | layer0_out[2955]);
    assign layer1_out[7090] = ~layer0_out[4251] | layer0_out[4252];
    assign layer1_out[7091] = ~layer0_out[1288] | layer0_out[1289];
    assign layer1_out[7092] = 1'b1;
    assign layer1_out[7093] = ~(layer0_out[6719] ^ layer0_out[6720]);
    assign layer1_out[7094] = ~(layer0_out[3746] | layer0_out[3747]);
    assign layer1_out[7095] = ~layer0_out[5090];
    assign layer1_out[7096] = ~(layer0_out[5815] | layer0_out[5816]);
    assign layer1_out[7097] = ~(layer0_out[7675] ^ layer0_out[7676]);
    assign layer1_out[7098] = layer0_out[1514] & ~layer0_out[1513];
    assign layer1_out[7099] = ~(layer0_out[4652] | layer0_out[4653]);
    assign layer1_out[7100] = ~layer0_out[4728];
    assign layer1_out[7101] = ~(layer0_out[4640] ^ layer0_out[4641]);
    assign layer1_out[7102] = layer0_out[3527] | layer0_out[3528];
    assign layer1_out[7103] = layer0_out[4378];
    assign layer1_out[7104] = layer0_out[3394] | layer0_out[3395];
    assign layer1_out[7105] = ~layer0_out[2137];
    assign layer1_out[7106] = ~layer0_out[1368];
    assign layer1_out[7107] = ~layer0_out[2004];
    assign layer1_out[7108] = ~(layer0_out[3236] | layer0_out[3237]);
    assign layer1_out[7109] = layer0_out[5805] & ~layer0_out[5804];
    assign layer1_out[7110] = ~layer0_out[3880] | layer0_out[3881];
    assign layer1_out[7111] = ~layer0_out[1663];
    assign layer1_out[7112] = ~layer0_out[3293];
    assign layer1_out[7113] = ~layer0_out[5030] | layer0_out[5029];
    assign layer1_out[7114] = layer0_out[2487] & ~layer0_out[2488];
    assign layer1_out[7115] = ~layer0_out[6015] | layer0_out[6014];
    assign layer1_out[7116] = 1'b1;
    assign layer1_out[7117] = ~layer0_out[6090];
    assign layer1_out[7118] = ~(layer0_out[896] & layer0_out[897]);
    assign layer1_out[7119] = ~(layer0_out[343] | layer0_out[344]);
    assign layer1_out[7120] = layer0_out[6098] & ~layer0_out[6097];
    assign layer1_out[7121] = layer0_out[6437] & ~layer0_out[6436];
    assign layer1_out[7122] = 1'b0;
    assign layer1_out[7123] = layer0_out[6738];
    assign layer1_out[7124] = ~layer0_out[5434] | layer0_out[5433];
    assign layer1_out[7125] = ~layer0_out[6232] | layer0_out[6233];
    assign layer1_out[7126] = ~layer0_out[829] | layer0_out[830];
    assign layer1_out[7127] = ~(layer0_out[3637] | layer0_out[3638]);
    assign layer1_out[7128] = ~layer0_out[5011];
    assign layer1_out[7129] = layer0_out[3006];
    assign layer1_out[7130] = layer0_out[800];
    assign layer1_out[7131] = layer0_out[5691] ^ layer0_out[5692];
    assign layer1_out[7132] = ~layer0_out[244] | layer0_out[245];
    assign layer1_out[7133] = ~layer0_out[617] | layer0_out[618];
    assign layer1_out[7134] = layer0_out[7523] ^ layer0_out[7524];
    assign layer1_out[7135] = layer0_out[2231];
    assign layer1_out[7136] = layer0_out[4099] & ~layer0_out[4100];
    assign layer1_out[7137] = ~layer0_out[2034];
    assign layer1_out[7138] = ~(layer0_out[2953] & layer0_out[2954]);
    assign layer1_out[7139] = ~layer0_out[7384];
    assign layer1_out[7140] = ~(layer0_out[1751] | layer0_out[1752]);
    assign layer1_out[7141] = layer0_out[2214] & layer0_out[2215];
    assign layer1_out[7142] = ~layer0_out[649];
    assign layer1_out[7143] = layer0_out[4257];
    assign layer1_out[7144] = layer0_out[5277] & ~layer0_out[5276];
    assign layer1_out[7145] = ~layer0_out[62];
    assign layer1_out[7146] = layer0_out[624] | layer0_out[625];
    assign layer1_out[7147] = layer0_out[2480] & ~layer0_out[2481];
    assign layer1_out[7148] = ~layer0_out[4328] | layer0_out[4327];
    assign layer1_out[7149] = layer0_out[7191];
    assign layer1_out[7150] = 1'b0;
    assign layer1_out[7151] = layer0_out[7518];
    assign layer1_out[7152] = layer0_out[1814] | layer0_out[1815];
    assign layer1_out[7153] = layer0_out[7119] ^ layer0_out[7120];
    assign layer1_out[7154] = ~(layer0_out[5086] ^ layer0_out[5087]);
    assign layer1_out[7155] = layer0_out[4639] & layer0_out[4640];
    assign layer1_out[7156] = ~layer0_out[7133] | layer0_out[7132];
    assign layer1_out[7157] = layer0_out[590] & layer0_out[591];
    assign layer1_out[7158] = ~layer0_out[6231] | layer0_out[6230];
    assign layer1_out[7159] = ~layer0_out[5972];
    assign layer1_out[7160] = ~(layer0_out[2693] & layer0_out[2694]);
    assign layer1_out[7161] = layer0_out[2131] & layer0_out[2132];
    assign layer1_out[7162] = ~layer0_out[6872] | layer0_out[6871];
    assign layer1_out[7163] = ~layer0_out[3905] | layer0_out[3906];
    assign layer1_out[7164] = ~layer0_out[3171] | layer0_out[3172];
    assign layer1_out[7165] = ~(layer0_out[7529] & layer0_out[7530]);
    assign layer1_out[7166] = layer0_out[936] & layer0_out[937];
    assign layer1_out[7167] = layer0_out[416];
    assign layer1_out[7168] = layer0_out[3064];
    assign layer1_out[7169] = ~layer0_out[6698] | layer0_out[6697];
    assign layer1_out[7170] = ~(layer0_out[4568] & layer0_out[4569]);
    assign layer1_out[7171] = ~(layer0_out[6686] ^ layer0_out[6687]);
    assign layer1_out[7172] = layer0_out[7003];
    assign layer1_out[7173] = layer0_out[6440] & layer0_out[6441];
    assign layer1_out[7174] = ~(layer0_out[3381] & layer0_out[3382]);
    assign layer1_out[7175] = ~(layer0_out[4330] | layer0_out[4331]);
    assign layer1_out[7176] = ~(layer0_out[6934] | layer0_out[6935]);
    assign layer1_out[7177] = ~layer0_out[2461];
    assign layer1_out[7178] = ~layer0_out[6638];
    assign layer1_out[7179] = 1'b0;
    assign layer1_out[7180] = layer0_out[1350] & layer0_out[1351];
    assign layer1_out[7181] = layer0_out[6223] | layer0_out[6224];
    assign layer1_out[7182] = 1'b0;
    assign layer1_out[7183] = ~layer0_out[6156] | layer0_out[6157];
    assign layer1_out[7184] = ~(layer0_out[655] & layer0_out[656]);
    assign layer1_out[7185] = layer0_out[4234] ^ layer0_out[4235];
    assign layer1_out[7186] = ~layer0_out[4994] | layer0_out[4995];
    assign layer1_out[7187] = layer0_out[493];
    assign layer1_out[7188] = ~layer0_out[3719];
    assign layer1_out[7189] = ~layer0_out[712];
    assign layer1_out[7190] = layer0_out[6779];
    assign layer1_out[7191] = layer0_out[4951];
    assign layer1_out[7192] = 1'b1;
    assign layer1_out[7193] = ~(layer0_out[2517] ^ layer0_out[2518]);
    assign layer1_out[7194] = ~layer0_out[7836];
    assign layer1_out[7195] = layer0_out[7797];
    assign layer1_out[7196] = ~(layer0_out[7649] | layer0_out[7650]);
    assign layer1_out[7197] = ~layer0_out[3520];
    assign layer1_out[7198] = layer0_out[5234] | layer0_out[5235];
    assign layer1_out[7199] = ~(layer0_out[7141] | layer0_out[7142]);
    assign layer1_out[7200] = layer0_out[1759] ^ layer0_out[1760];
    assign layer1_out[7201] = layer0_out[5682] | layer0_out[5683];
    assign layer1_out[7202] = layer0_out[6948] & ~layer0_out[6947];
    assign layer1_out[7203] = layer0_out[5429] & ~layer0_out[5430];
    assign layer1_out[7204] = ~(layer0_out[1765] | layer0_out[1766]);
    assign layer1_out[7205] = layer0_out[431] & ~layer0_out[430];
    assign layer1_out[7206] = layer0_out[54] & ~layer0_out[53];
    assign layer1_out[7207] = ~layer0_out[7206];
    assign layer1_out[7208] = layer0_out[5301];
    assign layer1_out[7209] = layer0_out[5901] | layer0_out[5902];
    assign layer1_out[7210] = ~layer0_out[4522] | layer0_out[4521];
    assign layer1_out[7211] = ~layer0_out[7826] | layer0_out[7825];
    assign layer1_out[7212] = layer0_out[5620];
    assign layer1_out[7213] = layer0_out[1934];
    assign layer1_out[7214] = layer0_out[6701] & ~layer0_out[6702];
    assign layer1_out[7215] = layer0_out[6583] ^ layer0_out[6584];
    assign layer1_out[7216] = ~(layer0_out[3834] | layer0_out[3835]);
    assign layer1_out[7217] = layer0_out[3259] | layer0_out[3260];
    assign layer1_out[7218] = ~(layer0_out[368] & layer0_out[369]);
    assign layer1_out[7219] = layer0_out[3356] & layer0_out[3357];
    assign layer1_out[7220] = ~(layer0_out[2906] & layer0_out[2907]);
    assign layer1_out[7221] = ~layer0_out[3195];
    assign layer1_out[7222] = layer0_out[708] & ~layer0_out[709];
    assign layer1_out[7223] = ~(layer0_out[5615] ^ layer0_out[5616]);
    assign layer1_out[7224] = layer0_out[7525] | layer0_out[7526];
    assign layer1_out[7225] = ~(layer0_out[6525] ^ layer0_out[6526]);
    assign layer1_out[7226] = ~layer0_out[779] | layer0_out[780];
    assign layer1_out[7227] = ~layer0_out[186] | layer0_out[185];
    assign layer1_out[7228] = ~(layer0_out[6992] | layer0_out[6993]);
    assign layer1_out[7229] = layer0_out[1691] & ~layer0_out[1692];
    assign layer1_out[7230] = ~(layer0_out[7886] | layer0_out[7887]);
    assign layer1_out[7231] = ~(layer0_out[7469] ^ layer0_out[7470]);
    assign layer1_out[7232] = 1'b1;
    assign layer1_out[7233] = ~layer0_out[3285] | layer0_out[3286];
    assign layer1_out[7234] = layer0_out[7413] & layer0_out[7414];
    assign layer1_out[7235] = 1'b1;
    assign layer1_out[7236] = layer0_out[675] ^ layer0_out[676];
    assign layer1_out[7237] = 1'b1;
    assign layer1_out[7238] = ~(layer0_out[1666] ^ layer0_out[1667]);
    assign layer1_out[7239] = ~layer0_out[2322];
    assign layer1_out[7240] = layer0_out[1699] & ~layer0_out[1700];
    assign layer1_out[7241] = layer0_out[1555];
    assign layer1_out[7242] = 1'b0;
    assign layer1_out[7243] = layer0_out[3540] | layer0_out[3541];
    assign layer1_out[7244] = ~(layer0_out[433] ^ layer0_out[434]);
    assign layer1_out[7245] = ~layer0_out[1525] | layer0_out[1526];
    assign layer1_out[7246] = layer0_out[716];
    assign layer1_out[7247] = layer0_out[4800];
    assign layer1_out[7248] = ~layer0_out[1722] | layer0_out[1723];
    assign layer1_out[7249] = 1'b0;
    assign layer1_out[7250] = layer0_out[1757];
    assign layer1_out[7251] = layer0_out[1293];
    assign layer1_out[7252] = ~(layer0_out[3524] | layer0_out[3525]);
    assign layer1_out[7253] = 1'b1;
    assign layer1_out[7254] = layer0_out[168] & layer0_out[169];
    assign layer1_out[7255] = layer0_out[4237] & ~layer0_out[4238];
    assign layer1_out[7256] = layer0_out[7745] ^ layer0_out[7746];
    assign layer1_out[7257] = layer0_out[5569] & ~layer0_out[5570];
    assign layer1_out[7258] = layer0_out[2558] ^ layer0_out[2559];
    assign layer1_out[7259] = ~(layer0_out[1088] | layer0_out[1089]);
    assign layer1_out[7260] = layer0_out[6942];
    assign layer1_out[7261] = 1'b0;
    assign layer1_out[7262] = ~layer0_out[2589] | layer0_out[2588];
    assign layer1_out[7263] = layer0_out[2795];
    assign layer1_out[7264] = ~layer0_out[2583] | layer0_out[2582];
    assign layer1_out[7265] = layer0_out[2354] | layer0_out[2355];
    assign layer1_out[7266] = ~(layer0_out[5800] | layer0_out[5801]);
    assign layer1_out[7267] = layer0_out[3220] & ~layer0_out[3219];
    assign layer1_out[7268] = ~layer0_out[3239];
    assign layer1_out[7269] = layer0_out[49] & ~layer0_out[50];
    assign layer1_out[7270] = layer0_out[6480] ^ layer0_out[6481];
    assign layer1_out[7271] = ~layer0_out[340] | layer0_out[341];
    assign layer1_out[7272] = ~layer0_out[6402];
    assign layer1_out[7273] = ~layer0_out[3306] | layer0_out[3305];
    assign layer1_out[7274] = layer0_out[976];
    assign layer1_out[7275] = ~layer0_out[4620];
    assign layer1_out[7276] = layer0_out[2123];
    assign layer1_out[7277] = ~layer0_out[7879];
    assign layer1_out[7278] = 1'b0;
    assign layer1_out[7279] = layer0_out[3078] ^ layer0_out[3079];
    assign layer1_out[7280] = layer0_out[7619] & layer0_out[7620];
    assign layer1_out[7281] = layer0_out[1798] & layer0_out[1799];
    assign layer1_out[7282] = layer0_out[7312];
    assign layer1_out[7283] = layer0_out[6095];
    assign layer1_out[7284] = ~layer0_out[3360] | layer0_out[3359];
    assign layer1_out[7285] = ~(layer0_out[409] ^ layer0_out[410]);
    assign layer1_out[7286] = ~layer0_out[1409] | layer0_out[1408];
    assign layer1_out[7287] = ~(layer0_out[375] & layer0_out[376]);
    assign layer1_out[7288] = ~(layer0_out[6611] | layer0_out[6612]);
    assign layer1_out[7289] = 1'b0;
    assign layer1_out[7290] = layer0_out[366] & ~layer0_out[367];
    assign layer1_out[7291] = ~layer0_out[4131] | layer0_out[4130];
    assign layer1_out[7292] = layer0_out[6214];
    assign layer1_out[7293] = layer0_out[7421];
    assign layer1_out[7294] = ~(layer0_out[6627] ^ layer0_out[6628]);
    assign layer1_out[7295] = ~(layer0_out[1746] | layer0_out[1747]);
    assign layer1_out[7296] = ~(layer0_out[4445] ^ layer0_out[4446]);
    assign layer1_out[7297] = ~layer0_out[7953];
    assign layer1_out[7298] = ~layer0_out[5599] | layer0_out[5598];
    assign layer1_out[7299] = layer0_out[7810] | layer0_out[7811];
    assign layer1_out[7300] = ~layer0_out[7593] | layer0_out[7592];
    assign layer1_out[7301] = ~(layer0_out[4454] | layer0_out[4455]);
    assign layer1_out[7302] = 1'b1;
    assign layer1_out[7303] = ~(layer0_out[699] | layer0_out[700]);
    assign layer1_out[7304] = 1'b1;
    assign layer1_out[7305] = ~(layer0_out[3704] | layer0_out[3705]);
    assign layer1_out[7306] = ~layer0_out[7735];
    assign layer1_out[7307] = layer0_out[3441] | layer0_out[3442];
    assign layer1_out[7308] = layer0_out[72];
    assign layer1_out[7309] = layer0_out[2797] ^ layer0_out[2798];
    assign layer1_out[7310] = 1'b1;
    assign layer1_out[7311] = ~layer0_out[7354];
    assign layer1_out[7312] = layer0_out[2689];
    assign layer1_out[7313] = ~layer0_out[7688] | layer0_out[7689];
    assign layer1_out[7314] = layer0_out[1107] | layer0_out[1108];
    assign layer1_out[7315] = layer0_out[6011] & ~layer0_out[6012];
    assign layer1_out[7316] = ~(layer0_out[90] & layer0_out[91]);
    assign layer1_out[7317] = layer0_out[5738];
    assign layer1_out[7318] = layer0_out[4141];
    assign layer1_out[7319] = 1'b1;
    assign layer1_out[7320] = ~layer0_out[6125];
    assign layer1_out[7321] = 1'b0;
    assign layer1_out[7322] = layer0_out[1180] ^ layer0_out[1181];
    assign layer1_out[7323] = layer0_out[4485];
    assign layer1_out[7324] = ~layer0_out[3356] | layer0_out[3355];
    assign layer1_out[7325] = ~layer0_out[6047] | layer0_out[6046];
    assign layer1_out[7326] = layer0_out[5555] & layer0_out[5556];
    assign layer1_out[7327] = ~layer0_out[1958] | layer0_out[1957];
    assign layer1_out[7328] = layer0_out[2760];
    assign layer1_out[7329] = layer0_out[3048] ^ layer0_out[3049];
    assign layer1_out[7330] = layer0_out[839];
    assign layer1_out[7331] = layer0_out[175] & ~layer0_out[176];
    assign layer1_out[7332] = ~(layer0_out[1259] ^ layer0_out[1260]);
    assign layer1_out[7333] = layer0_out[2981] & ~layer0_out[2982];
    assign layer1_out[7334] = layer0_out[6001] & layer0_out[6002];
    assign layer1_out[7335] = ~(layer0_out[7023] | layer0_out[7024]);
    assign layer1_out[7336] = ~layer0_out[1229];
    assign layer1_out[7337] = layer0_out[3225] | layer0_out[3226];
    assign layer1_out[7338] = layer0_out[5314];
    assign layer1_out[7339] = layer0_out[1586] & ~layer0_out[1585];
    assign layer1_out[7340] = layer0_out[2342];
    assign layer1_out[7341] = layer0_out[2480] & ~layer0_out[2479];
    assign layer1_out[7342] = 1'b1;
    assign layer1_out[7343] = layer0_out[1041];
    assign layer1_out[7344] = layer0_out[7920];
    assign layer1_out[7345] = 1'b0;
    assign layer1_out[7346] = layer0_out[1324] ^ layer0_out[1325];
    assign layer1_out[7347] = ~layer0_out[6192];
    assign layer1_out[7348] = ~layer0_out[4460] | layer0_out[4459];
    assign layer1_out[7349] = ~(layer0_out[257] | layer0_out[258]);
    assign layer1_out[7350] = layer0_out[2274] & ~layer0_out[2273];
    assign layer1_out[7351] = layer0_out[6865] | layer0_out[6866];
    assign layer1_out[7352] = layer0_out[5121] ^ layer0_out[5122];
    assign layer1_out[7353] = ~layer0_out[6161];
    assign layer1_out[7354] = 1'b0;
    assign layer1_out[7355] = ~(layer0_out[3931] & layer0_out[3932]);
    assign layer1_out[7356] = layer0_out[7645] & ~layer0_out[7644];
    assign layer1_out[7357] = ~layer0_out[3490];
    assign layer1_out[7358] = 1'b1;
    assign layer1_out[7359] = layer0_out[6179] & layer0_out[6180];
    assign layer1_out[7360] = 1'b1;
    assign layer1_out[7361] = layer0_out[3279] | layer0_out[3280];
    assign layer1_out[7362] = 1'b1;
    assign layer1_out[7363] = layer0_out[7900];
    assign layer1_out[7364] = layer0_out[4650] & ~layer0_out[4649];
    assign layer1_out[7365] = layer0_out[2077];
    assign layer1_out[7366] = ~(layer0_out[7532] ^ layer0_out[7533]);
    assign layer1_out[7367] = layer0_out[3062];
    assign layer1_out[7368] = ~(layer0_out[5168] ^ layer0_out[5169]);
    assign layer1_out[7369] = ~layer0_out[2865];
    assign layer1_out[7370] = ~layer0_out[743];
    assign layer1_out[7371] = ~layer0_out[4775];
    assign layer1_out[7372] = layer0_out[1336];
    assign layer1_out[7373] = ~(layer0_out[5709] | layer0_out[5710]);
    assign layer1_out[7374] = ~layer0_out[5601] | layer0_out[5600];
    assign layer1_out[7375] = ~layer0_out[23];
    assign layer1_out[7376] = layer0_out[249] & ~layer0_out[248];
    assign layer1_out[7377] = ~layer0_out[3954] | layer0_out[3953];
    assign layer1_out[7378] = layer0_out[3853] | layer0_out[3854];
    assign layer1_out[7379] = ~layer0_out[7098] | layer0_out[7099];
    assign layer1_out[7380] = ~(layer0_out[6441] ^ layer0_out[6442]);
    assign layer1_out[7381] = layer0_out[5649];
    assign layer1_out[7382] = 1'b0;
    assign layer1_out[7383] = layer0_out[3506] | layer0_out[3507];
    assign layer1_out[7384] = ~(layer0_out[5952] & layer0_out[5953]);
    assign layer1_out[7385] = layer0_out[4610];
    assign layer1_out[7386] = layer0_out[5836] ^ layer0_out[5837];
    assign layer1_out[7387] = ~layer0_out[1926] | layer0_out[1927];
    assign layer1_out[7388] = ~(layer0_out[3855] | layer0_out[3856]);
    assign layer1_out[7389] = layer0_out[2625];
    assign layer1_out[7390] = ~layer0_out[4669] | layer0_out[4668];
    assign layer1_out[7391] = ~layer0_out[4701];
    assign layer1_out[7392] = ~layer0_out[2738] | layer0_out[2737];
    assign layer1_out[7393] = layer0_out[2135] & ~layer0_out[2134];
    assign layer1_out[7394] = layer0_out[7796] & layer0_out[7797];
    assign layer1_out[7395] = layer0_out[4892] & ~layer0_out[4893];
    assign layer1_out[7396] = ~layer0_out[3399];
    assign layer1_out[7397] = ~(layer0_out[4904] | layer0_out[4905]);
    assign layer1_out[7398] = layer0_out[3412] & ~layer0_out[3411];
    assign layer1_out[7399] = 1'b1;
    assign layer1_out[7400] = layer0_out[530];
    assign layer1_out[7401] = layer0_out[716] & ~layer0_out[715];
    assign layer1_out[7402] = 1'b1;
    assign layer1_out[7403] = layer0_out[4829];
    assign layer1_out[7404] = ~layer0_out[3222];
    assign layer1_out[7405] = ~layer0_out[201];
    assign layer1_out[7406] = layer0_out[6595] & layer0_out[6596];
    assign layer1_out[7407] = layer0_out[756] & ~layer0_out[755];
    assign layer1_out[7408] = ~layer0_out[6278];
    assign layer1_out[7409] = layer0_out[4399] & ~layer0_out[4398];
    assign layer1_out[7410] = ~(layer0_out[468] ^ layer0_out[469]);
    assign layer1_out[7411] = layer0_out[5120] & ~layer0_out[5121];
    assign layer1_out[7412] = 1'b1;
    assign layer1_out[7413] = layer0_out[1418] & layer0_out[1419];
    assign layer1_out[7414] = layer0_out[3961] ^ layer0_out[3962];
    assign layer1_out[7415] = ~layer0_out[2667];
    assign layer1_out[7416] = layer0_out[1092] & ~layer0_out[1091];
    assign layer1_out[7417] = ~layer0_out[402];
    assign layer1_out[7418] = ~(layer0_out[4498] | layer0_out[4499]);
    assign layer1_out[7419] = ~layer0_out[7791];
    assign layer1_out[7420] = ~(layer0_out[6315] | layer0_out[6316]);
    assign layer1_out[7421] = layer0_out[1551] | layer0_out[1552];
    assign layer1_out[7422] = layer0_out[1482] ^ layer0_out[1483];
    assign layer1_out[7423] = layer0_out[3448] & ~layer0_out[3449];
    assign layer1_out[7424] = ~layer0_out[7194];
    assign layer1_out[7425] = ~layer0_out[5509] | layer0_out[5508];
    assign layer1_out[7426] = ~(layer0_out[1211] & layer0_out[1212]);
    assign layer1_out[7427] = ~layer0_out[679] | layer0_out[678];
    assign layer1_out[7428] = ~layer0_out[2912] | layer0_out[2913];
    assign layer1_out[7429] = layer0_out[7335] | layer0_out[7336];
    assign layer1_out[7430] = ~(layer0_out[6807] ^ layer0_out[6808]);
    assign layer1_out[7431] = ~(layer0_out[5913] ^ layer0_out[5914]);
    assign layer1_out[7432] = ~layer0_out[1609];
    assign layer1_out[7433] = ~layer0_out[4586] | layer0_out[4585];
    assign layer1_out[7434] = ~layer0_out[7318];
    assign layer1_out[7435] = ~(layer0_out[447] & layer0_out[448]);
    assign layer1_out[7436] = layer0_out[3182];
    assign layer1_out[7437] = ~layer0_out[6695];
    assign layer1_out[7438] = ~layer0_out[3189];
    assign layer1_out[7439] = ~(layer0_out[2748] | layer0_out[2749]);
    assign layer1_out[7440] = layer0_out[1558] | layer0_out[1559];
    assign layer1_out[7441] = layer0_out[1562] & ~layer0_out[1561];
    assign layer1_out[7442] = ~(layer0_out[3191] & layer0_out[3192]);
    assign layer1_out[7443] = ~layer0_out[372] | layer0_out[373];
    assign layer1_out[7444] = ~(layer0_out[5634] & layer0_out[5635]);
    assign layer1_out[7445] = layer0_out[1978] & ~layer0_out[1979];
    assign layer1_out[7446] = ~layer0_out[231];
    assign layer1_out[7447] = layer0_out[7668] & layer0_out[7669];
    assign layer1_out[7448] = ~layer0_out[2729] | layer0_out[2730];
    assign layer1_out[7449] = ~(layer0_out[5202] | layer0_out[5203]);
    assign layer1_out[7450] = ~(layer0_out[3832] & layer0_out[3833]);
    assign layer1_out[7451] = layer0_out[4];
    assign layer1_out[7452] = ~(layer0_out[2581] ^ layer0_out[2582]);
    assign layer1_out[7453] = layer0_out[947];
    assign layer1_out[7454] = ~layer0_out[192];
    assign layer1_out[7455] = ~(layer0_out[3755] | layer0_out[3756]);
    assign layer1_out[7456] = layer0_out[7470] & ~layer0_out[7471];
    assign layer1_out[7457] = ~layer0_out[2620] | layer0_out[2621];
    assign layer1_out[7458] = layer0_out[5539] & ~layer0_out[5540];
    assign layer1_out[7459] = ~(layer0_out[4810] & layer0_out[4811]);
    assign layer1_out[7460] = layer0_out[5451];
    assign layer1_out[7461] = ~layer0_out[3935];
    assign layer1_out[7462] = layer0_out[5550];
    assign layer1_out[7463] = layer0_out[3379] & layer0_out[3380];
    assign layer1_out[7464] = layer0_out[6541] ^ layer0_out[6542];
    assign layer1_out[7465] = layer0_out[7280] ^ layer0_out[7281];
    assign layer1_out[7466] = layer0_out[2349];
    assign layer1_out[7467] = layer0_out[853];
    assign layer1_out[7468] = ~layer0_out[4869];
    assign layer1_out[7469] = ~(layer0_out[2903] | layer0_out[2904]);
    assign layer1_out[7470] = 1'b0;
    assign layer1_out[7471] = ~layer0_out[7346] | layer0_out[7347];
    assign layer1_out[7472] = layer0_out[769] & ~layer0_out[768];
    assign layer1_out[7473] = ~layer0_out[2462];
    assign layer1_out[7474] = ~layer0_out[240] | layer0_out[239];
    assign layer1_out[7475] = layer0_out[2729];
    assign layer1_out[7476] = layer0_out[1708] | layer0_out[1709];
    assign layer1_out[7477] = layer0_out[2559] & ~layer0_out[2560];
    assign layer1_out[7478] = layer0_out[619];
    assign layer1_out[7479] = ~layer0_out[5338] | layer0_out[5337];
    assign layer1_out[7480] = ~layer0_out[2660];
    assign layer1_out[7481] = ~layer0_out[177];
    assign layer1_out[7482] = ~layer0_out[3097] | layer0_out[3096];
    assign layer1_out[7483] = layer0_out[6105] | layer0_out[6106];
    assign layer1_out[7484] = ~layer0_out[4329];
    assign layer1_out[7485] = ~layer0_out[6633] | layer0_out[6632];
    assign layer1_out[7486] = ~layer0_out[7575] | layer0_out[7576];
    assign layer1_out[7487] = ~layer0_out[1315] | layer0_out[1316];
    assign layer1_out[7488] = layer0_out[4340];
    assign layer1_out[7489] = layer0_out[119];
    assign layer1_out[7490] = 1'b0;
    assign layer1_out[7491] = layer0_out[2200] | layer0_out[2201];
    assign layer1_out[7492] = 1'b0;
    assign layer1_out[7493] = ~layer0_out[7673];
    assign layer1_out[7494] = 1'b0;
    assign layer1_out[7495] = ~layer0_out[4103] | layer0_out[4104];
    assign layer1_out[7496] = 1'b0;
    assign layer1_out[7497] = layer0_out[406] | layer0_out[407];
    assign layer1_out[7498] = layer0_out[3126] & ~layer0_out[3127];
    assign layer1_out[7499] = layer0_out[1600] & layer0_out[1601];
    assign layer1_out[7500] = layer0_out[2191] & ~layer0_out[2192];
    assign layer1_out[7501] = ~(layer0_out[2280] & layer0_out[2281]);
    assign layer1_out[7502] = layer0_out[4354] | layer0_out[4355];
    assign layer1_out[7503] = ~(layer0_out[2262] | layer0_out[2263]);
    assign layer1_out[7504] = ~layer0_out[1360] | layer0_out[1361];
    assign layer1_out[7505] = ~(layer0_out[5962] & layer0_out[5963]);
    assign layer1_out[7506] = ~layer0_out[6028];
    assign layer1_out[7507] = ~layer0_out[6432] | layer0_out[6431];
    assign layer1_out[7508] = layer0_out[1209] | layer0_out[1210];
    assign layer1_out[7509] = layer0_out[6313] & ~layer0_out[6314];
    assign layer1_out[7510] = ~(layer0_out[605] | layer0_out[606]);
    assign layer1_out[7511] = ~(layer0_out[2236] | layer0_out[2237]);
    assign layer1_out[7512] = layer0_out[2435] & layer0_out[2436];
    assign layer1_out[7513] = ~(layer0_out[6420] | layer0_out[6421]);
    assign layer1_out[7514] = ~(layer0_out[1439] & layer0_out[1440]);
    assign layer1_out[7515] = layer0_out[3153] & ~layer0_out[3152];
    assign layer1_out[7516] = ~(layer0_out[3322] & layer0_out[3323]);
    assign layer1_out[7517] = layer0_out[3351];
    assign layer1_out[7518] = ~(layer0_out[2525] & layer0_out[2526]);
    assign layer1_out[7519] = layer0_out[5817] & layer0_out[5818];
    assign layer1_out[7520] = ~layer0_out[542];
    assign layer1_out[7521] = ~(layer0_out[1522] & layer0_out[1523]);
    assign layer1_out[7522] = layer0_out[2338] | layer0_out[2339];
    assign layer1_out[7523] = ~layer0_out[4833];
    assign layer1_out[7524] = 1'b1;
    assign layer1_out[7525] = layer0_out[6770];
    assign layer1_out[7526] = ~layer0_out[2040];
    assign layer1_out[7527] = layer0_out[7633] & layer0_out[7634];
    assign layer1_out[7528] = layer0_out[4212] ^ layer0_out[4213];
    assign layer1_out[7529] = ~layer0_out[5094] | layer0_out[5095];
    assign layer1_out[7530] = ~layer0_out[5393];
    assign layer1_out[7531] = ~layer0_out[6063];
    assign layer1_out[7532] = layer0_out[2927] & layer0_out[2928];
    assign layer1_out[7533] = 1'b0;
    assign layer1_out[7534] = ~layer0_out[1230];
    assign layer1_out[7535] = layer0_out[5856] & layer0_out[5857];
    assign layer1_out[7536] = ~layer0_out[3452] | layer0_out[3451];
    assign layer1_out[7537] = ~layer0_out[7236];
    assign layer1_out[7538] = 1'b1;
    assign layer1_out[7539] = ~layer0_out[486] | layer0_out[487];
    assign layer1_out[7540] = 1'b1;
    assign layer1_out[7541] = layer0_out[5718];
    assign layer1_out[7542] = ~(layer0_out[1423] & layer0_out[1424]);
    assign layer1_out[7543] = ~layer0_out[347];
    assign layer1_out[7544] = layer0_out[2301] & ~layer0_out[2300];
    assign layer1_out[7545] = layer0_out[1593] & ~layer0_out[1594];
    assign layer1_out[7546] = ~layer0_out[3126];
    assign layer1_out[7547] = layer0_out[2536];
    assign layer1_out[7548] = layer0_out[3907] | layer0_out[3908];
    assign layer1_out[7549] = layer0_out[6560];
    assign layer1_out[7550] = layer0_out[6013] ^ layer0_out[6014];
    assign layer1_out[7551] = 1'b0;
    assign layer1_out[7552] = ~(layer0_out[1913] & layer0_out[1914]);
    assign layer1_out[7553] = ~(layer0_out[6487] ^ layer0_out[6488]);
    assign layer1_out[7554] = ~(layer0_out[7830] | layer0_out[7831]);
    assign layer1_out[7555] = layer0_out[2787];
    assign layer1_out[7556] = ~layer0_out[6418] | layer0_out[6417];
    assign layer1_out[7557] = ~layer0_out[2930];
    assign layer1_out[7558] = ~layer0_out[3390];
    assign layer1_out[7559] = layer0_out[5194] | layer0_out[5195];
    assign layer1_out[7560] = layer0_out[3766] & ~layer0_out[3765];
    assign layer1_out[7561] = layer0_out[6915];
    assign layer1_out[7562] = layer0_out[2122];
    assign layer1_out[7563] = 1'b1;
    assign layer1_out[7564] = ~layer0_out[156] | layer0_out[157];
    assign layer1_out[7565] = layer0_out[3325];
    assign layer1_out[7566] = ~(layer0_out[3715] | layer0_out[3716]);
    assign layer1_out[7567] = 1'b1;
    assign layer1_out[7568] = 1'b1;
    assign layer1_out[7569] = layer0_out[7279];
    assign layer1_out[7570] = ~layer0_out[2387] | layer0_out[2388];
    assign layer1_out[7571] = layer0_out[4385] ^ layer0_out[4386];
    assign layer1_out[7572] = layer0_out[4468] | layer0_out[4469];
    assign layer1_out[7573] = ~layer0_out[5578] | layer0_out[5577];
    assign layer1_out[7574] = ~(layer0_out[4004] | layer0_out[4005]);
    assign layer1_out[7575] = ~layer0_out[2902];
    assign layer1_out[7576] = ~layer0_out[164] | layer0_out[165];
    assign layer1_out[7577] = layer0_out[1821] | layer0_out[1822];
    assign layer1_out[7578] = layer0_out[6047] ^ layer0_out[6048];
    assign layer1_out[7579] = layer0_out[5807] & layer0_out[5808];
    assign layer1_out[7580] = layer0_out[427] | layer0_out[428];
    assign layer1_out[7581] = ~layer0_out[2841];
    assign layer1_out[7582] = layer0_out[501] & ~layer0_out[500];
    assign layer1_out[7583] = ~(layer0_out[916] & layer0_out[917]);
    assign layer1_out[7584] = layer0_out[3202];
    assign layer1_out[7585] = layer0_out[5694] | layer0_out[5695];
    assign layer1_out[7586] = layer0_out[6510];
    assign layer1_out[7587] = layer0_out[1404] | layer0_out[1405];
    assign layer1_out[7588] = ~(layer0_out[4592] | layer0_out[4593]);
    assign layer1_out[7589] = ~(layer0_out[4300] | layer0_out[4301]);
    assign layer1_out[7590] = layer0_out[1493];
    assign layer1_out[7591] = layer0_out[5492] & ~layer0_out[5491];
    assign layer1_out[7592] = layer0_out[7157] ^ layer0_out[7158];
    assign layer1_out[7593] = ~(layer0_out[4862] | layer0_out[4863]);
    assign layer1_out[7594] = ~layer0_out[4088];
    assign layer1_out[7595] = ~(layer0_out[4961] & layer0_out[4962]);
    assign layer1_out[7596] = layer0_out[1101];
    assign layer1_out[7597] = layer0_out[5876] | layer0_out[5877];
    assign layer1_out[7598] = layer0_out[6131] & ~layer0_out[6130];
    assign layer1_out[7599] = ~layer0_out[7117];
    assign layer1_out[7600] = ~layer0_out[5399] | layer0_out[5400];
    assign layer1_out[7601] = layer0_out[5066] & ~layer0_out[5065];
    assign layer1_out[7602] = layer0_out[6104] & layer0_out[6105];
    assign layer1_out[7603] = ~layer0_out[6318] | layer0_out[6319];
    assign layer1_out[7604] = layer0_out[4237];
    assign layer1_out[7605] = 1'b0;
    assign layer1_out[7606] = ~layer0_out[2911];
    assign layer1_out[7607] = layer0_out[7504] & layer0_out[7505];
    assign layer1_out[7608] = layer0_out[7522] & ~layer0_out[7523];
    assign layer1_out[7609] = layer0_out[199];
    assign layer1_out[7610] = layer0_out[4072];
    assign layer1_out[7611] = layer0_out[3319] & layer0_out[3320];
    assign layer1_out[7612] = layer0_out[7173] | layer0_out[7174];
    assign layer1_out[7613] = ~layer0_out[3169] | layer0_out[3168];
    assign layer1_out[7614] = layer0_out[2025] | layer0_out[2026];
    assign layer1_out[7615] = ~layer0_out[5359];
    assign layer1_out[7616] = ~layer0_out[3154];
    assign layer1_out[7617] = ~(layer0_out[7120] & layer0_out[7121]);
    assign layer1_out[7618] = ~layer0_out[745];
    assign layer1_out[7619] = layer0_out[7166] & ~layer0_out[7165];
    assign layer1_out[7620] = layer0_out[268] | layer0_out[269];
    assign layer1_out[7621] = layer0_out[864];
    assign layer1_out[7622] = ~layer0_out[5219];
    assign layer1_out[7623] = layer0_out[867] & layer0_out[868];
    assign layer1_out[7624] = layer0_out[3073];
    assign layer1_out[7625] = ~layer0_out[3762] | layer0_out[3763];
    assign layer1_out[7626] = layer0_out[2243];
    assign layer1_out[7627] = ~layer0_out[868] | layer0_out[869];
    assign layer1_out[7628] = layer0_out[6466];
    assign layer1_out[7629] = ~layer0_out[4187] | layer0_out[4186];
    assign layer1_out[7630] = layer0_out[3026] & ~layer0_out[3025];
    assign layer1_out[7631] = layer0_out[1719];
    assign layer1_out[7632] = ~layer0_out[4065];
    assign layer1_out[7633] = ~layer0_out[6570];
    assign layer1_out[7634] = layer0_out[5766];
    assign layer1_out[7635] = ~layer0_out[6935] | layer0_out[6936];
    assign layer1_out[7636] = layer0_out[329] & ~layer0_out[330];
    assign layer1_out[7637] = ~layer0_out[3405];
    assign layer1_out[7638] = layer0_out[1287] & ~layer0_out[1286];
    assign layer1_out[7639] = ~(layer0_out[4965] ^ layer0_out[4966]);
    assign layer1_out[7640] = layer0_out[3358] & layer0_out[3359];
    assign layer1_out[7641] = ~layer0_out[7197] | layer0_out[7196];
    assign layer1_out[7642] = ~layer0_out[4395];
    assign layer1_out[7643] = ~(layer0_out[1120] & layer0_out[1121]);
    assign layer1_out[7644] = 1'b1;
    assign layer1_out[7645] = 1'b0;
    assign layer1_out[7646] = ~(layer0_out[4611] ^ layer0_out[4612]);
    assign layer1_out[7647] = ~(layer0_out[3372] | layer0_out[3373]);
    assign layer1_out[7648] = layer0_out[2702];
    assign layer1_out[7649] = ~layer0_out[3348] | layer0_out[3347];
    assign layer1_out[7650] = layer0_out[122] & layer0_out[123];
    assign layer1_out[7651] = ~(layer0_out[5878] ^ layer0_out[5879]);
    assign layer1_out[7652] = ~layer0_out[6027];
    assign layer1_out[7653] = ~(layer0_out[7415] & layer0_out[7416]);
    assign layer1_out[7654] = ~layer0_out[4679];
    assign layer1_out[7655] = 1'b1;
    assign layer1_out[7656] = layer0_out[4818] & ~layer0_out[4817];
    assign layer1_out[7657] = layer0_out[6341];
    assign layer1_out[7658] = ~layer0_out[2712];
    assign layer1_out[7659] = layer0_out[7457];
    assign layer1_out[7660] = ~(layer0_out[5410] & layer0_out[5411]);
    assign layer1_out[7661] = ~(layer0_out[6472] & layer0_out[6473]);
    assign layer1_out[7662] = ~layer0_out[7902];
    assign layer1_out[7663] = layer0_out[1371] ^ layer0_out[1372];
    assign layer1_out[7664] = ~layer0_out[3859] | layer0_out[3858];
    assign layer1_out[7665] = ~layer0_out[2642] | layer0_out[2643];
    assign layer1_out[7666] = ~layer0_out[3198] | layer0_out[3199];
    assign layer1_out[7667] = ~(layer0_out[5816] | layer0_out[5817]);
    assign layer1_out[7668] = layer0_out[3086] ^ layer0_out[3087];
    assign layer1_out[7669] = layer0_out[6016] & layer0_out[6017];
    assign layer1_out[7670] = ~(layer0_out[7710] & layer0_out[7711]);
    assign layer1_out[7671] = ~layer0_out[6581];
    assign layer1_out[7672] = layer0_out[2575] & layer0_out[2576];
    assign layer1_out[7673] = ~layer0_out[5681];
    assign layer1_out[7674] = ~layer0_out[798] | layer0_out[797];
    assign layer1_out[7675] = ~layer0_out[3586] | layer0_out[3587];
    assign layer1_out[7676] = layer0_out[1341];
    assign layer1_out[7677] = ~(layer0_out[3037] & layer0_out[3038]);
    assign layer1_out[7678] = 1'b1;
    assign layer1_out[7679] = layer0_out[1615] & ~layer0_out[1614];
    assign layer1_out[7680] = ~layer0_out[4776] | layer0_out[4777];
    assign layer1_out[7681] = ~(layer0_out[3597] | layer0_out[3598]);
    assign layer1_out[7682] = ~(layer0_out[2715] ^ layer0_out[2716]);
    assign layer1_out[7683] = layer0_out[1170];
    assign layer1_out[7684] = ~layer0_out[2567];
    assign layer1_out[7685] = ~(layer0_out[2137] ^ layer0_out[2138]);
    assign layer1_out[7686] = ~layer0_out[18] | layer0_out[17];
    assign layer1_out[7687] = layer0_out[1933] & ~layer0_out[1932];
    assign layer1_out[7688] = 1'b0;
    assign layer1_out[7689] = ~layer0_out[4202];
    assign layer1_out[7690] = ~layer0_out[4225];
    assign layer1_out[7691] = ~(layer0_out[4993] & layer0_out[4994]);
    assign layer1_out[7692] = layer0_out[4510] | layer0_out[4511];
    assign layer1_out[7693] = layer0_out[4587] & ~layer0_out[4586];
    assign layer1_out[7694] = ~layer0_out[6531] | layer0_out[6530];
    assign layer1_out[7695] = ~(layer0_out[5119] & layer0_out[5120]);
    assign layer1_out[7696] = ~layer0_out[5437];
    assign layer1_out[7697] = ~layer0_out[1721];
    assign layer1_out[7698] = layer0_out[2380] | layer0_out[2381];
    assign layer1_out[7699] = layer0_out[5271];
    assign layer1_out[7700] = ~(layer0_out[2028] | layer0_out[2029]);
    assign layer1_out[7701] = ~layer0_out[5616] | layer0_out[5617];
    assign layer1_out[7702] = layer0_out[7321] | layer0_out[7322];
    assign layer1_out[7703] = 1'b0;
    assign layer1_out[7704] = layer0_out[785] & ~layer0_out[784];
    assign layer1_out[7705] = ~layer0_out[240] | layer0_out[241];
    assign layer1_out[7706] = layer0_out[6637];
    assign layer1_out[7707] = layer0_out[1015];
    assign layer1_out[7708] = ~(layer0_out[5195] | layer0_out[5196]);
    assign layer1_out[7709] = ~layer0_out[6461] | layer0_out[6462];
    assign layer1_out[7710] = ~layer0_out[4145];
    assign layer1_out[7711] = layer0_out[1524] | layer0_out[1525];
    assign layer1_out[7712] = 1'b0;
    assign layer1_out[7713] = ~layer0_out[7764];
    assign layer1_out[7714] = layer0_out[5870];
    assign layer1_out[7715] = 1'b1;
    assign layer1_out[7716] = layer0_out[6549] | layer0_out[6550];
    assign layer1_out[7717] = ~layer0_out[7927];
    assign layer1_out[7718] = ~layer0_out[7510];
    assign layer1_out[7719] = ~(layer0_out[178] ^ layer0_out[179]);
    assign layer1_out[7720] = layer0_out[5587] & layer0_out[5588];
    assign layer1_out[7721] = layer0_out[5386];
    assign layer1_out[7722] = ~layer0_out[1954] | layer0_out[1953];
    assign layer1_out[7723] = layer0_out[5850] & ~layer0_out[5849];
    assign layer1_out[7724] = layer0_out[6406] & ~layer0_out[6407];
    assign layer1_out[7725] = layer0_out[1266] & layer0_out[1267];
    assign layer1_out[7726] = layer0_out[3004] & ~layer0_out[3003];
    assign layer1_out[7727] = ~layer0_out[3396];
    assign layer1_out[7728] = 1'b1;
    assign layer1_out[7729] = ~layer0_out[4406];
    assign layer1_out[7730] = ~layer0_out[3124] | layer0_out[3123];
    assign layer1_out[7731] = layer0_out[6744] & layer0_out[6745];
    assign layer1_out[7732] = ~layer0_out[5663];
    assign layer1_out[7733] = ~layer0_out[320] | layer0_out[321];
    assign layer1_out[7734] = layer0_out[3414] & layer0_out[3415];
    assign layer1_out[7735] = ~layer0_out[1135] | layer0_out[1136];
    assign layer1_out[7736] = layer0_out[1014];
    assign layer1_out[7737] = ~(layer0_out[4037] & layer0_out[4038]);
    assign layer1_out[7738] = layer0_out[4938] | layer0_out[4939];
    assign layer1_out[7739] = layer0_out[5526] & layer0_out[5527];
    assign layer1_out[7740] = ~(layer0_out[6348] | layer0_out[6349]);
    assign layer1_out[7741] = ~(layer0_out[6620] | layer0_out[6621]);
    assign layer1_out[7742] = ~(layer0_out[154] | layer0_out[155]);
    assign layer1_out[7743] = ~layer0_out[2122] | layer0_out[2121];
    assign layer1_out[7744] = ~(layer0_out[485] & layer0_out[486]);
    assign layer1_out[7745] = layer0_out[3626] ^ layer0_out[3627];
    assign layer1_out[7746] = layer0_out[7556] | layer0_out[7557];
    assign layer1_out[7747] = layer0_out[1438] | layer0_out[1439];
    assign layer1_out[7748] = layer0_out[2287];
    assign layer1_out[7749] = layer0_out[1967];
    assign layer1_out[7750] = ~layer0_out[7555];
    assign layer1_out[7751] = layer0_out[7562];
    assign layer1_out[7752] = layer0_out[4871] & ~layer0_out[4870];
    assign layer1_out[7753] = ~(layer0_out[7348] ^ layer0_out[7349]);
    assign layer1_out[7754] = ~(layer0_out[3049] ^ layer0_out[3050]);
    assign layer1_out[7755] = 1'b1;
    assign layer1_out[7756] = layer0_out[3516] & ~layer0_out[3515];
    assign layer1_out[7757] = layer0_out[6700] & layer0_out[6701];
    assign layer1_out[7758] = ~layer0_out[301] | layer0_out[300];
    assign layer1_out[7759] = layer0_out[5096] & ~layer0_out[5097];
    assign layer1_out[7760] = ~(layer0_out[6298] | layer0_out[6299]);
    assign layer1_out[7761] = 1'b0;
    assign layer1_out[7762] = ~layer0_out[102];
    assign layer1_out[7763] = layer0_out[7492];
    assign layer1_out[7764] = layer0_out[2475];
    assign layer1_out[7765] = layer0_out[5032];
    assign layer1_out[7766] = layer0_out[1245] & ~layer0_out[1246];
    assign layer1_out[7767] = 1'b1;
    assign layer1_out[7768] = ~layer0_out[7398] | layer0_out[7399];
    assign layer1_out[7769] = layer0_out[2142];
    assign layer1_out[7770] = ~layer0_out[1905];
    assign layer1_out[7771] = ~(layer0_out[4411] | layer0_out[4412]);
    assign layer1_out[7772] = layer0_out[4160];
    assign layer1_out[7773] = ~layer0_out[2883] | layer0_out[2882];
    assign layer1_out[7774] = ~(layer0_out[6488] | layer0_out[6489]);
    assign layer1_out[7775] = layer0_out[3192] ^ layer0_out[3193];
    assign layer1_out[7776] = layer0_out[6225] | layer0_out[6226];
    assign layer1_out[7777] = ~layer0_out[3342];
    assign layer1_out[7778] = ~layer0_out[6606] | layer0_out[6605];
    assign layer1_out[7779] = ~layer0_out[5669];
    assign layer1_out[7780] = ~layer0_out[7555];
    assign layer1_out[7781] = ~layer0_out[2327];
    assign layer1_out[7782] = ~layer0_out[4101] | layer0_out[4100];
    assign layer1_out[7783] = 1'b0;
    assign layer1_out[7784] = 1'b0;
    assign layer1_out[7785] = layer0_out[2206] & layer0_out[2207];
    assign layer1_out[7786] = 1'b1;
    assign layer1_out[7787] = layer0_out[4996] & layer0_out[4997];
    assign layer1_out[7788] = layer0_out[6144] ^ layer0_out[6145];
    assign layer1_out[7789] = ~(layer0_out[4848] | layer0_out[4849]);
    assign layer1_out[7790] = ~layer0_out[6727];
    assign layer1_out[7791] = layer0_out[1332] & ~layer0_out[1333];
    assign layer1_out[7792] = layer0_out[3260] & layer0_out[3261];
    assign layer1_out[7793] = layer0_out[7176] | layer0_out[7177];
    assign layer1_out[7794] = ~layer0_out[2808];
    assign layer1_out[7795] = layer0_out[2192] & layer0_out[2193];
    assign layer1_out[7796] = ~(layer0_out[1186] | layer0_out[1187]);
    assign layer1_out[7797] = ~layer0_out[1042] | layer0_out[1043];
    assign layer1_out[7798] = ~layer0_out[7335];
    assign layer1_out[7799] = ~layer0_out[4577] | layer0_out[4576];
    assign layer1_out[7800] = ~(layer0_out[6568] & layer0_out[6569]);
    assign layer1_out[7801] = layer0_out[6879] & ~layer0_out[6880];
    assign layer1_out[7802] = ~layer0_out[651] | layer0_out[650];
    assign layer1_out[7803] = 1'b1;
    assign layer1_out[7804] = layer0_out[1330] | layer0_out[1331];
    assign layer1_out[7805] = ~(layer0_out[994] | layer0_out[995]);
    assign layer1_out[7806] = ~(layer0_out[3810] ^ layer0_out[3811]);
    assign layer1_out[7807] = layer0_out[4710];
    assign layer1_out[7808] = ~layer0_out[7983] | layer0_out[7982];
    assign layer1_out[7809] = ~layer0_out[7568];
    assign layer1_out[7810] = layer0_out[4076];
    assign layer1_out[7811] = layer0_out[2184];
    assign layer1_out[7812] = layer0_out[3827] & layer0_out[3828];
    assign layer1_out[7813] = ~layer0_out[4964];
    assign layer1_out[7814] = 1'b1;
    assign layer1_out[7815] = layer0_out[5637] | layer0_out[5638];
    assign layer1_out[7816] = layer0_out[6782];
    assign layer1_out[7817] = ~(layer0_out[2749] & layer0_out[2750]);
    assign layer1_out[7818] = ~layer0_out[4934];
    assign layer1_out[7819] = ~(layer0_out[1911] ^ layer0_out[1912]);
    assign layer1_out[7820] = layer0_out[6579] & ~layer0_out[6580];
    assign layer1_out[7821] = ~(layer0_out[3050] | layer0_out[3051]);
    assign layer1_out[7822] = ~(layer0_out[2161] | layer0_out[2162]);
    assign layer1_out[7823] = ~(layer0_out[7237] ^ layer0_out[7238]);
    assign layer1_out[7824] = layer0_out[7223] ^ layer0_out[7224];
    assign layer1_out[7825] = layer0_out[1788] | layer0_out[1789];
    assign layer1_out[7826] = layer0_out[4942] & layer0_out[4943];
    assign layer1_out[7827] = 1'b0;
    assign layer1_out[7828] = ~layer0_out[4409];
    assign layer1_out[7829] = 1'b1;
    assign layer1_out[7830] = layer0_out[1780] & ~layer0_out[1781];
    assign layer1_out[7831] = 1'b1;
    assign layer1_out[7832] = layer0_out[4222] & layer0_out[4223];
    assign layer1_out[7833] = ~layer0_out[6588] | layer0_out[6587];
    assign layer1_out[7834] = layer0_out[6262] & ~layer0_out[6263];
    assign layer1_out[7835] = layer0_out[752];
    assign layer1_out[7836] = 1'b1;
    assign layer1_out[7837] = layer0_out[2888];
    assign layer1_out[7838] = layer0_out[4813] & layer0_out[4814];
    assign layer1_out[7839] = ~layer0_out[1090];
    assign layer1_out[7840] = layer0_out[7338];
    assign layer1_out[7841] = ~layer0_out[4795];
    assign layer1_out[7842] = layer0_out[7285] | layer0_out[7286];
    assign layer1_out[7843] = layer0_out[7910] & ~layer0_out[7911];
    assign layer1_out[7844] = ~layer0_out[4308] | layer0_out[4309];
    assign layer1_out[7845] = ~layer0_out[1001];
    assign layer1_out[7846] = ~layer0_out[3471];
    assign layer1_out[7847] = layer0_out[923] ^ layer0_out[924];
    assign layer1_out[7848] = ~(layer0_out[7758] & layer0_out[7759]);
    assign layer1_out[7849] = layer0_out[7923];
    assign layer1_out[7850] = layer0_out[7564];
    assign layer1_out[7851] = ~layer0_out[5696] | layer0_out[5695];
    assign layer1_out[7852] = layer0_out[4980] & ~layer0_out[4979];
    assign layer1_out[7853] = layer0_out[2745] | layer0_out[2746];
    assign layer1_out[7854] = layer0_out[5081] | layer0_out[5082];
    assign layer1_out[7855] = ~layer0_out[2629];
    assign layer1_out[7856] = ~layer0_out[614] | layer0_out[615];
    assign layer1_out[7857] = ~(layer0_out[6378] & layer0_out[6379]);
    assign layer1_out[7858] = layer0_out[7725] & layer0_out[7726];
    assign layer1_out[7859] = ~layer0_out[3600];
    assign layer1_out[7860] = layer0_out[4986] | layer0_out[4987];
    assign layer1_out[7861] = 1'b0;
    assign layer1_out[7862] = layer0_out[7959];
    assign layer1_out[7863] = ~layer0_out[138] | layer0_out[139];
    assign layer1_out[7864] = layer0_out[4471] & ~layer0_out[4472];
    assign layer1_out[7865] = layer0_out[7973] & layer0_out[7974];
    assign layer1_out[7866] = layer0_out[6127];
    assign layer1_out[7867] = ~(layer0_out[4822] ^ layer0_out[4823]);
    assign layer1_out[7868] = layer0_out[6972] & ~layer0_out[6973];
    assign layer1_out[7869] = ~(layer0_out[1099] | layer0_out[1100]);
    assign layer1_out[7870] = 1'b1;
    assign layer1_out[7871] = layer0_out[6866] ^ layer0_out[6867];
    assign layer1_out[7872] = 1'b0;
    assign layer1_out[7873] = layer0_out[767] & ~layer0_out[768];
    assign layer1_out[7874] = 1'b1;
    assign layer1_out[7875] = ~layer0_out[667] | layer0_out[666];
    assign layer1_out[7876] = ~layer0_out[1231];
    assign layer1_out[7877] = ~layer0_out[3959];
    assign layer1_out[7878] = ~layer0_out[3224];
    assign layer1_out[7879] = layer0_out[7632];
    assign layer1_out[7880] = ~layer0_out[161];
    assign layer1_out[7881] = 1'b1;
    assign layer1_out[7882] = ~layer0_out[7814];
    assign layer1_out[7883] = ~layer0_out[5257] | layer0_out[5256];
    assign layer1_out[7884] = ~layer0_out[3714];
    assign layer1_out[7885] = layer0_out[903] & layer0_out[904];
    assign layer1_out[7886] = layer0_out[1381];
    assign layer1_out[7887] = ~layer0_out[3546];
    assign layer1_out[7888] = ~layer0_out[3640] | layer0_out[3639];
    assign layer1_out[7889] = ~(layer0_out[7857] | layer0_out[7858]);
    assign layer1_out[7890] = ~layer0_out[6435] | layer0_out[6436];
    assign layer1_out[7891] = layer0_out[1634];
    assign layer1_out[7892] = layer0_out[1886] & ~layer0_out[1885];
    assign layer1_out[7893] = layer0_out[4759] & layer0_out[4760];
    assign layer1_out[7894] = ~layer0_out[5749];
    assign layer1_out[7895] = ~layer0_out[5010];
    assign layer1_out[7896] = ~(layer0_out[1204] | layer0_out[1205]);
    assign layer1_out[7897] = ~layer0_out[2681];
    assign layer1_out[7898] = layer0_out[699] & ~layer0_out[698];
    assign layer1_out[7899] = layer0_out[530] ^ layer0_out[531];
    assign layer1_out[7900] = layer0_out[5583] & layer0_out[5584];
    assign layer1_out[7901] = ~layer0_out[6413] | layer0_out[6412];
    assign layer1_out[7902] = ~(layer0_out[5791] ^ layer0_out[5792]);
    assign layer1_out[7903] = ~layer0_out[3274] | layer0_out[3273];
    assign layer1_out[7904] = layer0_out[273];
    assign layer1_out[7905] = 1'b1;
    assign layer1_out[7906] = ~layer0_out[4157];
    assign layer1_out[7907] = ~(layer0_out[3280] & layer0_out[3281]);
    assign layer1_out[7908] = ~layer0_out[6801] | layer0_out[6802];
    assign layer1_out[7909] = layer0_out[3010];
    assign layer1_out[7910] = layer0_out[847];
    assign layer1_out[7911] = layer0_out[3719];
    assign layer1_out[7912] = layer0_out[3232];
    assign layer1_out[7913] = ~layer0_out[1774] | layer0_out[1773];
    assign layer1_out[7914] = layer0_out[1763] ^ layer0_out[1764];
    assign layer1_out[7915] = ~layer0_out[7763] | layer0_out[7762];
    assign layer1_out[7916] = ~(layer0_out[4975] & layer0_out[4976]);
    assign layer1_out[7917] = layer0_out[70] | layer0_out[71];
    assign layer1_out[7918] = layer0_out[4878] | layer0_out[4879];
    assign layer1_out[7919] = layer0_out[3670] & ~layer0_out[3671];
    assign layer1_out[7920] = layer0_out[160] & ~layer0_out[159];
    assign layer1_out[7921] = layer0_out[4750] | layer0_out[4751];
    assign layer1_out[7922] = ~layer0_out[4056];
    assign layer1_out[7923] = ~layer0_out[3213];
    assign layer1_out[7924] = layer0_out[2688] & ~layer0_out[2687];
    assign layer1_out[7925] = ~layer0_out[1094];
    assign layer1_out[7926] = ~layer0_out[6223] | layer0_out[6222];
    assign layer1_out[7927] = ~(layer0_out[6884] ^ layer0_out[6885]);
    assign layer1_out[7928] = ~layer0_out[4160];
    assign layer1_out[7929] = ~layer0_out[892];
    assign layer1_out[7930] = ~layer0_out[4247] | layer0_out[4248];
    assign layer1_out[7931] = layer0_out[4742] ^ layer0_out[4743];
    assign layer1_out[7932] = layer0_out[2899] & ~layer0_out[2898];
    assign layer1_out[7933] = layer0_out[127];
    assign layer1_out[7934] = ~layer0_out[1165];
    assign layer1_out[7935] = ~layer0_out[1107];
    assign layer1_out[7936] = ~layer0_out[3098] | layer0_out[3097];
    assign layer1_out[7937] = layer0_out[6827];
    assign layer1_out[7938] = layer0_out[7894] & ~layer0_out[7893];
    assign layer1_out[7939] = ~layer0_out[6763];
    assign layer1_out[7940] = layer0_out[5100];
    assign layer1_out[7941] = layer0_out[7268] ^ layer0_out[7269];
    assign layer1_out[7942] = layer0_out[5267];
    assign layer1_out[7943] = layer0_out[1597] | layer0_out[1598];
    assign layer1_out[7944] = layer0_out[7869] & ~layer0_out[7868];
    assign layer1_out[7945] = ~layer0_out[6290];
    assign layer1_out[7946] = layer0_out[5400];
    assign layer1_out[7947] = layer0_out[1395] & layer0_out[1396];
    assign layer1_out[7948] = layer0_out[3124] ^ layer0_out[3125];
    assign layer1_out[7949] = layer0_out[4764];
    assign layer1_out[7950] = layer0_out[2181] | layer0_out[2182];
    assign layer1_out[7951] = layer0_out[1317] & ~layer0_out[1318];
    assign layer1_out[7952] = layer0_out[4216] & ~layer0_out[4215];
    assign layer1_out[7953] = layer0_out[2747];
    assign layer1_out[7954] = ~layer0_out[1130];
    assign layer1_out[7955] = layer0_out[5478] & layer0_out[5479];
    assign layer1_out[7956] = layer0_out[2499] & ~layer0_out[2498];
    assign layer1_out[7957] = layer0_out[1008];
    assign layer1_out[7958] = layer0_out[6908];
    assign layer1_out[7959] = layer0_out[4563] & ~layer0_out[4562];
    assign layer1_out[7960] = ~(layer0_out[103] & layer0_out[104]);
    assign layer1_out[7961] = layer0_out[3084] & ~layer0_out[3085];
    assign layer1_out[7962] = 1'b0;
    assign layer1_out[7963] = 1'b1;
    assign layer1_out[7964] = ~layer0_out[5178];
    assign layer1_out[7965] = layer0_out[6750] | layer0_out[6751];
    assign layer1_out[7966] = layer0_out[4967];
    assign layer1_out[7967] = ~layer0_out[6007];
    assign layer1_out[7968] = ~layer0_out[6084] | layer0_out[6083];
    assign layer1_out[7969] = layer0_out[568] & ~layer0_out[569];
    assign layer1_out[7970] = layer0_out[6329] & ~layer0_out[6330];
    assign layer1_out[7971] = layer0_out[6137] & ~layer0_out[6136];
    assign layer1_out[7972] = layer0_out[7898];
    assign layer1_out[7973] = ~layer0_out[6854];
    assign layer1_out[7974] = layer0_out[834] ^ layer0_out[835];
    assign layer1_out[7975] = layer0_out[3956] & ~layer0_out[3957];
    assign layer1_out[7976] = layer0_out[3590] & ~layer0_out[3591];
    assign layer1_out[7977] = layer0_out[6055];
    assign layer1_out[7978] = ~(layer0_out[6277] & layer0_out[6278]);
    assign layer1_out[7979] = ~layer0_out[559];
    assign layer1_out[7980] = layer0_out[2502] & layer0_out[2503];
    assign layer1_out[7981] = ~layer0_out[6325];
    assign layer1_out[7982] = layer0_out[1990];
    assign layer1_out[7983] = ~layer0_out[5972];
    assign layer1_out[7984] = 1'b1;
    assign layer1_out[7985] = ~layer0_out[5318] | layer0_out[5317];
    assign layer1_out[7986] = layer0_out[172];
    assign layer1_out[7987] = ~(layer0_out[7105] | layer0_out[7106]);
    assign layer1_out[7988] = ~layer0_out[1688];
    assign layer1_out[7989] = ~layer0_out[4757] | layer0_out[4756];
    assign layer1_out[7990] = layer0_out[3417] | layer0_out[3418];
    assign layer1_out[7991] = layer0_out[4705];
    assign layer1_out[7992] = 1'b1;
    assign layer1_out[7993] = ~layer0_out[3336] | layer0_out[3335];
    assign layer1_out[7994] = ~(layer0_out[7793] | layer0_out[7794]);
    assign layer1_out[7995] = ~layer0_out[2343];
    assign layer1_out[7996] = ~layer0_out[3662] | layer0_out[3661];
    assign layer1_out[7997] = ~layer0_out[6307];
    assign layer1_out[7998] = ~layer0_out[4789] | layer0_out[4788];
    assign layer1_out[7999] = ~layer0_out[5905];
    assign layer2_out[0] = layer1_out[6798] & layer1_out[6799];
    assign layer2_out[1] = ~(layer1_out[1705] & layer1_out[1706]);
    assign layer2_out[2] = 1'b0;
    assign layer2_out[3] = layer1_out[6799];
    assign layer2_out[4] = ~layer1_out[4999] | layer1_out[4998];
    assign layer2_out[5] = ~layer1_out[2729] | layer1_out[2730];
    assign layer2_out[6] = layer1_out[2348];
    assign layer2_out[7] = 1'b0;
    assign layer2_out[8] = layer1_out[7939];
    assign layer2_out[9] = layer1_out[3397] & ~layer1_out[3398];
    assign layer2_out[10] = layer1_out[4167];
    assign layer2_out[11] = ~layer1_out[5831];
    assign layer2_out[12] = layer1_out[1431];
    assign layer2_out[13] = ~layer1_out[241] | layer1_out[242];
    assign layer2_out[14] = layer1_out[4546];
    assign layer2_out[15] = 1'b1;
    assign layer2_out[16] = layer1_out[1420] | layer1_out[1421];
    assign layer2_out[17] = ~layer1_out[6646];
    assign layer2_out[18] = layer1_out[7021] & ~layer1_out[7020];
    assign layer2_out[19] = layer1_out[4827];
    assign layer2_out[20] = ~layer1_out[4028];
    assign layer2_out[21] = layer1_out[4058];
    assign layer2_out[22] = ~layer1_out[639];
    assign layer2_out[23] = ~(layer1_out[654] ^ layer1_out[655]);
    assign layer2_out[24] = layer1_out[2152] & ~layer1_out[2151];
    assign layer2_out[25] = ~layer1_out[7476];
    assign layer2_out[26] = ~layer1_out[6361];
    assign layer2_out[27] = layer1_out[1986] & layer1_out[1987];
    assign layer2_out[28] = ~(layer1_out[1286] ^ layer1_out[1287]);
    assign layer2_out[29] = ~(layer1_out[7325] | layer1_out[7326]);
    assign layer2_out[30] = ~(layer1_out[6400] ^ layer1_out[6401]);
    assign layer2_out[31] = ~layer1_out[7745];
    assign layer2_out[32] = ~layer1_out[6430];
    assign layer2_out[33] = ~(layer1_out[7194] ^ layer1_out[7195]);
    assign layer2_out[34] = ~layer1_out[1891];
    assign layer2_out[35] = layer1_out[3733];
    assign layer2_out[36] = ~layer1_out[2520];
    assign layer2_out[37] = layer1_out[5291] | layer1_out[5292];
    assign layer2_out[38] = ~layer1_out[7320];
    assign layer2_out[39] = ~layer1_out[1877] | layer1_out[1876];
    assign layer2_out[40] = ~layer1_out[2301] | layer1_out[2302];
    assign layer2_out[41] = ~(layer1_out[721] & layer1_out[722]);
    assign layer2_out[42] = ~layer1_out[6665] | layer1_out[6664];
    assign layer2_out[43] = ~layer1_out[7462] | layer1_out[7463];
    assign layer2_out[44] = layer1_out[2354] & layer1_out[2355];
    assign layer2_out[45] = layer1_out[4456] | layer1_out[4457];
    assign layer2_out[46] = layer1_out[5990];
    assign layer2_out[47] = ~(layer1_out[2957] & layer1_out[2958]);
    assign layer2_out[48] = layer1_out[5977];
    assign layer2_out[49] = layer1_out[3111];
    assign layer2_out[50] = ~layer1_out[5119] | layer1_out[5120];
    assign layer2_out[51] = ~layer1_out[420] | layer1_out[421];
    assign layer2_out[52] = layer1_out[7430] & ~layer1_out[7431];
    assign layer2_out[53] = layer1_out[4197] & ~layer1_out[4196];
    assign layer2_out[54] = ~layer1_out[1042];
    assign layer2_out[55] = ~layer1_out[361];
    assign layer2_out[56] = ~layer1_out[5034];
    assign layer2_out[57] = layer1_out[4329] | layer1_out[4330];
    assign layer2_out[58] = layer1_out[1907] & ~layer1_out[1906];
    assign layer2_out[59] = layer1_out[75] & ~layer1_out[74];
    assign layer2_out[60] = layer1_out[5444] & layer1_out[5445];
    assign layer2_out[61] = ~layer1_out[2686] | layer1_out[2685];
    assign layer2_out[62] = layer1_out[2386] & ~layer1_out[2385];
    assign layer2_out[63] = ~layer1_out[4192];
    assign layer2_out[64] = ~(layer1_out[3782] ^ layer1_out[3783]);
    assign layer2_out[65] = ~(layer1_out[1019] ^ layer1_out[1020]);
    assign layer2_out[66] = layer1_out[2892];
    assign layer2_out[67] = 1'b0;
    assign layer2_out[68] = layer1_out[2413] | layer1_out[2414];
    assign layer2_out[69] = ~layer1_out[1010] | layer1_out[1011];
    assign layer2_out[70] = layer1_out[1548] & ~layer1_out[1547];
    assign layer2_out[71] = layer1_out[6924];
    assign layer2_out[72] = layer1_out[3658] & ~layer1_out[3659];
    assign layer2_out[73] = ~(layer1_out[7775] | layer1_out[7776]);
    assign layer2_out[74] = layer1_out[3826] & ~layer1_out[3827];
    assign layer2_out[75] = ~layer1_out[4656];
    assign layer2_out[76] = 1'b1;
    assign layer2_out[77] = layer1_out[2696];
    assign layer2_out[78] = layer1_out[1257] & layer1_out[1258];
    assign layer2_out[79] = layer1_out[5131] | layer1_out[5132];
    assign layer2_out[80] = layer1_out[6794];
    assign layer2_out[81] = ~layer1_out[1270] | layer1_out[1271];
    assign layer2_out[82] = layer1_out[2809];
    assign layer2_out[83] = ~layer1_out[426];
    assign layer2_out[84] = ~(layer1_out[3028] & layer1_out[3029]);
    assign layer2_out[85] = ~(layer1_out[1435] ^ layer1_out[1436]);
    assign layer2_out[86] = layer1_out[260] & ~layer1_out[261];
    assign layer2_out[87] = layer1_out[2919] | layer1_out[2920];
    assign layer2_out[88] = layer1_out[2875];
    assign layer2_out[89] = layer1_out[3333] | layer1_out[3334];
    assign layer2_out[90] = layer1_out[2358];
    assign layer2_out[91] = ~(layer1_out[45] & layer1_out[46]);
    assign layer2_out[92] = layer1_out[2831] & layer1_out[2832];
    assign layer2_out[93] = ~layer1_out[5833];
    assign layer2_out[94] = layer1_out[2330];
    assign layer2_out[95] = ~layer1_out[6907];
    assign layer2_out[96] = ~(layer1_out[39] & layer1_out[40]);
    assign layer2_out[97] = ~layer1_out[3612] | layer1_out[3613];
    assign layer2_out[98] = layer1_out[7431] | layer1_out[7432];
    assign layer2_out[99] = layer1_out[4188];
    assign layer2_out[100] = ~layer1_out[5459];
    assign layer2_out[101] = ~layer1_out[7159];
    assign layer2_out[102] = layer1_out[5340] | layer1_out[5341];
    assign layer2_out[103] = ~layer1_out[3446];
    assign layer2_out[104] = 1'b0;
    assign layer2_out[105] = ~layer1_out[2230] | layer1_out[2231];
    assign layer2_out[106] = layer1_out[6016];
    assign layer2_out[107] = ~layer1_out[4943];
    assign layer2_out[108] = layer1_out[4766] & layer1_out[4767];
    assign layer2_out[109] = ~(layer1_out[7476] | layer1_out[7477]);
    assign layer2_out[110] = layer1_out[6920] & layer1_out[6921];
    assign layer2_out[111] = ~layer1_out[7849];
    assign layer2_out[112] = ~layer1_out[6362];
    assign layer2_out[113] = ~(layer1_out[2530] ^ layer1_out[2531]);
    assign layer2_out[114] = ~layer1_out[7715] | layer1_out[7716];
    assign layer2_out[115] = ~(layer1_out[131] ^ layer1_out[132]);
    assign layer2_out[116] = ~layer1_out[703];
    assign layer2_out[117] = ~(layer1_out[7615] ^ layer1_out[7616]);
    assign layer2_out[118] = layer1_out[106];
    assign layer2_out[119] = layer1_out[4303] & ~layer1_out[4302];
    assign layer2_out[120] = ~layer1_out[5016];
    assign layer2_out[121] = layer1_out[7794] & layer1_out[7795];
    assign layer2_out[122] = 1'b1;
    assign layer2_out[123] = ~layer1_out[6157];
    assign layer2_out[124] = layer1_out[1797] & ~layer1_out[1798];
    assign layer2_out[125] = ~layer1_out[5294] | layer1_out[5295];
    assign layer2_out[126] = layer1_out[3962] & layer1_out[3963];
    assign layer2_out[127] = layer1_out[3215] & ~layer1_out[3214];
    assign layer2_out[128] = layer1_out[3428];
    assign layer2_out[129] = layer1_out[1429] | layer1_out[1430];
    assign layer2_out[130] = layer1_out[3211] | layer1_out[3212];
    assign layer2_out[131] = ~layer1_out[4947] | layer1_out[4946];
    assign layer2_out[132] = layer1_out[5553];
    assign layer2_out[133] = layer1_out[3498] | layer1_out[3499];
    assign layer2_out[134] = layer1_out[7638];
    assign layer2_out[135] = ~layer1_out[1556];
    assign layer2_out[136] = layer1_out[2218] ^ layer1_out[2219];
    assign layer2_out[137] = ~layer1_out[3591];
    assign layer2_out[138] = ~(layer1_out[770] ^ layer1_out[771]);
    assign layer2_out[139] = layer1_out[3897] & ~layer1_out[3896];
    assign layer2_out[140] = ~layer1_out[4749];
    assign layer2_out[141] = layer1_out[6615] ^ layer1_out[6616];
    assign layer2_out[142] = ~(layer1_out[1565] | layer1_out[1566]);
    assign layer2_out[143] = ~layer1_out[3483] | layer1_out[3482];
    assign layer2_out[144] = layer1_out[5929];
    assign layer2_out[145] = ~layer1_out[1087] | layer1_out[1088];
    assign layer2_out[146] = ~(layer1_out[4544] & layer1_out[4545]);
    assign layer2_out[147] = ~layer1_out[3373] | layer1_out[3372];
    assign layer2_out[148] = layer1_out[1313];
    assign layer2_out[149] = layer1_out[3769];
    assign layer2_out[150] = layer1_out[2647] ^ layer1_out[2648];
    assign layer2_out[151] = 1'b1;
    assign layer2_out[152] = ~layer1_out[4702];
    assign layer2_out[153] = layer1_out[4535];
    assign layer2_out[154] = layer1_out[6214];
    assign layer2_out[155] = 1'b1;
    assign layer2_out[156] = ~layer1_out[2939];
    assign layer2_out[157] = layer1_out[3582] & ~layer1_out[3581];
    assign layer2_out[158] = 1'b1;
    assign layer2_out[159] = ~layer1_out[4413];
    assign layer2_out[160] = ~layer1_out[1617];
    assign layer2_out[161] = ~layer1_out[3056];
    assign layer2_out[162] = layer1_out[234] & ~layer1_out[233];
    assign layer2_out[163] = layer1_out[4910] | layer1_out[4911];
    assign layer2_out[164] = layer1_out[5530] ^ layer1_out[5531];
    assign layer2_out[165] = layer1_out[5310];
    assign layer2_out[166] = layer1_out[2111] & ~layer1_out[2112];
    assign layer2_out[167] = ~layer1_out[4589];
    assign layer2_out[168] = ~layer1_out[1982] | layer1_out[1983];
    assign layer2_out[169] = layer1_out[3517] & ~layer1_out[3518];
    assign layer2_out[170] = layer1_out[5687] | layer1_out[5688];
    assign layer2_out[171] = ~(layer1_out[1772] & layer1_out[1773]);
    assign layer2_out[172] = ~(layer1_out[646] ^ layer1_out[647]);
    assign layer2_out[173] = ~layer1_out[5857];
    assign layer2_out[174] = ~layer1_out[312] | layer1_out[311];
    assign layer2_out[175] = layer1_out[989];
    assign layer2_out[176] = layer1_out[1875];
    assign layer2_out[177] = ~layer1_out[446];
    assign layer2_out[178] = ~(layer1_out[5197] ^ layer1_out[5198]);
    assign layer2_out[179] = ~layer1_out[5795];
    assign layer2_out[180] = ~(layer1_out[7713] & layer1_out[7714]);
    assign layer2_out[181] = layer1_out[7416] & layer1_out[7417];
    assign layer2_out[182] = layer1_out[3327] & layer1_out[3328];
    assign layer2_out[183] = layer1_out[5157];
    assign layer2_out[184] = layer1_out[876] & ~layer1_out[877];
    assign layer2_out[185] = layer1_out[1841] & ~layer1_out[1840];
    assign layer2_out[186] = ~(layer1_out[4863] | layer1_out[4864]);
    assign layer2_out[187] = layer1_out[6447];
    assign layer2_out[188] = ~(layer1_out[5092] & layer1_out[5093]);
    assign layer2_out[189] = layer1_out[4970];
    assign layer2_out[190] = ~layer1_out[3080];
    assign layer2_out[191] = layer1_out[5918] & ~layer1_out[5919];
    assign layer2_out[192] = layer1_out[2021];
    assign layer2_out[193] = layer1_out[3700] | layer1_out[3701];
    assign layer2_out[194] = ~(layer1_out[6590] & layer1_out[6591]);
    assign layer2_out[195] = layer1_out[7880];
    assign layer2_out[196] = ~layer1_out[2135];
    assign layer2_out[197] = ~layer1_out[4952];
    assign layer2_out[198] = ~layer1_out[5267];
    assign layer2_out[199] = 1'b0;
    assign layer2_out[200] = ~(layer1_out[6065] ^ layer1_out[6066]);
    assign layer2_out[201] = layer1_out[5623];
    assign layer2_out[202] = layer1_out[5481] & ~layer1_out[5482];
    assign layer2_out[203] = layer1_out[2702];
    assign layer2_out[204] = layer1_out[6718] | layer1_out[6719];
    assign layer2_out[205] = ~(layer1_out[4019] | layer1_out[4020]);
    assign layer2_out[206] = ~layer1_out[1483];
    assign layer2_out[207] = layer1_out[4520];
    assign layer2_out[208] = layer1_out[1511];
    assign layer2_out[209] = layer1_out[393] | layer1_out[394];
    assign layer2_out[210] = ~layer1_out[2700];
    assign layer2_out[211] = ~layer1_out[2215] | layer1_out[2216];
    assign layer2_out[212] = ~layer1_out[6134];
    assign layer2_out[213] = ~layer1_out[1904];
    assign layer2_out[214] = ~layer1_out[107];
    assign layer2_out[215] = layer1_out[1778];
    assign layer2_out[216] = layer1_out[2312] & ~layer1_out[2313];
    assign layer2_out[217] = ~(layer1_out[4230] ^ layer1_out[4231]);
    assign layer2_out[218] = 1'b0;
    assign layer2_out[219] = layer1_out[205] & ~layer1_out[206];
    assign layer2_out[220] = ~layer1_out[4414] | layer1_out[4415];
    assign layer2_out[221] = ~layer1_out[2535];
    assign layer2_out[222] = 1'b1;
    assign layer2_out[223] = ~layer1_out[748] | layer1_out[747];
    assign layer2_out[224] = ~layer1_out[3735] | layer1_out[3734];
    assign layer2_out[225] = layer1_out[4694] | layer1_out[4695];
    assign layer2_out[226] = layer1_out[3232] & ~layer1_out[3231];
    assign layer2_out[227] = layer1_out[7244] & ~layer1_out[7245];
    assign layer2_out[228] = layer1_out[2399];
    assign layer2_out[229] = layer1_out[581];
    assign layer2_out[230] = ~layer1_out[7337];
    assign layer2_out[231] = ~(layer1_out[2364] ^ layer1_out[2365]);
    assign layer2_out[232] = ~layer1_out[4954];
    assign layer2_out[233] = ~layer1_out[6414] | layer1_out[6415];
    assign layer2_out[234] = ~(layer1_out[2808] | layer1_out[2809]);
    assign layer2_out[235] = layer1_out[156] ^ layer1_out[157];
    assign layer2_out[236] = ~(layer1_out[7102] & layer1_out[7103]);
    assign layer2_out[237] = ~layer1_out[1755] | layer1_out[1754];
    assign layer2_out[238] = ~layer1_out[760] | layer1_out[759];
    assign layer2_out[239] = layer1_out[987];
    assign layer2_out[240] = ~(layer1_out[3914] & layer1_out[3915]);
    assign layer2_out[241] = ~(layer1_out[4858] ^ layer1_out[4859]);
    assign layer2_out[242] = ~layer1_out[6104];
    assign layer2_out[243] = ~layer1_out[6837];
    assign layer2_out[244] = layer1_out[49] ^ layer1_out[50];
    assign layer2_out[245] = ~layer1_out[7497];
    assign layer2_out[246] = ~layer1_out[5924] | layer1_out[5925];
    assign layer2_out[247] = ~layer1_out[4927];
    assign layer2_out[248] = layer1_out[6714];
    assign layer2_out[249] = ~(layer1_out[6600] ^ layer1_out[6601]);
    assign layer2_out[250] = layer1_out[3944] | layer1_out[3945];
    assign layer2_out[251] = ~layer1_out[1762] | layer1_out[1763];
    assign layer2_out[252] = ~layer1_out[1437];
    assign layer2_out[253] = 1'b0;
    assign layer2_out[254] = layer1_out[2150];
    assign layer2_out[255] = ~layer1_out[1466];
    assign layer2_out[256] = ~(layer1_out[7030] & layer1_out[7031]);
    assign layer2_out[257] = layer1_out[7308];
    assign layer2_out[258] = layer1_out[2702];
    assign layer2_out[259] = ~(layer1_out[7257] & layer1_out[7258]);
    assign layer2_out[260] = ~(layer1_out[3521] & layer1_out[3522]);
    assign layer2_out[261] = ~layer1_out[1128] | layer1_out[1129];
    assign layer2_out[262] = layer1_out[3485];
    assign layer2_out[263] = ~(layer1_out[1256] & layer1_out[1257]);
    assign layer2_out[264] = layer1_out[7651] & layer1_out[7652];
    assign layer2_out[265] = layer1_out[1461];
    assign layer2_out[266] = ~layer1_out[6421];
    assign layer2_out[267] = ~layer1_out[4361] | layer1_out[4362];
    assign layer2_out[268] = layer1_out[7881] & layer1_out[7882];
    assign layer2_out[269] = ~layer1_out[6900];
    assign layer2_out[270] = layer1_out[7031] & layer1_out[7032];
    assign layer2_out[271] = ~(layer1_out[5288] ^ layer1_out[5289]);
    assign layer2_out[272] = layer1_out[2380] & ~layer1_out[2379];
    assign layer2_out[273] = layer1_out[2599];
    assign layer2_out[274] = ~layer1_out[942];
    assign layer2_out[275] = ~(layer1_out[270] | layer1_out[271]);
    assign layer2_out[276] = layer1_out[5354] & layer1_out[5355];
    assign layer2_out[277] = layer1_out[4761] & ~layer1_out[4762];
    assign layer2_out[278] = ~(layer1_out[5867] ^ layer1_out[5868]);
    assign layer2_out[279] = ~layer1_out[2855];
    assign layer2_out[280] = layer1_out[718] & ~layer1_out[717];
    assign layer2_out[281] = ~layer1_out[3594] | layer1_out[3595];
    assign layer2_out[282] = ~(layer1_out[6463] ^ layer1_out[6464]);
    assign layer2_out[283] = layer1_out[5786] & ~layer1_out[5787];
    assign layer2_out[284] = ~layer1_out[3801];
    assign layer2_out[285] = ~layer1_out[2625];
    assign layer2_out[286] = layer1_out[3121];
    assign layer2_out[287] = layer1_out[1640] & ~layer1_out[1641];
    assign layer2_out[288] = ~layer1_out[832] | layer1_out[833];
    assign layer2_out[289] = ~layer1_out[6038];
    assign layer2_out[290] = layer1_out[1941];
    assign layer2_out[291] = layer1_out[4178] & layer1_out[4179];
    assign layer2_out[292] = ~layer1_out[2470];
    assign layer2_out[293] = layer1_out[5228];
    assign layer2_out[294] = layer1_out[4921];
    assign layer2_out[295] = layer1_out[346] & ~layer1_out[345];
    assign layer2_out[296] = ~(layer1_out[1344] & layer1_out[1345]);
    assign layer2_out[297] = ~(layer1_out[6782] | layer1_out[6783]);
    assign layer2_out[298] = ~layer1_out[6191];
    assign layer2_out[299] = ~layer1_out[441];
    assign layer2_out[300] = 1'b1;
    assign layer2_out[301] = layer1_out[3225];
    assign layer2_out[302] = ~layer1_out[4883];
    assign layer2_out[303] = 1'b1;
    assign layer2_out[304] = ~(layer1_out[1568] | layer1_out[1569]);
    assign layer2_out[305] = layer1_out[7510];
    assign layer2_out[306] = ~(layer1_out[5729] & layer1_out[5730]);
    assign layer2_out[307] = layer1_out[6258];
    assign layer2_out[308] = layer1_out[6496];
    assign layer2_out[309] = ~layer1_out[385] | layer1_out[386];
    assign layer2_out[310] = ~(layer1_out[2319] ^ layer1_out[2320]);
    assign layer2_out[311] = ~(layer1_out[1035] | layer1_out[1036]);
    assign layer2_out[312] = ~layer1_out[3266];
    assign layer2_out[313] = ~layer1_out[6230];
    assign layer2_out[314] = layer1_out[2479] & ~layer1_out[2480];
    assign layer2_out[315] = layer1_out[1472] ^ layer1_out[1473];
    assign layer2_out[316] = ~layer1_out[3422] | layer1_out[3423];
    assign layer2_out[317] = 1'b1;
    assign layer2_out[318] = ~layer1_out[2923];
    assign layer2_out[319] = ~(layer1_out[5887] ^ layer1_out[5888]);
    assign layer2_out[320] = ~(layer1_out[5542] & layer1_out[5543]);
    assign layer2_out[321] = layer1_out[7016] & ~layer1_out[7017];
    assign layer2_out[322] = layer1_out[6300] & ~layer1_out[6299];
    assign layer2_out[323] = layer1_out[2189];
    assign layer2_out[324] = layer1_out[1926];
    assign layer2_out[325] = layer1_out[6964] & ~layer1_out[6965];
    assign layer2_out[326] = layer1_out[378] & ~layer1_out[377];
    assign layer2_out[327] = ~layer1_out[1476] | layer1_out[1475];
    assign layer2_out[328] = layer1_out[228] & layer1_out[229];
    assign layer2_out[329] = ~(layer1_out[7932] | layer1_out[7933]);
    assign layer2_out[330] = ~(layer1_out[5353] | layer1_out[5354]);
    assign layer2_out[331] = layer1_out[4239] | layer1_out[4240];
    assign layer2_out[332] = 1'b1;
    assign layer2_out[333] = ~(layer1_out[6101] | layer1_out[6102]);
    assign layer2_out[334] = ~(layer1_out[6093] & layer1_out[6094]);
    assign layer2_out[335] = layer1_out[6044] & ~layer1_out[6045];
    assign layer2_out[336] = layer1_out[2567] ^ layer1_out[2568];
    assign layer2_out[337] = layer1_out[410] & ~layer1_out[409];
    assign layer2_out[338] = layer1_out[6677];
    assign layer2_out[339] = ~layer1_out[7580] | layer1_out[7581];
    assign layer2_out[340] = ~layer1_out[6488];
    assign layer2_out[341] = ~layer1_out[7216];
    assign layer2_out[342] = ~layer1_out[4475];
    assign layer2_out[343] = layer1_out[6554];
    assign layer2_out[344] = ~layer1_out[3710];
    assign layer2_out[345] = layer1_out[4088] & layer1_out[4089];
    assign layer2_out[346] = layer1_out[4465];
    assign layer2_out[347] = ~layer1_out[492];
    assign layer2_out[348] = ~layer1_out[3313];
    assign layer2_out[349] = layer1_out[5995];
    assign layer2_out[350] = ~layer1_out[4337] | layer1_out[4336];
    assign layer2_out[351] = ~layer1_out[5537] | layer1_out[5536];
    assign layer2_out[352] = layer1_out[3458] | layer1_out[3459];
    assign layer2_out[353] = layer1_out[516] & ~layer1_out[517];
    assign layer2_out[354] = layer1_out[2750];
    assign layer2_out[355] = layer1_out[1095] ^ layer1_out[1096];
    assign layer2_out[356] = ~layer1_out[4207] | layer1_out[4206];
    assign layer2_out[357] = layer1_out[5185];
    assign layer2_out[358] = ~layer1_out[2663];
    assign layer2_out[359] = layer1_out[1022] & ~layer1_out[1023];
    assign layer2_out[360] = ~layer1_out[1716] | layer1_out[1715];
    assign layer2_out[361] = ~(layer1_out[4425] & layer1_out[4426]);
    assign layer2_out[362] = layer1_out[765];
    assign layer2_out[363] = layer1_out[2228];
    assign layer2_out[364] = ~(layer1_out[2921] ^ layer1_out[2922]);
    assign layer2_out[365] = layer1_out[5978] ^ layer1_out[5979];
    assign layer2_out[366] = layer1_out[2825] & layer1_out[2826];
    assign layer2_out[367] = layer1_out[3064] & ~layer1_out[3065];
    assign layer2_out[368] = ~(layer1_out[869] | layer1_out[870]);
    assign layer2_out[369] = layer1_out[1758];
    assign layer2_out[370] = 1'b1;
    assign layer2_out[371] = ~layer1_out[954];
    assign layer2_out[372] = layer1_out[622] | layer1_out[623];
    assign layer2_out[373] = layer1_out[4556] & ~layer1_out[4557];
    assign layer2_out[374] = layer1_out[3711] & ~layer1_out[3710];
    assign layer2_out[375] = ~(layer1_out[4584] | layer1_out[4585]);
    assign layer2_out[376] = layer1_out[7855];
    assign layer2_out[377] = ~layer1_out[3759] | layer1_out[3760];
    assign layer2_out[378] = 1'b0;
    assign layer2_out[379] = ~layer1_out[4904] | layer1_out[4905];
    assign layer2_out[380] = ~layer1_out[3634];
    assign layer2_out[381] = layer1_out[7572];
    assign layer2_out[382] = ~layer1_out[1937] | layer1_out[1938];
    assign layer2_out[383] = ~layer1_out[564];
    assign layer2_out[384] = layer1_out[5947] ^ layer1_out[5948];
    assign layer2_out[385] = ~layer1_out[7933];
    assign layer2_out[386] = layer1_out[935] | layer1_out[936];
    assign layer2_out[387] = layer1_out[907];
    assign layer2_out[388] = layer1_out[3838] | layer1_out[3839];
    assign layer2_out[389] = layer1_out[752] | layer1_out[753];
    assign layer2_out[390] = ~(layer1_out[1358] | layer1_out[1359]);
    assign layer2_out[391] = layer1_out[2731] | layer1_out[2732];
    assign layer2_out[392] = ~layer1_out[1193];
    assign layer2_out[393] = ~layer1_out[2283] | layer1_out[2282];
    assign layer2_out[394] = ~layer1_out[4498] | layer1_out[4497];
    assign layer2_out[395] = layer1_out[5988] | layer1_out[5989];
    assign layer2_out[396] = layer1_out[3063];
    assign layer2_out[397] = layer1_out[1399] & ~layer1_out[1400];
    assign layer2_out[398] = layer1_out[4063] | layer1_out[4064];
    assign layer2_out[399] = ~layer1_out[6082] | layer1_out[6081];
    assign layer2_out[400] = 1'b1;
    assign layer2_out[401] = layer1_out[3670] | layer1_out[3671];
    assign layer2_out[402] = layer1_out[6426] & ~layer1_out[6425];
    assign layer2_out[403] = layer1_out[4625] | layer1_out[4626];
    assign layer2_out[404] = ~layer1_out[5325];
    assign layer2_out[405] = ~layer1_out[1769] | layer1_out[1770];
    assign layer2_out[406] = layer1_out[4424] | layer1_out[4425];
    assign layer2_out[407] = ~layer1_out[5528];
    assign layer2_out[408] = ~(layer1_out[6625] | layer1_out[6626]);
    assign layer2_out[409] = layer1_out[5316] ^ layer1_out[5317];
    assign layer2_out[410] = ~layer1_out[3904];
    assign layer2_out[411] = layer1_out[7845] & ~layer1_out[7846];
    assign layer2_out[412] = layer1_out[1274];
    assign layer2_out[413] = ~(layer1_out[5318] | layer1_out[5319]);
    assign layer2_out[414] = layer1_out[4042] & ~layer1_out[4041];
    assign layer2_out[415] = ~layer1_out[5776];
    assign layer2_out[416] = ~layer1_out[2232];
    assign layer2_out[417] = layer1_out[4160] & ~layer1_out[4159];
    assign layer2_out[418] = layer1_out[251];
    assign layer2_out[419] = ~layer1_out[5771];
    assign layer2_out[420] = layer1_out[7303] & ~layer1_out[7304];
    assign layer2_out[421] = ~(layer1_out[1469] ^ layer1_out[1470]);
    assign layer2_out[422] = ~(layer1_out[213] ^ layer1_out[214]);
    assign layer2_out[423] = 1'b1;
    assign layer2_out[424] = layer1_out[4139] & layer1_out[4140];
    assign layer2_out[425] = layer1_out[3149];
    assign layer2_out[426] = layer1_out[2688] & ~layer1_out[2687];
    assign layer2_out[427] = layer1_out[889];
    assign layer2_out[428] = layer1_out[3332] ^ layer1_out[3333];
    assign layer2_out[429] = ~layer1_out[7846] | layer1_out[7847];
    assign layer2_out[430] = layer1_out[4919];
    assign layer2_out[431] = ~layer1_out[4965];
    assign layer2_out[432] = ~(layer1_out[3229] & layer1_out[3230]);
    assign layer2_out[433] = layer1_out[4560];
    assign layer2_out[434] = ~layer1_out[6596] | layer1_out[6597];
    assign layer2_out[435] = ~(layer1_out[2295] | layer1_out[2296]);
    assign layer2_out[436] = layer1_out[6309];
    assign layer2_out[437] = layer1_out[1561] & layer1_out[1562];
    assign layer2_out[438] = ~layer1_out[1412] | layer1_out[1411];
    assign layer2_out[439] = ~(layer1_out[6953] & layer1_out[6954]);
    assign layer2_out[440] = ~(layer1_out[2549] & layer1_out[2550]);
    assign layer2_out[441] = layer1_out[7640] & ~layer1_out[7639];
    assign layer2_out[442] = layer1_out[6419] & layer1_out[6420];
    assign layer2_out[443] = layer1_out[6492] & ~layer1_out[6493];
    assign layer2_out[444] = layer1_out[1002] & ~layer1_out[1003];
    assign layer2_out[445] = 1'b0;
    assign layer2_out[446] = ~(layer1_out[1169] | layer1_out[1170]);
    assign layer2_out[447] = ~layer1_out[7204] | layer1_out[7203];
    assign layer2_out[448] = layer1_out[1572];
    assign layer2_out[449] = layer1_out[537];
    assign layer2_out[450] = ~(layer1_out[4348] ^ layer1_out[4349]);
    assign layer2_out[451] = layer1_out[4473];
    assign layer2_out[452] = ~(layer1_out[4874] & layer1_out[4875]);
    assign layer2_out[453] = layer1_out[1884];
    assign layer2_out[454] = ~(layer1_out[7731] | layer1_out[7732]);
    assign layer2_out[455] = ~layer1_out[2902] | layer1_out[2903];
    assign layer2_out[456] = ~layer1_out[2162] | layer1_out[2161];
    assign layer2_out[457] = layer1_out[6540] & layer1_out[6541];
    assign layer2_out[458] = ~layer1_out[3371] | layer1_out[3370];
    assign layer2_out[459] = ~(layer1_out[4013] ^ layer1_out[4014]);
    assign layer2_out[460] = ~(layer1_out[374] | layer1_out[375]);
    assign layer2_out[461] = layer1_out[6759];
    assign layer2_out[462] = layer1_out[7347] & ~layer1_out[7348];
    assign layer2_out[463] = layer1_out[7508] & ~layer1_out[7509];
    assign layer2_out[464] = 1'b1;
    assign layer2_out[465] = layer1_out[3417] & ~layer1_out[3416];
    assign layer2_out[466] = layer1_out[1343] & ~layer1_out[1344];
    assign layer2_out[467] = layer1_out[4505];
    assign layer2_out[468] = layer1_out[7095];
    assign layer2_out[469] = layer1_out[5849];
    assign layer2_out[470] = layer1_out[6456] & ~layer1_out[6455];
    assign layer2_out[471] = layer1_out[6179] & layer1_out[6180];
    assign layer2_out[472] = layer1_out[4499] & ~layer1_out[4498];
    assign layer2_out[473] = ~layer1_out[340];
    assign layer2_out[474] = ~(layer1_out[324] ^ layer1_out[325]);
    assign layer2_out[475] = layer1_out[4842] & layer1_out[4843];
    assign layer2_out[476] = ~(layer1_out[272] ^ layer1_out[273]);
    assign layer2_out[477] = layer1_out[6939];
    assign layer2_out[478] = layer1_out[605];
    assign layer2_out[479] = layer1_out[462];
    assign layer2_out[480] = ~(layer1_out[5216] ^ layer1_out[5217]);
    assign layer2_out[481] = layer1_out[6585] | layer1_out[6586];
    assign layer2_out[482] = layer1_out[845] & layer1_out[846];
    assign layer2_out[483] = layer1_out[3684];
    assign layer2_out[484] = ~layer1_out[6608];
    assign layer2_out[485] = layer1_out[7277];
    assign layer2_out[486] = ~layer1_out[6028];
    assign layer2_out[487] = 1'b0;
    assign layer2_out[488] = layer1_out[423] & ~layer1_out[422];
    assign layer2_out[489] = ~layer1_out[7882];
    assign layer2_out[490] = layer1_out[3865] & layer1_out[3866];
    assign layer2_out[491] = layer1_out[4591] | layer1_out[4592];
    assign layer2_out[492] = 1'b1;
    assign layer2_out[493] = ~layer1_out[7421] | layer1_out[7420];
    assign layer2_out[494] = layer1_out[2374];
    assign layer2_out[495] = ~layer1_out[4006];
    assign layer2_out[496] = ~layer1_out[6197] | layer1_out[6198];
    assign layer2_out[497] = layer1_out[29] & ~layer1_out[28];
    assign layer2_out[498] = 1'b0;
    assign layer2_out[499] = layer1_out[4275];
    assign layer2_out[500] = ~layer1_out[2581];
    assign layer2_out[501] = layer1_out[7871];
    assign layer2_out[502] = ~(layer1_out[7920] & layer1_out[7921]);
    assign layer2_out[503] = ~(layer1_out[4096] & layer1_out[4097]);
    assign layer2_out[504] = layer1_out[3838];
    assign layer2_out[505] = ~layer1_out[1033];
    assign layer2_out[506] = ~layer1_out[4813] | layer1_out[4814];
    assign layer2_out[507] = layer1_out[1531] & ~layer1_out[1530];
    assign layer2_out[508] = layer1_out[6854] & ~layer1_out[6853];
    assign layer2_out[509] = ~layer1_out[3614] | layer1_out[3613];
    assign layer2_out[510] = ~layer1_out[2587];
    assign layer2_out[511] = 1'b1;
    assign layer2_out[512] = layer1_out[2254];
    assign layer2_out[513] = ~layer1_out[811];
    assign layer2_out[514] = 1'b1;
    assign layer2_out[515] = ~layer1_out[5624];
    assign layer2_out[516] = ~(layer1_out[2148] | layer1_out[2149]);
    assign layer2_out[517] = ~layer1_out[2307] | layer1_out[2306];
    assign layer2_out[518] = layer1_out[3307] & ~layer1_out[3308];
    assign layer2_out[519] = ~(layer1_out[2716] | layer1_out[2717]);
    assign layer2_out[520] = ~layer1_out[3038];
    assign layer2_out[521] = layer1_out[7852] & layer1_out[7853];
    assign layer2_out[522] = layer1_out[5615];
    assign layer2_out[523] = ~layer1_out[5857];
    assign layer2_out[524] = ~layer1_out[7558];
    assign layer2_out[525] = layer1_out[51];
    assign layer2_out[526] = layer1_out[3511];
    assign layer2_out[527] = layer1_out[5606];
    assign layer2_out[528] = ~layer1_out[2182] | layer1_out[2181];
    assign layer2_out[529] = layer1_out[1863];
    assign layer2_out[530] = ~layer1_out[6395];
    assign layer2_out[531] = ~layer1_out[3843];
    assign layer2_out[532] = ~layer1_out[2350];
    assign layer2_out[533] = layer1_out[443];
    assign layer2_out[534] = ~layer1_out[6419];
    assign layer2_out[535] = layer1_out[2428];
    assign layer2_out[536] = ~layer1_out[2098] | layer1_out[2097];
    assign layer2_out[537] = layer1_out[4797];
    assign layer2_out[538] = 1'b1;
    assign layer2_out[539] = layer1_out[3363] & ~layer1_out[3362];
    assign layer2_out[540] = ~layer1_out[7329];
    assign layer2_out[541] = ~layer1_out[2344] | layer1_out[2343];
    assign layer2_out[542] = layer1_out[2971] ^ layer1_out[2972];
    assign layer2_out[543] = ~layer1_out[1952];
    assign layer2_out[544] = layer1_out[2187] & ~layer1_out[2188];
    assign layer2_out[545] = ~layer1_out[2929] | layer1_out[2930];
    assign layer2_out[546] = layer1_out[7904];
    assign layer2_out[547] = layer1_out[462] | layer1_out[463];
    assign layer2_out[548] = layer1_out[4] & layer1_out[5];
    assign layer2_out[549] = layer1_out[4903] & ~layer1_out[4902];
    assign layer2_out[550] = ~layer1_out[4656];
    assign layer2_out[551] = layer1_out[3444] | layer1_out[3445];
    assign layer2_out[552] = ~layer1_out[1516] | layer1_out[1515];
    assign layer2_out[553] = layer1_out[3421] | layer1_out[3422];
    assign layer2_out[554] = ~(layer1_out[1943] | layer1_out[1944]);
    assign layer2_out[555] = ~layer1_out[3216] | layer1_out[3217];
    assign layer2_out[556] = ~(layer1_out[3867] | layer1_out[3868]);
    assign layer2_out[557] = layer1_out[7066] & ~layer1_out[7065];
    assign layer2_out[558] = layer1_out[2828] & ~layer1_out[2827];
    assign layer2_out[559] = layer1_out[1298];
    assign layer2_out[560] = layer1_out[343];
    assign layer2_out[561] = ~(layer1_out[5221] ^ layer1_out[5222]);
    assign layer2_out[562] = layer1_out[2151] & ~layer1_out[2150];
    assign layer2_out[563] = ~layer1_out[5391];
    assign layer2_out[564] = ~layer1_out[7386];
    assign layer2_out[565] = layer1_out[5805] | layer1_out[5806];
    assign layer2_out[566] = ~layer1_out[2667] | layer1_out[2668];
    assign layer2_out[567] = ~(layer1_out[2252] | layer1_out[2253]);
    assign layer2_out[568] = ~layer1_out[6884];
    assign layer2_out[569] = layer1_out[5178] & ~layer1_out[5179];
    assign layer2_out[570] = ~layer1_out[7986];
    assign layer2_out[571] = layer1_out[1965] ^ layer1_out[1966];
    assign layer2_out[572] = ~(layer1_out[5188] & layer1_out[5189]);
    assign layer2_out[573] = ~layer1_out[3426];
    assign layer2_out[574] = layer1_out[4154] & ~layer1_out[4155];
    assign layer2_out[575] = layer1_out[5845] & ~layer1_out[5844];
    assign layer2_out[576] = ~(layer1_out[1059] | layer1_out[1060]);
    assign layer2_out[577] = 1'b1;
    assign layer2_out[578] = layer1_out[6863];
    assign layer2_out[579] = layer1_out[5965] & ~layer1_out[5966];
    assign layer2_out[580] = ~layer1_out[3271];
    assign layer2_out[581] = layer1_out[114] & ~layer1_out[115];
    assign layer2_out[582] = layer1_out[6030] ^ layer1_out[6031];
    assign layer2_out[583] = ~layer1_out[6442];
    assign layer2_out[584] = ~layer1_out[6803];
    assign layer2_out[585] = layer1_out[7736];
    assign layer2_out[586] = 1'b1;
    assign layer2_out[587] = layer1_out[4536] & layer1_out[4537];
    assign layer2_out[588] = layer1_out[3064] & ~layer1_out[3063];
    assign layer2_out[589] = ~layer1_out[7419];
    assign layer2_out[590] = ~(layer1_out[7184] & layer1_out[7185]);
    assign layer2_out[591] = ~layer1_out[748];
    assign layer2_out[592] = ~(layer1_out[81] & layer1_out[82]);
    assign layer2_out[593] = ~layer1_out[1506] | layer1_out[1505];
    assign layer2_out[594] = ~layer1_out[4855];
    assign layer2_out[595] = layer1_out[6326] & layer1_out[6327];
    assign layer2_out[596] = layer1_out[7480] & ~layer1_out[7479];
    assign layer2_out[597] = layer1_out[802] & ~layer1_out[803];
    assign layer2_out[598] = ~(layer1_out[7393] & layer1_out[7394]);
    assign layer2_out[599] = layer1_out[7850] & ~layer1_out[7851];
    assign layer2_out[600] = layer1_out[73];
    assign layer2_out[601] = ~layer1_out[6450];
    assign layer2_out[602] = layer1_out[5368];
    assign layer2_out[603] = ~(layer1_out[6744] | layer1_out[6745]);
    assign layer2_out[604] = ~layer1_out[1582];
    assign layer2_out[605] = ~layer1_out[96];
    assign layer2_out[606] = ~layer1_out[2645];
    assign layer2_out[607] = layer1_out[6979];
    assign layer2_out[608] = layer1_out[6649] & layer1_out[6650];
    assign layer2_out[609] = ~(layer1_out[297] & layer1_out[298]);
    assign layer2_out[610] = layer1_out[4609];
    assign layer2_out[611] = layer1_out[2548] & layer1_out[2549];
    assign layer2_out[612] = ~layer1_out[7790] | layer1_out[7791];
    assign layer2_out[613] = ~layer1_out[5160] | layer1_out[5161];
    assign layer2_out[614] = layer1_out[1023] ^ layer1_out[1024];
    assign layer2_out[615] = ~layer1_out[4631] | layer1_out[4632];
    assign layer2_out[616] = layer1_out[1104];
    assign layer2_out[617] = ~(layer1_out[3264] & layer1_out[3265]);
    assign layer2_out[618] = 1'b0;
    assign layer2_out[619] = 1'b1;
    assign layer2_out[620] = layer1_out[5921] & layer1_out[5922];
    assign layer2_out[621] = ~layer1_out[7910];
    assign layer2_out[622] = 1'b1;
    assign layer2_out[623] = ~layer1_out[6312] | layer1_out[6311];
    assign layer2_out[624] = layer1_out[4396] & ~layer1_out[4395];
    assign layer2_out[625] = ~layer1_out[4358] | layer1_out[4357];
    assign layer2_out[626] = ~(layer1_out[4437] | layer1_out[4438]);
    assign layer2_out[627] = ~layer1_out[4740] | layer1_out[4741];
    assign layer2_out[628] = ~layer1_out[5556];
    assign layer2_out[629] = ~layer1_out[1468] | layer1_out[1467];
    assign layer2_out[630] = ~layer1_out[7917];
    assign layer2_out[631] = 1'b1;
    assign layer2_out[632] = layer1_out[5176];
    assign layer2_out[633] = layer1_out[4667];
    assign layer2_out[634] = ~layer1_out[244];
    assign layer2_out[635] = ~layer1_out[489];
    assign layer2_out[636] = layer1_out[6252] & ~layer1_out[6251];
    assign layer2_out[637] = ~(layer1_out[606] & layer1_out[607]);
    assign layer2_out[638] = layer1_out[7027] ^ layer1_out[7028];
    assign layer2_out[639] = layer1_out[3598] & ~layer1_out[3599];
    assign layer2_out[640] = layer1_out[5246];
    assign layer2_out[641] = layer1_out[5974];
    assign layer2_out[642] = ~(layer1_out[7433] ^ layer1_out[7434]);
    assign layer2_out[643] = ~(layer1_out[3895] | layer1_out[3896]);
    assign layer2_out[644] = ~(layer1_out[6439] | layer1_out[6440]);
    assign layer2_out[645] = layer1_out[4637];
    assign layer2_out[646] = ~(layer1_out[5212] | layer1_out[5213]);
    assign layer2_out[647] = ~(layer1_out[3019] & layer1_out[3020]);
    assign layer2_out[648] = layer1_out[4247] ^ layer1_out[4248];
    assign layer2_out[649] = ~(layer1_out[55] & layer1_out[56]);
    assign layer2_out[650] = layer1_out[1190] ^ layer1_out[1191];
    assign layer2_out[651] = ~(layer1_out[2769] & layer1_out[2770]);
    assign layer2_out[652] = 1'b0;
    assign layer2_out[653] = layer1_out[6021] & ~layer1_out[6020];
    assign layer2_out[654] = layer1_out[3595] & layer1_out[3596];
    assign layer2_out[655] = ~layer1_out[4118];
    assign layer2_out[656] = layer1_out[4595];
    assign layer2_out[657] = layer1_out[4169];
    assign layer2_out[658] = ~layer1_out[254] | layer1_out[253];
    assign layer2_out[659] = 1'b0;
    assign layer2_out[660] = ~layer1_out[6819];
    assign layer2_out[661] = layer1_out[854] & layer1_out[855];
    assign layer2_out[662] = ~(layer1_out[4775] & layer1_out[4776]);
    assign layer2_out[663] = layer1_out[4060] & ~layer1_out[4059];
    assign layer2_out[664] = ~layer1_out[1793];
    assign layer2_out[665] = ~layer1_out[3897];
    assign layer2_out[666] = ~layer1_out[2482] | layer1_out[2483];
    assign layer2_out[667] = layer1_out[4282];
    assign layer2_out[668] = layer1_out[3179];
    assign layer2_out[669] = layer1_out[814] ^ layer1_out[815];
    assign layer2_out[670] = layer1_out[6286] & layer1_out[6287];
    assign layer2_out[671] = ~(layer1_out[6873] | layer1_out[6874]);
    assign layer2_out[672] = layer1_out[3368] & layer1_out[3369];
    assign layer2_out[673] = ~(layer1_out[2394] & layer1_out[2395]);
    assign layer2_out[674] = layer1_out[3988] & layer1_out[3989];
    assign layer2_out[675] = ~layer1_out[2425] | layer1_out[2426];
    assign layer2_out[676] = layer1_out[6856];
    assign layer2_out[677] = ~(layer1_out[6252] | layer1_out[6253]);
    assign layer2_out[678] = layer1_out[2620] & layer1_out[2621];
    assign layer2_out[679] = ~layer1_out[941] | layer1_out[942];
    assign layer2_out[680] = layer1_out[6911];
    assign layer2_out[681] = ~layer1_out[728] | layer1_out[729];
    assign layer2_out[682] = layer1_out[6053] & ~layer1_out[6054];
    assign layer2_out[683] = ~layer1_out[3955] | layer1_out[3954];
    assign layer2_out[684] = layer1_out[4698] & ~layer1_out[4697];
    assign layer2_out[685] = layer1_out[3873] & ~layer1_out[3874];
    assign layer2_out[686] = ~(layer1_out[2033] ^ layer1_out[2034]);
    assign layer2_out[687] = ~(layer1_out[3276] | layer1_out[3277]);
    assign layer2_out[688] = ~layer1_out[4244];
    assign layer2_out[689] = ~layer1_out[2595] | layer1_out[2594];
    assign layer2_out[690] = ~layer1_out[1184];
    assign layer2_out[691] = ~(layer1_out[7642] & layer1_out[7643]);
    assign layer2_out[692] = layer1_out[2671] & layer1_out[2672];
    assign layer2_out[693] = layer1_out[5200];
    assign layer2_out[694] = ~layer1_out[1806];
    assign layer2_out[695] = ~(layer1_out[7770] | layer1_out[7771]);
    assign layer2_out[696] = layer1_out[3949];
    assign layer2_out[697] = layer1_out[4407] ^ layer1_out[4408];
    assign layer2_out[698] = ~(layer1_out[1560] & layer1_out[1561]);
    assign layer2_out[699] = ~layer1_out[7663];
    assign layer2_out[700] = layer1_out[1220] | layer1_out[1221];
    assign layer2_out[701] = ~layer1_out[1545];
    assign layer2_out[702] = ~layer1_out[3304] | layer1_out[3303];
    assign layer2_out[703] = layer1_out[5699] & ~layer1_out[5700];
    assign layer2_out[704] = layer1_out[3622] | layer1_out[3623];
    assign layer2_out[705] = layer1_out[809] & ~layer1_out[808];
    assign layer2_out[706] = layer1_out[813] | layer1_out[814];
    assign layer2_out[707] = layer1_out[5709];
    assign layer2_out[708] = ~layer1_out[5048];
    assign layer2_out[709] = layer1_out[4390] & layer1_out[4391];
    assign layer2_out[710] = ~layer1_out[1831];
    assign layer2_out[711] = ~layer1_out[3780];
    assign layer2_out[712] = ~layer1_out[5375];
    assign layer2_out[713] = ~layer1_out[578] | layer1_out[577];
    assign layer2_out[714] = layer1_out[5655] & layer1_out[5656];
    assign layer2_out[715] = 1'b0;
    assign layer2_out[716] = layer1_out[5377] | layer1_out[5378];
    assign layer2_out[717] = layer1_out[4744] & layer1_out[4745];
    assign layer2_out[718] = ~(layer1_out[716] ^ layer1_out[717]);
    assign layer2_out[719] = layer1_out[1623] & ~layer1_out[1622];
    assign layer2_out[720] = ~(layer1_out[1384] ^ layer1_out[1385]);
    assign layer2_out[721] = ~layer1_out[7142];
    assign layer2_out[722] = ~layer1_out[724] | layer1_out[725];
    assign layer2_out[723] = layer1_out[1047] & ~layer1_out[1048];
    assign layer2_out[724] = layer1_out[5637];
    assign layer2_out[725] = layer1_out[412] & layer1_out[413];
    assign layer2_out[726] = layer1_out[2140] & layer1_out[2141];
    assign layer2_out[727] = ~layer1_out[2552];
    assign layer2_out[728] = 1'b1;
    assign layer2_out[729] = ~(layer1_out[4572] ^ layer1_out[4573]);
    assign layer2_out[730] = layer1_out[1867];
    assign layer2_out[731] = layer1_out[5535];
    assign layer2_out[732] = ~layer1_out[5254];
    assign layer2_out[733] = ~layer1_out[3672];
    assign layer2_out[734] = ~(layer1_out[3859] & layer1_out[3860]);
    assign layer2_out[735] = layer1_out[153] & ~layer1_out[154];
    assign layer2_out[736] = ~layer1_out[1977];
    assign layer2_out[737] = layer1_out[1260];
    assign layer2_out[738] = layer1_out[2511] & layer1_out[2512];
    assign layer2_out[739] = layer1_out[3501];
    assign layer2_out[740] = ~layer1_out[2587];
    assign layer2_out[741] = ~layer1_out[3121];
    assign layer2_out[742] = layer1_out[4085];
    assign layer2_out[743] = layer1_out[1302];
    assign layer2_out[744] = layer1_out[7286] & ~layer1_out[7287];
    assign layer2_out[745] = ~(layer1_out[6034] & layer1_out[6035]);
    assign layer2_out[746] = ~(layer1_out[7782] | layer1_out[7783]);
    assign layer2_out[747] = ~layer1_out[7049];
    assign layer2_out[748] = ~layer1_out[7083];
    assign layer2_out[749] = layer1_out[1027] & layer1_out[1028];
    assign layer2_out[750] = layer1_out[1711] ^ layer1_out[1712];
    assign layer2_out[751] = ~layer1_out[6960] | layer1_out[6959];
    assign layer2_out[752] = layer1_out[3204] & ~layer1_out[3203];
    assign layer2_out[753] = layer1_out[4607] & ~layer1_out[4606];
    assign layer2_out[754] = ~layer1_out[3328];
    assign layer2_out[755] = ~layer1_out[3424];
    assign layer2_out[756] = layer1_out[3140] & ~layer1_out[3141];
    assign layer2_out[757] = ~layer1_out[3979];
    assign layer2_out[758] = ~layer1_out[4820];
    assign layer2_out[759] = 1'b1;
    assign layer2_out[760] = ~layer1_out[5468];
    assign layer2_out[761] = layer1_out[3129] | layer1_out[3130];
    assign layer2_out[762] = ~layer1_out[1540];
    assign layer2_out[763] = ~(layer1_out[1609] & layer1_out[1610]);
    assign layer2_out[764] = layer1_out[5809] & ~layer1_out[5810];
    assign layer2_out[765] = layer1_out[87] & layer1_out[88];
    assign layer2_out[766] = layer1_out[5173] & ~layer1_out[5172];
    assign layer2_out[767] = ~layer1_out[3388];
    assign layer2_out[768] = ~layer1_out[3730];
    assign layer2_out[769] = layer1_out[6273] & ~layer1_out[6272];
    assign layer2_out[770] = ~layer1_out[7528];
    assign layer2_out[771] = ~(layer1_out[7445] | layer1_out[7446]);
    assign layer2_out[772] = ~(layer1_out[7337] & layer1_out[7338]);
    assign layer2_out[773] = layer1_out[7158] | layer1_out[7159];
    assign layer2_out[774] = layer1_out[5435] & layer1_out[5436];
    assign layer2_out[775] = ~(layer1_out[110] ^ layer1_out[111]);
    assign layer2_out[776] = ~layer1_out[1402] | layer1_out[1401];
    assign layer2_out[777] = ~layer1_out[738];
    assign layer2_out[778] = layer1_out[6804];
    assign layer2_out[779] = ~(layer1_out[5722] ^ layer1_out[5723]);
    assign layer2_out[780] = ~layer1_out[7007] | layer1_out[7008];
    assign layer2_out[781] = ~(layer1_out[147] | layer1_out[148]);
    assign layer2_out[782] = layer1_out[4642] & ~layer1_out[4641];
    assign layer2_out[783] = ~layer1_out[4177];
    assign layer2_out[784] = ~layer1_out[6804] | layer1_out[6803];
    assign layer2_out[785] = layer1_out[4466] ^ layer1_out[4467];
    assign layer2_out[786] = ~layer1_out[2734] | layer1_out[2733];
    assign layer2_out[787] = ~(layer1_out[2738] | layer1_out[2739]);
    assign layer2_out[788] = layer1_out[3950] & ~layer1_out[3951];
    assign layer2_out[789] = layer1_out[1633];
    assign layer2_out[790] = ~layer1_out[3688] | layer1_out[3687];
    assign layer2_out[791] = ~layer1_out[4078];
    assign layer2_out[792] = layer1_out[3340] & ~layer1_out[3339];
    assign layer2_out[793] = ~layer1_out[7118];
    assign layer2_out[794] = ~layer1_out[7768];
    assign layer2_out[795] = layer1_out[3276];
    assign layer2_out[796] = layer1_out[7291] & layer1_out[7292];
    assign layer2_out[797] = ~layer1_out[3697] | layer1_out[3696];
    assign layer2_out[798] = ~(layer1_out[7127] & layer1_out[7128]);
    assign layer2_out[799] = layer1_out[829] | layer1_out[830];
    assign layer2_out[800] = layer1_out[6871];
    assign layer2_out[801] = layer1_out[48] & layer1_out[49];
    assign layer2_out[802] = ~layer1_out[5557];
    assign layer2_out[803] = ~layer1_out[6396] | layer1_out[6397];
    assign layer2_out[804] = layer1_out[1361] & layer1_out[1362];
    assign layer2_out[805] = layer1_out[2284] & ~layer1_out[2283];
    assign layer2_out[806] = layer1_out[6880] & ~layer1_out[6879];
    assign layer2_out[807] = 1'b0;
    assign layer2_out[808] = ~layer1_out[5848] | layer1_out[5847];
    assign layer2_out[809] = layer1_out[2661];
    assign layer2_out[810] = ~layer1_out[4948] | layer1_out[4949];
    assign layer2_out[811] = layer1_out[2580];
    assign layer2_out[812] = ~layer1_out[4067];
    assign layer2_out[813] = layer1_out[5406];
    assign layer2_out[814] = layer1_out[6869] | layer1_out[6870];
    assign layer2_out[815] = layer1_out[5578];
    assign layer2_out[816] = layer1_out[7537];
    assign layer2_out[817] = ~layer1_out[5434];
    assign layer2_out[818] = layer1_out[22];
    assign layer2_out[819] = ~layer1_out[6470];
    assign layer2_out[820] = 1'b1;
    assign layer2_out[821] = layer1_out[1191];
    assign layer2_out[822] = layer1_out[6688] & ~layer1_out[6687];
    assign layer2_out[823] = layer1_out[5369] ^ layer1_out[5370];
    assign layer2_out[824] = layer1_out[109] & ~layer1_out[108];
    assign layer2_out[825] = ~layer1_out[5836];
    assign layer2_out[826] = layer1_out[2887];
    assign layer2_out[827] = layer1_out[1177] & layer1_out[1178];
    assign layer2_out[828] = layer1_out[3475] & ~layer1_out[3476];
    assign layer2_out[829] = layer1_out[225] ^ layer1_out[226];
    assign layer2_out[830] = layer1_out[2285] & layer1_out[2286];
    assign layer2_out[831] = ~layer1_out[3109];
    assign layer2_out[832] = ~layer1_out[5816] | layer1_out[5817];
    assign layer2_out[833] = layer1_out[7109];
    assign layer2_out[834] = ~(layer1_out[5049] | layer1_out[5050]);
    assign layer2_out[835] = layer1_out[927];
    assign layer2_out[836] = layer1_out[2300];
    assign layer2_out[837] = layer1_out[6845] & layer1_out[6846];
    assign layer2_out[838] = ~layer1_out[739];
    assign layer2_out[839] = layer1_out[1914] & ~layer1_out[1913];
    assign layer2_out[840] = ~layer1_out[7228] | layer1_out[7229];
    assign layer2_out[841] = layer1_out[3046] | layer1_out[3047];
    assign layer2_out[842] = ~(layer1_out[3153] | layer1_out[3154]);
    assign layer2_out[843] = ~(layer1_out[6310] ^ layer1_out[6311]);
    assign layer2_out[844] = ~(layer1_out[6598] ^ layer1_out[6599]);
    assign layer2_out[845] = ~(layer1_out[596] | layer1_out[597]);
    assign layer2_out[846] = layer1_out[5489] & layer1_out[5490];
    assign layer2_out[847] = ~layer1_out[7294];
    assign layer2_out[848] = layer1_out[4467];
    assign layer2_out[849] = layer1_out[1718] & ~layer1_out[1717];
    assign layer2_out[850] = layer1_out[7200];
    assign layer2_out[851] = layer1_out[5710] & layer1_out[5711];
    assign layer2_out[852] = ~layer1_out[5551] | layer1_out[5552];
    assign layer2_out[853] = ~(layer1_out[5766] & layer1_out[5767]);
    assign layer2_out[854] = layer1_out[3319] ^ layer1_out[3320];
    assign layer2_out[855] = layer1_out[2208];
    assign layer2_out[856] = ~(layer1_out[7211] & layer1_out[7212]);
    assign layer2_out[857] = 1'b1;
    assign layer2_out[858] = layer1_out[4037] & ~layer1_out[4036];
    assign layer2_out[859] = ~layer1_out[1771];
    assign layer2_out[860] = 1'b1;
    assign layer2_out[861] = layer1_out[6350];
    assign layer2_out[862] = ~layer1_out[1360];
    assign layer2_out[863] = layer1_out[3811] & ~layer1_out[3810];
    assign layer2_out[864] = 1'b0;
    assign layer2_out[865] = 1'b0;
    assign layer2_out[866] = layer1_out[7291];
    assign layer2_out[867] = layer1_out[5907] & ~layer1_out[5906];
    assign layer2_out[868] = layer1_out[7355];
    assign layer2_out[869] = layer1_out[4635];
    assign layer2_out[870] = ~layer1_out[4869] | layer1_out[4870];
    assign layer2_out[871] = ~layer1_out[1282] | layer1_out[1281];
    assign layer2_out[872] = layer1_out[4967] & layer1_out[4968];
    assign layer2_out[873] = layer1_out[2680] & ~layer1_out[2681];
    assign layer2_out[874] = ~layer1_out[3968];
    assign layer2_out[875] = ~(layer1_out[6473] & layer1_out[6474]);
    assign layer2_out[876] = layer1_out[276];
    assign layer2_out[877] = layer1_out[5155];
    assign layer2_out[878] = ~layer1_out[3258];
    assign layer2_out[879] = ~(layer1_out[432] ^ layer1_out[433]);
    assign layer2_out[880] = ~layer1_out[3701];
    assign layer2_out[881] = ~layer1_out[3025];
    assign layer2_out[882] = ~(layer1_out[3610] & layer1_out[3611]);
    assign layer2_out[883] = layer1_out[4076];
    assign layer2_out[884] = layer1_out[7071] & ~layer1_out[7070];
    assign layer2_out[885] = layer1_out[630];
    assign layer2_out[886] = layer1_out[7659] & ~layer1_out[7658];
    assign layer2_out[887] = ~layer1_out[6859];
    assign layer2_out[888] = ~layer1_out[429];
    assign layer2_out[889] = ~(layer1_out[1978] ^ layer1_out[1979]);
    assign layer2_out[890] = layer1_out[6129] & ~layer1_out[6130];
    assign layer2_out[891] = layer1_out[4208];
    assign layer2_out[892] = layer1_out[166] & ~layer1_out[165];
    assign layer2_out[893] = layer1_out[167] ^ layer1_out[168];
    assign layer2_out[894] = layer1_out[2976];
    assign layer2_out[895] = layer1_out[1260];
    assign layer2_out[896] = layer1_out[7786];
    assign layer2_out[897] = layer1_out[4950] & ~layer1_out[4951];
    assign layer2_out[898] = layer1_out[4165] | layer1_out[4166];
    assign layer2_out[899] = layer1_out[6329];
    assign layer2_out[900] = layer1_out[115] & layer1_out[116];
    assign layer2_out[901] = ~layer1_out[4350];
    assign layer2_out[902] = ~(layer1_out[478] & layer1_out[479]);
    assign layer2_out[903] = ~(layer1_out[7746] | layer1_out[7747]);
    assign layer2_out[904] = ~(layer1_out[4903] ^ layer1_out[4904]);
    assign layer2_out[905] = layer1_out[5002] & ~layer1_out[5003];
    assign layer2_out[906] = ~(layer1_out[3354] ^ layer1_out[3355]);
    assign layer2_out[907] = ~layer1_out[4872];
    assign layer2_out[908] = layer1_out[4354];
    assign layer2_out[909] = ~(layer1_out[6160] | layer1_out[6161]);
    assign layer2_out[910] = layer1_out[2920] & layer1_out[2921];
    assign layer2_out[911] = ~layer1_out[1121];
    assign layer2_out[912] = ~layer1_out[7112] | layer1_out[7111];
    assign layer2_out[913] = ~layer1_out[2597] | layer1_out[2596];
    assign layer2_out[914] = ~(layer1_out[2958] & layer1_out[2959]);
    assign layer2_out[915] = layer1_out[4982] & layer1_out[4983];
    assign layer2_out[916] = ~(layer1_out[3095] | layer1_out[3096]);
    assign layer2_out[917] = layer1_out[5940];
    assign layer2_out[918] = ~(layer1_out[4550] | layer1_out[4551]);
    assign layer2_out[919] = ~(layer1_out[7511] ^ layer1_out[7512]);
    assign layer2_out[920] = layer1_out[6130];
    assign layer2_out[921] = ~(layer1_out[7728] & layer1_out[7729]);
    assign layer2_out[922] = ~layer1_out[1763];
    assign layer2_out[923] = layer1_out[4741] ^ layer1_out[4742];
    assign layer2_out[924] = layer1_out[7525] & layer1_out[7526];
    assign layer2_out[925] = ~(layer1_out[1444] & layer1_out[1445]);
    assign layer2_out[926] = layer1_out[6285];
    assign layer2_out[927] = ~layer1_out[3142];
    assign layer2_out[928] = layer1_out[7012] | layer1_out[7013];
    assign layer2_out[929] = layer1_out[6882];
    assign layer2_out[930] = layer1_out[7068] & layer1_out[7069];
    assign layer2_out[931] = layer1_out[6914] & ~layer1_out[6915];
    assign layer2_out[932] = 1'b0;
    assign layer2_out[933] = layer1_out[5350];
    assign layer2_out[934] = 1'b0;
    assign layer2_out[935] = 1'b0;
    assign layer2_out[936] = ~layer1_out[939];
    assign layer2_out[937] = ~(layer1_out[2391] | layer1_out[2392]);
    assign layer2_out[938] = layer1_out[7286];
    assign layer2_out[939] = ~(layer1_out[5150] & layer1_out[5151]);
    assign layer2_out[940] = ~layer1_out[2259] | layer1_out[2260];
    assign layer2_out[941] = ~layer1_out[1478] | layer1_out[1477];
    assign layer2_out[942] = layer1_out[7614] & ~layer1_out[7615];
    assign layer2_out[943] = layer1_out[1354] | layer1_out[1355];
    assign layer2_out[944] = ~layer1_out[6105];
    assign layer2_out[945] = layer1_out[3586] & layer1_out[3587];
    assign layer2_out[946] = ~layer1_out[613];
    assign layer2_out[947] = 1'b0;
    assign layer2_out[948] = layer1_out[1370] & layer1_out[1371];
    assign layer2_out[949] = layer1_out[7609] & ~layer1_out[7610];
    assign layer2_out[950] = layer1_out[6481] & ~layer1_out[6482];
    assign layer2_out[951] = layer1_out[4330] & layer1_out[4331];
    assign layer2_out[952] = layer1_out[3661] | layer1_out[3662];
    assign layer2_out[953] = ~layer1_out[4911] | layer1_out[4912];
    assign layer2_out[954] = ~(layer1_out[4479] & layer1_out[4480]);
    assign layer2_out[955] = layer1_out[2977] & layer1_out[2978];
    assign layer2_out[956] = ~layer1_out[1835];
    assign layer2_out[957] = ~layer1_out[2039] | layer1_out[2038];
    assign layer2_out[958] = layer1_out[6952];
    assign layer2_out[959] = layer1_out[5909] & ~layer1_out[5910];
    assign layer2_out[960] = 1'b0;
    assign layer2_out[961] = layer1_out[235] & ~layer1_out[234];
    assign layer2_out[962] = layer1_out[1291] & layer1_out[1292];
    assign layer2_out[963] = layer1_out[707] | layer1_out[708];
    assign layer2_out[964] = ~layer1_out[5481];
    assign layer2_out[965] = layer1_out[606];
    assign layer2_out[966] = ~layer1_out[4945] | layer1_out[4944];
    assign layer2_out[967] = layer1_out[830] & ~layer1_out[831];
    assign layer2_out[968] = layer1_out[6329];
    assign layer2_out[969] = ~layer1_out[2960] | layer1_out[2959];
    assign layer2_out[970] = layer1_out[123];
    assign layer2_out[971] = ~layer1_out[2014] | layer1_out[2015];
    assign layer2_out[972] = layer1_out[173] & layer1_out[174];
    assign layer2_out[973] = layer1_out[3684] | layer1_out[3685];
    assign layer2_out[974] = layer1_out[5419] & layer1_out[5420];
    assign layer2_out[975] = ~layer1_out[3702];
    assign layer2_out[976] = layer1_out[3985];
    assign layer2_out[977] = ~layer1_out[6120];
    assign layer2_out[978] = 1'b1;
    assign layer2_out[979] = layer1_out[4549];
    assign layer2_out[980] = layer1_out[1649] | layer1_out[1650];
    assign layer2_out[981] = ~layer1_out[7829];
    assign layer2_out[982] = layer1_out[2493] | layer1_out[2494];
    assign layer2_out[983] = 1'b1;
    assign layer2_out[984] = layer1_out[1839];
    assign layer2_out[985] = ~(layer1_out[3345] ^ layer1_out[3346]);
    assign layer2_out[986] = ~layer1_out[7023];
    assign layer2_out[987] = layer1_out[4174];
    assign layer2_out[988] = ~(layer1_out[948] | layer1_out[949]);
    assign layer2_out[989] = layer1_out[4224] & ~layer1_out[4223];
    assign layer2_out[990] = layer1_out[2946] & layer1_out[2947];
    assign layer2_out[991] = ~(layer1_out[4095] & layer1_out[4096]);
    assign layer2_out[992] = ~(layer1_out[5719] | layer1_out[5720]);
    assign layer2_out[993] = layer1_out[7955] & ~layer1_out[7954];
    assign layer2_out[994] = layer1_out[6235];
    assign layer2_out[995] = ~(layer1_out[4069] ^ layer1_out[4070]);
    assign layer2_out[996] = layer1_out[3619] & ~layer1_out[3620];
    assign layer2_out[997] = layer1_out[670];
    assign layer2_out[998] = layer1_out[2472];
    assign layer2_out[999] = ~(layer1_out[1686] & layer1_out[1687]);
    assign layer2_out[1000] = ~layer1_out[452];
    assign layer2_out[1001] = ~layer1_out[7689];
    assign layer2_out[1002] = ~layer1_out[7821] | layer1_out[7822];
    assign layer2_out[1003] = ~layer1_out[1426] | layer1_out[1425];
    assign layer2_out[1004] = layer1_out[4588] & layer1_out[4589];
    assign layer2_out[1005] = ~layer1_out[3082];
    assign layer2_out[1006] = layer1_out[2435];
    assign layer2_out[1007] = layer1_out[2785];
    assign layer2_out[1008] = layer1_out[3145] | layer1_out[3146];
    assign layer2_out[1009] = ~layer1_out[7276];
    assign layer2_out[1010] = 1'b1;
    assign layer2_out[1011] = ~(layer1_out[3920] ^ layer1_out[3921]);
    assign layer2_out[1012] = layer1_out[6978];
    assign layer2_out[1013] = layer1_out[6541] ^ layer1_out[6542];
    assign layer2_out[1014] = ~layer1_out[7018];
    assign layer2_out[1015] = layer1_out[6180];
    assign layer2_out[1016] = ~layer1_out[7683];
    assign layer2_out[1017] = layer1_out[1013] & ~layer1_out[1012];
    assign layer2_out[1018] = layer1_out[7316] & ~layer1_out[7317];
    assign layer2_out[1019] = layer1_out[7357];
    assign layer2_out[1020] = ~(layer1_out[7997] & layer1_out[7998]);
    assign layer2_out[1021] = layer1_out[1900] & ~layer1_out[1899];
    assign layer2_out[1022] = 1'b0;
    assign layer2_out[1023] = ~layer1_out[2631] | layer1_out[2632];
    assign layer2_out[1024] = layer1_out[2804];
    assign layer2_out[1025] = layer1_out[2912] & ~layer1_out[2911];
    assign layer2_out[1026] = layer1_out[5413];
    assign layer2_out[1027] = layer1_out[1760];
    assign layer2_out[1028] = layer1_out[7449] | layer1_out[7450];
    assign layer2_out[1029] = layer1_out[543] | layer1_out[544];
    assign layer2_out[1030] = layer1_out[6043] & layer1_out[6044];
    assign layer2_out[1031] = ~layer1_out[5918];
    assign layer2_out[1032] = ~layer1_out[5306];
    assign layer2_out[1033] = layer1_out[4186] & ~layer1_out[4185];
    assign layer2_out[1034] = 1'b1;
    assign layer2_out[1035] = ~layer1_out[915] | layer1_out[914];
    assign layer2_out[1036] = ~(layer1_out[4418] | layer1_out[4419]);
    assign layer2_out[1037] = layer1_out[5801];
    assign layer2_out[1038] = ~layer1_out[5561];
    assign layer2_out[1039] = ~layer1_out[6536];
    assign layer2_out[1040] = layer1_out[3711] & layer1_out[3712];
    assign layer2_out[1041] = layer1_out[5987];
    assign layer2_out[1042] = ~layer1_out[7410] | layer1_out[7409];
    assign layer2_out[1043] = layer1_out[6567] & ~layer1_out[6566];
    assign layer2_out[1044] = layer1_out[6564] & ~layer1_out[6565];
    assign layer2_out[1045] = ~(layer1_out[5414] & layer1_out[5415]);
    assign layer2_out[1046] = ~(layer1_out[485] & layer1_out[486]);
    assign layer2_out[1047] = layer1_out[1638];
    assign layer2_out[1048] = layer1_out[2124];
    assign layer2_out[1049] = layer1_out[1119];
    assign layer2_out[1050] = ~layer1_out[7467];
    assign layer2_out[1051] = ~(layer1_out[440] & layer1_out[441]);
    assign layer2_out[1052] = layer1_out[2963] & ~layer1_out[2964];
    assign layer2_out[1053] = layer1_out[674] & ~layer1_out[675];
    assign layer2_out[1054] = layer1_out[2819] ^ layer1_out[2820];
    assign layer2_out[1055] = layer1_out[2648] | layer1_out[2649];
    assign layer2_out[1056] = layer1_out[6257] & ~layer1_out[6256];
    assign layer2_out[1057] = ~(layer1_out[1172] | layer1_out[1173]);
    assign layer2_out[1058] = ~layer1_out[1739] | layer1_out[1738];
    assign layer2_out[1059] = 1'b1;
    assign layer2_out[1060] = ~layer1_out[15];
    assign layer2_out[1061] = layer1_out[135] & layer1_out[136];
    assign layer2_out[1062] = layer1_out[3175] & ~layer1_out[3176];
    assign layer2_out[1063] = layer1_out[5575];
    assign layer2_out[1064] = layer1_out[1124];
    assign layer2_out[1065] = layer1_out[7812];
    assign layer2_out[1066] = 1'b0;
    assign layer2_out[1067] = ~(layer1_out[223] ^ layer1_out[224]);
    assign layer2_out[1068] = ~layer1_out[3560];
    assign layer2_out[1069] = ~layer1_out[7474] | layer1_out[7475];
    assign layer2_out[1070] = ~layer1_out[4817];
    assign layer2_out[1071] = layer1_out[6177];
    assign layer2_out[1072] = layer1_out[6784] ^ layer1_out[6785];
    assign layer2_out[1073] = ~layer1_out[5494];
    assign layer2_out[1074] = layer1_out[1589] & ~layer1_out[1590];
    assign layer2_out[1075] = layer1_out[4587] ^ layer1_out[4588];
    assign layer2_out[1076] = ~layer1_out[4193];
    assign layer2_out[1077] = layer1_out[7254];
    assign layer2_out[1078] = ~layer1_out[6512] | layer1_out[6513];
    assign layer2_out[1079] = layer1_out[7796] ^ layer1_out[7797];
    assign layer2_out[1080] = ~layer1_out[3194];
    assign layer2_out[1081] = layer1_out[566];
    assign layer2_out[1082] = ~(layer1_out[7175] & layer1_out[7176]);
    assign layer2_out[1083] = layer1_out[4854] | layer1_out[4855];
    assign layer2_out[1084] = ~layer1_out[6348];
    assign layer2_out[1085] = layer1_out[831] & ~layer1_out[832];
    assign layer2_out[1086] = ~(layer1_out[203] | layer1_out[204]);
    assign layer2_out[1087] = layer1_out[6037];
    assign layer2_out[1088] = ~layer1_out[71];
    assign layer2_out[1089] = ~layer1_out[2143];
    assign layer2_out[1090] = ~layer1_out[2527];
    assign layer2_out[1091] = ~layer1_out[2191];
    assign layer2_out[1092] = ~layer1_out[2462];
    assign layer2_out[1093] = ~layer1_out[4758];
    assign layer2_out[1094] = ~(layer1_out[3977] & layer1_out[3978]);
    assign layer2_out[1095] = ~layer1_out[6115] | layer1_out[6116];
    assign layer2_out[1096] = layer1_out[5628];
    assign layer2_out[1097] = layer1_out[1338] & ~layer1_out[1339];
    assign layer2_out[1098] = layer1_out[1998] | layer1_out[1999];
    assign layer2_out[1099] = layer1_out[961] | layer1_out[962];
    assign layer2_out[1100] = ~layer1_out[3808];
    assign layer2_out[1101] = ~layer1_out[4633];
    assign layer2_out[1102] = ~layer1_out[4522] | layer1_out[4521];
    assign layer2_out[1103] = ~layer1_out[293] | layer1_out[294];
    assign layer2_out[1104] = layer1_out[3536] | layer1_out[3537];
    assign layer2_out[1105] = ~layer1_out[5028] | layer1_out[5027];
    assign layer2_out[1106] = ~(layer1_out[5675] | layer1_out[5676]);
    assign layer2_out[1107] = ~layer1_out[5402];
    assign layer2_out[1108] = ~layer1_out[7279];
    assign layer2_out[1109] = layer1_out[542];
    assign layer2_out[1110] = ~layer1_out[1113];
    assign layer2_out[1111] = layer1_out[4176] & ~layer1_out[4175];
    assign layer2_out[1112] = layer1_out[4547] ^ layer1_out[4548];
    assign layer2_out[1113] = ~(layer1_out[5717] ^ layer1_out[5718]);
    assign layer2_out[1114] = ~layer1_out[5360];
    assign layer2_out[1115] = layer1_out[1407] & ~layer1_out[1406];
    assign layer2_out[1116] = ~(layer1_out[2627] | layer1_out[2628]);
    assign layer2_out[1117] = ~(layer1_out[753] | layer1_out[754]);
    assign layer2_out[1118] = layer1_out[7817] & ~layer1_out[7816];
    assign layer2_out[1119] = layer1_out[1596];
    assign layer2_out[1120] = ~layer1_out[5183];
    assign layer2_out[1121] = layer1_out[5790];
    assign layer2_out[1122] = layer1_out[4293] & ~layer1_out[4292];
    assign layer2_out[1123] = ~layer1_out[7520];
    assign layer2_out[1124] = layer1_out[1729];
    assign layer2_out[1125] = layer1_out[5621] | layer1_out[5622];
    assign layer2_out[1126] = layer1_out[6787] | layer1_out[6788];
    assign layer2_out[1127] = ~layer1_out[3488];
    assign layer2_out[1128] = ~layer1_out[4514];
    assign layer2_out[1129] = ~(layer1_out[7877] | layer1_out[7878]);
    assign layer2_out[1130] = ~(layer1_out[3541] ^ layer1_out[3542]);
    assign layer2_out[1131] = layer1_out[6944];
    assign layer2_out[1132] = ~layer1_out[4900] | layer1_out[4899];
    assign layer2_out[1133] = ~(layer1_out[2838] & layer1_out[2839]);
    assign layer2_out[1134] = ~(layer1_out[3674] ^ layer1_out[3675]);
    assign layer2_out[1135] = ~layer1_out[1256];
    assign layer2_out[1136] = ~layer1_out[2944];
    assign layer2_out[1137] = layer1_out[3678];
    assign layer2_out[1138] = ~layer1_out[4358];
    assign layer2_out[1139] = layer1_out[1660] & ~layer1_out[1659];
    assign layer2_out[1140] = ~(layer1_out[510] & layer1_out[511]);
    assign layer2_out[1141] = ~(layer1_out[5190] ^ layer1_out[5191]);
    assign layer2_out[1142] = ~layer1_out[1847];
    assign layer2_out[1143] = layer1_out[4401];
    assign layer2_out[1144] = ~(layer1_out[6582] | layer1_out[6583]);
    assign layer2_out[1145] = layer1_out[1027];
    assign layer2_out[1146] = layer1_out[5170];
    assign layer2_out[1147] = layer1_out[7902];
    assign layer2_out[1148] = 1'b0;
    assign layer2_out[1149] = layer1_out[1112] & ~layer1_out[1111];
    assign layer2_out[1150] = ~layer1_out[2483];
    assign layer2_out[1151] = ~layer1_out[4879] | layer1_out[4878];
    assign layer2_out[1152] = layer1_out[4398] | layer1_out[4399];
    assign layer2_out[1153] = ~(layer1_out[7473] & layer1_out[7474]);
    assign layer2_out[1154] = layer1_out[1326];
    assign layer2_out[1155] = layer1_out[2168];
    assign layer2_out[1156] = ~(layer1_out[3072] ^ layer1_out[3073]);
    assign layer2_out[1157] = 1'b1;
    assign layer2_out[1158] = ~(layer1_out[7576] & layer1_out[7577]);
    assign layer2_out[1159] = ~(layer1_out[5089] ^ layer1_out[5090]);
    assign layer2_out[1160] = ~layer1_out[5021];
    assign layer2_out[1161] = layer1_out[5447];
    assign layer2_out[1162] = layer1_out[5232] & ~layer1_out[5231];
    assign layer2_out[1163] = ~layer1_out[2510];
    assign layer2_out[1164] = layer1_out[3119];
    assign layer2_out[1165] = layer1_out[6657] & ~layer1_out[6656];
    assign layer2_out[1166] = ~layer1_out[1583];
    assign layer2_out[1167] = layer1_out[6283] & layer1_out[6284];
    assign layer2_out[1168] = ~layer1_out[2493] | layer1_out[2492];
    assign layer2_out[1169] = layer1_out[6041];
    assign layer2_out[1170] = layer1_out[2695];
    assign layer2_out[1171] = ~layer1_out[171];
    assign layer2_out[1172] = layer1_out[1209];
    assign layer2_out[1173] = ~layer1_out[6316];
    assign layer2_out[1174] = layer1_out[3583] & layer1_out[3584];
    assign layer2_out[1175] = layer1_out[7886] & ~layer1_out[7885];
    assign layer2_out[1176] = ~layer1_out[2192] | layer1_out[2193];
    assign layer2_out[1177] = layer1_out[4433] & ~layer1_out[4434];
    assign layer2_out[1178] = layer1_out[1008] | layer1_out[1009];
    assign layer2_out[1179] = layer1_out[2248];
    assign layer2_out[1180] = 1'b0;
    assign layer2_out[1181] = ~layer1_out[2339];
    assign layer2_out[1182] = 1'b0;
    assign layer2_out[1183] = ~layer1_out[5335] | layer1_out[5336];
    assign layer2_out[1184] = layer1_out[6774] & ~layer1_out[6775];
    assign layer2_out[1185] = ~layer1_out[6854];
    assign layer2_out[1186] = ~(layer1_out[3614] & layer1_out[3615]);
    assign layer2_out[1187] = layer1_out[5315] ^ layer1_out[5316];
    assign layer2_out[1188] = layer1_out[2478] & ~layer1_out[2479];
    assign layer2_out[1189] = layer1_out[1550];
    assign layer2_out[1190] = layer1_out[2512];
    assign layer2_out[1191] = ~(layer1_out[4611] & layer1_out[4612]);
    assign layer2_out[1192] = ~layer1_out[5299] | layer1_out[5298];
    assign layer2_out[1193] = ~(layer1_out[868] | layer1_out[869]);
    assign layer2_out[1194] = layer1_out[2221] ^ layer1_out[2222];
    assign layer2_out[1195] = layer1_out[6729] & layer1_out[6730];
    assign layer2_out[1196] = ~layer1_out[182];
    assign layer2_out[1197] = layer1_out[2364];
    assign layer2_out[1198] = layer1_out[4180] | layer1_out[4181];
    assign layer2_out[1199] = layer1_out[282] | layer1_out[283];
    assign layer2_out[1200] = layer1_out[6409];
    assign layer2_out[1201] = ~(layer1_out[6931] & layer1_out[6932]);
    assign layer2_out[1202] = layer1_out[1026] & ~layer1_out[1025];
    assign layer2_out[1203] = ~(layer1_out[7934] ^ layer1_out[7935]);
    assign layer2_out[1204] = ~layer1_out[6259] | layer1_out[6258];
    assign layer2_out[1205] = layer1_out[316];
    assign layer2_out[1206] = ~layer1_out[7403];
    assign layer2_out[1207] = ~layer1_out[557];
    assign layer2_out[1208] = layer1_out[4439] & layer1_out[4440];
    assign layer2_out[1209] = layer1_out[3781];
    assign layer2_out[1210] = ~layer1_out[1762];
    assign layer2_out[1211] = layer1_out[6062];
    assign layer2_out[1212] = ~layer1_out[6514];
    assign layer2_out[1213] = layer1_out[3332];
    assign layer2_out[1214] = ~layer1_out[7772] | layer1_out[7771];
    assign layer2_out[1215] = ~layer1_out[5153];
    assign layer2_out[1216] = layer1_out[3529] & ~layer1_out[3528];
    assign layer2_out[1217] = layer1_out[7460];
    assign layer2_out[1218] = layer1_out[3094];
    assign layer2_out[1219] = ~(layer1_out[5180] & layer1_out[5181]);
    assign layer2_out[1220] = ~layer1_out[5056] | layer1_out[5057];
    assign layer2_out[1221] = ~layer1_out[7676] | layer1_out[7677];
    assign layer2_out[1222] = ~layer1_out[2172] | layer1_out[2173];
    assign layer2_out[1223] = ~layer1_out[4236];
    assign layer2_out[1224] = layer1_out[2705] & ~layer1_out[2706];
    assign layer2_out[1225] = layer1_out[3377];
    assign layer2_out[1226] = ~layer1_out[2099];
    assign layer2_out[1227] = ~(layer1_out[3011] | layer1_out[3012]);
    assign layer2_out[1228] = layer1_out[3589] & layer1_out[3590];
    assign layer2_out[1229] = ~(layer1_out[5380] & layer1_out[5381]);
    assign layer2_out[1230] = ~layer1_out[4866];
    assign layer2_out[1231] = layer1_out[4484] & ~layer1_out[4483];
    assign layer2_out[1232] = layer1_out[4993] & layer1_out[4994];
    assign layer2_out[1233] = ~layer1_out[7394];
    assign layer2_out[1234] = ~(layer1_out[134] & layer1_out[135]);
    assign layer2_out[1235] = layer1_out[6461] & ~layer1_out[6462];
    assign layer2_out[1236] = layer1_out[1719] & layer1_out[1720];
    assign layer2_out[1237] = ~layer1_out[5003] | layer1_out[5004];
    assign layer2_out[1238] = ~layer1_out[3995] | layer1_out[3994];
    assign layer2_out[1239] = ~(layer1_out[7839] | layer1_out[7840]);
    assign layer2_out[1240] = ~layer1_out[5515] | layer1_out[5516];
    assign layer2_out[1241] = ~layer1_out[1655];
    assign layer2_out[1242] = layer1_out[5397] & ~layer1_out[5396];
    assign layer2_out[1243] = layer1_out[2086] | layer1_out[2087];
    assign layer2_out[1244] = ~layer1_out[4114] | layer1_out[4113];
    assign layer2_out[1245] = ~(layer1_out[5733] | layer1_out[5734]);
    assign layer2_out[1246] = ~layer1_out[2303];
    assign layer2_out[1247] = ~(layer1_out[5496] | layer1_out[5497]);
    assign layer2_out[1248] = layer1_out[3318];
    assign layer2_out[1249] = layer1_out[1635] & ~layer1_out[1634];
    assign layer2_out[1250] = ~layer1_out[7187] | layer1_out[7186];
    assign layer2_out[1251] = layer1_out[3840] & layer1_out[3841];
    assign layer2_out[1252] = layer1_out[2378];
    assign layer2_out[1253] = ~layer1_out[4254] | layer1_out[4255];
    assign layer2_out[1254] = ~layer1_out[7259] | layer1_out[7260];
    assign layer2_out[1255] = ~layer1_out[466];
    assign layer2_out[1256] = ~layer1_out[6052];
    assign layer2_out[1257] = ~layer1_out[6639] | layer1_out[6640];
    assign layer2_out[1258] = ~(layer1_out[3207] | layer1_out[3208]);
    assign layer2_out[1259] = layer1_out[6254] & layer1_out[6255];
    assign layer2_out[1260] = layer1_out[7223];
    assign layer2_out[1261] = layer1_out[5975] | layer1_out[5976];
    assign layer2_out[1262] = ~layer1_out[7379] | layer1_out[7380];
    assign layer2_out[1263] = ~layer1_out[4412] | layer1_out[4413];
    assign layer2_out[1264] = layer1_out[136] & layer1_out[137];
    assign layer2_out[1265] = layer1_out[4929] & ~layer1_out[4928];
    assign layer2_out[1266] = layer1_out[7335] ^ layer1_out[7336];
    assign layer2_out[1267] = ~layer1_out[1500];
    assign layer2_out[1268] = 1'b0;
    assign layer2_out[1269] = 1'b1;
    assign layer2_out[1270] = 1'b1;
    assign layer2_out[1271] = layer1_out[2102];
    assign layer2_out[1272] = ~layer1_out[4952];
    assign layer2_out[1273] = ~(layer1_out[4857] | layer1_out[4858]);
    assign layer2_out[1274] = ~layer1_out[5186] | layer1_out[5187];
    assign layer2_out[1275] = 1'b0;
    assign layer2_out[1276] = layer1_out[3048] | layer1_out[3049];
    assign layer2_out[1277] = layer1_out[1470] ^ layer1_out[1471];
    assign layer2_out[1278] = ~layer1_out[5305];
    assign layer2_out[1279] = layer1_out[2502] & layer1_out[2503];
    assign layer2_out[1280] = ~(layer1_out[5768] ^ layer1_out[5769]);
    assign layer2_out[1281] = layer1_out[4089];
    assign layer2_out[1282] = ~layer1_out[3411];
    assign layer2_out[1283] = ~layer1_out[7517] | layer1_out[7518];
    assign layer2_out[1284] = layer1_out[3162] & ~layer1_out[3163];
    assign layer2_out[1285] = layer1_out[6492] & ~layer1_out[6491];
    assign layer2_out[1286] = layer1_out[1306] & layer1_out[1307];
    assign layer2_out[1287] = layer1_out[6407] & ~layer1_out[6408];
    assign layer2_out[1288] = layer1_out[6277];
    assign layer2_out[1289] = layer1_out[6879];
    assign layer2_out[1290] = ~layer1_out[6186];
    assign layer2_out[1291] = layer1_out[209] & layer1_out[210];
    assign layer2_out[1292] = ~layer1_out[3724];
    assign layer2_out[1293] = layer1_out[3400] | layer1_out[3401];
    assign layer2_out[1294] = ~layer1_out[3561];
    assign layer2_out[1295] = ~(layer1_out[6875] | layer1_out[6876]);
    assign layer2_out[1296] = layer1_out[6822] & layer1_out[6823];
    assign layer2_out[1297] = ~(layer1_out[1923] & layer1_out[1924]);
    assign layer2_out[1298] = layer1_out[4201] & ~layer1_out[4202];
    assign layer2_out[1299] = ~layer1_out[5343];
    assign layer2_out[1300] = ~(layer1_out[5240] & layer1_out[5241]);
    assign layer2_out[1301] = ~layer1_out[3391] | layer1_out[3392];
    assign layer2_out[1302] = ~layer1_out[4601];
    assign layer2_out[1303] = layer1_out[7298] & layer1_out[7299];
    assign layer2_out[1304] = ~layer1_out[7625] | layer1_out[7626];
    assign layer2_out[1305] = layer1_out[1122] | layer1_out[1123];
    assign layer2_out[1306] = layer1_out[2021] & ~layer1_out[2020];
    assign layer2_out[1307] = ~layer1_out[3997];
    assign layer2_out[1308] = ~layer1_out[5235] | layer1_out[5234];
    assign layer2_out[1309] = ~(layer1_out[6306] & layer1_out[6307]);
    assign layer2_out[1310] = ~layer1_out[6417] | layer1_out[6416];
    assign layer2_out[1311] = layer1_out[7926];
    assign layer2_out[1312] = ~layer1_out[3809];
    assign layer2_out[1313] = layer1_out[2906];
    assign layer2_out[1314] = ~(layer1_out[7732] ^ layer1_out[7733]);
    assign layer2_out[1315] = layer1_out[5008];
    assign layer2_out[1316] = layer1_out[2590] ^ layer1_out[2591];
    assign layer2_out[1317] = ~layer1_out[7258] | layer1_out[7259];
    assign layer2_out[1318] = ~layer1_out[4135] | layer1_out[4136];
    assign layer2_out[1319] = ~(layer1_out[3456] ^ layer1_out[3457]);
    assign layer2_out[1320] = ~layer1_out[5049] | layer1_out[5048];
    assign layer2_out[1321] = ~layer1_out[5629] | layer1_out[5630];
    assign layer2_out[1322] = layer1_out[5149] & layer1_out[5150];
    assign layer2_out[1323] = ~layer1_out[7207];
    assign layer2_out[1324] = layer1_out[1170];
    assign layer2_out[1325] = ~layer1_out[212];
    assign layer2_out[1326] = layer1_out[7989];
    assign layer2_out[1327] = 1'b0;
    assign layer2_out[1328] = layer1_out[6374] & layer1_out[6375];
    assign layer2_out[1329] = ~layer1_out[1089] | layer1_out[1090];
    assign layer2_out[1330] = layer1_out[7408] & layer1_out[7409];
    assign layer2_out[1331] = layer1_out[1931] ^ layer1_out[1932];
    assign layer2_out[1332] = ~layer1_out[585];
    assign layer2_out[1333] = ~layer1_out[1814];
    assign layer2_out[1334] = ~(layer1_out[2255] & layer1_out[2256]);
    assign layer2_out[1335] = ~layer1_out[7719];
    assign layer2_out[1336] = layer1_out[1646] | layer1_out[1647];
    assign layer2_out[1337] = ~(layer1_out[7726] | layer1_out[7727]);
    assign layer2_out[1338] = layer1_out[4398];
    assign layer2_out[1339] = layer1_out[1437] & layer1_out[1438];
    assign layer2_out[1340] = ~layer1_out[656];
    assign layer2_out[1341] = 1'b0;
    assign layer2_out[1342] = ~layer1_out[6279];
    assign layer2_out[1343] = ~(layer1_out[5372] & layer1_out[5373]);
    assign layer2_out[1344] = layer1_out[2996] | layer1_out[2997];
    assign layer2_out[1345] = layer1_out[371] & ~layer1_out[372];
    assign layer2_out[1346] = ~layer1_out[6655];
    assign layer2_out[1347] = layer1_out[6986] | layer1_out[6987];
    assign layer2_out[1348] = ~layer1_out[660];
    assign layer2_out[1349] = ~layer1_out[2501];
    assign layer2_out[1350] = layer1_out[6061];
    assign layer2_out[1351] = layer1_out[4932];
    assign layer2_out[1352] = layer1_out[3659] | layer1_out[3660];
    assign layer2_out[1353] = layer1_out[6940];
    assign layer2_out[1354] = layer1_out[2896] ^ layer1_out[2897];
    assign layer2_out[1355] = layer1_out[2797] & ~layer1_out[2796];
    assign layer2_out[1356] = ~layer1_out[4503];
    assign layer2_out[1357] = layer1_out[2401] & layer1_out[2402];
    assign layer2_out[1358] = layer1_out[2614] & ~layer1_out[2613];
    assign layer2_out[1359] = ~layer1_out[821];
    assign layer2_out[1360] = layer1_out[147] & ~layer1_out[146];
    assign layer2_out[1361] = ~layer1_out[5032] | layer1_out[5031];
    assign layer2_out[1362] = ~(layer1_out[3741] & layer1_out[3742]);
    assign layer2_out[1363] = ~(layer1_out[6593] | layer1_out[6594]);
    assign layer2_out[1364] = ~layer1_out[4063];
    assign layer2_out[1365] = layer1_out[4038];
    assign layer2_out[1366] = layer1_out[7422];
    assign layer2_out[1367] = ~layer1_out[7407];
    assign layer2_out[1368] = layer1_out[6612];
    assign layer2_out[1369] = ~layer1_out[278] | layer1_out[279];
    assign layer2_out[1370] = ~(layer1_out[3516] & layer1_out[3517]);
    assign layer2_out[1371] = ~layer1_out[5431] | layer1_out[5432];
    assign layer2_out[1372] = layer1_out[2275] & ~layer1_out[2276];
    assign layer2_out[1373] = layer1_out[5032] | layer1_out[5033];
    assign layer2_out[1374] = layer1_out[517];
    assign layer2_out[1375] = ~(layer1_out[1786] ^ layer1_out[1787]);
    assign layer2_out[1376] = layer1_out[5919] ^ layer1_out[5920];
    assign layer2_out[1377] = ~layer1_out[7261];
    assign layer2_out[1378] = ~layer1_out[1520];
    assign layer2_out[1379] = ~layer1_out[6159];
    assign layer2_out[1380] = ~(layer1_out[1774] ^ layer1_out[1775]);
    assign layer2_out[1381] = ~(layer1_out[5257] ^ layer1_out[5258]);
    assign layer2_out[1382] = layer1_out[1764] & layer1_out[1765];
    assign layer2_out[1383] = ~layer1_out[3665];
    assign layer2_out[1384] = layer1_out[3807];
    assign layer2_out[1385] = ~(layer1_out[3875] | layer1_out[3876]);
    assign layer2_out[1386] = ~layer1_out[2268];
    assign layer2_out[1387] = layer1_out[296] ^ layer1_out[297];
    assign layer2_out[1388] = ~layer1_out[6581];
    assign layer2_out[1389] = layer1_out[3506] & layer1_out[3507];
    assign layer2_out[1390] = ~layer1_out[6707];
    assign layer2_out[1391] = layer1_out[1962] & ~layer1_out[1961];
    assign layer2_out[1392] = layer1_out[7121] ^ layer1_out[7122];
    assign layer2_out[1393] = ~(layer1_out[5574] ^ layer1_out[5575]);
    assign layer2_out[1394] = ~layer1_out[4183];
    assign layer2_out[1395] = layer1_out[529] & ~layer1_out[530];
    assign layer2_out[1396] = ~layer1_out[2673] | layer1_out[2674];
    assign layer2_out[1397] = ~(layer1_out[3866] ^ layer1_out[3867]);
    assign layer2_out[1398] = ~layer1_out[4236];
    assign layer2_out[1399] = ~(layer1_out[143] | layer1_out[144]);
    assign layer2_out[1400] = layer1_out[7939] & ~layer1_out[7940];
    assign layer2_out[1401] = ~(layer1_out[7451] | layer1_out[7452]);
    assign layer2_out[1402] = layer1_out[5866] & ~layer1_out[5865];
    assign layer2_out[1403] = layer1_out[5568] & ~layer1_out[5569];
    assign layer2_out[1404] = ~layer1_out[4937] | layer1_out[4936];
    assign layer2_out[1405] = ~(layer1_out[7477] & layer1_out[7478]);
    assign layer2_out[1406] = ~(layer1_out[4554] | layer1_out[4555]);
    assign layer2_out[1407] = layer1_out[5778] & ~layer1_out[5777];
    assign layer2_out[1408] = ~layer1_out[2605];
    assign layer2_out[1409] = ~layer1_out[3467];
    assign layer2_out[1410] = layer1_out[6290] & ~layer1_out[6289];
    assign layer2_out[1411] = layer1_out[2960] & layer1_out[2961];
    assign layer2_out[1412] = ~layer1_out[2753];
    assign layer2_out[1413] = layer1_out[1412] & layer1_out[1413];
    assign layer2_out[1414] = ~layer1_out[6432];
    assign layer2_out[1415] = ~(layer1_out[7530] & layer1_out[7531]);
    assign layer2_out[1416] = layer1_out[7889] & layer1_out[7890];
    assign layer2_out[1417] = layer1_out[129] | layer1_out[130];
    assign layer2_out[1418] = layer1_out[2406] | layer1_out[2407];
    assign layer2_out[1419] = layer1_out[4109] & ~layer1_out[4110];
    assign layer2_out[1420] = ~layer1_out[2975];
    assign layer2_out[1421] = ~layer1_out[523];
    assign layer2_out[1422] = ~layer1_out[545];
    assign layer2_out[1423] = layer1_out[4344];
    assign layer2_out[1424] = ~layer1_out[4809] | layer1_out[4810];
    assign layer2_out[1425] = layer1_out[4039] & ~layer1_out[4040];
    assign layer2_out[1426] = ~(layer1_out[4021] & layer1_out[4022]);
    assign layer2_out[1427] = layer1_out[424] ^ layer1_out[425];
    assign layer2_out[1428] = 1'b0;
    assign layer2_out[1429] = layer1_out[2196];
    assign layer2_out[1430] = layer1_out[1963];
    assign layer2_out[1431] = 1'b0;
    assign layer2_out[1432] = ~(layer1_out[5388] & layer1_out[5389]);
    assign layer2_out[1433] = layer1_out[5206] | layer1_out[5207];
    assign layer2_out[1434] = ~layer1_out[131];
    assign layer2_out[1435] = layer1_out[389] | layer1_out[390];
    assign layer2_out[1436] = layer1_out[5526] & ~layer1_out[5525];
    assign layer2_out[1437] = ~layer1_out[3978];
    assign layer2_out[1438] = layer1_out[2798];
    assign layer2_out[1439] = layer1_out[1894];
    assign layer2_out[1440] = layer1_out[3320];
    assign layer2_out[1441] = ~(layer1_out[2463] & layer1_out[2464]);
    assign layer2_out[1442] = ~(layer1_out[874] | layer1_out[875]);
    assign layer2_out[1443] = layer1_out[2019] | layer1_out[2020];
    assign layer2_out[1444] = ~layer1_out[4116];
    assign layer2_out[1445] = ~(layer1_out[6453] ^ layer1_out[6454]);
    assign layer2_out[1446] = ~layer1_out[6714] | layer1_out[6713];
    assign layer2_out[1447] = layer1_out[7722];
    assign layer2_out[1448] = ~(layer1_out[2193] ^ layer1_out[2194]);
    assign layer2_out[1449] = layer1_out[778];
    assign layer2_out[1450] = ~layer1_out[7161];
    assign layer2_out[1451] = layer1_out[1413] | layer1_out[1414];
    assign layer2_out[1452] = ~layer1_out[911];
    assign layer2_out[1453] = ~layer1_out[6370] | layer1_out[6371];
    assign layer2_out[1454] = ~layer1_out[6300];
    assign layer2_out[1455] = ~layer1_out[6283] | layer1_out[6282];
    assign layer2_out[1456] = 1'b1;
    assign layer2_out[1457] = layer1_out[4705];
    assign layer2_out[1458] = layer1_out[3707];
    assign layer2_out[1459] = ~layer1_out[4215] | layer1_out[4214];
    assign layer2_out[1460] = layer1_out[5073] & ~layer1_out[5072];
    assign layer2_out[1461] = ~layer1_out[3366];
    assign layer2_out[1462] = 1'b1;
    assign layer2_out[1463] = layer1_out[549] & layer1_out[550];
    assign layer2_out[1464] = ~(layer1_out[3512] & layer1_out[3513]);
    assign layer2_out[1465] = ~layer1_out[5704];
    assign layer2_out[1466] = ~layer1_out[5076];
    assign layer2_out[1467] = layer1_out[3380] | layer1_out[3381];
    assign layer2_out[1468] = layer1_out[3737] | layer1_out[3738];
    assign layer2_out[1469] = layer1_out[2670] & layer1_out[2671];
    assign layer2_out[1470] = ~layer1_out[1760];
    assign layer2_out[1471] = layer1_out[6908] | layer1_out[6909];
    assign layer2_out[1472] = layer1_out[1874];
    assign layer2_out[1473] = layer1_out[3563];
    assign layer2_out[1474] = layer1_out[5671];
    assign layer2_out[1475] = ~layer1_out[4477];
    assign layer2_out[1476] = layer1_out[2824];
    assign layer2_out[1477] = ~layer1_out[6438];
    assign layer2_out[1478] = ~layer1_out[4269];
    assign layer2_out[1479] = layer1_out[3395];
    assign layer2_out[1480] = layer1_out[4411];
    assign layer2_out[1481] = ~layer1_out[4680];
    assign layer2_out[1482] = layer1_out[1063] & ~layer1_out[1062];
    assign layer2_out[1483] = ~layer1_out[7173] | layer1_out[7174];
    assign layer2_out[1484] = layer1_out[2732] & layer1_out[2733];
    assign layer2_out[1485] = layer1_out[4986] & ~layer1_out[4985];
    assign layer2_out[1486] = ~(layer1_out[5751] & layer1_out[5752]);
    assign layer2_out[1487] = layer1_out[1795] | layer1_out[1796];
    assign layer2_out[1488] = layer1_out[3277];
    assign layer2_out[1489] = 1'b1;
    assign layer2_out[1490] = ~layer1_out[7252];
    assign layer2_out[1491] = layer1_out[5438] & ~layer1_out[5437];
    assign layer2_out[1492] = ~layer1_out[4138];
    assign layer2_out[1493] = layer1_out[4737];
    assign layer2_out[1494] = ~layer1_out[2291];
    assign layer2_out[1495] = layer1_out[7425] & ~layer1_out[7424];
    assign layer2_out[1496] = ~(layer1_out[863] | layer1_out[864]);
    assign layer2_out[1497] = ~(layer1_out[6616] & layer1_out[6617]);
    assign layer2_out[1498] = ~layer1_out[335];
    assign layer2_out[1499] = layer1_out[2356];
    assign layer2_out[1500] = layer1_out[1927];
    assign layer2_out[1501] = layer1_out[5547];
    assign layer2_out[1502] = layer1_out[2576] ^ layer1_out[2577];
    assign layer2_out[1503] = ~(layer1_out[3629] & layer1_out[3630]);
    assign layer2_out[1504] = ~(layer1_out[2755] & layer1_out[2756]);
    assign layer2_out[1505] = layer1_out[3966];
    assign layer2_out[1506] = ~layer1_out[2164] | layer1_out[2163];
    assign layer2_out[1507] = layer1_out[7806] & ~layer1_out[7807];
    assign layer2_out[1508] = layer1_out[99] ^ layer1_out[100];
    assign layer2_out[1509] = layer1_out[877] & ~layer1_out[878];
    assign layer2_out[1510] = layer1_out[3200] | layer1_out[3201];
    assign layer2_out[1511] = layer1_out[1990] & layer1_out[1991];
    assign layer2_out[1512] = ~(layer1_out[1387] & layer1_out[1388]);
    assign layer2_out[1513] = layer1_out[553] ^ layer1_out[554];
    assign layer2_out[1514] = layer1_out[1015] & layer1_out[1016];
    assign layer2_out[1515] = layer1_out[4551] & ~layer1_out[4552];
    assign layer2_out[1516] = ~layer1_out[75];
    assign layer2_out[1517] = layer1_out[7627] | layer1_out[7628];
    assign layer2_out[1518] = ~layer1_out[2004];
    assign layer2_out[1519] = ~(layer1_out[5064] & layer1_out[5065]);
    assign layer2_out[1520] = layer1_out[865] & layer1_out[866];
    assign layer2_out[1521] = layer1_out[1848];
    assign layer2_out[1522] = ~layer1_out[431];
    assign layer2_out[1523] = ~layer1_out[5158];
    assign layer2_out[1524] = ~layer1_out[1104] | layer1_out[1103];
    assign layer2_out[1525] = layer1_out[6723];
    assign layer2_out[1526] = ~(layer1_out[4447] | layer1_out[4448]);
    assign layer2_out[1527] = layer1_out[6889] & ~layer1_out[6890];
    assign layer2_out[1528] = layer1_out[4130];
    assign layer2_out[1529] = layer1_out[35] | layer1_out[36];
    assign layer2_out[1530] = layer1_out[3557] & ~layer1_out[3558];
    assign layer2_out[1531] = ~layer1_out[3615] | layer1_out[3616];
    assign layer2_out[1532] = ~layer1_out[5870] | layer1_out[5869];
    assign layer2_out[1533] = layer1_out[768];
    assign layer2_out[1534] = ~(layer1_out[3386] & layer1_out[3387]);
    assign layer2_out[1535] = layer1_out[6898];
    assign layer2_out[1536] = ~(layer1_out[3261] ^ layer1_out[3262]);
    assign layer2_out[1537] = layer1_out[2584] & ~layer1_out[2583];
    assign layer2_out[1538] = layer1_out[7937];
    assign layer2_out[1539] = ~layer1_out[6027] | layer1_out[6028];
    assign layer2_out[1540] = ~layer1_out[6467];
    assign layer2_out[1541] = ~layer1_out[6007];
    assign layer2_out[1542] = layer1_out[5251];
    assign layer2_out[1543] = ~(layer1_out[904] | layer1_out[905]);
    assign layer2_out[1544] = ~(layer1_out[4064] | layer1_out[4065]);
    assign layer2_out[1545] = layer1_out[2423] & layer1_out[2424];
    assign layer2_out[1546] = layer1_out[4585] & ~layer1_out[4586];
    assign layer2_out[1547] = layer1_out[7926] & layer1_out[7927];
    assign layer2_out[1548] = layer1_out[2455];
    assign layer2_out[1549] = ~layer1_out[3637];
    assign layer2_out[1550] = layer1_out[6383] ^ layer1_out[6384];
    assign layer2_out[1551] = layer1_out[926] & layer1_out[927];
    assign layer2_out[1552] = layer1_out[4430] & ~layer1_out[4429];
    assign layer2_out[1553] = layer1_out[883] | layer1_out[884];
    assign layer2_out[1554] = ~layer1_out[5979];
    assign layer2_out[1555] = 1'b1;
    assign layer2_out[1556] = ~layer1_out[5250];
    assign layer2_out[1557] = layer1_out[6607];
    assign layer2_out[1558] = ~layer1_out[5579] | layer1_out[5578];
    assign layer2_out[1559] = layer1_out[7873];
    assign layer2_out[1560] = layer1_out[2037] & ~layer1_out[2038];
    assign layer2_out[1561] = 1'b0;
    assign layer2_out[1562] = ~layer1_out[76] | layer1_out[77];
    assign layer2_out[1563] = ~(layer1_out[7168] | layer1_out[7169]);
    assign layer2_out[1564] = layer1_out[7061] ^ layer1_out[7062];
    assign layer2_out[1565] = layer1_out[7949];
    assign layer2_out[1566] = layer1_out[4394] ^ layer1_out[4395];
    assign layer2_out[1567] = layer1_out[3099] | layer1_out[3100];
    assign layer2_out[1568] = layer1_out[5594] & layer1_out[5595];
    assign layer2_out[1569] = ~layer1_out[4542];
    assign layer2_out[1570] = ~(layer1_out[2102] | layer1_out[2103]);
    assign layer2_out[1571] = ~(layer1_out[4128] | layer1_out[4129]);
    assign layer2_out[1572] = layer1_out[1987] & ~layer1_out[1988];
    assign layer2_out[1573] = 1'b1;
    assign layer2_out[1574] = layer1_out[2186];
    assign layer2_out[1575] = ~layer1_out[7205];
    assign layer2_out[1576] = ~(layer1_out[4257] | layer1_out[4258]);
    assign layer2_out[1577] = layer1_out[7093] & ~layer1_out[7094];
    assign layer2_out[1578] = 1'b0;
    assign layer2_out[1579] = layer1_out[5992] ^ layer1_out[5993];
    assign layer2_out[1580] = ~(layer1_out[3651] | layer1_out[3652]);
    assign layer2_out[1581] = ~layer1_out[7310] | layer1_out[7311];
    assign layer2_out[1582] = layer1_out[567] | layer1_out[568];
    assign layer2_out[1583] = 1'b0;
    assign layer2_out[1584] = ~layer1_out[1692] | layer1_out[1691];
    assign layer2_out[1585] = layer1_out[3409];
    assign layer2_out[1586] = layer1_out[641] | layer1_out[642];
    assign layer2_out[1587] = layer1_out[2773];
    assign layer2_out[1588] = 1'b0;
    assign layer2_out[1589] = layer1_out[660] & ~layer1_out[661];
    assign layer2_out[1590] = ~layer1_out[6181] | layer1_out[6182];
    assign layer2_out[1591] = ~layer1_out[3708];
    assign layer2_out[1592] = ~layer1_out[7718];
    assign layer2_out[1593] = layer1_out[1997];
    assign layer2_out[1594] = layer1_out[6353] & layer1_out[6354];
    assign layer2_out[1595] = ~(layer1_out[859] & layer1_out[860]);
    assign layer2_out[1596] = layer1_out[3570] | layer1_out[3571];
    assign layer2_out[1597] = ~layer1_out[5400];
    assign layer2_out[1598] = 1'b1;
    assign layer2_out[1599] = ~layer1_out[3930];
    assign layer2_out[1600] = ~(layer1_out[4194] | layer1_out[4195]);
    assign layer2_out[1601] = ~(layer1_out[5012] & layer1_out[5013]);
    assign layer2_out[1602] = ~layer1_out[6336] | layer1_out[6337];
    assign layer2_out[1603] = layer1_out[881] & ~layer1_out[880];
    assign layer2_out[1604] = ~layer1_out[6762];
    assign layer2_out[1605] = layer1_out[5684] ^ layer1_out[5685];
    assign layer2_out[1606] = ~layer1_out[3245] | layer1_out[3246];
    assign layer2_out[1607] = layer1_out[6301] & ~layer1_out[6302];
    assign layer2_out[1608] = ~layer1_out[5522];
    assign layer2_out[1609] = layer1_out[2928];
    assign layer2_out[1610] = layer1_out[3721];
    assign layer2_out[1611] = ~(layer1_out[1887] | layer1_out[1888]);
    assign layer2_out[1612] = layer1_out[2695] & ~layer1_out[2694];
    assign layer2_out[1613] = layer1_out[2266] | layer1_out[2267];
    assign layer2_out[1614] = layer1_out[1934] & ~layer1_out[1935];
    assign layer2_out[1615] = layer1_out[3765] & layer1_out[3766];
    assign layer2_out[1616] = layer1_out[1240] | layer1_out[1241];
    assign layer2_out[1617] = layer1_out[1611] & ~layer1_out[1610];
    assign layer2_out[1618] = layer1_out[3045] & ~layer1_out[3044];
    assign layer2_out[1619] = layer1_out[3993] & ~layer1_out[3994];
    assign layer2_out[1620] = layer1_out[4169];
    assign layer2_out[1621] = ~(layer1_out[7840] & layer1_out[7841]);
    assign layer2_out[1622] = layer1_out[7701];
    assign layer2_out[1623] = ~layer1_out[6339];
    assign layer2_out[1624] = ~layer1_out[3627];
    assign layer2_out[1625] = layer1_out[1973] | layer1_out[1974];
    assign layer2_out[1626] = layer1_out[4142];
    assign layer2_out[1627] = layer1_out[7429] & ~layer1_out[7428];
    assign layer2_out[1628] = ~layer1_out[0];
    assign layer2_out[1629] = layer1_out[4186] & ~layer1_out[4187];
    assign layer2_out[1630] = layer1_out[1896] & layer1_out[1897];
    assign layer2_out[1631] = layer1_out[6226];
    assign layer2_out[1632] = ~layer1_out[3174];
    assign layer2_out[1633] = layer1_out[4094] & ~layer1_out[4093];
    assign layer2_out[1634] = ~layer1_out[211] | layer1_out[212];
    assign layer2_out[1635] = ~(layer1_out[3242] & layer1_out[3243]);
    assign layer2_out[1636] = layer1_out[1645] & ~layer1_out[1646];
    assign layer2_out[1637] = layer1_out[5840];
    assign layer2_out[1638] = layer1_out[7105] & ~layer1_out[7106];
    assign layer2_out[1639] = ~layer1_out[7052];
    assign layer2_out[1640] = ~(layer1_out[5897] ^ layer1_out[5898]);
    assign layer2_out[1641] = layer1_out[5510] & ~layer1_out[5511];
    assign layer2_out[1642] = ~layer1_out[2917];
    assign layer2_out[1643] = layer1_out[4303] & layer1_out[4304];
    assign layer2_out[1644] = layer1_out[1195];
    assign layer2_out[1645] = layer1_out[404] ^ layer1_out[405];
    assign layer2_out[1646] = ~layer1_out[3844];
    assign layer2_out[1647] = ~layer1_out[2007];
    assign layer2_out[1648] = ~layer1_out[993] | layer1_out[994];
    assign layer2_out[1649] = ~(layer1_out[3248] | layer1_out[3249]);
    assign layer2_out[1650] = layer1_out[3474];
    assign layer2_out[1651] = layer1_out[6568];
    assign layer2_out[1652] = ~layer1_out[5456];
    assign layer2_out[1653] = 1'b1;
    assign layer2_out[1654] = layer1_out[6189];
    assign layer2_out[1655] = layer1_out[2286];
    assign layer2_out[1656] = ~layer1_out[1300];
    assign layer2_out[1657] = ~(layer1_out[5600] ^ layer1_out[5601]);
    assign layer2_out[1658] = ~layer1_out[7120];
    assign layer2_out[1659] = layer1_out[5247] & ~layer1_out[5246];
    assign layer2_out[1660] = layer1_out[169] | layer1_out[170];
    assign layer2_out[1661] = ~layer1_out[7671] | layer1_out[7672];
    assign layer2_out[1662] = layer1_out[5913] ^ layer1_out[5914];
    assign layer2_out[1663] = layer1_out[484] ^ layer1_out[485];
    assign layer2_out[1664] = layer1_out[7654];
    assign layer2_out[1665] = layer1_out[7110] & layer1_out[7111];
    assign layer2_out[1666] = ~layer1_out[6964];
    assign layer2_out[1667] = 1'b1;
    assign layer2_out[1668] = ~layer1_out[6047] | layer1_out[6048];
    assign layer2_out[1669] = layer1_out[6254];
    assign layer2_out[1670] = ~(layer1_out[5937] ^ layer1_out[5938]);
    assign layer2_out[1671] = layer1_out[6856];
    assign layer2_out[1672] = layer1_out[6445] | layer1_out[6446];
    assign layer2_out[1673] = layer1_out[1938] & layer1_out[1939];
    assign layer2_out[1674] = layer1_out[4604] & layer1_out[4605];
    assign layer2_out[1675] = ~layer1_out[2878];
    assign layer2_out[1676] = layer1_out[3924];
    assign layer2_out[1677] = layer1_out[7722] & ~layer1_out[7723];
    assign layer2_out[1678] = ~layer1_out[15] | layer1_out[16];
    assign layer2_out[1679] = layer1_out[332];
    assign layer2_out[1680] = layer1_out[982] | layer1_out[983];
    assign layer2_out[1681] = 1'b0;
    assign layer2_out[1682] = layer1_out[1336];
    assign layer2_out[1683] = ~layer1_out[1708] | layer1_out[1707];
    assign layer2_out[1684] = ~layer1_out[7920];
    assign layer2_out[1685] = 1'b1;
    assign layer2_out[1686] = ~layer1_out[415];
    assign layer2_out[1687] = layer1_out[763] & ~layer1_out[764];
    assign layer2_out[1688] = layer1_out[5460];
    assign layer2_out[1689] = ~(layer1_out[5490] & layer1_out[5491]);
    assign layer2_out[1690] = layer1_out[3638];
    assign layer2_out[1691] = layer1_out[1329] & layer1_out[1330];
    assign layer2_out[1692] = ~layer1_out[6777] | layer1_out[6776];
    assign layer2_out[1693] = ~layer1_out[5124] | layer1_out[5125];
    assign layer2_out[1694] = layer1_out[133];
    assign layer2_out[1695] = layer1_out[6662];
    assign layer2_out[1696] = layer1_out[3778] & ~layer1_out[3777];
    assign layer2_out[1697] = layer1_out[5530];
    assign layer2_out[1698] = 1'b0;
    assign layer2_out[1699] = layer1_out[5789];
    assign layer2_out[1700] = layer1_out[2454];
    assign layer2_out[1701] = ~layer1_out[3015];
    assign layer2_out[1702] = layer1_out[598] ^ layer1_out[599];
    assign layer2_out[1703] = ~layer1_out[4595];
    assign layer2_out[1704] = layer1_out[2206] & ~layer1_out[2207];
    assign layer2_out[1705] = ~layer1_out[1732] | layer1_out[1733];
    assign layer2_out[1706] = layer1_out[7506];
    assign layer2_out[1707] = ~layer1_out[7227];
    assign layer2_out[1708] = ~layer1_out[4525] | layer1_out[4524];
    assign layer2_out[1709] = ~layer1_out[2486];
    assign layer2_out[1710] = layer1_out[934] & ~layer1_out[933];
    assign layer2_out[1711] = layer1_out[3184];
    assign layer2_out[1712] = layer1_out[3154] | layer1_out[3155];
    assign layer2_out[1713] = ~layer1_out[5878];
    assign layer2_out[1714] = 1'b0;
    assign layer2_out[1715] = 1'b0;
    assign layer2_out[1716] = layer1_out[6772] ^ layer1_out[6773];
    assign layer2_out[1717] = layer1_out[7541];
    assign layer2_out[1718] = ~layer1_out[6270];
    assign layer2_out[1719] = ~(layer1_out[4043] ^ layer1_out[4044]);
    assign layer2_out[1720] = layer1_out[6715];
    assign layer2_out[1721] = layer1_out[2719] & layer1_out[2720];
    assign layer2_out[1722] = layer1_out[816];
    assign layer2_out[1723] = ~(layer1_out[2173] | layer1_out[2174]);
    assign layer2_out[1724] = layer1_out[7478] & layer1_out[7479];
    assign layer2_out[1725] = layer1_out[3831] & ~layer1_out[3832];
    assign layer2_out[1726] = ~layer1_out[7815];
    assign layer2_out[1727] = layer1_out[4320];
    assign layer2_out[1728] = layer1_out[4324] ^ layer1_out[4325];
    assign layer2_out[1729] = layer1_out[3143] & ~layer1_out[3144];
    assign layer2_out[1730] = 1'b1;
    assign layer2_out[1731] = ~(layer1_out[6705] & layer1_out[6706]);
    assign layer2_out[1732] = ~(layer1_out[1393] | layer1_out[1394]);
    assign layer2_out[1733] = ~layer1_out[1609] | layer1_out[1608];
    assign layer2_out[1734] = layer1_out[4220];
    assign layer2_out[1735] = layer1_out[528] | layer1_out[529];
    assign layer2_out[1736] = layer1_out[1432] & layer1_out[1433];
    assign layer2_out[1737] = layer1_out[1811] & ~layer1_out[1812];
    assign layer2_out[1738] = ~(layer1_out[5043] & layer1_out[5044]);
    assign layer2_out[1739] = ~layer1_out[7272] | layer1_out[7273];
    assign layer2_out[1740] = layer1_out[4159] & ~layer1_out[4158];
    assign layer2_out[1741] = ~layer1_out[4181];
    assign layer2_out[1742] = ~(layer1_out[7003] | layer1_out[7004]);
    assign layer2_out[1743] = layer1_out[7546] ^ layer1_out[7547];
    assign layer2_out[1744] = ~(layer1_out[2746] | layer1_out[2747]);
    assign layer2_out[1745] = ~layer1_out[3092] | layer1_out[3093];
    assign layer2_out[1746] = ~layer1_out[7508];
    assign layer2_out[1747] = layer1_out[3980] | layer1_out[3981];
    assign layer2_out[1748] = ~(layer1_out[2791] ^ layer1_out[2792]);
    assign layer2_out[1749] = layer1_out[3543];
    assign layer2_out[1750] = ~(layer1_out[7720] | layer1_out[7721]);
    assign layer2_out[1751] = layer1_out[5117];
    assign layer2_out[1752] = layer1_out[6220] & ~layer1_out[6219];
    assign layer2_out[1753] = ~(layer1_out[403] & layer1_out[404]);
    assign layer2_out[1754] = layer1_out[137];
    assign layer2_out[1755] = layer1_out[2136];
    assign layer2_out[1756] = layer1_out[5965] & ~layer1_out[5964];
    assign layer2_out[1757] = layer1_out[6577] & ~layer1_out[6576];
    assign layer2_out[1758] = ~(layer1_out[68] & layer1_out[69]);
    assign layer2_out[1759] = ~layer1_out[3077] | layer1_out[3076];
    assign layer2_out[1760] = ~(layer1_out[2967] & layer1_out[2968]);
    assign layer2_out[1761] = layer1_out[1058] & ~layer1_out[1057];
    assign layer2_out[1762] = ~(layer1_out[2623] & layer1_out[2624]);
    assign layer2_out[1763] = layer1_out[944] & ~layer1_out[943];
    assign layer2_out[1764] = ~layer1_out[1394];
    assign layer2_out[1765] = ~(layer1_out[2284] & layer1_out[2285]);
    assign layer2_out[1766] = ~layer1_out[331] | layer1_out[330];
    assign layer2_out[1767] = ~(layer1_out[36] ^ layer1_out[37]);
    assign layer2_out[1768] = layer1_out[4471] ^ layer1_out[4472];
    assign layer2_out[1769] = layer1_out[6457] & ~layer1_out[6456];
    assign layer2_out[1770] = layer1_out[6092];
    assign layer2_out[1771] = layer1_out[5533];
    assign layer2_out[1772] = layer1_out[5063] ^ layer1_out[5064];
    assign layer2_out[1773] = layer1_out[368] & ~layer1_out[367];
    assign layer2_out[1774] = layer1_out[844];
    assign layer2_out[1775] = ~(layer1_out[53] | layer1_out[54]);
    assign layer2_out[1776] = layer1_out[6906];
    assign layer2_out[1777] = layer1_out[3960] & ~layer1_out[3961];
    assign layer2_out[1778] = layer1_out[5389] | layer1_out[5390];
    assign layer2_out[1779] = layer1_out[3824] & ~layer1_out[3823];
    assign layer2_out[1780] = ~layer1_out[6786] | layer1_out[6785];
    assign layer2_out[1781] = layer1_out[4751] & layer1_out[4752];
    assign layer2_out[1782] = layer1_out[3420] & ~layer1_out[3419];
    assign layer2_out[1783] = 1'b0;
    assign layer2_out[1784] = layer1_out[5884] & ~layer1_out[5883];
    assign layer2_out[1785] = ~layer1_out[4768] | layer1_out[4769];
    assign layer2_out[1786] = 1'b1;
    assign layer2_out[1787] = layer1_out[3228] ^ layer1_out[3229];
    assign layer2_out[1788] = ~layer1_out[7149];
    assign layer2_out[1789] = ~layer1_out[2074];
    assign layer2_out[1790] = layer1_out[6368];
    assign layer2_out[1791] = layer1_out[7653] & ~layer1_out[7652];
    assign layer2_out[1792] = layer1_out[4622] & ~layer1_out[4621];
    assign layer2_out[1793] = layer1_out[4867] & layer1_out[4868];
    assign layer2_out[1794] = ~layer1_out[4234] | layer1_out[4233];
    assign layer2_out[1795] = ~layer1_out[1373] | layer1_out[1374];
    assign layer2_out[1796] = ~(layer1_out[981] ^ layer1_out[982]);
    assign layer2_out[1797] = layer1_out[3019] & ~layer1_out[3018];
    assign layer2_out[1798] = layer1_out[7122] & layer1_out[7123];
    assign layer2_out[1799] = layer1_out[7976] & ~layer1_out[7977];
    assign layer2_out[1800] = ~(layer1_out[5450] & layer1_out[5451]);
    assign layer2_out[1801] = ~(layer1_out[5130] | layer1_out[5131]);
    assign layer2_out[1802] = ~layer1_out[5713] | layer1_out[5712];
    assign layer2_out[1803] = ~layer1_out[4711] | layer1_out[4712];
    assign layer2_out[1804] = layer1_out[5868] | layer1_out[5869];
    assign layer2_out[1805] = ~layer1_out[505] | layer1_out[506];
    assign layer2_out[1806] = layer1_out[6746] ^ layer1_out[6747];
    assign layer2_out[1807] = ~(layer1_out[4889] | layer1_out[4890]);
    assign layer2_out[1808] = ~layer1_out[3786];
    assign layer2_out[1809] = ~layer1_out[7451] | layer1_out[7450];
    assign layer2_out[1810] = ~layer1_out[1651] | layer1_out[1650];
    assign layer2_out[1811] = layer1_out[449] ^ layer1_out[450];
    assign layer2_out[1812] = layer1_out[7913] & ~layer1_out[7912];
    assign layer2_out[1813] = ~layer1_out[7682] | layer1_out[7681];
    assign layer2_out[1814] = ~layer1_out[4894] | layer1_out[4895];
    assign layer2_out[1815] = ~layer1_out[1924];
    assign layer2_out[1816] = ~layer1_out[1935];
    assign layer2_out[1817] = layer1_out[7280];
    assign layer2_out[1818] = layer1_out[7221] & ~layer1_out[7222];
    assign layer2_out[1819] = ~(layer1_out[760] ^ layer1_out[761]);
    assign layer2_out[1820] = layer1_out[2202] | layer1_out[2203];
    assign layer2_out[1821] = ~(layer1_out[2937] & layer1_out[2938]);
    assign layer2_out[1822] = layer1_out[4338] & ~layer1_out[4339];
    assign layer2_out[1823] = layer1_out[1283] & layer1_out[1284];
    assign layer2_out[1824] = layer1_out[3349] & layer1_out[3350];
    assign layer2_out[1825] = layer1_out[2804];
    assign layer2_out[1826] = layer1_out[2789] | layer1_out[2790];
    assign layer2_out[1827] = ~layer1_out[2175];
    assign layer2_out[1828] = layer1_out[3804] & ~layer1_out[3805];
    assign layer2_out[1829] = 1'b1;
    assign layer2_out[1830] = layer1_out[78] & ~layer1_out[77];
    assign layer2_out[1831] = ~layer1_out[5743];
    assign layer2_out[1832] = layer1_out[3288];
    assign layer2_out[1833] = layer1_out[6068];
    assign layer2_out[1834] = ~layer1_out[997];
    assign layer2_out[1835] = layer1_out[5070] & layer1_out[5071];
    assign layer2_out[1836] = layer1_out[355] | layer1_out[356];
    assign layer2_out[1837] = layer1_out[7406] ^ layer1_out[7407];
    assign layer2_out[1838] = layer1_out[7888];
    assign layer2_out[1839] = ~layer1_out[5240];
    assign layer2_out[1840] = layer1_out[3021] & ~layer1_out[3020];
    assign layer2_out[1841] = layer1_out[4391] | layer1_out[4392];
    assign layer2_out[1842] = layer1_out[4964];
    assign layer2_out[1843] = layer1_out[755];
    assign layer2_out[1844] = ~layer1_out[1525];
    assign layer2_out[1845] = ~layer1_out[5656];
    assign layer2_out[1846] = ~(layer1_out[4482] & layer1_out[4483]);
    assign layer2_out[1847] = ~layer1_out[3247];
    assign layer2_out[1848] = ~(layer1_out[7229] & layer1_out[7230]);
    assign layer2_out[1849] = ~layer1_out[2040] | layer1_out[2039];
    assign layer2_out[1850] = layer1_out[5724];
    assign layer2_out[1851] = ~layer1_out[3548];
    assign layer2_out[1852] = layer1_out[184];
    assign layer2_out[1853] = layer1_out[5564] & ~layer1_out[5563];
    assign layer2_out[1854] = layer1_out[4227] | layer1_out[4228];
    assign layer2_out[1855] = layer1_out[7366] & ~layer1_out[7365];
    assign layer2_out[1856] = ~(layer1_out[2412] | layer1_out[2413]);
    assign layer2_out[1857] = layer1_out[262];
    assign layer2_out[1858] = ~layer1_out[4075];
    assign layer2_out[1859] = layer1_out[3873] & ~layer1_out[3872];
    assign layer2_out[1860] = layer1_out[2028];
    assign layer2_out[1861] = layer1_out[4385];
    assign layer2_out[1862] = ~(layer1_out[3021] ^ layer1_out[3022]);
    assign layer2_out[1863] = layer1_out[475] | layer1_out[476];
    assign layer2_out[1864] = layer1_out[5018] & ~layer1_out[5019];
    assign layer2_out[1865] = 1'b1;
    assign layer2_out[1866] = ~(layer1_out[6135] | layer1_out[6136]);
    assign layer2_out[1867] = ~(layer1_out[853] ^ layer1_out[854]);
    assign layer2_out[1868] = ~layer1_out[7295] | layer1_out[7294];
    assign layer2_out[1869] = ~layer1_out[1867] | layer1_out[1866];
    assign layer2_out[1870] = layer1_out[7042] & layer1_out[7043];
    assign layer2_out[1871] = layer1_out[4694];
    assign layer2_out[1872] = layer1_out[774];
    assign layer2_out[1873] = 1'b0;
    assign layer2_out[1874] = 1'b1;
    assign layer2_out[1875] = ~layer1_out[4987];
    assign layer2_out[1876] = ~(layer1_out[5242] & layer1_out[5243]);
    assign layer2_out[1877] = layer1_out[6820] & layer1_out[6821];
    assign layer2_out[1878] = ~layer1_out[2851];
    assign layer2_out[1879] = ~layer1_out[3282];
    assign layer2_out[1880] = layer1_out[6969];
    assign layer2_out[1881] = ~layer1_out[6655] | layer1_out[6654];
    assign layer2_out[1882] = layer1_out[5225] & ~layer1_out[5224];
    assign layer2_out[1883] = ~layer1_out[1957] | layer1_out[1956];
    assign layer2_out[1884] = ~(layer1_out[6158] & layer1_out[6159]);
    assign layer2_out[1885] = layer1_out[1414];
    assign layer2_out[1886] = ~(layer1_out[6334] & layer1_out[6335]);
    assign layer2_out[1887] = layer1_out[3682];
    assign layer2_out[1888] = layer1_out[680] | layer1_out[681];
    assign layer2_out[1889] = layer1_out[2388] & ~layer1_out[2389];
    assign layer2_out[1890] = layer1_out[2599] & layer1_out[2600];
    assign layer2_out[1891] = ~(layer1_out[5079] & layer1_out[5080]);
    assign layer2_out[1892] = ~layer1_out[1702];
    assign layer2_out[1893] = layer1_out[2492];
    assign layer2_out[1894] = ~layer1_out[4151] | layer1_out[4152];
    assign layer2_out[1895] = layer1_out[2324] & ~layer1_out[2323];
    assign layer2_out[1896] = 1'b1;
    assign layer2_out[1897] = ~layer1_out[7202] | layer1_out[7201];
    assign layer2_out[1898] = layer1_out[222];
    assign layer2_out[1899] = layer1_out[4509];
    assign layer2_out[1900] = layer1_out[3256] & layer1_out[3257];
    assign layer2_out[1901] = layer1_out[6379];
    assign layer2_out[1902] = layer1_out[6970] & ~layer1_out[6971];
    assign layer2_out[1903] = ~(layer1_out[2345] & layer1_out[2346]);
    assign layer2_out[1904] = ~layer1_out[1244] | layer1_out[1243];
    assign layer2_out[1905] = layer1_out[363] & ~layer1_out[362];
    assign layer2_out[1906] = ~(layer1_out[5520] | layer1_out[5521]);
    assign layer2_out[1907] = ~(layer1_out[6275] ^ layer1_out[6276]);
    assign layer2_out[1908] = 1'b0;
    assign layer2_out[1909] = ~layer1_out[908] | layer1_out[909];
    assign layer2_out[1910] = ~(layer1_out[5235] & layer1_out[5236]);
    assign layer2_out[1911] = layer1_out[6610] ^ layer1_out[6611];
    assign layer2_out[1912] = ~layer1_out[4328];
    assign layer2_out[1913] = ~(layer1_out[2751] | layer1_out[2752]);
    assign layer2_out[1914] = ~layer1_out[3430];
    assign layer2_out[1915] = layer1_out[3589];
    assign layer2_out[1916] = ~(layer1_out[7691] ^ layer1_out[7692]);
    assign layer2_out[1917] = ~layer1_out[3036];
    assign layer2_out[1918] = ~(layer1_out[3402] & layer1_out[3403]);
    assign layer2_out[1919] = layer1_out[5286] & ~layer1_out[5287];
    assign layer2_out[1920] = layer1_out[5163];
    assign layer2_out[1921] = ~layer1_out[5297];
    assign layer2_out[1922] = ~layer1_out[6050] | layer1_out[6049];
    assign layer2_out[1923] = ~layer1_out[7052];
    assign layer2_out[1924] = layer1_out[2727] & ~layer1_out[2728];
    assign layer2_out[1925] = layer1_out[6634] & layer1_out[6635];
    assign layer2_out[1926] = layer1_out[3238];
    assign layer2_out[1927] = ~layer1_out[3508];
    assign layer2_out[1928] = 1'b0;
    assign layer2_out[1929] = ~(layer1_out[1154] | layer1_out[1155]);
    assign layer2_out[1930] = ~layer1_out[3953];
    assign layer2_out[1931] = ~(layer1_out[698] ^ layer1_out[699]);
    assign layer2_out[1932] = layer1_out[6097] ^ layer1_out[6098];
    assign layer2_out[1933] = ~layer1_out[5057] | layer1_out[5058];
    assign layer2_out[1934] = layer1_out[7528];
    assign layer2_out[1935] = layer1_out[1910] | layer1_out[1911];
    assign layer2_out[1936] = 1'b1;
    assign layer2_out[1937] = layer1_out[3085];
    assign layer2_out[1938] = ~(layer1_out[5932] & layer1_out[5933]);
    assign layer2_out[1939] = ~layer1_out[3652] | layer1_out[3653];
    assign layer2_out[1940] = layer1_out[3514];
    assign layer2_out[1941] = ~layer1_out[5565];
    assign layer2_out[1942] = ~(layer1_out[7656] | layer1_out[7657]);
    assign layer2_out[1943] = layer1_out[5960];
    assign layer2_out[1944] = layer1_out[186] | layer1_out[187];
    assign layer2_out[1945] = ~(layer1_out[1102] ^ layer1_out[1103]);
    assign layer2_out[1946] = layer1_out[5933] & ~layer1_out[5934];
    assign layer2_out[1947] = layer1_out[5459] & layer1_out[5460];
    assign layer2_out[1948] = layer1_out[6426];
    assign layer2_out[1949] = ~layer1_out[5621] | layer1_out[5620];
    assign layer2_out[1950] = layer1_out[2198];
    assign layer2_out[1951] = layer1_out[1844];
    assign layer2_out[1952] = ~layer1_out[6060];
    assign layer2_out[1953] = ~layer1_out[863];
    assign layer2_out[1954] = layer1_out[5367] & layer1_out[5368];
    assign layer2_out[1955] = ~(layer1_out[6327] & layer1_out[6328]);
    assign layer2_out[1956] = layer1_out[410];
    assign layer2_out[1957] = layer1_out[7387] | layer1_out[7388];
    assign layer2_out[1958] = layer1_out[2477] & layer1_out[2478];
    assign layer2_out[1959] = 1'b1;
    assign layer2_out[1960] = ~(layer1_out[7464] | layer1_out[7465]);
    assign layer2_out[1961] = layer1_out[3530];
    assign layer2_out[1962] = layer1_out[3999];
    assign layer2_out[1963] = layer1_out[10];
    assign layer2_out[1964] = ~layer1_out[489];
    assign layer2_out[1965] = layer1_out[304] | layer1_out[305];
    assign layer2_out[1966] = layer1_out[3968];
    assign layer2_out[1967] = layer1_out[2765] & ~layer1_out[2764];
    assign layer2_out[1968] = ~layer1_out[7750];
    assign layer2_out[1969] = ~(layer1_out[7980] ^ layer1_out[7981]);
    assign layer2_out[1970] = layer1_out[3884] | layer1_out[3885];
    assign layer2_out[1971] = ~layer1_out[3091];
    assign layer2_out[1972] = layer1_out[4294] & ~layer1_out[4295];
    assign layer2_out[1973] = ~layer1_out[6892] | layer1_out[6891];
    assign layer2_out[1974] = layer1_out[6574];
    assign layer2_out[1975] = layer1_out[3428] & ~layer1_out[3427];
    assign layer2_out[1976] = ~(layer1_out[3945] & layer1_out[3946]);
    assign layer2_out[1977] = layer1_out[601] & ~layer1_out[602];
    assign layer2_out[1978] = layer1_out[1725] & ~layer1_out[1724];
    assign layer2_out[1979] = layer1_out[6260];
    assign layer2_out[1980] = layer1_out[7860];
    assign layer2_out[1981] = layer1_out[7577] & ~layer1_out[7578];
    assign layer2_out[1982] = layer1_out[2035] & layer1_out[2036];
    assign layer2_out[1983] = layer1_out[1714];
    assign layer2_out[1984] = layer1_out[7458] & ~layer1_out[7457];
    assign layer2_out[1985] = layer1_out[2490];
    assign layer2_out[1986] = ~(layer1_out[3441] & layer1_out[3442]);
    assign layer2_out[1987] = ~layer1_out[7411] | layer1_out[7412];
    assign layer2_out[1988] = layer1_out[7974];
    assign layer2_out[1989] = layer1_out[7292] & layer1_out[7293];
    assign layer2_out[1990] = layer1_out[3158];
    assign layer2_out[1991] = layer1_out[7993] ^ layer1_out[7994];
    assign layer2_out[1992] = layer1_out[3186] & layer1_out[3187];
    assign layer2_out[1993] = layer1_out[7593] | layer1_out[7594];
    assign layer2_out[1994] = 1'b1;
    assign layer2_out[1995] = 1'b1;
    assign layer2_out[1996] = layer1_out[2855];
    assign layer2_out[1997] = layer1_out[340];
    assign layer2_out[1998] = ~layer1_out[3171];
    assign layer2_out[1999] = ~layer1_out[3908];
    assign layer2_out[2000] = layer1_out[7282] | layer1_out[7283];
    assign layer2_out[2001] = layer1_out[4648];
    assign layer2_out[2002] = layer1_out[5504];
    assign layer2_out[2003] = ~layer1_out[7411] | layer1_out[7410];
    assign layer2_out[2004] = layer1_out[917] & ~layer1_out[916];
    assign layer2_out[2005] = 1'b0;
    assign layer2_out[2006] = layer1_out[4897] & ~layer1_out[4896];
    assign layer2_out[2007] = layer1_out[1285] & layer1_out[1286];
    assign layer2_out[2008] = ~layer1_out[2592];
    assign layer2_out[2009] = layer1_out[3604] & ~layer1_out[3605];
    assign layer2_out[2010] = layer1_out[5233] | layer1_out[5234];
    assign layer2_out[2011] = 1'b0;
    assign layer2_out[2012] = layer1_out[2677] & ~layer1_out[2676];
    assign layer2_out[2013] = ~layer1_out[4473] | layer1_out[4472];
    assign layer2_out[2014] = ~layer1_out[3678] | layer1_out[3679];
    assign layer2_out[2015] = layer1_out[4583] & ~layer1_out[4582];
    assign layer2_out[2016] = layer1_out[733] | layer1_out[734];
    assign layer2_out[2017] = ~layer1_out[2961];
    assign layer2_out[2018] = ~(layer1_out[7686] | layer1_out[7687]);
    assign layer2_out[2019] = ~layer1_out[6344] | layer1_out[6345];
    assign layer2_out[2020] = ~layer1_out[7234];
    assign layer2_out[2021] = layer1_out[5262] & ~layer1_out[5261];
    assign layer2_out[2022] = ~layer1_out[7397];
    assign layer2_out[2023] = layer1_out[4721];
    assign layer2_out[2024] = ~layer1_out[4238] | layer1_out[4239];
    assign layer2_out[2025] = ~(layer1_out[7055] | layer1_out[7056]);
    assign layer2_out[2026] = layer1_out[4439];
    assign layer2_out[2027] = layer1_out[1315];
    assign layer2_out[2028] = ~(layer1_out[695] ^ layer1_out[696]);
    assign layer2_out[2029] = layer1_out[3490] | layer1_out[3491];
    assign layer2_out[2030] = ~layer1_out[1918] | layer1_out[1917];
    assign layer2_out[2031] = ~layer1_out[2668];
    assign layer2_out[2032] = ~(layer1_out[4980] & layer1_out[4981]);
    assign layer2_out[2033] = ~(layer1_out[190] | layer1_out[191]);
    assign layer2_out[2034] = layer1_out[1449];
    assign layer2_out[2035] = ~(layer1_out[5905] ^ layer1_out[5906]);
    assign layer2_out[2036] = layer1_out[971] & ~layer1_out[972];
    assign layer2_out[2037] = 1'b0;
    assign layer2_out[2038] = layer1_out[714];
    assign layer2_out[2039] = layer1_out[7928];
    assign layer2_out[2040] = layer1_out[900];
    assign layer2_out[2041] = ~layer1_out[7674];
    assign layer2_out[2042] = layer1_out[919] & ~layer1_out[918];
    assign layer2_out[2043] = 1'b0;
    assign layer2_out[2044] = ~(layer1_out[3916] | layer1_out[3917]);
    assign layer2_out[2045] = ~layer1_out[3038];
    assign layer2_out[2046] = ~layer1_out[5177] | layer1_out[5178];
    assign layer2_out[2047] = layer1_out[4404] ^ layer1_out[4405];
    assign layer2_out[2048] = layer1_out[238] & ~layer1_out[239];
    assign layer2_out[2049] = ~(layer1_out[3367] & layer1_out[3368]);
    assign layer2_out[2050] = 1'b0;
    assign layer2_out[2051] = layer1_out[7494] ^ layer1_out[7495];
    assign layer2_out[2052] = layer1_out[2261] & ~layer1_out[2262];
    assign layer2_out[2053] = ~layer1_out[4489] | layer1_out[4488];
    assign layer2_out[2054] = layer1_out[5166];
    assign layer2_out[2055] = ~layer1_out[3526] | layer1_out[3525];
    assign layer2_out[2056] = ~layer1_out[838] | layer1_out[839];
    assign layer2_out[2057] = layer1_out[5612] | layer1_out[5613];
    assign layer2_out[2058] = ~layer1_out[2564] | layer1_out[2563];
    assign layer2_out[2059] = ~(layer1_out[3561] ^ layer1_out[3562]);
    assign layer2_out[2060] = layer1_out[5126] & layer1_out[5127];
    assign layer2_out[2061] = layer1_out[7552];
    assign layer2_out[2062] = layer1_out[5116];
    assign layer2_out[2063] = 1'b0;
    assign layer2_out[2064] = ~layer1_out[1950];
    assign layer2_out[2065] = ~layer1_out[1597];
    assign layer2_out[2066] = ~(layer1_out[5914] | layer1_out[5915]);
    assign layer2_out[2067] = ~(layer1_out[7075] & layer1_out[7076]);
    assign layer2_out[2068] = layer1_out[3744] | layer1_out[3745];
    assign layer2_out[2069] = layer1_out[1278] & layer1_out[1279];
    assign layer2_out[2070] = layer1_out[5151];
    assign layer2_out[2071] = layer1_out[6246] & ~layer1_out[6245];
    assign layer2_out[2072] = ~layer1_out[391];
    assign layer2_out[2073] = layer1_out[3278] & layer1_out[3279];
    assign layer2_out[2074] = layer1_out[5538] & ~layer1_out[5537];
    assign layer2_out[2075] = layer1_out[6595];
    assign layer2_out[2076] = layer1_out[1511] & layer1_out[1512];
    assign layer2_out[2077] = ~layer1_out[4722];
    assign layer2_out[2078] = layer1_out[3426] | layer1_out[3427];
    assign layer2_out[2079] = layer1_out[2833];
    assign layer2_out[2080] = ~layer1_out[2091];
    assign layer2_out[2081] = layer1_out[4228] & ~layer1_out[4229];
    assign layer2_out[2082] = ~layer1_out[6406] | layer1_out[6405];
    assign layer2_out[2083] = ~layer1_out[5192];
    assign layer2_out[2084] = 1'b1;
    assign layer2_out[2085] = layer1_out[4978];
    assign layer2_out[2086] = ~layer1_out[5107];
    assign layer2_out[2087] = layer1_out[4295] | layer1_out[4296];
    assign layer2_out[2088] = ~layer1_out[3053];
    assign layer2_out[2089] = ~layer1_out[2966] | layer1_out[2967];
    assign layer2_out[2090] = ~(layer1_out[6342] & layer1_out[6343]);
    assign layer2_out[2091] = layer1_out[481] | layer1_out[482];
    assign layer2_out[2092] = ~(layer1_out[3135] ^ layer1_out[3136]);
    assign layer2_out[2093] = layer1_out[5374];
    assign layer2_out[2094] = layer1_out[2953] & layer1_out[2954];
    assign layer2_out[2095] = layer1_out[4834] | layer1_out[4835];
    assign layer2_out[2096] = ~layer1_out[5353] | layer1_out[5352];
    assign layer2_out[2097] = layer1_out[3430];
    assign layer2_out[2098] = layer1_out[2745] & ~layer1_out[2744];
    assign layer2_out[2099] = ~layer1_out[5675];
    assign layer2_out[2100] = layer1_out[2373];
    assign layer2_out[2101] = ~(layer1_out[579] | layer1_out[580]);
    assign layer2_out[2102] = layer1_out[7180] ^ layer1_out[7181];
    assign layer2_out[2103] = layer1_out[5747] & ~layer1_out[5748];
    assign layer2_out[2104] = layer1_out[3167] & ~layer1_out[3166];
    assign layer2_out[2105] = ~(layer1_out[184] ^ layer1_out[185]);
    assign layer2_out[2106] = ~layer1_out[7566] | layer1_out[7567];
    assign layer2_out[2107] = ~layer1_out[6851] | layer1_out[6852];
    assign layer2_out[2108] = layer1_out[5837] & ~layer1_out[5838];
    assign layer2_out[2109] = layer1_out[4158] & ~layer1_out[4157];
    assign layer2_out[2110] = layer1_out[6516] & layer1_out[6517];
    assign layer2_out[2111] = layer1_out[1251] & ~layer1_out[1250];
    assign layer2_out[2112] = ~(layer1_out[3252] | layer1_out[3253]);
    assign layer2_out[2113] = layer1_out[668] ^ layer1_out[669];
    assign layer2_out[2114] = layer1_out[2305];
    assign layer2_out[2115] = ~(layer1_out[480] | layer1_out[481]);
    assign layer2_out[2116] = layer1_out[2544] | layer1_out[2545];
    assign layer2_out[2117] = layer1_out[3774] | layer1_out[3775];
    assign layer2_out[2118] = layer1_out[7672] | layer1_out[7673];
    assign layer2_out[2119] = layer1_out[5361] ^ layer1_out[5362];
    assign layer2_out[2120] = ~layer1_out[347] | layer1_out[346];
    assign layer2_out[2121] = layer1_out[7368] & ~layer1_out[7367];
    assign layer2_out[2122] = ~(layer1_out[7403] | layer1_out[7404]);
    assign layer2_out[2123] = layer1_out[998] | layer1_out[999];
    assign layer2_out[2124] = ~layer1_out[4373];
    assign layer2_out[2125] = layer1_out[651] & layer1_out[652];
    assign layer2_out[2126] = ~layer1_out[998] | layer1_out[997];
    assign layer2_out[2127] = layer1_out[5394] & ~layer1_out[5393];
    assign layer2_out[2128] = ~layer1_out[587] | layer1_out[588];
    assign layer2_out[2129] = layer1_out[4405] | layer1_out[4406];
    assign layer2_out[2130] = layer1_out[7367] & ~layer1_out[7366];
    assign layer2_out[2131] = layer1_out[1969] & ~layer1_out[1970];
    assign layer2_out[2132] = ~layer1_out[5601];
    assign layer2_out[2133] = 1'b1;
    assign layer2_out[2134] = ~layer1_out[2058];
    assign layer2_out[2135] = ~layer1_out[7055] | layer1_out[7054];
    assign layer2_out[2136] = ~layer1_out[3657] | layer1_out[3656];
    assign layer2_out[2137] = layer1_out[1289] & ~layer1_out[1288];
    assign layer2_out[2138] = ~layer1_out[2643] | layer1_out[2642];
    assign layer2_out[2139] = ~layer1_out[3497];
    assign layer2_out[2140] = layer1_out[3801];
    assign layer2_out[2141] = layer1_out[7134];
    assign layer2_out[2142] = ~layer1_out[1517];
    assign layer2_out[2143] = layer1_out[7271] & layer1_out[7272];
    assign layer2_out[2144] = layer1_out[6909];
    assign layer2_out[2145] = layer1_out[6514] & ~layer1_out[6513];
    assign layer2_out[2146] = layer1_out[1661] & ~layer1_out[1662];
    assign layer2_out[2147] = ~layer1_out[1601];
    assign layer2_out[2148] = ~layer1_out[7221];
    assign layer2_out[2149] = ~layer1_out[7281] | layer1_out[7282];
    assign layer2_out[2150] = ~layer1_out[4599];
    assign layer2_out[2151] = layer1_out[3343] & ~layer1_out[3344];
    assign layer2_out[2152] = ~layer1_out[591];
    assign layer2_out[2153] = ~(layer1_out[3529] ^ layer1_out[3530]);
    assign layer2_out[2154] = layer1_out[1299] & ~layer1_out[1298];
    assign layer2_out[2155] = layer1_out[1712] & ~layer1_out[1713];
    assign layer2_out[2156] = layer1_out[125];
    assign layer2_out[2157] = layer1_out[155] & ~layer1_out[156];
    assign layer2_out[2158] = ~(layer1_out[7370] | layer1_out[7371]);
    assign layer2_out[2159] = ~layer1_out[4153];
    assign layer2_out[2160] = ~layer1_out[3220];
    assign layer2_out[2161] = ~layer1_out[5470] | layer1_out[5471];
    assign layer2_out[2162] = 1'b1;
    assign layer2_out[2163] = ~layer1_out[1013];
    assign layer2_out[2164] = ~(layer1_out[6877] | layer1_out[6878]);
    assign layer2_out[2165] = ~layer1_out[4602] | layer1_out[4601];
    assign layer2_out[2166] = layer1_out[2795];
    assign layer2_out[2167] = layer1_out[4842] & ~layer1_out[4841];
    assign layer2_out[2168] = ~layer1_out[7320];
    assign layer2_out[2169] = layer1_out[7982];
    assign layer2_out[2170] = ~(layer1_out[6708] ^ layer1_out[6709]);
    assign layer2_out[2171] = ~layer1_out[4316] | layer1_out[4317];
    assign layer2_out[2172] = ~(layer1_out[312] | layer1_out[313]);
    assign layer2_out[2173] = layer1_out[406] | layer1_out[407];
    assign layer2_out[2174] = ~(layer1_out[7251] ^ layer1_out[7252]);
    assign layer2_out[2175] = layer1_out[1903] | layer1_out[1904];
    assign layer2_out[2176] = layer1_out[6098] & ~layer1_out[6099];
    assign layer2_out[2177] = ~(layer1_out[6663] & layer1_out[6664]);
    assign layer2_out[2178] = layer1_out[7238];
    assign layer2_out[2179] = ~layer1_out[6872] | layer1_out[6873];
    assign layer2_out[2180] = layer1_out[1905] & ~layer1_out[1906];
    assign layer2_out[2181] = ~layer1_out[4348];
    assign layer2_out[2182] = layer1_out[3074];
    assign layer2_out[2183] = ~layer1_out[6546];
    assign layer2_out[2184] = ~layer1_out[4679] | layer1_out[4678];
    assign layer2_out[2185] = ~layer1_out[5670] | layer1_out[5669];
    assign layer2_out[2186] = layer1_out[5360];
    assign layer2_out[2187] = ~layer1_out[7012];
    assign layer2_out[2188] = layer1_out[4971];
    assign layer2_out[2189] = layer1_out[5384] & layer1_out[5385];
    assign layer2_out[2190] = layer1_out[1944] & layer1_out[1945];
    assign layer2_out[2191] = 1'b0;
    assign layer2_out[2192] = ~layer1_out[1943];
    assign layer2_out[2193] = layer1_out[3400] & ~layer1_out[3399];
    assign layer2_out[2194] = ~layer1_out[5025];
    assign layer2_out[2195] = 1'b0;
    assign layer2_out[2196] = ~(layer1_out[3533] & layer1_out[3534]);
    assign layer2_out[2197] = layer1_out[6183] & ~layer1_out[6182];
    assign layer2_out[2198] = ~(layer1_out[3226] ^ layer1_out[3227]);
    assign layer2_out[2199] = layer1_out[2210] & ~layer1_out[2209];
    assign layer2_out[2200] = ~(layer1_out[2106] & layer1_out[2107]);
    assign layer2_out[2201] = layer1_out[4995] & layer1_out[4996];
    assign layer2_out[2202] = 1'b0;
    assign layer2_out[2203] = layer1_out[4225] ^ layer1_out[4226];
    assign layer2_out[2204] = layer1_out[6448] | layer1_out[6449];
    assign layer2_out[2205] = ~layer1_out[3965];
    assign layer2_out[2206] = ~layer1_out[6972];
    assign layer2_out[2207] = layer1_out[4761];
    assign layer2_out[2208] = layer1_out[1156];
    assign layer2_out[2209] = layer1_out[5525] & ~layer1_out[5524];
    assign layer2_out[2210] = layer1_out[6736] | layer1_out[6737];
    assign layer2_out[2211] = ~layer1_out[1569];
    assign layer2_out[2212] = ~(layer1_out[4262] & layer1_out[4263]);
    assign layer2_out[2213] = layer1_out[6680];
    assign layer2_out[2214] = layer1_out[4502] & ~layer1_out[4503];
    assign layer2_out[2215] = ~layer1_out[7300];
    assign layer2_out[2216] = layer1_out[4836] & ~layer1_out[4837];
    assign layer2_out[2217] = layer1_out[3169] & layer1_out[3170];
    assign layer2_out[2218] = layer1_out[1923];
    assign layer2_out[2219] = ~layer1_out[1450];
    assign layer2_out[2220] = ~layer1_out[3817] | layer1_out[3816];
    assign layer2_out[2221] = ~layer1_out[4219];
    assign layer2_out[2222] = ~(layer1_out[1069] & layer1_out[1070]);
    assign layer2_out[2223] = layer1_out[1694];
    assign layer2_out[2224] = layer1_out[6993] & ~layer1_out[6994];
    assign layer2_out[2225] = layer1_out[2059] | layer1_out[2060];
    assign layer2_out[2226] = ~layer1_out[644] | layer1_out[643];
    assign layer2_out[2227] = ~layer1_out[6662] | layer1_out[6663];
    assign layer2_out[2228] = layer1_out[1814];
    assign layer2_out[2229] = ~layer1_out[7807] | layer1_out[7808];
    assign layer2_out[2230] = layer1_out[6573] & ~layer1_out[6572];
    assign layer2_out[2231] = layer1_out[980] ^ layer1_out[981];
    assign layer2_out[2232] = layer1_out[2715] | layer1_out[2716];
    assign layer2_out[2233] = layer1_out[6913] & ~layer1_out[6912];
    assign layer2_out[2234] = ~layer1_out[7694] | layer1_out[7693];
    assign layer2_out[2235] = ~layer1_out[5343];
    assign layer2_out[2236] = ~layer1_out[5579];
    assign layer2_out[2237] = ~(layer1_out[2474] | layer1_out[2475]);
    assign layer2_out[2238] = layer1_out[4696] | layer1_out[4697];
    assign layer2_out[2239] = layer1_out[7799];
    assign layer2_out[2240] = layer1_out[866];
    assign layer2_out[2241] = layer1_out[3312];
    assign layer2_out[2242] = ~layer1_out[5973] | layer1_out[5972];
    assign layer2_out[2243] = ~layer1_out[2003] | layer1_out[2002];
    assign layer2_out[2244] = layer1_out[99];
    assign layer2_out[2245] = layer1_out[6000];
    assign layer2_out[2246] = layer1_out[7891] & ~layer1_out[7892];
    assign layer2_out[2247] = ~(layer1_out[2375] | layer1_out[2376]);
    assign layer2_out[2248] = ~layer1_out[2724] | layer1_out[2723];
    assign layer2_out[2249] = layer1_out[1594];
    assign layer2_out[2250] = layer1_out[4018] & ~layer1_out[4017];
    assign layer2_out[2251] = ~(layer1_out[7274] & layer1_out[7275]);
    assign layer2_out[2252] = ~(layer1_out[6168] & layer1_out[6169]);
    assign layer2_out[2253] = ~layer1_out[4448];
    assign layer2_out[2254] = ~layer1_out[280] | layer1_out[281];
    assign layer2_out[2255] = layer1_out[5218] & layer1_out[5219];
    assign layer2_out[2256] = layer1_out[5608] & ~layer1_out[5607];
    assign layer2_out[2257] = layer1_out[397];
    assign layer2_out[2258] = layer1_out[2737] | layer1_out[2738];
    assign layer2_out[2259] = layer1_out[1642] & ~layer1_out[1643];
    assign layer2_out[2260] = ~layer1_out[1116] | layer1_out[1115];
    assign layer2_out[2261] = layer1_out[1948] & layer1_out[1949];
    assign layer2_out[2262] = 1'b1;
    assign layer2_out[2263] = layer1_out[6363] & ~layer1_out[6364];
    assign layer2_out[2264] = ~(layer1_out[6721] ^ layer1_out[6722]);
    assign layer2_out[2265] = layer1_out[3871] & ~layer1_out[3872];
    assign layer2_out[2266] = ~layer1_out[6522];
    assign layer2_out[2267] = ~(layer1_out[1237] & layer1_out[1238]);
    assign layer2_out[2268] = ~(layer1_out[3963] ^ layer1_out[3964]);
    assign layer2_out[2269] = ~(layer1_out[4259] & layer1_out[4260]);
    assign layer2_out[2270] = ~(layer1_out[1251] & layer1_out[1252]);
    assign layer2_out[2271] = ~(layer1_out[5259] ^ layer1_out[5260]);
    assign layer2_out[2272] = ~(layer1_out[934] | layer1_out[935]);
    assign layer2_out[2273] = ~layer1_out[4409];
    assign layer2_out[2274] = layer1_out[7167];
    assign layer2_out[2275] = layer1_out[4101] & ~layer1_out[4100];
    assign layer2_out[2276] = layer1_out[1880] & ~layer1_out[1881];
    assign layer2_out[2277] = layer1_out[6848] & layer1_out[6849];
    assign layer2_out[2278] = ~(layer1_out[3001] | layer1_out[3002]);
    assign layer2_out[2279] = layer1_out[7380];
    assign layer2_out[2280] = ~layer1_out[2835];
    assign layer2_out[2281] = ~(layer1_out[932] | layer1_out[933]);
    assign layer2_out[2282] = ~(layer1_out[5487] ^ layer1_out[5488]);
    assign layer2_out[2283] = layer1_out[7749] & layer1_out[7750];
    assign layer2_out[2284] = layer1_out[952];
    assign layer2_out[2285] = layer1_out[5106] & ~layer1_out[5105];
    assign layer2_out[2286] = ~(layer1_out[1100] | layer1_out[1101]);
    assign layer2_out[2287] = layer1_out[1692] | layer1_out[1693];
    assign layer2_out[2288] = layer1_out[5658];
    assign layer2_out[2289] = ~layer1_out[7248];
    assign layer2_out[2290] = layer1_out[5289] & ~layer1_out[5290];
    assign layer2_out[2291] = layer1_out[2725];
    assign layer2_out[2292] = layer1_out[4149] & ~layer1_out[4150];
    assign layer2_out[2293] = layer1_out[2857] & ~layer1_out[2858];
    assign layer2_out[2294] = layer1_out[5725];
    assign layer2_out[2295] = ~layer1_out[5385];
    assign layer2_out[2296] = ~(layer1_out[6539] & layer1_out[6540]);
    assign layer2_out[2297] = ~layer1_out[1036];
    assign layer2_out[2298] = ~layer1_out[5764];
    assign layer2_out[2299] = 1'b0;
    assign layer2_out[2300] = layer1_out[5955] & layer1_out[5956];
    assign layer2_out[2301] = layer1_out[2264] & layer1_out[2265];
    assign layer2_out[2302] = ~layer1_out[4309];
    assign layer2_out[2303] = 1'b0;
    assign layer2_out[2304] = ~layer1_out[946] | layer1_out[947];
    assign layer2_out[2305] = ~layer1_out[7749] | layer1_out[7748];
    assign layer2_out[2306] = layer1_out[870] | layer1_out[871];
    assign layer2_out[2307] = ~(layer1_out[1076] | layer1_out[1077]);
    assign layer2_out[2308] = ~(layer1_out[4905] & layer1_out[4906]);
    assign layer2_out[2309] = layer1_out[6953] & ~layer1_out[6952];
    assign layer2_out[2310] = ~layer1_out[1183] | layer1_out[1182];
    assign layer2_out[2311] = layer1_out[3899] & ~layer1_out[3898];
    assign layer2_out[2312] = layer1_out[4649] | layer1_out[4650];
    assign layer2_out[2313] = ~(layer1_out[3126] | layer1_out[3127]);
    assign layer2_out[2314] = 1'b1;
    assign layer2_out[2315] = ~(layer1_out[1898] | layer1_out[1899]);
    assign layer2_out[2316] = layer1_out[2690];
    assign layer2_out[2317] = ~layer1_out[5665];
    assign layer2_out[2318] = layer1_out[1308];
    assign layer2_out[2319] = layer1_out[1289] & ~layer1_out[1290];
    assign layer2_out[2320] = layer1_out[6398];
    assign layer2_out[2321] = ~layer1_out[5644];
    assign layer2_out[2322] = ~layer1_out[3676];
    assign layer2_out[2323] = layer1_out[1807] & ~layer1_out[1808];
    assign layer2_out[2324] = ~layer1_out[5458];
    assign layer2_out[2325] = layer1_out[1950];
    assign layer2_out[2326] = layer1_out[5456] & ~layer1_out[5457];
    assign layer2_out[2327] = 1'b1;
    assign layer2_out[2328] = layer1_out[7818] | layer1_out[7819];
    assign layer2_out[2329] = ~(layer1_out[5653] ^ layer1_out[5654]);
    assign layer2_out[2330] = layer1_out[4906] ^ layer1_out[4907];
    assign layer2_out[2331] = ~layer1_out[6228];
    assign layer2_out[2332] = layer1_out[5512];
    assign layer2_out[2333] = ~layer1_out[5617];
    assign layer2_out[2334] = layer1_out[2978] & ~layer1_out[2979];
    assign layer2_out[2335] = ~layer1_out[7698];
    assign layer2_out[2336] = 1'b1;
    assign layer2_out[2337] = layer1_out[2446] | layer1_out[2447];
    assign layer2_out[2338] = layer1_out[1629];
    assign layer2_out[2339] = ~layer1_out[1690];
    assign layer2_out[2340] = ~layer1_out[1810];
    assign layer2_out[2341] = ~layer1_out[782] | layer1_out[781];
    assign layer2_out[2342] = ~layer1_out[5781] | layer1_out[5782];
    assign layer2_out[2343] = ~(layer1_out[405] | layer1_out[406]);
    assign layer2_out[2344] = layer1_out[6866] | layer1_out[6867];
    assign layer2_out[2345] = 1'b0;
    assign layer2_out[2346] = layer1_out[195] & ~layer1_out[194];
    assign layer2_out[2347] = layer1_out[4318] & layer1_out[4319];
    assign layer2_out[2348] = layer1_out[124] & ~layer1_out[123];
    assign layer2_out[2349] = ~layer1_out[7585];
    assign layer2_out[2350] = ~layer1_out[3729];
    assign layer2_out[2351] = ~layer1_out[2536] | layer1_out[2535];
    assign layer2_out[2352] = 1'b1;
    assign layer2_out[2353] = ~layer1_out[3757];
    assign layer2_out[2354] = layer1_out[7600] & ~layer1_out[7601];
    assign layer2_out[2355] = layer1_out[250] & layer1_out[251];
    assign layer2_out[2356] = layer1_out[4256] ^ layer1_out[4257];
    assign layer2_out[2357] = ~layer1_out[7725];
    assign layer2_out[2358] = ~layer1_out[3463];
    assign layer2_out[2359] = layer1_out[5320] | layer1_out[5321];
    assign layer2_out[2360] = ~layer1_out[1464];
    assign layer2_out[2361] = layer1_out[3936] & ~layer1_out[3937];
    assign layer2_out[2362] = layer1_out[1564] & layer1_out[1565];
    assign layer2_out[2363] = ~layer1_out[3832];
    assign layer2_out[2364] = ~layer1_out[2050];
    assign layer2_out[2365] = ~(layer1_out[402] & layer1_out[403]);
    assign layer2_out[2366] = 1'b1;
    assign layer2_out[2367] = layer1_out[1442] | layer1_out[1443];
    assign layer2_out[2368] = layer1_out[2762] | layer1_out[2763];
    assign layer2_out[2369] = ~layer1_out[6152];
    assign layer2_out[2370] = ~layer1_out[4288] | layer1_out[4289];
    assign layer2_out[2371] = ~(layer1_out[3285] ^ layer1_out[3286]);
    assign layer2_out[2372] = 1'b1;
    assign layer2_out[2373] = layer1_out[7770] & ~layer1_out[7769];
    assign layer2_out[2374] = layer1_out[4388];
    assign layer2_out[2375] = ~(layer1_out[7089] & layer1_out[7090]);
    assign layer2_out[2376] = layer1_out[2322] & layer1_out[2323];
    assign layer2_out[2377] = 1'b0;
    assign layer2_out[2378] = ~(layer1_out[3040] | layer1_out[3041]);
    assign layer2_out[2379] = ~(layer1_out[6022] | layer1_out[6023]);
    assign layer2_out[2380] = ~layer1_out[6955];
    assign layer2_out[2381] = ~layer1_out[4049] | layer1_out[4050];
    assign layer2_out[2382] = ~layer1_out[350] | layer1_out[351];
    assign layer2_out[2383] = layer1_out[1981] | layer1_out[1982];
    assign layer2_out[2384] = ~layer1_out[898] | layer1_out[899];
    assign layer2_out[2385] = ~layer1_out[6457] | layer1_out[6458];
    assign layer2_out[2386] = ~layer1_out[2513] | layer1_out[2514];
    assign layer2_out[2387] = layer1_out[871];
    assign layer2_out[2388] = layer1_out[3052] & ~layer1_out[3053];
    assign layer2_out[2389] = layer1_out[560];
    assign layer2_out[2390] = ~layer1_out[1625];
    assign layer2_out[2391] = ~layer1_out[319] | layer1_out[320];
    assign layer2_out[2392] = ~layer1_out[3086] | layer1_out[3085];
    assign layer2_out[2393] = ~layer1_out[3379];
    assign layer2_out[2394] = layer1_out[2869] ^ layer1_out[2870];
    assign layer2_out[2395] = layer1_out[584] ^ layer1_out[585];
    assign layer2_out[2396] = ~layer1_out[6179] | layer1_out[6178];
    assign layer2_out[2397] = layer1_out[958] & ~layer1_out[959];
    assign layer2_out[2398] = layer1_out[4244] | layer1_out[4245];
    assign layer2_out[2399] = layer1_out[2637];
    assign layer2_out[2400] = layer1_out[6667];
    assign layer2_out[2401] = layer1_out[3098] & ~layer1_out[3097];
    assign layer2_out[2402] = ~layer1_out[6749];
    assign layer2_out[2403] = 1'b0;
    assign layer2_out[2404] = layer1_out[5482] ^ layer1_out[5483];
    assign layer2_out[2405] = layer1_out[82] & layer1_out[83];
    assign layer2_out[2406] = ~(layer1_out[1946] | layer1_out[1947]);
    assign layer2_out[2407] = layer1_out[2778];
    assign layer2_out[2408] = layer1_out[4258] & layer1_out[4259];
    assign layer2_out[2409] = layer1_out[3881];
    assign layer2_out[2410] = layer1_out[377] & ~layer1_out[376];
    assign layer2_out[2411] = layer1_out[163];
    assign layer2_out[2412] = layer1_out[6652] & ~layer1_out[6651];
    assign layer2_out[2413] = ~layer1_out[7317] | layer1_out[7318];
    assign layer2_out[2414] = ~layer1_out[2274];
    assign layer2_out[2415] = layer1_out[3471] & ~layer1_out[3472];
    assign layer2_out[2416] = layer1_out[1808] ^ layer1_out[1809];
    assign layer2_out[2417] = ~(layer1_out[1549] | layer1_out[1550]);
    assign layer2_out[2418] = layer1_out[3470];
    assign layer2_out[2419] = layer1_out[3374] & ~layer1_out[3373];
    assign layer2_out[2420] = layer1_out[5526];
    assign layer2_out[2421] = layer1_out[2930] & ~layer1_out[2931];
    assign layer2_out[2422] = layer1_out[2209] & ~layer1_out[2208];
    assign layer2_out[2423] = layer1_out[6464] ^ layer1_out[6465];
    assign layer2_out[2424] = ~layer1_out[1698];
    assign layer2_out[2425] = layer1_out[4389];
    assign layer2_out[2426] = ~(layer1_out[157] | layer1_out[158]);
    assign layer2_out[2427] = ~layer1_out[4454] | layer1_out[4455];
    assign layer2_out[2428] = layer1_out[6246] & layer1_out[6247];
    assign layer2_out[2429] = ~layer1_out[2746] | layer1_out[2745];
    assign layer2_out[2430] = layer1_out[2703] & layer1_out[2704];
    assign layer2_out[2431] = layer1_out[6154];
    assign layer2_out[2432] = layer1_out[5855] | layer1_out[5856];
    assign layer2_out[2433] = layer1_out[51] & ~layer1_out[52];
    assign layer2_out[2434] = layer1_out[1459];
    assign layer2_out[2435] = ~layer1_out[850] | layer1_out[851];
    assign layer2_out[2436] = layer1_out[5591];
    assign layer2_out[2437] = ~layer1_out[313];
    assign layer2_out[2438] = ~layer1_out[4309] | layer1_out[4310];
    assign layer2_out[2439] = ~(layer1_out[2182] ^ layer1_out[2183]);
    assign layer2_out[2440] = layer1_out[2858] ^ layer1_out[2859];
    assign layer2_out[2441] = ~layer1_out[6574];
    assign layer2_out[2442] = layer1_out[2080] | layer1_out[2081];
    assign layer2_out[2443] = ~layer1_out[1700];
    assign layer2_out[2444] = layer1_out[6542] ^ layer1_out[6543];
    assign layer2_out[2445] = layer1_out[6536] & layer1_out[6537];
    assign layer2_out[2446] = layer1_out[6399] | layer1_out[6400];
    assign layer2_out[2447] = layer1_out[4099];
    assign layer2_out[2448] = layer1_out[133];
    assign layer2_out[2449] = layer1_out[1399];
    assign layer2_out[2450] = ~layer1_out[236] | layer1_out[237];
    assign layer2_out[2451] = ~layer1_out[5736];
    assign layer2_out[2452] = ~layer1_out[4045];
    assign layer2_out[2453] = layer1_out[4253] & layer1_out[4254];
    assign layer2_out[2454] = layer1_out[2949] | layer1_out[2950];
    assign layer2_out[2455] = layer1_out[5118] & ~layer1_out[5119];
    assign layer2_out[2456] = ~layer1_out[2437];
    assign layer2_out[2457] = layer1_out[68] & ~layer1_out[67];
    assign layer2_out[2458] = ~layer1_out[1585];
    assign layer2_out[2459] = ~layer1_out[1612];
    assign layer2_out[2460] = ~layer1_out[611];
    assign layer2_out[2461] = layer1_out[7999];
    assign layer2_out[2462] = layer1_out[1830];
    assign layer2_out[2463] = layer1_out[5599];
    assign layer2_out[2464] = ~layer1_out[6285];
    assign layer2_out[2465] = ~layer1_out[2989];
    assign layer2_out[2466] = layer1_out[5013];
    assign layer2_out[2467] = layer1_out[6904];
    assign layer2_out[2468] = layer1_out[3361] & ~layer1_out[3362];
    assign layer2_out[2469] = layer1_out[7648] & layer1_out[7649];
    assign layer2_out[2470] = ~(layer1_out[4826] | layer1_out[4827]);
    assign layer2_out[2471] = ~layer1_out[7139];
    assign layer2_out[2472] = ~layer1_out[5570] | layer1_out[5569];
    assign layer2_out[2473] = ~(layer1_out[989] | layer1_out[990]);
    assign layer2_out[2474] = ~layer1_out[5087];
    assign layer2_out[2475] = layer1_out[6830] & ~layer1_out[6831];
    assign layer2_out[2476] = ~(layer1_out[3221] ^ layer1_out[3222]);
    assign layer2_out[2477] = layer1_out[5760] & ~layer1_out[5759];
    assign layer2_out[2478] = ~(layer1_out[6618] & layer1_out[6619]);
    assign layer2_out[2479] = layer1_out[7678] & ~layer1_out[7679];
    assign layer2_out[2480] = layer1_out[7036] ^ layer1_out[7037];
    assign layer2_out[2481] = layer1_out[7931] & ~layer1_out[7930];
    assign layer2_out[2482] = layer1_out[5785] & layer1_out[5786];
    assign layer2_out[2483] = ~layer1_out[4941];
    assign layer2_out[2484] = layer1_out[740] | layer1_out[741];
    assign layer2_out[2485] = ~layer1_out[4513];
    assign layer2_out[2486] = ~layer1_out[3645] | layer1_out[3646];
    assign layer2_out[2487] = layer1_out[4739] & ~layer1_out[4738];
    assign layer2_out[2488] = layer1_out[6231] ^ layer1_out[6232];
    assign layer2_out[2489] = ~(layer1_out[5948] | layer1_out[5949]);
    assign layer2_out[2490] = layer1_out[1238] & layer1_out[1239];
    assign layer2_out[2491] = ~layer1_out[6599];
    assign layer2_out[2492] = layer1_out[6270] & ~layer1_out[6269];
    assign layer2_out[2493] = ~(layer1_out[4107] ^ layer1_out[4108]);
    assign layer2_out[2494] = ~layer1_out[3181];
    assign layer2_out[2495] = ~layer1_out[6264];
    assign layer2_out[2496] = ~layer1_out[3571] | layer1_out[3572];
    assign layer2_out[2497] = ~layer1_out[6604] | layer1_out[6605];
    assign layer2_out[2498] = ~layer1_out[1079];
    assign layer2_out[2499] = layer1_out[4057] & ~layer1_out[4056];
    assign layer2_out[2500] = layer1_out[4073] ^ layer1_out[4074];
    assign layer2_out[2501] = ~layer1_out[5982];
    assign layer2_out[2502] = 1'b1;
    assign layer2_out[2503] = ~layer1_out[4444];
    assign layer2_out[2504] = layer1_out[5671];
    assign layer2_out[2505] = ~layer1_out[214] | layer1_out[215];
    assign layer2_out[2506] = layer1_out[126];
    assign layer2_out[2507] = layer1_out[7402] & ~layer1_out[7401];
    assign layer2_out[2508] = layer1_out[3692];
    assign layer2_out[2509] = ~(layer1_out[1368] | layer1_out[1369]);
    assign layer2_out[2510] = layer1_out[5609] & ~layer1_out[5610];
    assign layer2_out[2511] = layer1_out[4579] & ~layer1_out[4578];
    assign layer2_out[2512] = ~layer1_out[3350];
    assign layer2_out[2513] = layer1_out[1780];
    assign layer2_out[2514] = ~layer1_out[593];
    assign layer2_out[2515] = ~layer1_out[4529] | layer1_out[4528];
    assign layer2_out[2516] = layer1_out[1802];
    assign layer2_out[2517] = layer1_out[4700] ^ layer1_out[4701];
    assign layer2_out[2518] = layer1_out[4241] & layer1_out[4242];
    assign layer2_out[2519] = ~layer1_out[6936] | layer1_out[6937];
    assign layer2_out[2520] = layer1_out[7151];
    assign layer2_out[2521] = layer1_out[1115] & ~layer1_out[1114];
    assign layer2_out[2522] = ~(layer1_out[881] ^ layer1_out[882]);
    assign layer2_out[2523] = ~(layer1_out[3210] & layer1_out[3211]);
    assign layer2_out[2524] = layer1_out[3822] & ~layer1_out[3821];
    assign layer2_out[2525] = ~layer1_out[5866];
    assign layer2_out[2526] = ~layer1_out[7153];
    assign layer2_out[2527] = ~layer1_out[4747] | layer1_out[4746];
    assign layer2_out[2528] = 1'b1;
    assign layer2_out[2529] = ~layer1_out[3263];
    assign layer2_out[2530] = ~layer1_out[3956] | layer1_out[3957];
    assign layer2_out[2531] = layer1_out[7001] | layer1_out[7002];
    assign layer2_out[2532] = layer1_out[4616] & ~layer1_out[4617];
    assign layer2_out[2533] = ~layer1_out[7983];
    assign layer2_out[2534] = ~(layer1_out[569] & layer1_out[570]);
    assign layer2_out[2535] = layer1_out[3928] ^ layer1_out[3929];
    assign layer2_out[2536] = layer1_out[1155] & layer1_out[1156];
    assign layer2_out[2537] = ~layer1_out[589];
    assign layer2_out[2538] = 1'b1;
    assign layer2_out[2539] = layer1_out[5634] & ~layer1_out[5633];
    assign layer2_out[2540] = layer1_out[7328];
    assign layer2_out[2541] = ~layer1_out[1740];
    assign layer2_out[2542] = ~(layer1_out[2107] & layer1_out[2108]);
    assign layer2_out[2543] = layer1_out[6726];
    assign layer2_out[2544] = 1'b1;
    assign layer2_out[2545] = layer1_out[3698] ^ layer1_out[3699];
    assign layer2_out[2546] = layer1_out[4602] | layer1_out[4603];
    assign layer2_out[2547] = layer1_out[6186] & ~layer1_out[6185];
    assign layer2_out[2548] = layer1_out[7080];
    assign layer2_out[2549] = layer1_out[7552];
    assign layer2_out[2550] = layer1_out[5731];
    assign layer2_out[2551] = layer1_out[885];
    assign layer2_out[2552] = ~(layer1_out[4276] & layer1_out[4277]);
    assign layer2_out[2553] = ~layer1_out[2717] | layer1_out[2718];
    assign layer2_out[2554] = layer1_out[6842];
    assign layer2_out[2555] = layer1_out[6115] & ~layer1_out[6114];
    assign layer2_out[2556] = ~(layer1_out[7506] & layer1_out[7507]);
    assign layer2_out[2557] = 1'b1;
    assign layer2_out[2558] = layer1_out[1537] & layer1_out[1538];
    assign layer2_out[2559] = layer1_out[7906] | layer1_out[7907];
    assign layer2_out[2560] = ~(layer1_out[5553] & layer1_out[5554]);
    assign layer2_out[2561] = layer1_out[6475] & layer1_out[6476];
    assign layer2_out[2562] = layer1_out[2292] & ~layer1_out[2291];
    assign layer2_out[2563] = ~(layer1_out[391] & layer1_out[392]);
    assign layer2_out[2564] = ~(layer1_out[1032] | layer1_out[1033]);
    assign layer2_out[2565] = ~layer1_out[7032];
    assign layer2_out[2566] = ~(layer1_out[59] ^ layer1_out[60]);
    assign layer2_out[2567] = ~(layer1_out[3412] & layer1_out[3413]);
    assign layer2_out[2568] = ~layer1_out[3546];
    assign layer2_out[2569] = 1'b0;
    assign layer2_out[2570] = ~(layer1_out[3033] ^ layer1_out[3034]);
    assign layer2_out[2571] = layer1_out[4553];
    assign layer2_out[2572] = layer1_out[4633] & layer1_out[4634];
    assign layer2_out[2573] = ~layer1_out[629] | layer1_out[630];
    assign layer2_out[2574] = layer1_out[465] | layer1_out[466];
    assign layer2_out[2575] = layer1_out[1637] ^ layer1_out[1638];
    assign layer2_out[2576] = ~layer1_out[4648];
    assign layer2_out[2577] = layer1_out[3791] & layer1_out[3792];
    assign layer2_out[2578] = layer1_out[1126];
    assign layer2_out[2579] = layer1_out[619] & layer1_out[620];
    assign layer2_out[2580] = layer1_out[7072];
    assign layer2_out[2581] = ~layer1_out[366];
    assign layer2_out[2582] = ~(layer1_out[6504] ^ layer1_out[6505]);
    assign layer2_out[2583] = layer1_out[7077] | layer1_out[7078];
    assign layer2_out[2584] = ~layer1_out[3847];
    assign layer2_out[2585] = 1'b1;
    assign layer2_out[2586] = layer1_out[5836];
    assign layer2_out[2587] = layer1_out[6754];
    assign layer2_out[2588] = layer1_out[2224] & ~layer1_out[2223];
    assign layer2_out[2589] = layer1_out[34] & ~layer1_out[35];
    assign layer2_out[2590] = 1'b1;
    assign layer2_out[2591] = layer1_out[3842] | layer1_out[3843];
    assign layer2_out[2592] = ~layer1_out[3920];
    assign layer2_out[2593] = layer1_out[5573] ^ layer1_out[5574];
    assign layer2_out[2594] = layer1_out[6633] ^ layer1_out[6634];
    assign layer2_out[2595] = ~layer1_out[2782];
    assign layer2_out[2596] = 1'b1;
    assign layer2_out[2597] = layer1_out[1507] & ~layer1_out[1508];
    assign layer2_out[2598] = 1'b1;
    assign layer2_out[2599] = layer1_out[3549] ^ layer1_out[3550];
    assign layer2_out[2600] = layer1_out[25] & ~layer1_out[24];
    assign layer2_out[2601] = ~(layer1_out[5376] ^ layer1_out[5377]);
    assign layer2_out[2602] = layer1_out[7312] | layer1_out[7313];
    assign layer2_out[2603] = layer1_out[7067] ^ layer1_out[7068];
    assign layer2_out[2604] = layer1_out[7697] & ~layer1_out[7696];
    assign layer2_out[2605] = ~(layer1_out[3998] | layer1_out[3999]);
    assign layer2_out[2606] = ~layer1_out[7404];
    assign layer2_out[2607] = ~layer1_out[1621];
    assign layer2_out[2608] = layer1_out[3439] & ~layer1_out[3438];
    assign layer2_out[2609] = layer1_out[1200];
    assign layer2_out[2610] = ~layer1_out[6675] | layer1_out[6674];
    assign layer2_out[2611] = layer1_out[4299];
    assign layer2_out[2612] = layer1_out[5095] & ~layer1_out[5096];
    assign layer2_out[2613] = layer1_out[521] & ~layer1_out[522];
    assign layer2_out[2614] = layer1_out[3556];
    assign layer2_out[2615] = layer1_out[6386];
    assign layer2_out[2616] = ~(layer1_out[3108] | layer1_out[3109]);
    assign layer2_out[2617] = layer1_out[5823];
    assign layer2_out[2618] = layer1_out[7353] & ~layer1_out[7352];
    assign layer2_out[2619] = layer1_out[846] ^ layer1_out[847];
    assign layer2_out[2620] = layer1_out[5791];
    assign layer2_out[2621] = layer1_out[5694];
    assign layer2_out[2622] = layer1_out[3665];
    assign layer2_out[2623] = ~layer1_out[4814];
    assign layer2_out[2624] = ~layer1_out[5958];
    assign layer2_out[2625] = layer1_out[7522] & layer1_out[7523];
    assign layer2_out[2626] = layer1_out[3477] & ~layer1_out[3478];
    assign layer2_out[2627] = layer1_out[5210];
    assign layer2_out[2628] = ~layer1_out[551];
    assign layer2_out[2629] = layer1_out[4795] & ~layer1_out[4796];
    assign layer2_out[2630] = layer1_out[4707] | layer1_out[4708];
    assign layer2_out[2631] = ~layer1_out[5561];
    assign layer2_out[2632] = ~layer1_out[1495];
    assign layer2_out[2633] = layer1_out[3885] & ~layer1_out[3886];
    assign layer2_out[2634] = layer1_out[7697] & layer1_out[7698];
    assign layer2_out[2635] = ~layer1_out[5509];
    assign layer2_out[2636] = ~layer1_out[2652] | layer1_out[2651];
    assign layer2_out[2637] = ~(layer1_out[6893] ^ layer1_out[6894]);
    assign layer2_out[2638] = layer1_out[5784] & layer1_out[5785];
    assign layer2_out[2639] = layer1_out[4493];
    assign layer2_out[2640] = layer1_out[1510];
    assign layer2_out[2641] = ~(layer1_out[3088] ^ layer1_out[3089]);
    assign layer2_out[2642] = ~(layer1_out[27] ^ layer1_out[28]);
    assign layer2_out[2643] = ~(layer1_out[4226] & layer1_out[4227]);
    assign layer2_out[2644] = layer1_out[5686];
    assign layer2_out[2645] = layer1_out[2093] & ~layer1_out[2094];
    assign layer2_out[2646] = layer1_out[741] & ~layer1_out[742];
    assign layer2_out[2647] = ~layer1_out[4734];
    assign layer2_out[2648] = ~(layer1_out[2726] & layer1_out[2727]);
    assign layer2_out[2649] = ~layer1_out[3621];
    assign layer2_out[2650] = ~layer1_out[3306] | layer1_out[3307];
    assign layer2_out[2651] = layer1_out[1731];
    assign layer2_out[2652] = layer1_out[5201];
    assign layer2_out[2653] = layer1_out[7935] & ~layer1_out[7936];
    assign layer2_out[2654] = ~(layer1_out[2144] | layer1_out[2145]);
    assign layer2_out[2655] = layer1_out[3875];
    assign layer2_out[2656] = layer1_out[921] ^ layer1_out[922];
    assign layer2_out[2657] = layer1_out[800] & layer1_out[801];
    assign layer2_out[2658] = layer1_out[7212] | layer1_out[7213];
    assign layer2_out[2659] = ~layer1_out[4917];
    assign layer2_out[2660] = ~layer1_out[5000];
    assign layer2_out[2661] = layer1_out[7950] & ~layer1_out[7951];
    assign layer2_out[2662] = ~layer1_out[5991] | layer1_out[5992];
    assign layer2_out[2663] = layer1_out[7484] & layer1_out[7485];
    assign layer2_out[2664] = ~layer1_out[7800];
    assign layer2_out[2665] = ~layer1_out[7516];
    assign layer2_out[2666] = ~(layer1_out[5491] | layer1_out[5492]);
    assign layer2_out[2667] = layer1_out[6752] & ~layer1_out[6753];
    assign layer2_out[2668] = 1'b1;
    assign layer2_out[2669] = ~(layer1_out[1671] ^ layer1_out[1672]);
    assign layer2_out[2670] = layer1_out[6603] | layer1_out[6604];
    assign layer2_out[2671] = layer1_out[6177] & layer1_out[6178];
    assign layer2_out[2672] = ~layer1_out[5823];
    assign layer2_out[2673] = ~(layer1_out[5262] ^ layer1_out[5263]);
    assign layer2_out[2674] = layer1_out[7123] & layer1_out[7124];
    assign layer2_out[2675] = ~(layer1_out[320] & layer1_out[321]);
    assign layer2_out[2676] = layer1_out[4942] & ~layer1_out[4943];
    assign layer2_out[2677] = ~layer1_out[5971] | layer1_out[5970];
    assign layer2_out[2678] = ~(layer1_out[7660] | layer1_out[7661]);
    assign layer2_out[2679] = layer1_out[6094] & layer1_out[6095];
    assign layer2_out[2680] = layer1_out[7038] & ~layer1_out[7037];
    assign layer2_out[2681] = layer1_out[6281] & layer1_out[6282];
    assign layer2_out[2682] = layer1_out[2078] | layer1_out[2079];
    assign layer2_out[2683] = layer1_out[7713];
    assign layer2_out[2684] = ~layer1_out[6009];
    assign layer2_out[2685] = layer1_out[4742] ^ layer1_out[4743];
    assign layer2_out[2686] = layer1_out[4924] & ~layer1_out[4925];
    assign layer2_out[2687] = ~layer1_out[4031] | layer1_out[4032];
    assign layer2_out[2688] = ~(layer1_out[7612] ^ layer1_out[7613]);
    assign layer2_out[2689] = layer1_out[5271] | layer1_out[5272];
    assign layer2_out[2690] = layer1_out[3083] ^ layer1_out[3084];
    assign layer2_out[2691] = ~layer1_out[3184] | layer1_out[3185];
    assign layer2_out[2692] = layer1_out[447];
    assign layer2_out[2693] = layer1_out[3746] & ~layer1_out[3747];
    assign layer2_out[2694] = ~layer1_out[179];
    assign layer2_out[2695] = ~(layer1_out[5716] | layer1_out[5717]);
    assign layer2_out[2696] = layer1_out[4204];
    assign layer2_out[2697] = layer1_out[6403] ^ layer1_out[6404];
    assign layer2_out[2698] = ~layer1_out[3802];
    assign layer2_out[2699] = layer1_out[5312] & ~layer1_out[5313];
    assign layer2_out[2700] = ~layer1_out[5779];
    assign layer2_out[2701] = layer1_out[5667] & ~layer1_out[5666];
    assign layer2_out[2702] = ~(layer1_out[3799] | layer1_out[3800]);
    assign layer2_out[2703] = ~layer1_out[5826];
    assign layer2_out[2704] = layer1_out[3342] | layer1_out[3343];
    assign layer2_out[2705] = 1'b0;
    assign layer2_out[2706] = layer1_out[7897];
    assign layer2_out[2707] = layer1_out[2178] & ~layer1_out[2177];
    assign layer2_out[2708] = ~layer1_out[7764];
    assign layer2_out[2709] = layer1_out[6849] & layer1_out[6850];
    assign layer2_out[2710] = ~(layer1_out[4190] & layer1_out[4191]);
    assign layer2_out[2711] = ~(layer1_out[4541] | layer1_out[4542]);
    assign layer2_out[2712] = ~layer1_out[5999];
    assign layer2_out[2713] = ~layer1_out[7180];
    assign layer2_out[2714] = layer1_out[4489] & layer1_out[4490];
    assign layer2_out[2715] = ~layer1_out[6343];
    assign layer2_out[2716] = layer1_out[5913] & ~layer1_out[5912];
    assign layer2_out[2717] = ~(layer1_out[1842] | layer1_out[1843]);
    assign layer2_out[2718] = ~layer1_out[3345];
    assign layer2_out[2719] = 1'b0;
    assign layer2_out[2720] = layer1_out[4189] & layer1_out[4190];
    assign layer2_out[2721] = ~layer1_out[4107];
    assign layer2_out[2722] = layer1_out[6057] & ~layer1_out[6056];
    assign layer2_out[2723] = ~layer1_out[4807] | layer1_out[4808];
    assign layer2_out[2724] = layer1_out[6946];
    assign layer2_out[2725] = layer1_out[1567] ^ layer1_out[1568];
    assign layer2_out[2726] = ~layer1_out[6103] | layer1_out[6102];
    assign layer2_out[2727] = layer1_out[5086] ^ layer1_out[5087];
    assign layer2_out[2728] = layer1_out[5800];
    assign layer2_out[2729] = ~layer1_out[2113] | layer1_out[2112];
    assign layer2_out[2730] = layer1_out[6817];
    assign layer2_out[2731] = ~layer1_out[6800] | layer1_out[6801];
    assign layer2_out[2732] = layer1_out[4337];
    assign layer2_out[2733] = layer1_out[5303] & ~layer1_out[5304];
    assign layer2_out[2734] = 1'b0;
    assign layer2_out[2735] = layer1_out[4852];
    assign layer2_out[2736] = layer1_out[7680] & layer1_out[7681];
    assign layer2_out[2737] = layer1_out[5044] ^ layer1_out[5045];
    assign layer2_out[2738] = ~layer1_out[6033];
    assign layer2_out[2739] = layer1_out[6155];
    assign layer2_out[2740] = ~layer1_out[6606] | layer1_out[6605];
    assign layer2_out[2741] = layer1_out[1465];
    assign layer2_out[2742] = layer1_out[295];
    assign layer2_out[2743] = layer1_out[6754] & ~layer1_out[6753];
    assign layer2_out[2744] = layer1_out[2507] ^ layer1_out[2508];
    assign layer2_out[2745] = layer1_out[1720] | layer1_out[1721];
    assign layer2_out[2746] = ~layer1_out[2108];
    assign layer2_out[2747] = layer1_out[6524];
    assign layer2_out[2748] = 1'b1;
    assign layer2_out[2749] = layer1_out[4854] & ~layer1_out[4853];
    assign layer2_out[2750] = ~layer1_out[826];
    assign layer2_out[2751] = 1'b1;
    assign layer2_out[2752] = ~(layer1_out[3891] & layer1_out[3892]);
    assign layer2_out[2753] = ~(layer1_out[6459] & layer1_out[6460]);
    assign layer2_out[2754] = ~layer1_out[502] | layer1_out[501];
    assign layer2_out[2755] = ~(layer1_out[7486] & layer1_out[7487]);
    assign layer2_out[2756] = ~layer1_out[3957];
    assign layer2_out[2757] = layer1_out[1790];
    assign layer2_out[2758] = ~(layer1_out[5692] ^ layer1_out[5693]);
    assign layer2_out[2759] = layer1_out[4787];
    assign layer2_out[2760] = ~(layer1_out[2686] ^ layer1_out[2687]);
    assign layer2_out[2761] = layer1_out[3309];
    assign layer2_out[2762] = layer1_out[2523] & layer1_out[2524];
    assign layer2_out[2763] = layer1_out[6808] & ~layer1_out[6809];
    assign layer2_out[2764] = ~layer1_out[43];
    assign layer2_out[2765] = layer1_out[4920];
    assign layer2_out[2766] = layer1_out[6587] | layer1_out[6588];
    assign layer2_out[2767] = layer1_out[3714] & layer1_out[3715];
    assign layer2_out[2768] = layer1_out[7376];
    assign layer2_out[2769] = layer1_out[5844];
    assign layer2_out[2770] = layer1_out[3956] & ~layer1_out[3955];
    assign layer2_out[2771] = ~layer1_out[1818];
    assign layer2_out[2772] = layer1_out[1109] & layer1_out[1110];
    assign layer2_out[2773] = ~(layer1_out[7521] | layer1_out[7522]);
    assign layer2_out[2774] = ~(layer1_out[2915] ^ layer1_out[2916]);
    assign layer2_out[2775] = layer1_out[4445] & ~layer1_out[4446];
    assign layer2_out[2776] = layer1_out[542];
    assign layer2_out[2777] = layer1_out[6079];
    assign layer2_out[2778] = ~layer1_out[7378];
    assign layer2_out[2779] = layer1_out[4243];
    assign layer2_out[2780] = layer1_out[2905];
    assign layer2_out[2781] = ~layer1_out[7071];
    assign layer2_out[2782] = layer1_out[1253] & ~layer1_out[1252];
    assign layer2_out[2783] = 1'b0;
    assign layer2_out[2784] = layer1_out[232] & ~layer1_out[233];
    assign layer2_out[2785] = layer1_out[7963];
    assign layer2_out[2786] = layer1_out[4579] & ~layer1_out[4580];
    assign layer2_out[2787] = layer1_out[7168];
    assign layer2_out[2788] = ~layer1_out[3128];
    assign layer2_out[2789] = layer1_out[2659];
    assign layer2_out[2790] = ~layer1_out[6068];
    assign layer2_out[2791] = layer1_out[2377];
    assign layer2_out[2792] = ~layer1_out[4488] | layer1_out[4487];
    assign layer2_out[2793] = layer1_out[4954];
    assign layer2_out[2794] = layer1_out[1682] ^ layer1_out[1683];
    assign layer2_out[2795] = ~layer1_out[7472] | layer1_out[7471];
    assign layer2_out[2796] = ~layer1_out[5750];
    assign layer2_out[2797] = ~(layer1_out[7707] & layer1_out[7708]);
    assign layer2_out[2798] = layer1_out[4494] & ~layer1_out[4495];
    assign layer2_out[2799] = ~layer1_out[2015];
    assign layer2_out[2800] = layer1_out[5438];
    assign layer2_out[2801] = ~layer1_out[1892] | layer1_out[1891];
    assign layer2_out[2802] = ~(layer1_out[6755] | layer1_out[6756]);
    assign layer2_out[2803] = ~layer1_out[4431] | layer1_out[4432];
    assign layer2_out[2804] = ~layer1_out[692];
    assign layer2_out[2805] = ~layer1_out[1146];
    assign layer2_out[2806] = layer1_out[1536];
    assign layer2_out[2807] = ~layer1_out[7602] | layer1_out[7601];
    assign layer2_out[2808] = layer1_out[472];
    assign layer2_out[2809] = ~layer1_out[2305];
    assign layer2_out[2810] = layer1_out[2363] & ~layer1_out[2362];
    assign layer2_out[2811] = ~layer1_out[1620];
    assign layer2_out[2812] = ~layer1_out[7902];
    assign layer2_out[2813] = ~layer1_out[758];
    assign layer2_out[2814] = layer1_out[860] | layer1_out[861];
    assign layer2_out[2815] = ~layer1_out[6167] | layer1_out[6168];
    assign layer2_out[2816] = layer1_out[498] & layer1_out[499];
    assign layer2_out[2817] = layer1_out[3771] | layer1_out[3772];
    assign layer2_out[2818] = ~layer1_out[7980] | layer1_out[7979];
    assign layer2_out[2819] = ~layer1_out[7921];
    assign layer2_out[2820] = layer1_out[3895] & ~layer1_out[3894];
    assign layer2_out[2821] = layer1_out[7455] ^ layer1_out[7456];
    assign layer2_out[2822] = ~layer1_out[2174] | layer1_out[2175];
    assign layer2_out[2823] = ~layer1_out[2999];
    assign layer2_out[2824] = ~(layer1_out[1457] & layer1_out[1458]);
    assign layer2_out[2825] = ~layer1_out[6661] | layer1_out[6660];
    assign layer2_out[2826] = layer1_out[5854];
    assign layer2_out[2827] = ~layer1_out[4629];
    assign layer2_out[2828] = ~layer1_out[5264] | layer1_out[5265];
    assign layer2_out[2829] = layer1_out[1093] & ~layer1_out[1094];
    assign layer2_out[2830] = layer1_out[4143] & layer1_out[4144];
    assign layer2_out[2831] = layer1_out[7883] & ~layer1_out[7884];
    assign layer2_out[2832] = layer1_out[465] & ~layer1_out[464];
    assign layer2_out[2833] = layer1_out[3905];
    assign layer2_out[2834] = ~layer1_out[2844] | layer1_out[2843];
    assign layer2_out[2835] = layer1_out[1077];
    assign layer2_out[2836] = ~layer1_out[2918] | layer1_out[2917];
    assign layer2_out[2837] = ~(layer1_out[283] & layer1_out[284]);
    assign layer2_out[2838] = layer1_out[3230];
    assign layer2_out[2839] = layer1_out[4798] & ~layer1_out[4799];
    assign layer2_out[2840] = layer1_out[1159] | layer1_out[1160];
    assign layer2_out[2841] = layer1_out[3068] & ~layer1_out[3067];
    assign layer2_out[2842] = ~layer1_out[3170] | layer1_out[3171];
    assign layer2_out[2843] = layer1_out[3102];
    assign layer2_out[2844] = layer1_out[5210];
    assign layer2_out[2845] = ~layer1_out[3820];
    assign layer2_out[2846] = ~(layer1_out[1461] & layer1_out[1462]);
    assign layer2_out[2847] = ~(layer1_out[2189] ^ layer1_out[2190]);
    assign layer2_out[2848] = ~layer1_out[1349];
    assign layer2_out[2849] = layer1_out[5545];
    assign layer2_out[2850] = layer1_out[3187];
    assign layer2_out[2851] = layer1_out[6414];
    assign layer2_out[2852] = 1'b0;
    assign layer2_out[2853] = ~layer1_out[1397];
    assign layer2_out[2854] = ~layer1_out[2577];
    assign layer2_out[2855] = ~(layer1_out[7867] & layer1_out[7868]);
    assign layer2_out[2856] = ~(layer1_out[2405] | layer1_out[2406]);
    assign layer2_out[2857] = layer1_out[3969] & layer1_out[3970];
    assign layer2_out[2858] = layer1_out[1164] & layer1_out[1165];
    assign layer2_out[2859] = layer1_out[2353];
    assign layer2_out[2860] = layer1_out[4299];
    assign layer2_out[2861] = layer1_out[7811] ^ layer1_out[7812];
    assign layer2_out[2862] = layer1_out[1572] ^ layer1_out[1573];
    assign layer2_out[2863] = ~layer1_out[102];
    assign layer2_out[2864] = ~layer1_out[6121];
    assign layer2_out[2865] = layer1_out[7331] | layer1_out[7332];
    assign layer2_out[2866] = layer1_out[5323] & ~layer1_out[5324];
    assign layer2_out[2867] = 1'b1;
    assign layer2_out[2868] = ~(layer1_out[400] | layer1_out[401]);
    assign layer2_out[2869] = ~(layer1_out[6242] | layer1_out[6243]);
    assign layer2_out[2870] = layer1_out[6105] | layer1_out[6106];
    assign layer2_out[2871] = ~layer1_out[6732];
    assign layer2_out[2872] = ~(layer1_out[4333] & layer1_out[4334]);
    assign layer2_out[2873] = layer1_out[6151];
    assign layer2_out[2874] = layer1_out[2756] & ~layer1_out[2757];
    assign layer2_out[2875] = layer1_out[1708];
    assign layer2_out[2876] = ~layer1_out[2584] | layer1_out[2585];
    assign layer2_out[2877] = ~(layer1_out[5204] & layer1_out[5205]);
    assign layer2_out[2878] = layer1_out[2382];
    assign layer2_out[2879] = ~layer1_out[5277] | layer1_out[5276];
    assign layer2_out[2880] = layer1_out[3579];
    assign layer2_out[2881] = layer1_out[5757];
    assign layer2_out[2882] = ~layer1_out[6017] | layer1_out[6018];
    assign layer2_out[2883] = ~layer1_out[2925];
    assign layer2_out[2884] = ~layer1_out[7230] | layer1_out[7231];
    assign layer2_out[2885] = ~(layer1_out[3111] | layer1_out[3112]);
    assign layer2_out[2886] = ~layer1_out[4767] | layer1_out[4768];
    assign layer2_out[2887] = layer1_out[1314] | layer1_out[1315];
    assign layer2_out[2888] = layer1_out[4083] | layer1_out[4084];
    assign layer2_out[2889] = ~layer1_out[5411];
    assign layer2_out[2890] = 1'b0;
    assign layer2_out[2891] = layer1_out[6250] & ~layer1_out[6251];
    assign layer2_out[2892] = ~layer1_out[5484] | layer1_out[5483];
    assign layer2_out[2893] = ~(layer1_out[6054] ^ layer1_out[6055]);
    assign layer2_out[2894] = layer1_out[6211];
    assign layer2_out[2895] = layer1_out[4712] ^ layer1_out[4713];
    assign layer2_out[2896] = ~layer1_out[3511];
    assign layer2_out[2897] = ~(layer1_out[3848] ^ layer1_out[3849]);
    assign layer2_out[2898] = layer1_out[5473];
    assign layer2_out[2899] = ~layer1_out[2931];
    assign layer2_out[2900] = ~(layer1_out[1402] | layer1_out[1403]);
    assign layer2_out[2901] = ~(layer1_out[6767] & layer1_out[6768]);
    assign layer2_out[2902] = ~layer1_out[4914];
    assign layer2_out[2903] = ~(layer1_out[5878] ^ layer1_out[5879]);
    assign layer2_out[2904] = ~layer1_out[5163] | layer1_out[5164];
    assign layer2_out[2905] = ~layer1_out[4724] | layer1_out[4723];
    assign layer2_out[2906] = ~layer1_out[7760];
    assign layer2_out[2907] = ~layer1_out[4745];
    assign layer2_out[2908] = layer1_out[3102];
    assign layer2_out[2909] = layer1_out[2999] & layer1_out[3000];
    assign layer2_out[2910] = layer1_out[3220] & layer1_out[3221];
    assign layer2_out[2911] = layer1_out[5679];
    assign layer2_out[2912] = layer1_out[5205];
    assign layer2_out[2913] = ~layer1_out[3593];
    assign layer2_out[2914] = ~layer1_out[353];
    assign layer2_out[2915] = layer1_out[276];
    assign layer2_out[2916] = ~layer1_out[5448] | layer1_out[5447];
    assign layer2_out[2917] = ~(layer1_out[5807] & layer1_out[5808]);
    assign layer2_out[2918] = layer1_out[1452];
    assign layer2_out[2919] = ~layer1_out[6588] | layer1_out[6589];
    assign layer2_out[2920] = ~(layer1_out[3096] | layer1_out[3097]);
    assign layer2_out[2921] = ~layer1_out[1176] | layer1_out[1177];
    assign layer2_out[2922] = layer1_out[6774];
    assign layer2_out[2923] = layer1_out[4977] ^ layer1_out[4978];
    assign layer2_out[2924] = ~layer1_out[6564] | layer1_out[6563];
    assign layer2_out[2925] = layer1_out[1239] | layer1_out[1240];
    assign layer2_out[2926] = layer1_out[960];
    assign layer2_out[2927] = layer1_out[3539] ^ layer1_out[3540];
    assign layer2_out[2928] = layer1_out[1835] & ~layer1_out[1836];
    assign layer2_out[2929] = layer1_out[6806] | layer1_out[6807];
    assign layer2_out[2930] = layer1_out[4047] | layer1_out[4048];
    assign layer2_out[2931] = ~layer1_out[2812];
    assign layer2_out[2932] = ~layer1_out[4773] | layer1_out[4772];
    assign layer2_out[2933] = ~layer1_out[5137];
    assign layer2_out[2934] = ~(layer1_out[1333] & layer1_out[1334]);
    assign layer2_out[2935] = ~layer1_out[2268];
    assign layer2_out[2936] = layer1_out[1518] & layer1_out[1519];
    assign layer2_out[2937] = ~(layer1_out[5304] | layer1_out[5305]);
    assign layer2_out[2938] = ~layer1_out[3481];
    assign layer2_out[2939] = ~layer1_out[3389];
    assign layer2_out[2940] = ~(layer1_out[6062] | layer1_out[6063]);
    assign layer2_out[2941] = layer1_out[5260];
    assign layer2_out[2942] = layer1_out[4669] & ~layer1_out[4670];
    assign layer2_out[2943] = layer1_out[4177] & ~layer1_out[4176];
    assign layer2_out[2944] = ~(layer1_out[7649] | layer1_out[7650]);
    assign layer2_out[2945] = ~(layer1_out[3197] & layer1_out[3198]);
    assign layer2_out[2946] = layer1_out[2697] | layer1_out[2698];
    assign layer2_out[2947] = ~layer1_out[4719];
    assign layer2_out[2948] = layer1_out[1068] & ~layer1_out[1069];
    assign layer2_out[2949] = ~layer1_out[7485] | layer1_out[7486];
    assign layer2_out[2950] = layer1_out[4685];
    assign layer2_out[2951] = layer1_out[4908] & layer1_out[4909];
    assign layer2_out[2952] = layer1_out[6932];
    assign layer2_out[2953] = layer1_out[5042] & ~layer1_out[5041];
    assign layer2_out[2954] = layer1_out[7183] | layer1_out[7184];
    assign layer2_out[2955] = layer1_out[7105] & ~layer1_out[7104];
    assign layer2_out[2956] = ~(layer1_out[555] & layer1_out[556]);
    assign layer2_out[2957] = layer1_out[6905] & ~layer1_out[6906];
    assign layer2_out[2958] = ~(layer1_out[3086] | layer1_out[3087]);
    assign layer2_out[2959] = ~layer1_out[3552];
    assign layer2_out[2960] = ~layer1_out[5593] | layer1_out[5592];
    assign layer2_out[2961] = ~layer1_out[2480];
    assign layer2_out[2962] = ~layer1_out[5251] | layer1_out[5252];
    assign layer2_out[2963] = layer1_out[1570] & layer1_out[1571];
    assign layer2_out[2964] = ~layer1_out[4119] | layer1_out[4118];
    assign layer2_out[2965] = ~layer1_out[2736];
    assign layer2_out[2966] = layer1_out[5110] & ~layer1_out[5111];
    assign layer2_out[2967] = ~layer1_out[2542];
    assign layer2_out[2968] = ~(layer1_out[5387] & layer1_out[5388]);
    assign layer2_out[2969] = ~(layer1_out[5806] ^ layer1_out[5807]);
    assign layer2_out[2970] = layer1_out[18] | layer1_out[19];
    assign layer2_out[2971] = ~layer1_out[6892] | layer1_out[6893];
    assign layer2_out[2972] = layer1_out[6788];
    assign layer2_out[2973] = layer1_out[995] | layer1_out[996];
    assign layer2_out[2974] = layer1_out[5219] | layer1_out[5220];
    assign layer2_out[2975] = ~(layer1_out[4501] & layer1_out[4502]);
    assign layer2_out[2976] = ~layer1_out[3797] | layer1_out[3796];
    assign layer2_out[2977] = ~layer1_out[2681] | layer1_out[2682];
    assign layer2_out[2978] = ~(layer1_out[3646] ^ layer1_out[3647]);
    assign layer2_out[2979] = ~layer1_out[4115] | layer1_out[4116];
    assign layer2_out[2980] = ~layer1_out[7825] | layer1_out[7824];
    assign layer2_out[2981] = layer1_out[608] & ~layer1_out[607];
    assign layer2_out[2982] = layer1_out[7608] ^ layer1_out[7609];
    assign layer2_out[2983] = layer1_out[3662] & layer1_out[3663];
    assign layer2_out[2984] = ~layer1_out[5283] | layer1_out[5284];
    assign layer2_out[2985] = ~layer1_out[5990];
    assign layer2_out[2986] = layer1_out[5937];
    assign layer2_out[2987] = layer1_out[4321];
    assign layer2_out[2988] = ~(layer1_out[2031] | layer1_out[2032]);
    assign layer2_out[2989] = layer1_out[4971];
    assign layer2_out[2990] = ~(layer1_out[1953] | layer1_out[1954]);
    assign layer2_out[2991] = layer1_out[7459] & ~layer1_out[7460];
    assign layer2_out[2992] = ~layer1_out[2776] | layer1_out[2775];
    assign layer2_out[2993] = ~layer1_out[3289];
    assign layer2_out[2994] = layer1_out[7135];
    assign layer2_out[2995] = ~layer1_out[2410] | layer1_out[2411];
    assign layer2_out[2996] = ~(layer1_out[5543] ^ layer1_out[5544]);
    assign layer2_out[2997] = ~(layer1_out[1261] & layer1_out[1262]);
    assign layer2_out[2998] = ~layer1_out[2403] | layer1_out[2402];
    assign layer2_out[2999] = ~(layer1_out[4374] & layer1_out[4375]);
    assign layer2_out[3000] = ~layer1_out[2336] | layer1_out[2335];
    assign layer2_out[3001] = layer1_out[1748] & ~layer1_out[1749];
    assign layer2_out[3002] = ~layer1_out[1546];
    assign layer2_out[3003] = ~(layer1_out[2141] & layer1_out[2142]);
    assign layer2_out[3004] = layer1_out[2734] & ~layer1_out[2735];
    assign layer2_out[3005] = ~layer1_out[3609];
    assign layer2_out[3006] = layer1_out[4219] & layer1_out[4220];
    assign layer2_out[3007] = 1'b1;
    assign layer2_out[3008] = 1'b0;
    assign layer2_out[3009] = ~layer1_out[6035];
    assign layer2_out[3010] = layer1_out[7970];
    assign layer2_out[3011] = layer1_out[5039] & ~layer1_out[5040];
    assign layer2_out[3012] = layer1_out[6298];
    assign layer2_out[3013] = ~layer1_out[1341];
    assign layer2_out[3014] = ~(layer1_out[5922] | layer1_out[5923]);
    assign layer2_out[3015] = ~layer1_out[5684];
    assign layer2_out[3016] = layer1_out[7643];
    assign layer2_out[3017] = 1'b1;
    assign layer2_out[3018] = ~layer1_out[5771] | layer1_out[5772];
    assign layer2_out[3019] = layer1_out[6482] | layer1_out[6483];
    assign layer2_out[3020] = ~layer1_out[7884];
    assign layer2_out[3021] = layer1_out[7376] & layer1_out[7377];
    assign layer2_out[3022] = layer1_out[3] & layer1_out[4];
    assign layer2_out[3023] = layer1_out[2656];
    assign layer2_out[3024] = layer1_out[7427];
    assign layer2_out[3025] = 1'b1;
    assign layer2_out[3026] = ~(layer1_out[5715] & layer1_out[5716]);
    assign layer2_out[3027] = 1'b0;
    assign layer2_out[3028] = ~layer1_out[7444];
    assign layer2_out[3029] = ~layer1_out[171];
    assign layer2_out[3030] = ~layer1_out[714];
    assign layer2_out[3031] = ~layer1_out[2540];
    assign layer2_out[3032] = layer1_out[1895] & ~layer1_out[1896];
    assign layer2_out[3033] = ~layer1_out[1053];
    assign layer2_out[3034] = layer1_out[4754] & ~layer1_out[4753];
    assign layer2_out[3035] = ~layer1_out[7774];
    assign layer2_out[3036] = ~layer1_out[6919];
    assign layer2_out[3037] = ~(layer1_out[3208] ^ layer1_out[3209]);
    assign layer2_out[3038] = layer1_out[95] & ~layer1_out[94];
    assign layer2_out[3039] = ~(layer1_out[1804] ^ layer1_out[1805]);
    assign layer2_out[3040] = layer1_out[4314] | layer1_out[4315];
    assign layer2_out[3041] = ~(layer1_out[1683] ^ layer1_out[1684]);
    assign layer2_out[3042] = ~layer1_out[5605];
    assign layer2_out[3043] = layer1_out[2989];
    assign layer2_out[3044] = layer1_out[2817] & ~layer1_out[2818];
    assign layer2_out[3045] = ~layer1_out[2878] | layer1_out[2877];
    assign layer2_out[3046] = layer1_out[4939] & ~layer1_out[4938];
    assign layer2_out[3047] = ~layer1_out[1933] | layer1_out[1932];
    assign layer2_out[3048] = 1'b0;
    assign layer2_out[3049] = ~(layer1_out[7809] | layer1_out[7810]);
    assign layer2_out[3050] = ~(layer1_out[7005] | layer1_out[7006]);
    assign layer2_out[3051] = ~layer1_out[7927];
    assign layer2_out[3052] = layer1_out[7868] & ~layer1_out[7869];
    assign layer2_out[3053] = layer1_out[2660] | layer1_out[2661];
    assign layer2_out[3054] = layer1_out[4719] ^ layer1_out[4720];
    assign layer2_out[3055] = layer1_out[3940] & layer1_out[3941];
    assign layer2_out[3056] = ~layer1_out[4543];
    assign layer2_out[3057] = layer1_out[7570] | layer1_out[7571];
    assign layer2_out[3058] = layer1_out[1473] & ~layer1_out[1474];
    assign layer2_out[3059] = ~layer1_out[3690] | layer1_out[3691];
    assign layer2_out[3060] = ~(layer1_out[3853] ^ layer1_out[3854]);
    assign layer2_out[3061] = layer1_out[7480] & ~layer1_out[7481];
    assign layer2_out[3062] = 1'b0;
    assign layer2_out[3063] = ~layer1_out[719];
    assign layer2_out[3064] = layer1_out[1507] & ~layer1_out[1506];
    assign layer2_out[3065] = ~layer1_out[3382];
    assign layer2_out[3066] = ~layer1_out[6500];
    assign layer2_out[3067] = layer1_out[2994];
    assign layer2_out[3068] = ~(layer1_out[756] & layer1_out[757]);
    assign layer2_out[3069] = layer1_out[7412] & layer1_out[7413];
    assign layer2_out[3070] = ~(layer1_out[2495] & layer1_out[2496]);
    assign layer2_out[3071] = ~layer1_out[7758];
    assign layer2_out[3072] = 1'b0;
    assign layer2_out[3073] = 1'b1;
    assign layer2_out[3074] = layer1_out[5416] | layer1_out[5417];
    assign layer2_out[3075] = 1'b1;
    assign layer2_out[3076] = layer1_out[6216];
    assign layer2_out[3077] = layer1_out[6966];
    assign layer2_out[3078] = layer1_out[6237] & layer1_out[6238];
    assign layer2_out[3079] = ~(layer1_out[343] ^ layer1_out[344]);
    assign layer2_out[3080] = layer1_out[386] | layer1_out[387];
    assign layer2_out[3081] = ~layer1_out[903];
    assign layer2_out[3082] = layer1_out[7614];
    assign layer2_out[3083] = layer1_out[1690] & layer1_out[1691];
    assign layer2_out[3084] = layer1_out[1541];
    assign layer2_out[3085] = layer1_out[5983] & ~layer1_out[5984];
    assign layer2_out[3086] = ~(layer1_out[7624] | layer1_out[7625]);
    assign layer2_out[3087] = ~layer1_out[5112];
    assign layer2_out[3088] = 1'b1;
    assign layer2_out[3089] = ~layer1_out[5052];
    assign layer2_out[3090] = layer1_out[1526];
    assign layer2_out[3091] = layer1_out[4845] & ~layer1_out[4844];
    assign layer2_out[3092] = layer1_out[4434] | layer1_out[4435];
    assign layer2_out[3093] = layer1_out[1714];
    assign layer2_out[3094] = ~layer1_out[1664] | layer1_out[1665];
    assign layer2_out[3095] = layer1_out[7790] & ~layer1_out[7789];
    assign layer2_out[3096] = layer1_out[3584] ^ layer1_out[3585];
    assign layer2_out[3097] = ~(layer1_out[5593] & layer1_out[5594]);
    assign layer2_out[3098] = layer1_out[4460] & ~layer1_out[4459];
    assign layer2_out[3099] = layer1_out[791];
    assign layer2_out[3100] = ~layer1_out[3699];
    assign layer2_out[3101] = layer1_out[5238] & ~layer1_out[5239];
    assign layer2_out[3102] = ~layer1_out[4332];
    assign layer2_out[3103] = ~layer1_out[2122];
    assign layer2_out[3104] = 1'b1;
    assign layer2_out[3105] = layer1_out[5498];
    assign layer2_out[3106] = ~layer1_out[3682];
    assign layer2_out[3107] = ~(layer1_out[3879] ^ layer1_out[3880]);
    assign layer2_out[3108] = layer1_out[6238];
    assign layer2_out[3109] = ~layer1_out[5615] | layer1_out[5616];
    assign layer2_out[3110] = ~(layer1_out[3113] | layer1_out[3114]);
    assign layer2_out[3111] = ~layer1_out[4048];
    assign layer2_out[3112] = ~layer1_out[417];
    assign layer2_out[3113] = ~layer1_out[6638] | layer1_out[6637];
    assign layer2_out[3114] = ~layer1_out[6673] | layer1_out[6674];
    assign layer2_out[3115] = ~(layer1_out[7591] & layer1_out[7592]);
    assign layer2_out[3116] = ~layer1_out[2924] | layer1_out[2923];
    assign layer2_out[3117] = layer1_out[7267];
    assign layer2_out[3118] = ~(layer1_out[1351] ^ layer1_out[1352]);
    assign layer2_out[3119] = 1'b0;
    assign layer2_out[3120] = ~(layer1_out[6339] | layer1_out[6340]);
    assign layer2_out[3121] = 1'b1;
    assign layer2_out[3122] = ~layer1_out[5597] | layer1_out[5596];
    assign layer2_out[3123] = ~layer1_out[6950] | layer1_out[6949];
    assign layer2_out[3124] = ~layer1_out[6002];
    assign layer2_out[3125] = ~layer1_out[6348] | layer1_out[6349];
    assign layer2_out[3126] = ~layer1_out[3072] | layer1_out[3071];
    assign layer2_out[3127] = layer1_out[26] | layer1_out[27];
    assign layer2_out[3128] = layer1_out[3195] & layer1_out[3196];
    assign layer2_out[3129] = layer1_out[2619] & layer1_out[2620];
    assign layer2_out[3130] = ~layer1_out[6204];
    assign layer2_out[3131] = ~(layer1_out[4692] & layer1_out[4693]);
    assign layer2_out[3132] = ~layer1_out[4019] | layer1_out[4018];
    assign layer2_out[3133] = layer1_out[985] | layer1_out[986];
    assign layer2_out[3134] = layer1_out[4873] & ~layer1_out[4874];
    assign layer2_out[3135] = ~layer1_out[1122] | layer1_out[1121];
    assign layer2_out[3136] = 1'b0;
    assign layer2_out[3137] = layer1_out[1378];
    assign layer2_out[3138] = ~layer1_out[2222];
    assign layer2_out[3139] = layer1_out[1140] | layer1_out[1141];
    assign layer2_out[3140] = ~layer1_out[6915] | layer1_out[6916];
    assign layer2_out[3141] = ~layer1_out[4792] | layer1_out[4791];
    assign layer2_out[3142] = layer1_out[1471] & ~layer1_out[1472];
    assign layer2_out[3143] = layer1_out[4210];
    assign layer2_out[3144] = 1'b0;
    assign layer2_out[3145] = ~(layer1_out[3253] ^ layer1_out[3254]);
    assign layer2_out[3146] = ~layer1_out[2027];
    assign layer2_out[3147] = ~layer1_out[7975];
    assign layer2_out[3148] = layer1_out[2677];
    assign layer2_out[3149] = layer1_out[5626];
    assign layer2_out[3150] = 1'b0;
    assign layer2_out[3151] = layer1_out[6834] & ~layer1_out[6833];
    assign layer2_out[3152] = ~(layer1_out[7447] | layer1_out[7448]);
    assign layer2_out[3153] = ~(layer1_out[4161] | layer1_out[4162]);
    assign layer2_out[3154] = 1'b0;
    assign layer2_out[3155] = ~layer1_out[3044] | layer1_out[3043];
    assign layer2_out[3156] = ~layer1_out[1628];
    assign layer2_out[3157] = ~layer1_out[5704];
    assign layer2_out[3158] = layer1_out[2404];
    assign layer2_out[3159] = ~layer1_out[3670];
    assign layer2_out[3160] = layer1_out[4568] | layer1_out[4569];
    assign layer2_out[3161] = ~layer1_out[5324];
    assign layer2_out[3162] = ~layer1_out[6304];
    assign layer2_out[3163] = layer1_out[4533];
    assign layer2_out[3164] = ~layer1_out[3852] | layer1_out[3853];
    assign layer2_out[3165] = layer1_out[6562] & ~layer1_out[6561];
    assign layer2_out[3166] = layer1_out[5395] | layer1_out[5396];
    assign layer2_out[3167] = layer1_out[4522] ^ layer1_out[4523];
    assign layer2_out[3168] = layer1_out[7436];
    assign layer2_out[3169] = layer1_out[5139];
    assign layer2_out[3170] = layer1_out[5938] | layer1_out[5939];
    assign layer2_out[3171] = layer1_out[6840];
    assign layer2_out[3172] = layer1_out[7365] & ~layer1_out[7364];
    assign layer2_out[3173] = layer1_out[6359] & ~layer1_out[6360];
    assign layer2_out[3174] = ~(layer1_out[6428] & layer1_out[6429]);
    assign layer2_out[3175] = 1'b1;
    assign layer2_out[3176] = ~layer1_out[2739];
    assign layer2_out[3177] = layer1_out[862];
    assign layer2_out[3178] = layer1_out[690];
    assign layer2_out[3179] = ~(layer1_out[7084] | layer1_out[7085]);
    assign layer2_out[3180] = ~(layer1_out[5277] | layer1_out[5278]);
    assign layer2_out[3181] = ~layer1_out[3667] | layer1_out[3666];
    assign layer2_out[3182] = ~layer1_out[7198] | layer1_out[7197];
    assign layer2_out[3183] = layer1_out[1776];
    assign layer2_out[3184] = 1'b1;
    assign layer2_out[3185] = layer1_out[3739] | layer1_out[3740];
    assign layer2_out[3186] = ~layer1_out[5887] | layer1_out[5886];
    assign layer2_out[3187] = ~(layer1_out[6581] ^ layer1_out[6582]);
    assign layer2_out[3188] = ~layer1_out[4033];
    assign layer2_out[3189] = layer1_out[4120];
    assign layer2_out[3190] = layer1_out[7206] & layer1_out[7207];
    assign layer2_out[3191] = layer1_out[4521] & ~layer1_out[4520];
    assign layer2_out[3192] = layer1_out[2030] ^ layer1_out[2031];
    assign layer2_out[3193] = layer1_out[2054] | layer1_out[2055];
    assign layer2_out[3194] = layer1_out[6199] & ~layer1_out[6200];
    assign layer2_out[3195] = ~layer1_out[1838] | layer1_out[1837];
    assign layer2_out[3196] = layer1_out[2884] & ~layer1_out[2885];
    assign layer2_out[3197] = ~layer1_out[3827] | layer1_out[3828];
    assign layer2_out[3198] = ~(layer1_out[520] ^ layer1_out[521]);
    assign layer2_out[3199] = ~layer1_out[3876];
    assign layer2_out[3200] = ~(layer1_out[2640] & layer1_out[2641]);
    assign layer2_out[3201] = ~(layer1_out[3243] ^ layer1_out[3244]);
    assign layer2_out[3202] = ~layer1_out[5465] | layer1_out[5464];
    assign layer2_out[3203] = ~layer1_out[5635] | layer1_out[5634];
    assign layer2_out[3204] = ~layer1_out[5051];
    assign layer2_out[3205] = ~layer1_out[6402];
    assign layer2_out[3206] = layer1_out[4235] & ~layer1_out[4234];
    assign layer2_out[3207] = ~(layer1_out[7498] | layer1_out[7499]);
    assign layer2_out[3208] = ~layer1_out[6423];
    assign layer2_out[3209] = ~(layer1_out[644] & layer1_out[645]);
    assign layer2_out[3210] = layer1_out[5539] & layer1_out[5540];
    assign layer2_out[3211] = ~layer1_out[6214];
    assign layer2_out[3212] = ~layer1_out[6539] | layer1_out[6538];
    assign layer2_out[3213] = ~layer1_out[577];
    assign layer2_out[3214] = ~layer1_out[5517];
    assign layer2_out[3215] = ~layer1_out[2876];
    assign layer2_out[3216] = layer1_out[4427] & layer1_out[4428];
    assign layer2_out[3217] = ~layer1_out[1248];
    assign layer2_out[3218] = layer1_out[6575] & layer1_out[6576];
    assign layer2_out[3219] = ~layer1_out[218];
    assign layer2_out[3220] = ~layer1_out[7008];
    assign layer2_out[3221] = ~(layer1_out[5488] ^ layer1_out[5489]);
    assign layer2_out[3222] = ~(layer1_out[6224] & layer1_out[6225]);
    assign layer2_out[3223] = ~layer1_out[7172];
    assign layer2_out[3224] = layer1_out[1678];
    assign layer2_out[3225] = layer1_out[7472] | layer1_out[7473];
    assign layer2_out[3226] = layer1_out[2365] ^ layer1_out[2366];
    assign layer2_out[3227] = layer1_out[5740] & ~layer1_out[5739];
    assign layer2_out[3228] = layer1_out[256];
    assign layer2_out[3229] = ~layer1_out[5726] | layer1_out[5727];
    assign layer2_out[3230] = 1'b0;
    assign layer2_out[3231] = layer1_out[4529] | layer1_out[4530];
    assign layer2_out[3232] = layer1_out[5832];
    assign layer2_out[3233] = layer1_out[7255];
    assign layer2_out[3234] = layer1_out[7442];
    assign layer2_out[3235] = layer1_out[5680];
    assign layer2_out[3236] = layer1_out[3456];
    assign layer2_out[3237] = layer1_out[7994] | layer1_out[7995];
    assign layer2_out[3238] = layer1_out[1853] ^ layer1_out[1854];
    assign layer2_out[3239] = layer1_out[1236] | layer1_out[1237];
    assign layer2_out[3240] = ~(layer1_out[1356] | layer1_out[1357]);
    assign layer2_out[3241] = ~(layer1_out[1884] | layer1_out[1885]);
    assign layer2_out[3242] = ~(layer1_out[2510] | layer1_out[2511]);
    assign layer2_out[3243] = ~layer1_out[5120] | layer1_out[5121];
    assign layer2_out[3244] = layer1_out[6631] & ~layer1_out[6630];
    assign layer2_out[3245] = layer1_out[5518] | layer1_out[5519];
    assign layer2_out[3246] = layer1_out[1053] & ~layer1_out[1052];
    assign layer2_out[3247] = ~layer1_out[2926] | layer1_out[2925];
    assign layer2_out[3248] = layer1_out[336] | layer1_out[337];
    assign layer2_out[3249] = ~layer1_out[7440] | layer1_out[7439];
    assign layer2_out[3250] = layer1_out[1768];
    assign layer2_out[3251] = layer1_out[6951] & ~layer1_out[6950];
    assign layer2_out[3252] = layer1_out[5220];
    assign layer2_out[3253] = layer1_out[2611] & ~layer1_out[2610];
    assign layer2_out[3254] = layer1_out[2826] | layer1_out[2827];
    assign layer2_out[3255] = ~layer1_out[6032];
    assign layer2_out[3256] = ~layer1_out[6546] | layer1_out[6547];
    assign layer2_out[3257] = layer1_out[4384];
    assign layer2_out[3258] = 1'b0;
    assign layer2_out[3259] = layer1_out[5214] & layer1_out[5215];
    assign layer2_out[3260] = ~layer1_out[5202];
    assign layer2_out[3261] = layer1_out[2249];
    assign layer2_out[3262] = ~layer1_out[2537] | layer1_out[2536];
    assign layer2_out[3263] = ~(layer1_out[4285] | layer1_out[4286]);
    assign layer2_out[3264] = layer1_out[7370];
    assign layer2_out[3265] = ~layer1_out[7044];
    assign layer2_out[3266] = ~layer1_out[6981];
    assign layer2_out[3267] = layer1_out[3592];
    assign layer2_out[3268] = ~layer1_out[7262];
    assign layer2_out[3269] = ~layer1_out[819] | layer1_out[820];
    assign layer2_out[3270] = ~layer1_out[566];
    assign layer2_out[3271] = ~layer1_out[4431] | layer1_out[4430];
    assign layer2_out[3272] = ~(layer1_out[1962] ^ layer1_out[1963]);
    assign layer2_out[3273] = layer1_out[1606] & ~layer1_out[1607];
    assign layer2_out[3274] = layer1_out[17];
    assign layer2_out[3275] = ~(layer1_out[7863] & layer1_out[7864]);
    assign layer2_out[3276] = ~layer1_out[3450] | layer1_out[3449];
    assign layer2_out[3277] = ~(layer1_out[5237] | layer1_out[5238]);
    assign layer2_out[3278] = ~layer1_out[2646];
    assign layer2_out[3279] = layer1_out[3751] & ~layer1_out[3750];
    assign layer2_out[3280] = 1'b0;
    assign layer2_out[3281] = ~(layer1_out[1407] | layer1_out[1408]);
    assign layer2_out[3282] = 1'b1;
    assign layer2_out[3283] = layer1_out[1557] | layer1_out[1558];
    assign layer2_out[3284] = ~layer1_out[5854];
    assign layer2_out[3285] = ~layer1_out[6808] | layer1_out[6807];
    assign layer2_out[3286] = layer1_out[7191];
    assign layer2_out[3287] = ~layer1_out[5061] | layer1_out[5062];
    assign layer2_out[3288] = layer1_out[6205];
    assign layer2_out[3289] = layer1_out[5486] & ~layer1_out[5485];
    assign layer2_out[3290] = ~layer1_out[3554] | layer1_out[3553];
    assign layer2_out[3291] = ~(layer1_out[6882] & layer1_out[6883]);
    assign layer2_out[3292] = ~layer1_out[1631] | layer1_out[1632];
    assign layer2_out[3293] = layer1_out[2254] & ~layer1_out[2255];
    assign layer2_out[3294] = ~layer1_out[4567] | layer1_out[4568];
    assign layer2_out[3295] = ~(layer1_out[4773] & layer1_out[4774]);
    assign layer2_out[3296] = ~layer1_out[138];
    assign layer2_out[3297] = layer1_out[4009];
    assign layer2_out[3298] = ~layer1_out[7515];
    assign layer2_out[3299] = layer1_out[6001] ^ layer1_out[6002];
    assign layer2_out[3300] = ~(layer1_out[4237] ^ layer1_out[4238]);
    assign layer2_out[3301] = layer1_out[7712] & ~layer1_out[7711];
    assign layer2_out[3302] = 1'b0;
    assign layer2_out[3303] = ~layer1_out[6682];
    assign layer2_out[3304] = 1'b0;
    assign layer2_out[3305] = layer1_out[280] & ~layer1_out[279];
    assign layer2_out[3306] = layer1_out[7054];
    assign layer2_out[3307] = ~(layer1_out[7398] & layer1_out[7399]);
    assign layer2_out[3308] = ~layer1_out[1559];
    assign layer2_out[3309] = ~(layer1_out[6057] & layer1_out[6058]);
    assign layer2_out[3310] = layer1_out[5897];
    assign layer2_out[3311] = layer1_out[3233];
    assign layer2_out[3312] = layer1_out[5433];
    assign layer2_out[3313] = ~layer1_out[7324];
    assign layer2_out[3314] = layer1_out[1229] & ~layer1_out[1230];
    assign layer2_out[3315] = layer1_out[1711];
    assign layer2_out[3316] = ~layer1_out[6591] | layer1_out[6592];
    assign layer2_out[3317] = ~(layer1_out[4812] & layer1_out[4813]);
    assign layer2_out[3318] = layer1_out[193];
    assign layer2_out[3319] = layer1_out[7400];
    assign layer2_out[3320] = ~layer1_out[7624] | layer1_out[7623];
    assign layer2_out[3321] = layer1_out[6494] ^ layer1_out[6495];
    assign layer2_out[3322] = ~(layer1_out[4800] & layer1_out[4801]);
    assign layer2_out[3323] = ~layer1_out[6679];
    assign layer2_out[3324] = layer1_out[2836] ^ layer1_out[2837];
    assign layer2_out[3325] = ~(layer1_out[329] ^ layer1_out[330]);
    assign layer2_out[3326] = layer1_out[5194];
    assign layer2_out[3327] = ~layer1_out[4440];
    assign layer2_out[3328] = ~layer1_out[3505];
    assign layer2_out[3329] = 1'b1;
    assign layer2_out[3330] = ~(layer1_out[1214] ^ layer1_out[1215]);
    assign layer2_out[3331] = ~(layer1_out[149] ^ layer1_out[150]);
    assign layer2_out[3332] = 1'b0;
    assign layer2_out[3333] = ~layer1_out[1222];
    assign layer2_out[3334] = ~layer1_out[7739];
    assign layer2_out[3335] = ~layer1_out[6850] | layer1_out[6851];
    assign layer2_out[3336] = layer1_out[7263] & layer1_out[7264];
    assign layer2_out[3337] = ~(layer1_out[5187] & layer1_out[5188]);
    assign layer2_out[3338] = layer1_out[5705];
    assign layer2_out[3339] = ~(layer1_out[4114] ^ layer1_out[4115]);
    assign layer2_out[3340] = layer1_out[4686] & layer1_out[4687];
    assign layer2_out[3341] = ~layer1_out[3522];
    assign layer2_out[3342] = layer1_out[6372];
    assign layer2_out[3343] = ~(layer1_out[947] ^ layer1_out[948]);
    assign layer2_out[3344] = ~(layer1_out[2260] ^ layer1_out[2261]);
    assign layer2_out[3345] = ~layer1_out[2636] | layer1_out[2635];
    assign layer2_out[3346] = layer1_out[2807];
    assign layer2_out[3347] = ~(layer1_out[1078] & layer1_out[1079]);
    assign layer2_out[3348] = ~layer1_out[7876] | layer1_out[7875];
    assign layer2_out[3349] = layer1_out[3573] & layer1_out[3574];
    assign layer2_out[3350] = layer1_out[4983];
    assign layer2_out[3351] = ~layer1_out[5796] | layer1_out[5797];
    assign layer2_out[3352] = ~layer1_out[1535];
    assign layer2_out[3353] = ~(layer1_out[381] & layer1_out[382]);
    assign layer2_out[3354] = ~layer1_out[6968];
    assign layer2_out[3355] = ~(layer1_out[894] ^ layer1_out[895]);
    assign layer2_out[3356] = layer1_out[4432];
    assign layer2_out[3357] = layer1_out[3479];
    assign layer2_out[3358] = ~layer1_out[487];
    assign layer2_out[3359] = ~layer1_out[5364];
    assign layer2_out[3360] = layer1_out[4051] ^ layer1_out[4052];
    assign layer2_out[3361] = layer1_out[3261];
    assign layer2_out[3362] = layer1_out[7359];
    assign layer2_out[3363] = layer1_out[310];
    assign layer2_out[3364] = ~(layer1_out[4758] ^ layer1_out[4759]);
    assign layer2_out[3365] = ~layer1_out[32] | layer1_out[33];
    assign layer2_out[3366] = layer1_out[5900];
    assign layer2_out[3367] = ~(layer1_out[2811] ^ layer1_out[2812]);
    assign layer2_out[3368] = ~(layer1_out[610] & layer1_out[611]);
    assign layer2_out[3369] = ~layer1_out[2460];
    assign layer2_out[3370] = layer1_out[176];
    assign layer2_out[3371] = layer1_out[6955] | layer1_out[6956];
    assign layer2_out[3372] = ~(layer1_out[5727] & layer1_out[5728]);
    assign layer2_out[3373] = ~layer1_out[2684];
    assign layer2_out[3374] = ~(layer1_out[6111] & layer1_out[6112]);
    assign layer2_out[3375] = layer1_out[7064] & ~layer1_out[7065];
    assign layer2_out[3376] = layer1_out[2881];
    assign layer2_out[3377] = ~(layer1_out[4659] & layer1_out[4660]);
    assign layer2_out[3378] = ~layer1_out[7145];
    assign layer2_out[3379] = 1'b1;
    assign layer2_out[3380] = ~(layer1_out[5876] & layer1_out[5877]);
    assign layer2_out[3381] = layer1_out[5736];
    assign layer2_out[3382] = layer1_out[6629] ^ layer1_out[6630];
    assign layer2_out[3383] = layer1_out[2853];
    assign layer2_out[3384] = layer1_out[6941];
    assign layer2_out[3385] = ~layer1_out[7842];
    assign layer2_out[3386] = layer1_out[929];
    assign layer2_out[3387] = ~layer1_out[823] | layer1_out[824];
    assign layer2_out[3388] = layer1_out[5926] ^ layer1_out[5927];
    assign layer2_out[3389] = ~layer1_out[2954];
    assign layer2_out[3390] = layer1_out[6667] & layer1_out[6668];
    assign layer2_out[3391] = layer1_out[7441];
    assign layer2_out[3392] = layer1_out[3893] ^ layer1_out[3894];
    assign layer2_out[3393] = ~layer1_out[2014];
    assign layer2_out[3394] = ~(layer1_out[7391] ^ layer1_out[7392]);
    assign layer2_out[3395] = layer1_out[6085];
    assign layer2_out[3396] = layer1_out[5272] & layer1_out[5273];
    assign layer2_out[3397] = ~(layer1_out[5792] ^ layer1_out[5793]);
    assign layer2_out[3398] = ~layer1_out[243] | layer1_out[242];
    assign layer2_out[3399] = ~layer1_out[3360] | layer1_out[3359];
    assign layer2_out[3400] = layer1_out[1448] & layer1_out[1449];
    assign layer2_out[3401] = ~layer1_out[1188];
    assign layer2_out[3402] = layer1_out[5135] & ~layer1_out[5134];
    assign layer2_out[3403] = layer1_out[4876];
    assign layer2_out[3404] = layer1_out[159] & layer1_out[160];
    assign layer2_out[3405] = ~layer1_out[4282] | layer1_out[4281];
    assign layer2_out[3406] = layer1_out[5603] ^ layer1_out[5604];
    assign layer2_out[3407] = ~(layer1_out[1676] ^ layer1_out[1677]);
    assign layer2_out[3408] = layer1_out[3609];
    assign layer2_out[3409] = layer1_out[4422] & layer1_out[4423];
    assign layer2_out[3410] = ~layer1_out[1305];
    assign layer2_out[3411] = layer1_out[5103];
    assign layer2_out[3412] = ~(layer1_out[7859] & layer1_out[7860]);
    assign layer2_out[3413] = layer1_out[1090] ^ layer1_out[1091];
    assign layer2_out[3414] = ~(layer1_out[7841] ^ layer1_out[7842]);
    assign layer2_out[3415] = ~(layer1_out[6895] & layer1_out[6896]);
    assign layer2_out[3416] = ~layer1_out[6537];
    assign layer2_out[3417] = layer1_out[3157] & ~layer1_out[3156];
    assign layer2_out[3418] = layer1_out[4840] & ~layer1_out[4839];
    assign layer2_out[3419] = ~(layer1_out[3755] & layer1_out[3756]);
    assign layer2_out[3420] = layer1_out[3631];
    assign layer2_out[3421] = ~layer1_out[4638];
    assign layer2_out[3422] = layer1_out[204];
    assign layer2_out[3423] = ~layer1_out[6508] | layer1_out[6507];
    assign layer2_out[3424] = layer1_out[739];
    assign layer2_out[3425] = 1'b1;
    assign layer2_out[3426] = layer1_out[6827] | layer1_out[6828];
    assign layer2_out[3427] = layer1_out[3569] & ~layer1_out[3570];
    assign layer2_out[3428] = ~(layer1_out[479] | layer1_out[480]);
    assign layer2_out[3429] = layer1_out[6140] & layer1_out[6141];
    assign layer2_out[3430] = ~layer1_out[2602] | layer1_out[2603];
    assign layer2_out[3431] = layer1_out[5738] & ~layer1_out[5737];
    assign layer2_out[3432] = ~layer1_out[1041];
    assign layer2_out[3433] = layer1_out[2657] & layer1_out[2658];
    assign layer2_out[3434] = ~layer1_out[3703] | layer1_out[3704];
    assign layer2_out[3435] = ~layer1_out[7685];
    assign layer2_out[3436] = ~(layer1_out[6741] & layer1_out[6742]);
    assign layer2_out[3437] = ~(layer1_out[867] & layer1_out[868]);
    assign layer2_out[3438] = layer1_out[5321];
    assign layer2_out[3439] = ~layer1_out[766];
    assign layer2_out[3440] = layer1_out[6363] & ~layer1_out[6362];
    assign layer2_out[3441] = layer1_out[4470];
    assign layer2_out[3442] = ~layer1_out[286];
    assign layer2_out[3443] = layer1_out[3324] | layer1_out[3325];
    assign layer2_out[3444] = layer1_out[1411] & ~layer1_out[1410];
    assign layer2_out[3445] = ~(layer1_out[4120] & layer1_out[4121]);
    assign layer2_out[3446] = layer1_out[1552] & ~layer1_out[1551];
    assign layer2_out[3447] = ~layer1_out[4400] | layer1_out[4401];
    assign layer2_out[3448] = ~(layer1_out[4716] & layer1_out[4717]);
    assign layer2_out[3449] = layer1_out[1521] & ~layer1_out[1520];
    assign layer2_out[3450] = layer1_out[5547];
    assign layer2_out[3451] = ~layer1_out[3436];
    assign layer2_out[3452] = ~layer1_out[7040] | layer1_out[7041];
    assign layer2_out[3453] = ~layer1_out[4709];
    assign layer2_out[3454] = ~(layer1_out[755] & layer1_out[756]);
    assign layer2_out[3455] = layer1_out[2220] | layer1_out[2221];
    assign layer2_out[3456] = layer1_out[4011] & layer1_out[4012];
    assign layer2_out[3457] = ~layer1_out[628];
    assign layer2_out[3458] = ~(layer1_out[1481] | layer1_out[1482]);
    assign layer2_out[3459] = 1'b0;
    assign layer2_out[3460] = ~layer1_out[4044];
    assign layer2_out[3461] = layer1_out[7300] & ~layer1_out[7299];
    assign layer2_out[3462] = layer1_out[7233] & ~layer1_out[7232];
    assign layer2_out[3463] = layer1_out[4831] | layer1_out[4832];
    assign layer2_out[3464] = layer1_out[7062];
    assign layer2_out[3465] = layer1_out[2326] & ~layer1_out[2325];
    assign layer2_out[3466] = layer1_out[1620] & ~layer1_out[1619];
    assign layer2_out[3467] = ~layer1_out[66];
    assign layer2_out[3468] = layer1_out[7162] & layer1_out[7163];
    assign layer2_out[3469] = ~layer1_out[3449];
    assign layer2_out[3470] = layer1_out[5872];
    assign layer2_out[3471] = layer1_out[6814] | layer1_out[6815];
    assign layer2_out[3472] = layer1_out[6824] | layer1_out[6825];
    assign layer2_out[3473] = layer1_out[2280];
    assign layer2_out[3474] = layer1_out[2985] | layer1_out[2986];
    assign layer2_out[3475] = ~layer1_out[4333] | layer1_out[4332];
    assign layer2_out[3476] = ~layer1_out[4222];
    assign layer2_out[3477] = ~(layer1_out[2720] | layer1_out[2721]);
    assign layer2_out[3478] = ~layer1_out[2741];
    assign layer2_out[3479] = ~layer1_out[2919];
    assign layer2_out[3480] = layer1_out[1382] & layer1_out[1383];
    assign layer2_out[3481] = layer1_out[209];
    assign layer2_out[3482] = ~(layer1_out[5053] ^ layer1_out[5054]);
    assign layer2_out[3483] = ~layer1_out[1148] | layer1_out[1147];
    assign layer2_out[3484] = ~layer1_out[2844];
    assign layer2_out[3485] = ~layer1_out[6142] | layer1_out[6143];
    assign layer2_out[3486] = ~(layer1_out[2204] | layer1_out[2205]);
    assign layer2_out[3487] = layer1_out[4212] & ~layer1_out[4211];
    assign layer2_out[3488] = layer1_out[7955] & ~layer1_out[7956];
    assign layer2_out[3489] = ~layer1_out[7774];
    assign layer2_out[3490] = ~(layer1_out[2862] ^ layer1_out[2863]);
    assign layer2_out[3491] = ~layer1_out[3750];
    assign layer2_out[3492] = layer1_out[930] & layer1_out[931];
    assign layer2_out[3493] = ~(layer1_out[539] & layer1_out[540]);
    assign layer2_out[3494] = ~layer1_out[4278] | layer1_out[4279];
    assign layer2_out[3495] = ~layer1_out[7491];
    assign layer2_out[3496] = layer1_out[765] & layer1_out[766];
    assign layer2_out[3497] = 1'b1;
    assign layer2_out[3498] = layer1_out[5096] & layer1_out[5097];
    assign layer2_out[3499] = layer1_out[3754] & layer1_out[3755];
    assign layer2_out[3500] = layer1_out[3763];
    assign layer2_out[3501] = layer1_out[5931];
    assign layer2_out[3502] = layer1_out[1101] & layer1_out[1102];
    assign layer2_out[3503] = ~layer1_out[1184];
    assign layer2_out[3504] = layer1_out[5];
    assign layer2_out[3505] = ~(layer1_out[3100] & layer1_out[3101]);
    assign layer2_out[3506] = layer1_out[3310] & layer1_out[3311];
    assign layer2_out[3507] = ~(layer1_out[3564] | layer1_out[3565]);
    assign layer2_out[3508] = ~(layer1_out[7739] & layer1_out[7740]);
    assign layer2_out[3509] = layer1_out[1885];
    assign layer2_out[3510] = ~(layer1_out[4991] ^ layer1_out[4992]);
    assign layer2_out[3511] = layer1_out[4122] | layer1_out[4123];
    assign layer2_out[3512] = layer1_out[6500];
    assign layer2_out[3513] = layer1_out[7634] & ~layer1_out[7635];
    assign layer2_out[3514] = layer1_out[5408] | layer1_out[5409];
    assign layer2_out[3515] = layer1_out[7503] | layer1_out[7504];
    assign layer2_out[3516] = ~layer1_out[6210] | layer1_out[6209];
    assign layer2_out[3517] = layer1_out[828];
    assign layer2_out[3518] = 1'b0;
    assign layer2_out[3519] = layer1_out[1784] & ~layer1_out[1783];
    assign layer2_out[3520] = ~(layer1_out[3899] & layer1_out[3900]);
    assign layer2_out[3521] = 1'b1;
    assign layer2_out[3522] = ~layer1_out[554];
    assign layer2_out[3523] = ~layer1_out[7970];
    assign layer2_out[3524] = ~(layer1_out[2214] ^ layer1_out[2215]);
    assign layer2_out[3525] = layer1_out[2770];
    assign layer2_out[3526] = ~(layer1_out[2893] ^ layer1_out[2894]);
    assign layer2_out[3527] = layer1_out[7250];
    assign layer2_out[3528] = ~layer1_out[7005];
    assign layer2_out[3529] = layer1_out[7330];
    assign layer2_out[3530] = layer1_out[499] & layer1_out[500];
    assign layer2_out[3531] = layer1_out[4273] & ~layer1_out[4272];
    assign layer2_out[3532] = layer1_out[2659] & ~layer1_out[2658];
    assign layer2_out[3533] = layer1_out[1186] & ~layer1_out[1185];
    assign layer2_out[3534] = layer1_out[4493] & ~layer1_out[4494];
    assign layer2_out[3535] = ~layer1_out[6517] | layer1_out[6518];
    assign layer2_out[3536] = layer1_out[1439];
    assign layer2_out[3537] = layer1_out[348] & ~layer1_out[349];
    assign layer2_out[3538] = layer1_out[1980];
    assign layer2_out[3539] = ~layer1_out[230] | layer1_out[229];
    assign layer2_out[3540] = layer1_out[5629] & ~layer1_out[5628];
    assign layer2_out[3541] = layer1_out[3725] & ~layer1_out[3724];
    assign layer2_out[3542] = ~layer1_out[2360];
    assign layer2_out[3543] = layer1_out[7880];
    assign layer2_out[3544] = ~layer1_out[3953] | layer1_out[3954];
    assign layer2_out[3545] = layer1_out[784];
    assign layer2_out[3546] = layer1_out[2062];
    assign layer2_out[3547] = layer1_out[3280] | layer1_out[3281];
    assign layer2_out[3548] = ~(layer1_out[7987] & layer1_out[7988]);
    assign layer2_out[3549] = layer1_out[2783] ^ layer1_out[2784];
    assign layer2_out[3550] = ~(layer1_out[6638] ^ layer1_out[6639]);
    assign layer2_out[3551] = layer1_out[2943];
    assign layer2_out[3552] = layer1_out[6725] & ~layer1_out[6724];
    assign layer2_out[3553] = layer1_out[4843];
    assign layer2_out[3554] = layer1_out[62] | layer1_out[63];
    assign layer2_out[3555] = ~layer1_out[6917];
    assign layer2_out[3556] = ~layer1_out[1367] | layer1_out[1366];
    assign layer2_out[3557] = layer1_out[1922];
    assign layer2_out[3558] = 1'b1;
    assign layer2_out[3559] = ~(layer1_out[711] & layer1_out[712]);
    assign layer2_out[3560] = layer1_out[7125] & ~layer1_out[7124];
    assign layer2_out[3561] = ~layer1_out[6795];
    assign layer2_out[3562] = layer1_out[7483] ^ layer1_out[7484];
    assign layer2_out[3563] = layer1_out[4880];
    assign layer2_out[3564] = layer1_out[654];
    assign layer2_out[3565] = layer1_out[2636] & ~layer1_out[2637];
    assign layer2_out[3566] = ~layer1_out[4097];
    assign layer2_out[3567] = layer1_out[2799] & layer1_out[2800];
    assign layer2_out[3568] = layer1_out[6797] & ~layer1_out[6798];
    assign layer2_out[3569] = ~(layer1_out[3830] & layer1_out[3831]);
    assign layer2_out[3570] = ~layer1_out[6111];
    assign layer2_out[3571] = ~(layer1_out[3030] ^ layer1_out[3031]);
    assign layer2_out[3572] = layer1_out[2469];
    assign layer2_out[3573] = layer1_out[7706] & ~layer1_out[7707];
    assign layer2_out[3574] = layer1_out[5366];
    assign layer2_out[3575] = layer1_out[5236] | layer1_out[5237];
    assign layer2_out[3576] = ~layer1_out[7339] | layer1_out[7338];
    assign layer2_out[3577] = ~(layer1_out[1566] & layer1_out[1567]);
    assign layer2_out[3578] = ~layer1_out[4815];
    assign layer2_out[3579] = ~(layer1_out[4571] ^ layer1_out[4572]);
    assign layer2_out[3580] = layer1_out[3523];
    assign layer2_out[3581] = layer1_out[4925] | layer1_out[4926];
    assign layer2_out[3582] = layer1_out[3826];
    assign layer2_out[3583] = ~(layer1_out[458] | layer1_out[459]);
    assign layer2_out[3584] = layer1_out[2171];
    assign layer2_out[3585] = layer1_out[3941] | layer1_out[3942];
    assign layer2_out[3586] = ~layer1_out[3296] | layer1_out[3295];
    assign layer2_out[3587] = layer1_out[5779] & ~layer1_out[5778];
    assign layer2_out[3588] = layer1_out[439] & layer1_out[440];
    assign layer2_out[3589] = ~layer1_out[2814] | layer1_out[2815];
    assign layer2_out[3590] = layer1_out[979] | layer1_out[980];
    assign layer2_out[3591] = layer1_out[2560] & layer1_out[2561];
    assign layer2_out[3592] = layer1_out[1060] | layer1_out[1061];
    assign layer2_out[3593] = layer1_out[4575] & layer1_out[4576];
    assign layer2_out[3594] = layer1_out[2962] ^ layer1_out[2963];
    assign layer2_out[3595] = layer1_out[6847];
    assign layer2_out[3596] = ~layer1_out[3981];
    assign layer2_out[3597] = ~(layer1_out[6756] | layer1_out[6757]);
    assign layer2_out[3598] = layer1_out[3647];
    assign layer2_out[3599] = ~layer1_out[6440] | layer1_out[6441];
    assign layer2_out[3600] = layer1_out[2395] | layer1_out[2396];
    assign layer2_out[3601] = layer1_out[4421] ^ layer1_out[4422];
    assign layer2_out[3602] = layer1_out[7964] & ~layer1_out[7965];
    assign layer2_out[3603] = ~layer1_out[3576];
    assign layer2_out[3604] = ~(layer1_out[6719] ^ layer1_out[6720]);
    assign layer2_out[3605] = layer1_out[7205] & ~layer1_out[7204];
    assign layer2_out[3606] = layer1_out[2662] & ~layer1_out[2663];
    assign layer2_out[3607] = layer1_out[1512];
    assign layer2_out[3608] = layer1_out[4360];
    assign layer2_out[3609] = layer1_out[5256] & ~layer1_out[5257];
    assign layer2_out[3610] = ~layer1_out[4793];
    assign layer2_out[3611] = layer1_out[559];
    assign layer2_out[3612] = layer1_out[5927];
    assign layer2_out[3613] = ~layer1_out[2699];
    assign layer2_out[3614] = ~(layer1_out[3273] & layer1_out[3274]);
    assign layer2_out[3615] = ~layer1_out[6217];
    assign layer2_out[3616] = ~layer1_out[4539];
    assign layer2_out[3617] = layer1_out[395] ^ layer1_out[396];
    assign layer2_out[3618] = layer1_out[3374] ^ layer1_out[3375];
    assign layer2_out[3619] = ~layer1_out[1773] | layer1_out[1774];
    assign layer2_out[3620] = 1'b1;
    assign layer2_out[3621] = layer1_out[2342];
    assign layer2_out[3622] = layer1_out[6994] & layer1_out[6995];
    assign layer2_out[3623] = layer1_out[2530] & ~layer1_out[2529];
    assign layer2_out[3624] = ~layer1_out[6814];
    assign layer2_out[3625] = ~layer1_out[7553] | layer1_out[7554];
    assign layer2_out[3626] = ~(layer1_out[5365] | layer1_out[5366]);
    assign layer2_out[3627] = layer1_out[4646] & ~layer1_out[4645];
    assign layer2_out[3628] = 1'b0;
    assign layer2_out[3629] = ~(layer1_out[4900] | layer1_out[4901]);
    assign layer2_out[3630] = layer1_out[5203] | layer1_out[5204];
    assign layer2_out[3631] = ~layer1_out[6972] | layer1_out[6973];
    assign layer2_out[3632] = 1'b1;
    assign layer2_out[3633] = layer1_out[3649] & ~layer1_out[3648];
    assign layer2_out[3634] = ~layer1_out[7456];
    assign layer2_out[3635] = ~layer1_out[5359];
    assign layer2_out[3636] = ~layer1_out[7638] | layer1_out[7637];
    assign layer2_out[3637] = ~layer1_out[2991];
    assign layer2_out[3638] = layer1_out[1671];
    assign layer2_out[3639] = layer1_out[2543] & layer1_out[2544];
    assign layer2_out[3640] = ~(layer1_out[2666] ^ layer1_out[2667]);
    assign layer2_out[3641] = 1'b1;
    assign layer2_out[3642] = ~layer1_out[563] | layer1_out[564];
    assign layer2_out[3643] = layer1_out[4291] & ~layer1_out[4290];
    assign layer2_out[3644] = layer1_out[4218];
    assign layer2_out[3645] = layer1_out[1199];
    assign layer2_out[3646] = ~layer1_out[7743] | layer1_out[7742];
    assign layer2_out[3647] = 1'b1;
    assign layer2_out[3648] = layer1_out[2675] & ~layer1_out[2674];
    assign layer2_out[3649] = ~layer1_out[4683] | layer1_out[4682];
    assign layer2_out[3650] = layer1_out[3013];
    assign layer2_out[3651] = layer1_out[1335] & ~layer1_out[1334];
    assign layer2_out[3652] = ~layer1_out[4008];
    assign layer2_out[3653] = layer1_out[2103] ^ layer1_out[2104];
    assign layer2_out[3654] = layer1_out[5500] & ~layer1_out[5499];
    assign layer2_out[3655] = ~layer1_out[5610];
    assign layer2_out[3656] = layer1_out[1974];
    assign layer2_out[3657] = layer1_out[7430] & ~layer1_out[7429];
    assign layer2_out[3658] = ~(layer1_out[1148] | layer1_out[1149]);
    assign layer2_out[3659] = layer1_out[5680];
    assign layer2_out[3660] = ~(layer1_out[4586] ^ layer1_out[4587]);
    assign layer2_out[3661] = layer1_out[5346] & layer1_out[5347];
    assign layer2_out[3662] = ~layer1_out[965] | layer1_out[964];
    assign layer2_out[3663] = layer1_out[7967];
    assign layer2_out[3664] = layer1_out[3355] & layer1_out[3356];
    assign layer2_out[3665] = layer1_out[4862];
    assign layer2_out[3666] = ~(layer1_out[2912] & layer1_out[2913]);
    assign layer2_out[3667] = ~layer1_out[7737] | layer1_out[7736];
    assign layer2_out[3668] = ~(layer1_out[5586] | layer1_out[5587]);
    assign layer2_out[3669] = ~layer1_out[5824] | layer1_out[5825];
    assign layer2_out[3670] = layer1_out[2368];
    assign layer2_out[3671] = layer1_out[5582];
    assign layer2_out[3672] = layer1_out[3061];
    assign layer2_out[3673] = ~(layer1_out[6569] | layer1_out[6570]);
    assign layer2_out[3674] = layer1_out[235];
    assign layer2_out[3675] = ~layer1_out[2050];
    assign layer2_out[3676] = ~layer1_out[5062];
    assign layer2_out[3677] = ~(layer1_out[1130] | layer1_out[1131]);
    assign layer2_out[3678] = ~(layer1_out[7695] & layer1_out[7696]);
    assign layer2_out[3679] = ~layer1_out[349];
    assign layer2_out[3680] = layer1_out[1751];
    assign layer2_out[3681] = layer1_out[6968] | layer1_out[6969];
    assign layer2_out[3682] = layer1_out[7731];
    assign layer2_out[3683] = ~(layer1_out[3518] & layer1_out[3519]);
    assign layer2_out[3684] = ~(layer1_out[852] ^ layer1_out[853]);
    assign layer2_out[3685] = layer1_out[1524] & ~layer1_out[1523];
    assign layer2_out[3686] = layer1_out[2873] ^ layer1_out[2874];
    assign layer2_out[3687] = 1'b1;
    assign layer2_out[3688] = layer1_out[6087];
    assign layer2_out[3689] = layer1_out[662];
    assign layer2_out[3690] = layer1_out[202];
    assign layer2_out[3691] = layer1_out[1227] ^ layer1_out[1228];
    assign layer2_out[3692] = ~layer1_out[5164] | layer1_out[5165];
    assign layer2_out[3693] = layer1_out[7468];
    assign layer2_out[3694] = ~(layer1_out[2601] | layer1_out[2602]);
    assign layer2_out[3695] = layer1_out[4576] & layer1_out[4577];
    assign layer2_out[3696] = ~(layer1_out[6166] | layer1_out[6167]);
    assign layer2_out[3697] = ~(layer1_out[7659] ^ layer1_out[7660]);
    assign layer2_out[3698] = layer1_out[3150] | layer1_out[3151];
    assign layer2_out[3699] = layer1_out[514];
    assign layer2_out[3700] = layer1_out[1386];
    assign layer2_out[3701] = ~layer1_out[4015] | layer1_out[4014];
    assign layer2_out[3702] = ~layer1_out[3605];
    assign layer2_out[3703] = 1'b0;
    assign layer2_out[3704] = ~layer1_out[3795];
    assign layer2_out[3705] = 1'b0;
    assign layer2_out[3706] = ~(layer1_out[4717] ^ layer1_out[4718]);
    assign layer2_out[3707] = ~layer1_out[4512];
    assign layer2_out[3708] = ~(layer1_out[7119] | layer1_out[7120]);
    assign layer2_out[3709] = ~layer1_out[4002];
    assign layer2_out[3710] = ~layer1_out[7244] | layer1_out[7243];
    assign layer2_out[3711] = ~layer1_out[3667];
    assign layer2_out[3712] = ~layer1_out[648] | layer1_out[647];
    assign layer2_out[3713] = ~layer1_out[6929];
    assign layer2_out[3714] = layer1_out[2329];
    assign layer2_out[3715] = layer1_out[2179] ^ layer1_out[2180];
    assign layer2_out[3716] = layer1_out[2515] & ~layer1_out[2516];
    assign layer2_out[3717] = ~(layer1_out[6230] | layer1_out[6231]);
    assign layer2_out[3718] = ~layer1_out[7689] | layer1_out[7690];
    assign layer2_out[3719] = ~layer1_out[6680] | layer1_out[6679];
    assign layer2_out[3720] = layer1_out[4105];
    assign layer2_out[3721] = ~layer1_out[5859] | layer1_out[5860];
    assign layer2_out[3722] = layer1_out[7373] & layer1_out[7374];
    assign layer2_out[3723] = ~layer1_out[1503];
    assign layer2_out[3724] = ~layer1_out[3327] | layer1_out[3326];
    assign layer2_out[3725] = ~(layer1_out[2048] ^ layer1_out[2049]);
    assign layer2_out[3726] = layer1_out[3022] & ~layer1_out[3023];
    assign layer2_out[3727] = layer1_out[1188] & layer1_out[1189];
    assign layer2_out[3728] = ~layer1_out[2609];
    assign layer2_out[3729] = ~layer1_out[2089] | layer1_out[2088];
    assign layer2_out[3730] = layer1_out[5573] & ~layer1_out[5572];
    assign layer2_out[3731] = layer1_out[6983];
    assign layer2_out[3732] = ~layer1_out[1317];
    assign layer2_out[3733] = layer1_out[31];
    assign layer2_out[3734] = ~layer1_out[5590] | layer1_out[5591];
    assign layer2_out[3735] = ~layer1_out[6070] | layer1_out[6069];
    assign layer2_out[3736] = layer1_out[2256];
    assign layer2_out[3737] = ~(layer1_out[3878] & layer1_out[3879]);
    assign layer2_out[3738] = ~layer1_out[5800] | layer1_out[5799];
    assign layer2_out[3739] = layer1_out[4642] & layer1_out[4643];
    assign layer2_out[3740] = ~(layer1_out[6319] & layer1_out[6320]);
    assign layer2_out[3741] = layer1_out[216];
    assign layer2_out[3742] = ~(layer1_out[4739] & layer1_out[4740]);
    assign layer2_out[3743] = layer1_out[1823];
    assign layer2_out[3744] = layer1_out[246] | layer1_out[247];
    assign layer2_out[3745] = ~layer1_out[1928] | layer1_out[1929];
    assign layer2_out[3746] = layer1_out[3212] & ~layer1_out[3213];
    assign layer2_out[3747] = ~layer1_out[1264];
    assign layer2_out[3748] = ~(layer1_out[5308] | layer1_out[5309]);
    assign layer2_out[3749] = ~layer1_out[2941];
    assign layer2_out[3750] = ~layer1_out[3251];
    assign layer2_out[3751] = layer1_out[2979];
    assign layer2_out[3752] = ~layer1_out[5912];
    assign layer2_out[3753] = 1'b1;
    assign layer2_out[3754] = layer1_out[6825] & layer1_out[6826];
    assign layer2_out[3755] = 1'b1;
    assign layer2_out[3756] = ~layer1_out[1092];
    assign layer2_out[3757] = layer1_out[2713] & ~layer1_out[2714];
    assign layer2_out[3758] = layer1_out[6694] | layer1_out[6695];
    assign layer2_out[3759] = layer1_out[4687] | layer1_out[4688];
    assign layer2_out[3760] = ~(layer1_out[2160] & layer1_out[2161]);
    assign layer2_out[3761] = layer1_out[7535] & ~layer1_out[7534];
    assign layer2_out[3762] = ~(layer1_out[5328] ^ layer1_out[5329]);
    assign layer2_out[3763] = ~layer1_out[7791] | layer1_out[7792];
    assign layer2_out[3764] = ~layer1_out[4996];
    assign layer2_out[3765] = ~(layer1_out[2447] | layer1_out[2448]);
    assign layer2_out[3766] = layer1_out[3434];
    assign layer2_out[3767] = layer1_out[1044];
    assign layer2_out[3768] = ~layer1_out[6248];
    assign layer2_out[3769] = ~layer1_out[799];
    assign layer2_out[3770] = layer1_out[4731];
    assign layer2_out[3771] = 1'b1;
    assign layer2_out[3772] = layer1_out[4461] & ~layer1_out[4460];
    assign layer2_out[3773] = layer1_out[4715];
    assign layer2_out[3774] = ~layer1_out[3686];
    assign layer2_out[3775] = ~(layer1_out[6725] & layer1_out[6726]);
    assign layer2_out[3776] = layer1_out[2678] & layer1_out[2679];
    assign layer2_out[3777] = layer1_out[7889];
    assign layer2_out[3778] = ~layer1_out[1433];
    assign layer2_out[3779] = layer1_out[1740];
    assign layer2_out[3780] = layer1_out[6811];
    assign layer2_out[3781] = 1'b0;
    assign layer2_out[3782] = layer1_out[2377];
    assign layer2_out[3783] = ~layer1_out[1141] | layer1_out[1142];
    assign layer2_out[3784] = layer1_out[7010] | layer1_out[7011];
    assign layer2_out[3785] = ~layer1_out[2509];
    assign layer2_out[3786] = ~(layer1_out[1822] | layer1_out[1823]);
    assign layer2_out[3787] = layer1_out[6116] & ~layer1_out[6117];
    assign layer2_out[3788] = layer1_out[2195] & ~layer1_out[2194];
    assign layer2_out[3789] = layer1_out[4756] & ~layer1_out[4755];
    assign layer2_out[3790] = layer1_out[5009] | layer1_out[5010];
    assign layer2_out[3791] = ~layer1_out[6091] | layer1_out[6090];
    assign layer2_out[3792] = layer1_out[2830];
    assign layer2_out[3793] = layer1_out[2366] | layer1_out[2367];
    assign layer2_out[3794] = ~layer1_out[800];
    assign layer2_out[3795] = layer1_out[2155] & layer1_out[2156];
    assign layer2_out[3796] = layer1_out[3776];
    assign layer2_out[3797] = layer1_out[6771] | layer1_out[6772];
    assign layer2_out[3798] = ~layer1_out[804];
    assign layer2_out[3799] = ~(layer1_out[1527] ^ layer1_out[1528]);
    assign layer2_out[3800] = layer1_out[3846];
    assign layer2_out[3801] = layer1_out[4197];
    assign layer2_out[3802] = layer1_out[4779] & layer1_out[4780];
    assign layer2_out[3803] = ~layer1_out[6485] | layer1_out[6486];
    assign layer2_out[3804] = ~layer1_out[645];
    assign layer2_out[3805] = layer1_out[7351] | layer1_out[7352];
    assign layer2_out[3806] = layer1_out[7795] ^ layer1_out[7796];
    assign layer2_out[3807] = layer1_out[4403] | layer1_out[4404];
    assign layer2_out[3808] = ~layer1_out[6038] | layer1_out[6039];
    assign layer2_out[3809] = ~(layer1_out[4570] & layer1_out[4571]);
    assign layer2_out[3810] = ~layer1_out[4495] | layer1_out[4496];
    assign layer2_out[3811] = layer1_out[5141] ^ layer1_out[5142];
    assign layer2_out[3812] = layer1_out[1495] | layer1_out[1496];
    assign layer2_out[3813] = ~(layer1_out[4732] | layer1_out[4733]);
    assign layer2_out[3814] = layer1_out[149];
    assign layer2_out[3815] = ~layer1_out[1592] | layer1_out[1593];
    assign layer2_out[3816] = layer1_out[6288];
    assign layer2_out[3817] = layer1_out[3763] & layer1_out[3764];
    assign layer2_out[3818] = layer1_out[2006];
    assign layer2_out[3819] = layer1_out[5864];
    assign layer2_out[3820] = layer1_out[6124];
    assign layer2_out[3821] = ~(layer1_out[4068] & layer1_out[4069]);
    assign layer2_out[3822] = ~layer1_out[2113];
    assign layer2_out[3823] = layer1_out[4930];
    assign layer2_out[3824] = ~layer1_out[3687];
    assign layer2_out[3825] = layer1_out[2028];
    assign layer2_out[3826] = 1'b0;
    assign layer2_out[3827] = ~layer1_out[2719] | layer1_out[2718];
    assign layer2_out[3828] = ~layer1_out[5885];
    assign layer2_out[3829] = ~layer1_out[252] | layer1_out[253];
    assign layer2_out[3830] = ~(layer1_out[5951] | layer1_out[5952]);
    assign layer2_out[3831] = layer1_out[4296] ^ layer1_out[4297];
    assign layer2_out[3832] = ~(layer1_out[3047] | layer1_out[3048]);
    assign layer2_out[3833] = 1'b0;
    assign layer2_out[3834] = layer1_out[6050] & ~layer1_out[6051];
    assign layer2_out[3835] = layer1_out[6415];
    assign layer2_out[3836] = layer1_out[664];
    assign layer2_out[3837] = ~(layer1_out[7395] & layer1_out[7396]);
    assign layer2_out[3838] = layer1_out[4072] | layer1_out[4073];
    assign layer2_out[3839] = ~(layer1_out[1454] | layer1_out[1455]);
    assign layer2_out[3840] = ~layer1_out[3500];
    assign layer2_out[3841] = layer1_out[1854] & layer1_out[1855];
    assign layer2_out[3842] = layer1_out[2585] & ~layer1_out[2586];
    assign layer2_out[3843] = layer1_out[2300] & ~layer1_out[2299];
    assign layer2_out[3844] = layer1_out[6367] | layer1_out[6368];
    assign layer2_out[3845] = layer1_out[5420] & layer1_out[5421];
    assign layer2_out[3846] = ~layer1_out[3181];
    assign layer2_out[3847] = ~layer1_out[3376];
    assign layer2_out[3848] = ~layer1_out[92];
    assign layer2_out[3849] = layer1_out[1254] & layer1_out[1255];
    assign layer2_out[3850] = ~layer1_out[5002];
    assign layer2_out[3851] = ~layer1_out[199] | layer1_out[198];
    assign layer2_out[3852] = layer1_out[7130];
    assign layer2_out[3853] = layer1_out[6404] | layer1_out[6405];
    assign layer2_out[3854] = layer1_out[1639] & layer1_out[1640];
    assign layer2_out[3855] = ~layer1_out[4525] | layer1_out[4526];
    assign layer2_out[3856] = ~layer1_out[3526] | layer1_out[3527];
    assign layer2_out[3857] = ~layer1_out[6840] | layer1_out[6839];
    assign layer2_out[3858] = layer1_out[7857] & ~layer1_out[7858];
    assign layer2_out[3859] = layer1_out[1085];
    assign layer2_out[3860] = ~layer1_out[5840] | layer1_out[5841];
    assign layer2_out[3861] = ~layer1_out[6074];
    assign layer2_out[3862] = ~layer1_out[1780];
    assign layer2_out[3863] = layer1_out[696] & ~layer1_out[697];
    assign layer2_out[3864] = layer1_out[6148] ^ layer1_out[6149];
    assign layer2_out[3865] = layer1_out[6880] & ~layer1_out[6881];
    assign layer2_out[3866] = layer1_out[1582];
    assign layer2_out[3867] = layer1_out[6929] & ~layer1_out[6928];
    assign layer2_out[3868] = layer1_out[3413] & ~layer1_out[3414];
    assign layer2_out[3869] = layer1_out[4662];
    assign layer2_out[3870] = layer1_out[5067] & ~layer1_out[5066];
    assign layer2_out[3871] = ~layer1_out[6295];
    assign layer2_out[3872] = layer1_out[3983];
    assign layer2_out[3873] = layer1_out[341];
    assign layer2_out[3874] = 1'b0;
    assign layer2_out[3875] = layer1_out[6403] & ~layer1_out[6402];
    assign layer2_out[3876] = ~layer1_out[7558];
    assign layer2_out[3877] = ~layer1_out[7641] | layer1_out[7640];
    assign layer2_out[3878] = layer1_out[1658] | layer1_out[1659];
    assign layer2_out[3879] = layer1_out[1882] ^ layer1_out[1883];
    assign layer2_out[3880] = ~layer1_out[2034];
    assign layer2_out[3881] = ~layer1_out[3806];
    assign layer2_out[3882] = 1'b1;
    assign layer2_out[3883] = ~(layer1_out[1870] & layer1_out[1871]);
    assign layer2_out[3884] = 1'b0;
    assign layer2_out[3885] = layer1_out[890] & layer1_out[891];
    assign layer2_out[3886] = ~(layer1_out[4665] | layer1_out[4666]);
    assign layer2_out[3887] = ~layer1_out[7417];
    assign layer2_out[3888] = ~layer1_out[7603];
    assign layer2_out[3889] = layer1_out[1812] & ~layer1_out[1813];
    assign layer2_out[3890] = layer1_out[6449];
    assign layer2_out[3891] = layer1_out[7137] & layer1_out[7138];
    assign layer2_out[3892] = ~layer1_out[5652] | layer1_out[5651];
    assign layer2_out[3893] = ~layer1_out[3165];
    assign layer2_out[3894] = layer1_out[380];
    assign layer2_out[3895] = ~layer1_out[7313];
    assign layer2_out[3896] = layer1_out[6341] | layer1_out[6342];
    assign layer2_out[3897] = ~(layer1_out[3833] | layer1_out[3834]);
    assign layer2_out[3898] = layer1_out[3961];
    assign layer2_out[3899] = ~layer1_out[5929];
    assign layer2_out[3900] = layer1_out[4000];
    assign layer2_out[3901] = ~layer1_out[971];
    assign layer2_out[3902] = ~(layer1_out[7013] | layer1_out[7014]);
    assign layer2_out[3903] = ~layer1_out[5082];
    assign layer2_out[3904] = 1'b1;
    assign layer2_out[3905] = ~layer1_out[2615];
    assign layer2_out[3906] = layer1_out[1267] ^ layer1_out[1268];
    assign layer2_out[3907] = ~(layer1_out[2317] | layer1_out[2318]);
    assign layer2_out[3908] = ~layer1_out[3352];
    assign layer2_out[3909] = layer1_out[4785] ^ layer1_out[4786];
    assign layer2_out[3910] = layer1_out[7825] & ~layer1_out[7826];
    assign layer2_out[3911] = ~layer1_out[2474];
    assign layer2_out[3912] = ~(layer1_out[5548] | layer1_out[5549]);
    assign layer2_out[3913] = ~(layer1_out[473] | layer1_out[474]);
    assign layer2_out[3914] = layer1_out[7185] & ~layer1_out[7186];
    assign layer2_out[3915] = layer1_out[3765] & ~layer1_out[3764];
    assign layer2_out[3916] = ~layer1_out[4386] | layer1_out[4387];
    assign layer2_out[3917] = ~layer1_out[2288];
    assign layer2_out[3918] = layer1_out[5454];
    assign layer2_out[3919] = layer1_out[3294] & ~layer1_out[3293];
    assign layer2_out[3920] = layer1_out[5379];
    assign layer2_out[3921] = ~layer1_out[3466] | layer1_out[3465];
    assign layer2_out[3922] = layer1_out[6503] & ~layer1_out[6504];
    assign layer2_out[3923] = ~(layer1_out[4313] | layer1_out[4314]);
    assign layer2_out[3924] = ~layer1_out[3943];
    assign layer2_out[3925] = ~layer1_out[1439];
    assign layer2_out[3926] = 1'b1;
    assign layer2_out[3927] = 1'b0;
    assign layer2_out[3928] = ~layer1_out[2829] | layer1_out[2828];
    assign layer2_out[3929] = ~layer1_out[6192] | layer1_out[6193];
    assign layer2_out[3930] = layer1_out[4561] | layer1_out[4562];
    assign layer2_out[3931] = ~layer1_out[910];
    assign layer2_out[3932] = layer1_out[4213] & layer1_out[4214];
    assign layer2_out[3933] = 1'b0;
    assign layer2_out[3934] = ~(layer1_out[1552] ^ layer1_out[1553]);
    assign layer2_out[3935] = ~(layer1_out[676] & layer1_out[677]);
    assign layer2_out[3936] = ~layer1_out[1318];
    assign layer2_out[3937] = ~layer1_out[6317];
    assign layer2_out[3938] = ~(layer1_out[3457] ^ layer1_out[3458]);
    assign layer2_out[3939] = layer1_out[5161] & ~layer1_out[5162];
    assign layer2_out[3940] = layer1_out[3315];
    assign layer2_out[3941] = layer1_out[6041] ^ layer1_out[6042];
    assign layer2_out[3942] = ~(layer1_out[1616] & layer1_out[1617]);
    assign layer2_out[3943] = layer1_out[3118];
    assign layer2_out[3944] = ~(layer1_out[7164] ^ layer1_out[7165]);
    assign layer2_out[3945] = ~layer1_out[1941];
    assign layer2_out[3946] = ~(layer1_out[5916] ^ layer1_out[5917]);
    assign layer2_out[3947] = ~layer1_out[1848];
    assign layer2_out[3948] = ~layer1_out[3132] | layer1_out[3131];
    assign layer2_out[3949] = ~layer1_out[3209];
    assign layer2_out[3950] = layer1_out[4361];
    assign layer2_out[3951] = layer1_out[3854] & layer1_out[3855];
    assign layer2_out[3952] = layer1_out[1225] & ~layer1_out[1226];
    assign layer2_out[3953] = layer1_out[1353];
    assign layer2_out[3954] = ~layer1_out[2589];
    assign layer2_out[3955] = ~layer1_out[4635];
    assign layer2_out[3956] = layer1_out[6364] ^ layer1_out[6365];
    assign layer2_out[3957] = layer1_out[955] & ~layer1_out[954];
    assign layer2_out[3958] = ~layer1_out[329] | layer1_out[328];
    assign layer2_out[3959] = layer1_out[3204] & ~layer1_out[3205];
    assign layer2_out[3960] = ~layer1_out[4188] | layer1_out[4187];
    assign layer2_out[3961] = ~layer1_out[6669];
    assign layer2_out[3962] = layer1_out[3132] & ~layer1_out[3133];
    assign layer2_out[3963] = ~layer1_out[2329];
    assign layer2_out[3964] = ~layer1_out[2270] | layer1_out[2271];
    assign layer2_out[3965] = layer1_out[4794];
    assign layer2_out[3966] = layer1_out[937] ^ layer1_out[938];
    assign layer2_out[3967] = 1'b1;
    assign layer2_out[3968] = 1'b1;
    assign layer2_out[3969] = layer1_out[7837] & layer1_out[7838];
    assign layer2_out[3970] = ~layer1_out[6202];
    assign layer2_out[3971] = ~layer1_out[6747] | layer1_out[6748];
    assign layer2_out[3972] = layer1_out[5462] & ~layer1_out[5461];
    assign layer2_out[3973] = ~layer1_out[4832] | layer1_out[4833];
    assign layer2_out[3974] = layer1_out[2538];
    assign layer2_out[3975] = layer1_out[513] | layer1_out[514];
    assign layer2_out[3976] = ~layer1_out[4727];
    assign layer2_out[3977] = ~layer1_out[525];
    assign layer2_out[3978] = ~(layer1_out[333] ^ layer1_out[334]);
    assign layer2_out[3979] = ~(layer1_out[903] & layer1_out[904]);
    assign layer2_out[3980] = layer1_out[1205];
    assign layer2_out[3981] = layer1_out[2448] & layer1_out[2449];
    assign layer2_out[3982] = layer1_out[4039];
    assign layer2_out[3983] = layer1_out[7634] & ~layer1_out[7633];
    assign layer2_out[3984] = ~(layer1_out[5580] ^ layer1_out[5581]);
    assign layer2_out[3985] = layer1_out[510];
    assign layer2_out[3986] = ~layer1_out[4524];
    assign layer2_out[3987] = layer1_out[4677] & ~layer1_out[4676];
    assign layer2_out[3988] = layer1_out[1094] | layer1_out[1095];
    assign layer2_out[3989] = layer1_out[4964];
    assign layer2_out[3990] = ~layer1_out[1151] | layer1_out[1150];
    assign layer2_out[3991] = ~(layer1_out[7567] | layer1_out[7568]);
    assign layer2_out[3992] = ~layer1_out[2423];
    assign layer2_out[3993] = layer1_out[1249] | layer1_out[1250];
    assign layer2_out[3994] = layer1_out[298] & ~layer1_out[299];
    assign layer2_out[3995] = layer1_out[3023];
    assign layer2_out[3996] = ~layer1_out[7821] | layer1_out[7820];
    assign layer2_out[3997] = layer1_out[1058];
    assign layer2_out[3998] = layer1_out[5428];
    assign layer2_out[3999] = layer1_out[6704] & ~layer1_out[6703];
    assign layer2_out[4000] = ~layer1_out[5936];
    assign layer2_out[4001] = layer1_out[6595] | layer1_out[6596];
    assign layer2_out[4002] = layer1_out[6425];
    assign layer2_out[4003] = layer1_out[1816];
    assign layer2_out[4004] = layer1_out[3748];
    assign layer2_out[4005] = ~(layer1_out[2224] & layer1_out[2225]);
    assign layer2_out[4006] = ~layer1_out[1897];
    assign layer2_out[4007] = layer1_out[2349] ^ layer1_out[2350];
    assign layer2_out[4008] = layer1_out[4803] & ~layer1_out[4804];
    assign layer2_out[4009] = layer1_out[5810] ^ layer1_out[5811];
    assign layer2_out[4010] = ~(layer1_out[1679] & layer1_out[1680]);
    assign layer2_out[4011] = ~layer1_out[3959] | layer1_out[3960];
    assign layer2_out[4012] = layer1_out[1405];
    assign layer2_out[4013] = ~(layer1_out[3055] & layer1_out[3056]);
    assign layer2_out[4014] = ~(layer1_out[7063] & layer1_out[7064]);
    assign layer2_out[4015] = 1'b0;
    assign layer2_out[4016] = layer1_out[3137] & layer1_out[3138];
    assign layer2_out[4017] = layer1_out[3483] & layer1_out[3484];
    assign layer2_out[4018] = layer1_out[3669];
    assign layer2_out[4019] = layer1_out[3531];
    assign layer2_out[4020] = ~(layer1_out[834] & layer1_out[835]);
    assign layer2_out[4021] = layer1_out[7541];
    assign layer2_out[4022] = ~(layer1_out[7073] & layer1_out[7074]);
    assign layer2_out[4023] = ~(layer1_out[4674] | layer1_out[4675]);
    assign layer2_out[4024] = ~(layer1_out[3990] | layer1_out[3991]);
    assign layer2_out[4025] = 1'b0;
    assign layer2_out[4026] = ~(layer1_out[745] & layer1_out[746]);
    assign layer2_out[4027] = layer1_out[4143];
    assign layer2_out[4028] = ~layer1_out[6123];
    assign layer2_out[4029] = ~(layer1_out[3105] ^ layer1_out[3106]);
    assign layer2_out[4030] = 1'b1;
    assign layer2_out[4031] = layer1_out[5190];
    assign layer2_out[4032] = layer1_out[1858] & layer1_out[1859];
    assign layer2_out[4033] = ~layer1_out[4479] | layer1_out[4478];
    assign layer2_out[4034] = ~layer1_out[7684];
    assign layer2_out[4035] = ~layer1_out[4516] | layer1_out[4515];
    assign layer2_out[4036] = layer1_out[4539] & ~layer1_out[4540];
    assign layer2_out[4037] = ~(layer1_out[5545] & layer1_out[5546]);
    assign layer2_out[4038] = ~layer1_out[4700];
    assign layer2_out[4039] = layer1_out[6227];
    assign layer2_out[4040] = layer1_out[2472];
    assign layer2_out[4041] = ~layer1_out[6692] | layer1_out[6693];
    assign layer2_out[4042] = ~(layer1_out[1287] & layer1_out[1288]);
    assign layer2_out[4043] = layer1_out[2700];
    assign layer2_out[4044] = ~(layer1_out[7024] ^ layer1_out[7025]);
    assign layer2_out[4045] = ~layer1_out[4624];
    assign layer2_out[4046] = layer1_out[4087];
    assign layer2_out[4047] = 1'b1;
    assign layer2_out[4048] = layer1_out[2525] ^ layer1_out[2526];
    assign layer2_out[4049] = ~(layer1_out[3849] | layer1_out[3850]);
    assign layer2_out[4050] = layer1_out[3418] & layer1_out[3419];
    assign layer2_out[4051] = layer1_out[5089];
    assign layer2_out[4052] = layer1_out[152] & layer1_out[153];
    assign layer2_out[4053] = 1'b1;
    assign layer2_out[4054] = layer1_out[158];
    assign layer2_out[4055] = ~layer1_out[535] | layer1_out[534];
    assign layer2_out[4056] = layer1_out[2768] & layer1_out[2769];
    assign layer2_out[4057] = layer1_out[2776] & layer1_out[2777];
    assign layer2_out[4058] = layer1_out[2888];
    assign layer2_out[4059] = layer1_out[5268] | layer1_out[5269];
    assign layer2_out[4060] = layer1_out[6466] & ~layer1_out[6467];
    assign layer2_out[4061] = layer1_out[2165];
    assign layer2_out[4062] = ~layer1_out[4915] | layer1_out[4916];
    assign layer2_out[4063] = layer1_out[7109] & ~layer1_out[7108];
    assign layer2_out[4064] = ~(layer1_out[4650] & layer1_out[4651]);
    assign layer2_out[4065] = ~(layer1_out[3616] ^ layer1_out[3617]);
    assign layer2_out[4066] = ~(layer1_out[6422] ^ layer1_out[6423]);
    assign layer2_out[4067] = ~layer1_out[1349];
    assign layer2_out[4068] = ~layer1_out[2047] | layer1_out[2048];
    assign layer2_out[4069] = 1'b0;
    assign layer2_out[4070] = ~layer1_out[7368] | layer1_out[7369];
    assign layer2_out[4071] = layer1_out[5941];
    assign layer2_out[4072] = layer1_out[2631];
    assign layer2_out[4073] = ~layer1_out[777];
    assign layer2_out[4074] = layer1_out[4221] ^ layer1_out[4222];
    assign layer2_out[4075] = 1'b1;
    assign layer2_out[4076] = layer1_out[2843];
    assign layer2_out[4077] = layer1_out[60];
    assign layer2_out[4078] = 1'b0;
    assign layer2_out[4079] = ~(layer1_out[7378] & layer1_out[7379]);
    assign layer2_out[4080] = ~layer1_out[3727];
    assign layer2_out[4081] = ~(layer1_out[4090] ^ layer1_out[4091]);
    assign layer2_out[4082] = layer1_out[1491];
    assign layer2_out[4083] = layer1_out[4496];
    assign layer2_out[4084] = layer1_out[4627];
    assign layer2_out[4085] = ~layer1_out[5721] | layer1_out[5720];
    assign layer2_out[4086] = ~layer1_out[4891];
    assign layer2_out[4087] = ~layer1_out[1341];
    assign layer2_out[4088] = 1'b0;
    assign layer2_out[4089] = ~layer1_out[2707] | layer1_out[2708];
    assign layer2_out[4090] = layer1_out[7459];
    assign layer2_out[4091] = 1'b1;
    assign layer2_out[4092] = ~layer1_out[4024];
    assign layer2_out[4093] = 1'b0;
    assign layer2_out[4094] = ~(layer1_out[1295] & layer1_out[1296]);
    assign layer2_out[4095] = ~(layer1_out[139] ^ layer1_out[140]);
    assign layer2_out[4096] = layer1_out[4691] ^ layer1_out[4692];
    assign layer2_out[4097] = ~layer1_out[7190];
    assign layer2_out[4098] = layer1_out[1669] & ~layer1_out[1670];
    assign layer2_out[4099] = layer1_out[2644];
    assign layer2_out[4100] = ~layer1_out[2465] | layer1_out[2466];
    assign layer2_out[4101] = ~(layer1_out[546] | layer1_out[547]);
    assign layer2_out[4102] = 1'b0;
    assign layer2_out[4103] = ~layer1_out[4016];
    assign layer2_out[4104] = layer1_out[3174];
    assign layer2_out[4105] = ~layer1_out[2849] | layer1_out[2848];
    assign layer2_out[4106] = layer1_out[5226];
    assign layer2_out[4107] = ~(layer1_out[7598] & layer1_out[7599]);
    assign layer2_out[4108] = layer1_out[7074];
    assign layer2_out[4109] = ~(layer1_out[3268] ^ layer1_out[3269]);
    assign layer2_out[4110] = layer1_out[2654];
    assign layer2_out[4111] = layer1_out[2895];
    assign layer2_out[4112] = layer1_out[2860] & layer1_out[2861];
    assign layer2_out[4113] = layer1_out[3147];
    assign layer2_out[4114] = layer1_out[1845] ^ layer1_out[1846];
    assign layer2_out[4115] = layer1_out[7058] & layer1_out[7059];
    assign layer2_out[4116] = ~layer1_out[1187];
    assign layer2_out[4117] = ~(layer1_out[5985] ^ layer1_out[5986]);
    assign layer2_out[4118] = layer1_out[4618] | layer1_out[4619];
    assign layer2_out[4119] = ~(layer1_out[4060] & layer1_out[4061]);
    assign layer2_out[4120] = ~layer1_out[7346] | layer1_out[7347];
    assign layer2_out[4121] = layer1_out[5292] & layer1_out[5293];
    assign layer2_out[4122] = layer1_out[3032];
    assign layer2_out[4123] = layer1_out[1491];
    assign layer2_out[4124] = layer1_out[1607];
    assign layer2_out[4125] = ~layer1_out[5066];
    assign layer2_out[4126] = layer1_out[5467];
    assign layer2_out[4127] = layer1_out[1983] ^ layer1_out[1984];
    assign layer2_out[4128] = layer1_out[7622] & ~layer1_out[7623];
    assign layer2_out[4129] = ~layer1_out[2969] | layer1_out[2970];
    assign layer2_out[4130] = ~layer1_out[3651] | layer1_out[3650];
    assign layer2_out[4131] = layer1_out[1601] & ~layer1_out[1600];
    assign layer2_out[4132] = ~(layer1_out[7219] ^ layer1_out[7220]);
    assign layer2_out[4133] = layer1_out[1205] ^ layer1_out[1206];
    assign layer2_out[4134] = layer1_out[6724];
    assign layer2_out[4135] = ~(layer1_out[3507] ^ layer1_out[3508]);
    assign layer2_out[4136] = ~layer1_out[2308];
    assign layer2_out[4137] = ~layer1_out[5753];
    assign layer2_out[4138] = layer1_out[116] ^ layer1_out[117];
    assign layer2_out[4139] = layer1_out[2987];
    assign layer2_out[4140] = layer1_out[4748];
    assign layer2_out[4141] = layer1_out[1231];
    assign layer2_out[4142] = ~layer1_out[4901];
    assign layer2_out[4143] = ~layer1_out[3654] | layer1_out[3655];
    assign layer2_out[4144] = ~(layer1_out[4164] & layer1_out[4165]);
    assign layer2_out[4145] = layer1_out[2438] | layer1_out[2439];
    assign layer2_out[4146] = ~layer1_out[3134];
    assign layer2_out[4147] = ~layer1_out[6928] | layer1_out[6927];
    assign layer2_out[4148] = layer1_out[1049] & layer1_out[1050];
    assign layer2_out[4149] = ~layer1_out[7303];
    assign layer2_out[4150] = layer1_out[1072] & ~layer1_out[1071];
    assign layer2_out[4151] = 1'b1;
    assign layer2_out[4152] = ~layer1_out[5614];
    assign layer2_out[4153] = ~layer1_out[1678] | layer1_out[1679];
    assign layer2_out[4154] = layer1_out[4268];
    assign layer2_out[4155] = layer1_out[2315] | layer1_out[2316];
    assign layer2_out[4156] = ~layer1_out[562];
    assign layer2_out[4157] = ~layer1_out[3452];
    assign layer2_out[4158] = ~(layer1_out[5817] ^ layer1_out[5818]);
    assign layer2_out[4159] = ~layer1_out[1280];
    assign layer2_out[4160] = ~(layer1_out[6136] | layer1_out[6137]);
    assign layer2_out[4161] = layer1_out[327];
    assign layer2_out[4162] = ~layer1_out[5302];
    assign layer2_out[4163] = ~layer1_out[3825] | layer1_out[3824];
    assign layer2_out[4164] = ~layer1_out[1624];
    assign layer2_out[4165] = layer1_out[1919] & ~layer1_out[1918];
    assign layer2_out[4166] = layer1_out[6931] & ~layer1_out[6930];
    assign layer2_out[4167] = layer1_out[3193] ^ layer1_out[3194];
    assign layer2_out[4168] = ~(layer1_out[3039] | layer1_out[3040]);
    assign layer2_out[4169] = layer1_out[3502] & layer1_out[3503];
    assign layer2_out[4170] = ~layer1_out[6845];
    assign layer2_out[4171] = layer1_out[4790] & layer1_out[4791];
    assign layer2_out[4172] = layer1_out[7425] | layer1_out[7426];
    assign layer2_out[4173] = ~layer1_out[2551];
    assign layer2_out[4174] = ~layer1_out[745] | layer1_out[744];
    assign layer2_out[4175] = ~(layer1_out[7911] ^ layer1_out[7912]);
    assign layer2_out[4176] = 1'b0;
    assign layer2_out[4177] = ~layer1_out[2317];
    assign layer2_out[4178] = layer1_out[7223] ^ layer1_out[7224];
    assign layer2_out[4179] = layer1_out[6861];
    assign layer2_out[4180] = ~(layer1_out[5440] & layer1_out[5441]);
    assign layer2_out[4181] = layer1_out[6739] & ~layer1_out[6740];
    assign layer2_out[4182] = layer1_out[5825] & layer1_out[5826];
    assign layer2_out[4183] = ~layer1_out[503];
    assign layer2_out[4184] = layer1_out[1505] & ~layer1_out[1504];
    assign layer2_out[4185] = ~layer1_out[5755];
    assign layer2_out[4186] = ~(layer1_out[3337] | layer1_out[3338]);
    assign layer2_out[4187] = ~(layer1_out[7350] | layer1_out[7351]);
    assign layer2_out[4188] = layer1_out[3717];
    assign layer2_out[4189] = layer1_out[4241];
    assign layer2_out[4190] = ~layer1_out[609] | layer1_out[610];
    assign layer2_out[4191] = layer1_out[6015];
    assign layer2_out[4192] = ~(layer1_out[4947] ^ layer1_out[4948]);
    assign layer2_out[4193] = layer1_out[2554];
    assign layer2_out[4194] = ~layer1_out[220] | layer1_out[219];
    assign layer2_out[4195] = ~layer1_out[4074];
    assign layer2_out[4196] = layer1_out[4311] | layer1_out[4312];
    assign layer2_out[4197] = layer1_out[2908];
    assign layer2_out[4198] = layer1_out[2559];
    assign layer2_out[4199] = layer1_out[2766];
    assign layer2_out[4200] = layer1_out[6443] & layer1_out[6444];
    assign layer2_out[4201] = layer1_out[6026] & ~layer1_out[6025];
    assign layer2_out[4202] = layer1_out[3030] & ~layer1_out[3029];
    assign layer2_out[4203] = layer1_out[292] | layer1_out[293];
    assign layer2_out[4204] = layer1_out[6735];
    assign layer2_out[4205] = ~layer1_out[4620] | layer1_out[4621];
    assign layer2_out[4206] = layer1_out[2418] & ~layer1_out[2419];
    assign layer2_out[4207] = ~layer1_out[7915] | layer1_out[7914];
    assign layer2_out[4208] = ~(layer1_out[2075] | layer1_out[2076]);
    assign layer2_out[4209] = ~(layer1_out[6430] | layer1_out[6431]);
    assign layer2_out[4210] = layer1_out[3586];
    assign layer2_out[4211] = 1'b0;
    assign layer2_out[4212] = layer1_out[4955];
    assign layer2_out[4213] = ~layer1_out[5973] | layer1_out[5974];
    assign layer2_out[4214] = layer1_out[4160];
    assign layer2_out[4215] = layer1_out[6728];
    assign layer2_out[4216] = ~layer1_out[5502];
    assign layer2_out[4217] = ~(layer1_out[61] & layer1_out[62]);
    assign layer2_out[4218] = ~(layer1_out[849] & layer1_out[850]);
    assign layer2_out[4219] = layer1_out[7] & ~layer1_out[8];
    assign layer2_out[4220] = layer1_out[7918] | layer1_out[7919];
    assign layer2_out[4221] = ~layer1_out[240];
    assign layer2_out[4222] = layer1_out[10];
    assign layer2_out[4223] = ~layer1_out[3958] | layer1_out[3959];
    assign layer2_out[4224] = layer1_out[97] | layer1_out[98];
    assign layer2_out[4225] = ~layer1_out[7651];
    assign layer2_out[4226] = layer1_out[6530];
    assign layer2_out[4227] = ~layer1_out[5649] | layer1_out[5648];
    assign layer2_out[4228] = layer1_out[2574] & ~layer1_out[2573];
    assign layer2_out[4229] = layer1_out[4092];
    assign layer2_out[4230] = ~layer1_out[199] | layer1_out[200];
    assign layer2_out[4231] = ~layer1_out[6207] | layer1_out[6208];
    assign layer2_out[4232] = ~(layer1_out[3168] | layer1_out[3169]);
    assign layer2_out[4233] = ~layer1_out[6511];
    assign layer2_out[4234] = layer1_out[4680] & layer1_out[4681];
    assign layer2_out[4235] = ~layer1_out[4725] | layer1_out[4724];
    assign layer2_out[4236] = ~(layer1_out[84] | layer1_out[85]);
    assign layer2_out[4237] = ~layer1_out[6108] | layer1_out[6109];
    assign layer2_out[4238] = layer1_out[1216];
    assign layer2_out[4239] = ~layer1_out[945];
    assign layer2_out[4240] = layer1_out[6975] | layer1_out[6976];
    assign layer2_out[4241] = ~(layer1_out[2604] ^ layer1_out[2605]);
    assign layer2_out[4242] = layer1_out[4709] & ~layer1_out[4710];
    assign layer2_out[4243] = ~layer1_out[4285];
    assign layer2_out[4244] = ~layer1_out[3383];
    assign layer2_out[4245] = layer1_out[5500] ^ layer1_out[5501];
    assign layer2_out[4246] = layer1_out[3241];
    assign layer2_out[4247] = ~layer1_out[1989];
    assign layer2_out[4248] = ~layer1_out[194] | layer1_out[193];
    assign layer2_out[4249] = layer1_out[1129] | layer1_out[1130];
    assign layer2_out[4250] = layer1_out[4888];
    assign layer2_out[4251] = ~layer1_out[54];
    assign layer2_out[4252] = ~layer1_out[3973];
    assign layer2_out[4253] = ~layer1_out[5892];
    assign layer2_out[4254] = ~layer1_out[2356] | layer1_out[2357];
    assign layer2_out[4255] = layer1_out[3839];
    assign layer2_out[4256] = layer1_out[2129] & ~layer1_out[2128];
    assign layer2_out[4257] = layer1_out[2419];
    assign layer2_out[4258] = layer1_out[185];
    assign layer2_out[4259] = layer1_out[6710];
    assign layer2_out[4260] = layer1_out[2935];
    assign layer2_out[4261] = layer1_out[2125] & layer1_out[2126];
    assign layer2_out[4262] = layer1_out[5372];
    assign layer2_out[4263] = ~layer1_out[7873];
    assign layer2_out[4264] = layer1_out[4552] & layer1_out[4553];
    assign layer2_out[4265] = ~layer1_out[1380];
    assign layer2_out[4266] = layer1_out[573] ^ layer1_out[574];
    assign layer2_out[4267] = ~layer1_out[7050];
    assign layer2_out[4268] = ~(layer1_out[2042] | layer1_out[2043]);
    assign layer2_out[4269] = ~layer1_out[600];
    assign layer2_out[4270] = layer1_out[2003] | layer1_out[2004];
    assign layer2_out[4271] = ~layer1_out[6805];
    assign layer2_out[4272] = layer1_out[4173] & ~layer1_out[4174];
    assign layer2_out[4273] = 1'b1;
    assign layer2_out[4274] = layer1_out[5901];
    assign layer2_out[4275] = layer1_out[2873] & ~layer1_out[2872];
    assign layer2_out[4276] = layer1_out[6924];
    assign layer2_out[4277] = ~layer1_out[3569];
    assign layer2_out[4278] = ~layer1_out[6901];
    assign layer2_out[4279] = layer1_out[1745] & ~layer1_out[1746];
    assign layer2_out[4280] = 1'b1;
    assign layer2_out[4281] = ~layer1_out[6234];
    assign layer2_out[4282] = layer1_out[2071];
    assign layer2_out[4283] = ~(layer1_out[3012] | layer1_out[3013]);
    assign layer2_out[4284] = layer1_out[1685] | layer1_out[1686];
    assign layer2_out[4285] = layer1_out[1596];
    assign layer2_out[4286] = layer1_out[5379] | layer1_out[5380];
    assign layer2_out[4287] = layer1_out[25] & layer1_out[26];
    assign layer2_out[4288] = ~(layer1_out[382] ^ layer1_out[383]);
    assign layer2_out[4289] = layer1_out[1642];
    assign layer2_out[4290] = layer1_out[4399] | layer1_out[4400];
    assign layer2_out[4291] = layer1_out[6195];
    assign layer2_out[4292] = ~layer1_out[5798] | layer1_out[5799];
    assign layer2_out[4293] = ~layer1_out[2412];
    assign layer2_out[4294] = layer1_out[5197];
    assign layer2_out[4295] = ~layer1_out[2603] | layer1_out[2604];
    assign layer2_out[4296] = layer1_out[1422];
    assign layer2_out[4297] = ~layer1_out[7831] | layer1_out[7830];
    assign layer2_out[4298] = layer1_out[451] ^ layer1_out[452];
    assign layer2_out[4299] = layer1_out[448] & layer1_out[449];
    assign layer2_out[4300] = ~(layer1_out[4393] ^ layer1_out[4394]);
    assign layer2_out[4301] = ~layer1_out[7537];
    assign layer2_out[4302] = layer1_out[3128] & ~layer1_out[3127];
    assign layer2_out[4303] = ~(layer1_out[1580] ^ layer1_out[1581]);
    assign layer2_out[4304] = layer1_out[2794];
    assign layer2_out[4305] = ~layer1_out[5796];
    assign layer2_out[4306] = ~(layer1_out[4133] | layer1_out[4134]);
    assign layer2_out[4307] = layer1_out[5492] & layer1_out[5493];
    assign layer2_out[4308] = ~layer1_out[992] | layer1_out[993];
    assign layer2_out[4309] = layer1_out[4459];
    assign layer2_out[4310] = ~layer1_out[7718];
    assign layer2_out[4311] = layer1_out[6391];
    assign layer2_out[4312] = ~layer1_out[3183];
    assign layer2_out[4313] = ~layer1_out[4466];
    assign layer2_out[4314] = layer1_out[2476] & ~layer1_out[2477];
    assign layer2_out[4315] = layer1_out[1108];
    assign layer2_out[4316] = 1'b1;
    assign layer2_out[4317] = layer1_out[6306];
    assign layer2_out[4318] = ~(layer1_out[1199] & layer1_out[1200]);
    assign layer2_out[4319] = layer1_out[4616];
    assign layer2_out[4320] = 1'b1;
    assign layer2_out[4321] = layer1_out[5142] & layer1_out[5143];
    assign layer2_out[4322] = layer1_out[2484] & ~layer1_out[2485];
    assign layer2_out[4323] = layer1_out[7046] & ~layer1_out[7045];
    assign layer2_out[4324] = ~layer1_out[183];
    assign layer2_out[4325] = ~layer1_out[1081] | layer1_out[1080];
    assign layer2_out[4326] = ~layer1_out[715];
    assign layer2_out[4327] = ~layer1_out[731] | layer1_out[730];
    assign layer2_out[4328] = layer1_out[6925] & layer1_out[6926];
    assign layer2_out[4329] = ~layer1_out[5317] | layer1_out[5318];
    assign layer2_out[4330] = ~layer1_out[7406] | layer1_out[7405];
    assign layer2_out[4331] = layer1_out[4081];
    assign layer2_out[4332] = ~layer1_out[7740];
    assign layer2_out[4333] = layer1_out[959];
    assign layer2_out[4334] = layer1_out[4411] & ~layer1_out[4410];
    assign layer2_out[4335] = ~(layer1_out[6052] & layer1_out[6053]);
    assign layer2_out[4336] = layer1_out[2883] & ~layer1_out[2884];
    assign layer2_out[4337] = ~layer1_out[7218] | layer1_out[7217];
    assign layer2_out[4338] = ~(layer1_out[1024] & layer1_out[1025]);
    assign layer2_out[4339] = layer1_out[5946];
    assign layer2_out[4340] = layer1_out[4351] | layer1_out[4352];
    assign layer2_out[4341] = ~layer1_out[2666];
    assign layer2_out[4342] = layer1_out[7631];
    assign layer2_out[4343] = layer1_out[1176];
    assign layer2_out[4344] = layer1_out[2272] | layer1_out[2273];
    assign layer2_out[4345] = ~(layer1_out[1828] ^ layer1_out[1829]);
    assign layer2_out[4346] = ~layer1_out[7003] | layer1_out[7002];
    assign layer2_out[4347] = ~layer1_out[3635];
    assign layer2_out[4348] = ~layer1_out[420];
    assign layer2_out[4349] = layer1_out[1408];
    assign layer2_out[4350] = ~layer1_out[5602] | layer1_out[5603];
    assign layer2_out[4351] = layer1_out[7022];
    assign layer2_out[4352] = ~layer1_out[2987];
    assign layer2_out[4353] = ~layer1_out[4922];
    assign layer2_out[4354] = layer1_out[2684] & layer1_out[2685];
    assign layer2_out[4355] = ~layer1_out[7573];
    assign layer2_out[4356] = layer1_out[7226] & ~layer1_out[7225];
    assign layer2_out[4357] = ~layer1_out[6351] | layer1_out[6350];
    assign layer2_out[4358] = ~layer1_out[2180] | layer1_out[2181];
    assign layer2_out[4359] = ~layer1_out[3199];
    assign layer2_out[4360] = ~layer1_out[7438] | layer1_out[7437];
    assign layer2_out[4361] = layer1_out[3391] & ~layer1_out[3390];
    assign layer2_out[4362] = ~layer1_out[5646];
    assign layer2_out[4363] = ~(layer1_out[113] | layer1_out[114]);
    assign layer2_out[4364] = layer1_out[7908] & ~layer1_out[7907];
    assign layer2_out[4365] = ~(layer1_out[5668] & layer1_out[5669]);
    assign layer2_out[4366] = ~layer1_out[6477] | layer1_out[6478];
    assign layer2_out[4367] = layer1_out[1603] & ~layer1_out[1602];
    assign layer2_out[4368] = ~(layer1_out[7960] | layer1_out[7961]);
    assign layer2_out[4369] = 1'b0;
    assign layer2_out[4370] = ~layer1_out[2524] | layer1_out[2525];
    assign layer2_out[4371] = layer1_out[1917];
    assign layer2_out[4372] = layer1_out[695];
    assign layer2_out[4373] = layer1_out[5266] | layer1_out[5267];
    assign layer2_out[4374] = layer1_out[1851];
    assign layer2_out[4375] = ~(layer1_out[6096] | layer1_out[6097]);
    assign layer2_out[4376] = ~layer1_out[7798];
    assign layer2_out[4377] = layer1_out[7144];
    assign layer2_out[4378] = ~layer1_out[2013] | layer1_out[2012];
    assign layer2_out[4379] = layer1_out[4145];
    assign layer2_out[4380] = layer1_out[5035];
    assign layer2_out[4381] = layer1_out[5666] & ~layer1_out[5665];
    assign layer2_out[4382] = layer1_out[2486] & ~layer1_out[2485];
    assign layer2_out[4383] = layer1_out[2597];
    assign layer2_out[4384] = layer1_out[2876] | layer1_out[2877];
    assign layer2_out[4385] = ~(layer1_out[5093] ^ layer1_out[5094]);
    assign layer2_out[4386] = layer1_out[2546] & ~layer1_out[2545];
    assign layer2_out[4387] = ~layer1_out[6692];
    assign layer2_out[4388] = ~(layer1_out[1360] ^ layer1_out[1361]);
    assign layer2_out[4389] = layer1_out[3070] & layer1_out[3071];
    assign layer2_out[4390] = ~layer1_out[5728];
    assign layer2_out[4391] = ~layer1_out[4456] | layer1_out[4455];
    assign layer2_out[4392] = 1'b0;
    assign layer2_out[4393] = ~layer1_out[3939];
    assign layer2_out[4394] = ~layer1_out[4512] | layer1_out[4513];
    assign layer2_out[4395] = layer1_out[3409];
    assign layer2_out[4396] = ~layer1_out[1097];
    assign layer2_out[4397] = layer1_out[5375];
    assign layer2_out[4398] = ~(layer1_out[7817] | layer1_out[7818]);
    assign layer2_out[4399] = ~layer1_out[3000];
    assign layer2_out[4400] = ~layer1_out[2390];
    assign layer2_out[4401] = layer1_out[2407] & ~layer1_out[2408];
    assign layer2_out[4402] = layer1_out[6477];
    assign layer2_out[4403] = ~(layer1_out[6685] ^ layer1_out[6686]);
    assign layer2_out[4404] = ~layer1_out[807];
    assign layer2_out[4405] = layer1_out[6642] & ~layer1_out[6643];
    assign layer2_out[4406] = ~layer1_out[1878];
    assign layer2_out[4407] = ~layer1_out[3122];
    assign layer2_out[4408] = layer1_out[1175];
    assign layer2_out[4409] = ~layer1_out[6389];
    assign layer2_out[4410] = ~layer1_out[2761];
    assign layer2_out[4411] = ~layer1_out[5172];
    assign layer2_out[4412] = layer1_out[5505] & ~layer1_out[5506];
    assign layer2_out[4413] = ~layer1_out[2252];
    assign layer2_out[4414] = layer1_out[1513];
    assign layer2_out[4415] = ~(layer1_out[3321] | layer1_out[3322]);
    assign layer2_out[4416] = ~layer1_out[1826] | layer1_out[1825];
    assign layer2_out[4417] = ~(layer1_out[5075] & layer1_out[5076]);
    assign layer2_out[4418] = 1'b1;
    assign layer2_out[4419] = ~layer1_out[1966] | layer1_out[1967];
    assign layer2_out[4420] = ~(layer1_out[4997] ^ layer1_out[4998]);
    assign layer2_out[4421] = 1'b0;
    assign layer2_out[4422] = ~layer1_out[2841];
    assign layer2_out[4423] = ~(layer1_out[621] & layer1_out[622]);
    assign layer2_out[4424] = ~layer1_out[3338] | layer1_out[3339];
    assign layer2_out[4425] = ~(layer1_out[5667] & layer1_out[5668]);
    assign layer2_out[4426] = ~layer1_out[750];
    assign layer2_out[4427] = layer1_out[3552] | layer1_out[3553];
    assign layer2_out[4428] = layer1_out[413] ^ layer1_out[414];
    assign layer2_out[4429] = layer1_out[1093];
    assign layer2_out[4430] = 1'b0;
    assign layer2_out[4431] = ~layer1_out[5551];
    assign layer2_out[4432] = layer1_out[2654] & ~layer1_out[2653];
    assign layer2_out[4433] = layer1_out[839] ^ layer1_out[840];
    assign layer2_out[4434] = ~layer1_out[4485] | layer1_out[4484];
    assign layer2_out[4435] = ~layer1_out[6463];
    assign layer2_out[4436] = ~layer1_out[4920];
    assign layer2_out[4437] = ~(layer1_out[6358] | layer1_out[6359]);
    assign layer2_out[4438] = ~(layer1_out[2] | layer1_out[3]);
    assign layer2_out[4439] = layer1_out[1242] & ~layer1_out[1243];
    assign layer2_out[4440] = layer1_out[2506] & layer1_out[2507];
    assign layer2_out[4441] = layer1_out[792];
    assign layer2_out[4442] = ~layer1_out[6691];
    assign layer2_out[4443] = ~layer1_out[1615];
    assign layer2_out[4444] = layer1_out[1274];
    assign layer2_out[4445] = ~layer1_out[6544];
    assign layer2_out[4446] = ~layer1_out[2444];
    assign layer2_out[4447] = layer1_out[6324] & ~layer1_out[6323];
    assign layer2_out[4448] = layer1_out[6174];
    assign layer2_out[4449] = layer1_out[6709] & layer1_out[6710];
    assign layer2_out[4450] = ~layer1_out[906];
    assign layer2_out[4451] = layer1_out[2708] | layer1_out[2709];
    assign layer2_out[4452] = ~(layer1_out[1347] | layer1_out[1348]);
    assign layer2_out[4453] = ~(layer1_out[2278] & layer1_out[2279]);
    assign layer2_out[4454] = ~layer1_out[513];
    assign layer2_out[4455] = ~(layer1_out[4022] | layer1_out[4023]);
    assign layer2_out[4456] = ~layer1_out[4356];
    assign layer2_out[4457] = layer1_out[6976] ^ layer1_out[6977];
    assign layer2_out[4458] = layer1_out[6079] & layer1_out[6080];
    assign layer2_out[4459] = ~layer1_out[7446];
    assign layer2_out[4460] = layer1_out[7307];
    assign layer2_out[4461] = ~layer1_out[4809] | layer1_out[4808];
    assign layer2_out[4462] = layer1_out[7931] | layer1_out[7932];
    assign layer2_out[4463] = layer1_out[7276] & ~layer1_out[7275];
    assign layer2_out[4464] = layer1_out[3783] | layer1_out[3784];
    assign layer2_out[4465] = layer1_out[5890];
    assign layer2_out[4466] = layer1_out[65];
    assign layer2_out[4467] = layer1_out[840] ^ layer1_out[841];
    assign layer2_out[4468] = ~layer1_out[6484] | layer1_out[6483];
    assign layer2_out[4469] = ~(layer1_out[3294] ^ layer1_out[3295]);
    assign layer2_out[4470] = ~layer1_out[1113] | layer1_out[1114];
    assign layer2_out[4471] = layer1_out[5961] | layer1_out[5962];
    assign layer2_out[4472] = layer1_out[3334] & layer1_out[3335];
    assign layer2_out[4473] = ~layer1_out[7039];
    assign layer2_out[4474] = layer1_out[2099] | layer1_out[2100];
    assign layer2_out[4475] = ~layer1_out[2712];
    assign layer2_out[4476] = layer1_out[5967] | layer1_out[5968];
    assign layer2_out[4477] = ~(layer1_out[4683] ^ layer1_out[4684]);
    assign layer2_out[4478] = ~layer1_out[5627] | layer1_out[5626];
    assign layer2_out[4479] = ~layer1_out[1197] | layer1_out[1196];
    assign layer2_out[4480] = layer1_out[7305] | layer1_out[7306];
    assign layer2_out[4481] = ~layer1_out[4113] | layer1_out[4112];
    assign layer2_out[4482] = ~(layer1_out[3322] & layer1_out[3323]);
    assign layer2_out[4483] = ~layer1_out[7250];
    assign layer2_out[4484] = ~layer1_out[1743] | layer1_out[1742];
    assign layer2_out[4485] = layer1_out[240];
    assign layer2_out[4486] = layer1_out[6077] | layer1_out[6078];
    assign layer2_out[4487] = ~layer1_out[4755] | layer1_out[4754];
    assign layer2_out[4488] = layer1_out[3851];
    assign layer2_out[4489] = ~layer1_out[7183] | layer1_out[7182];
    assign layer2_out[4490] = layer1_out[6933] & layer1_out[6934];
    assign layer2_out[4491] = layer1_out[2781];
    assign layer2_out[4492] = ~layer1_out[4031] | layer1_out[4030];
    assign layer2_out[4493] = ~layer1_out[3237] | layer1_out[3236];
    assign layer2_out[4494] = 1'b0;
    assign layer2_out[4495] = ~(layer1_out[1266] & layer1_out[1267]);
    assign layer2_out[4496] = layer1_out[434] ^ layer1_out[435];
    assign layer2_out[4497] = ~layer1_out[1048] | layer1_out[1049];
    assign layer2_out[4498] = layer1_out[3436];
    assign layer2_out[4499] = ~layer1_out[5638];
    assign layer2_out[4500] = layer1_out[2327] & ~layer1_out[2326];
    assign layer2_out[4501] = ~layer1_out[4706];
    assign layer2_out[4502] = layer1_out[6571] & ~layer1_out[6570];
    assign layer2_out[4503] = layer1_out[751] & ~layer1_out[752];
    assign layer2_out[4504] = layer1_out[2993] | layer1_out[2994];
    assign layer2_out[4505] = layer1_out[5326] ^ layer1_out[5327];
    assign layer2_out[4506] = ~(layer1_out[6262] & layer1_out[6263]);
    assign layer2_out[4507] = ~(layer1_out[742] | layer1_out[743]);
    assign layer2_out[4508] = ~(layer1_out[5790] & layer1_out[5791]);
    assign layer2_out[4509] = layer1_out[2867];
    assign layer2_out[4510] = layer1_out[6648];
    assign layer2_out[4511] = layer1_out[4750];
    assign layer2_out[4512] = ~layer1_out[1657];
    assign layer2_out[4513] = layer1_out[4975];
    assign layer2_out[4514] = ~layer1_out[5141] | layer1_out[5140];
    assign layer2_out[4515] = ~layer1_out[7015];
    assign layer2_out[4516] = layer1_out[1050];
    assign layer2_out[4517] = layer1_out[526];
    assign layer2_out[4518] = layer1_out[1118];
    assign layer2_out[4519] = ~(layer1_out[2497] & layer1_out[2498]);
    assign layer2_out[4520] = layer1_out[1841] & layer1_out[1842];
    assign layer2_out[4521] = layer1_out[6129];
    assign layer2_out[4522] = ~layer1_out[6262];
    assign layer2_out[4523] = layer1_out[3366];
    assign layer2_out[4524] = ~(layer1_out[2186] | layer1_out[2187]);
    assign layer2_out[4525] = layer1_out[6011];
    assign layer2_out[4526] = ~layer1_out[5672] | layer1_out[5673];
    assign layer2_out[4527] = layer1_out[1776] & layer1_out[1777];
    assign layer2_out[4528] = ~(layer1_out[6118] ^ layer1_out[6119]);
    assign layer2_out[4529] = layer1_out[4409] | layer1_out[4410];
    assign layer2_out[4530] = layer1_out[3882];
    assign layer2_out[4531] = layer1_out[6490] | layer1_out[6491];
    assign layer2_out[4532] = layer1_out[3947];
    assign layer2_out[4533] = layer1_out[1375] | layer1_out[1376];
    assign layer2_out[4534] = ~layer1_out[5950];
    assign layer2_out[4535] = ~(layer1_out[5834] & layer1_out[5835]);
    assign layer2_out[4536] = ~(layer1_out[3513] ^ layer1_out[3514]);
    assign layer2_out[4537] = ~(layer1_out[2334] | layer1_out[2335]);
    assign layer2_out[4538] = 1'b0;
    assign layer2_out[4539] = layer1_out[5635] | layer1_out[5636];
    assign layer2_out[4540] = ~layer1_out[6957] | layer1_out[6958];
    assign layer2_out[4541] = layer1_out[4797];
    assign layer2_out[4542] = layer1_out[1901] & ~layer1_out[1900];
    assign layer2_out[4543] = layer1_out[1005];
    assign layer2_out[4544] = ~layer1_out[4013] | layer1_out[4012];
    assign layer2_out[4545] = ~(layer1_out[4094] & layer1_out[4095]);
    assign layer2_out[4546] = ~(layer1_out[4733] ^ layer1_out[4734]);
    assign layer2_out[4547] = ~(layer1_out[7238] & layer1_out[7239]);
    assign layer2_out[4548] = 1'b0;
    assign layer2_out[4549] = ~(layer1_out[7803] | layer1_out[7804]);
    assign layer2_out[4550] = ~layer1_out[2271];
    assign layer2_out[4551] = ~layer1_out[4253];
    assign layer2_out[4552] = layer1_out[3459] ^ layer1_out[3460];
    assign layer2_out[4553] = ~layer1_out[4509] | layer1_out[4508];
    assign layer2_out[4554] = layer1_out[6769] & ~layer1_out[6768];
    assign layer2_out[4555] = layer1_out[706] & layer1_out[707];
    assign layer2_out[4556] = ~layer1_out[4415];
    assign layer2_out[4557] = ~layer1_out[6897] | layer1_out[6898];
    assign layer2_out[4558] = ~(layer1_out[4317] | layer1_out[4318]);
    assign layer2_out[4559] = layer1_out[6839];
    assign layer2_out[4560] = ~(layer1_out[4071] | layer1_out[4072]);
    assign layer2_out[4561] = ~layer1_out[5643];
    assign layer2_out[4562] = layer1_out[3971] & layer1_out[3972];
    assign layer2_out[4563] = 1'b0;
    assign layer2_out[4564] = layer1_out[1914];
    assign layer2_out[4565] = layer1_out[1340];
    assign layer2_out[4566] = layer1_out[7604] ^ layer1_out[7605];
    assign layer2_out[4567] = layer1_out[1667];
    assign layer2_out[4568] = layer1_out[6086];
    assign layer2_out[4569] = ~(layer1_out[6592] | layer1_out[6593]);
    assign layer2_out[4570] = ~layer1_out[4147] | layer1_out[4146];
    assign layer2_out[4571] = layer1_out[7059] & ~layer1_out[7060];
    assign layer2_out[4572] = ~layer1_out[2046];
    assign layer2_out[4573] = ~(layer1_out[4268] & layer1_out[4269]);
    assign layer2_out[4574] = layer1_out[4198] & ~layer1_out[4199];
    assign layer2_out[4575] = ~layer1_out[457] | layer1_out[456];
    assign layer2_out[4576] = layer1_out[3218] | layer1_out[3219];
    assign layer2_out[4577] = layer1_out[5600];
    assign layer2_out[4578] = layer1_out[1409] & layer1_out[1410];
    assign layer2_out[4579] = ~layer1_out[6435];
    assign layer2_out[4580] = ~(layer1_out[1168] & layer1_out[1169]);
    assign layer2_out[4581] = ~layer1_out[4973];
    assign layer2_out[4582] = 1'b1;
    assign layer2_out[4583] = layer1_out[3587] & ~layer1_out[3588];
    assign layer2_out[4584] = ~(layer1_out[3026] & layer1_out[3027]);
    assign layer2_out[4585] = layer1_out[1483] ^ layer1_out[1484];
    assign layer2_out[4586] = layer1_out[4500] & ~layer1_out[4501];
    assign layer2_out[4587] = layer1_out[693] & ~layer1_out[694];
    assign layer2_out[4588] = layer1_out[1687] & layer1_out[1688];
    assign layer2_out[4589] = layer1_out[6748] & ~layer1_out[6749];
    assign layer2_out[4590] = ~layer1_out[4469] | layer1_out[4468];
    assign layer2_out[4591] = ~layer1_out[44];
    assign layer2_out[4592] = layer1_out[7898] ^ layer1_out[7899];
    assign layer2_out[4593] = ~layer1_out[2928] | layer1_out[2929];
    assign layer2_out[4594] = ~layer1_out[4940];
    assign layer2_out[4595] = layer1_out[4370] ^ layer1_out[4371];
    assign layer2_out[4596] = ~(layer1_out[6997] & layer1_out[6998]);
    assign layer2_out[4597] = layer1_out[1040];
    assign layer2_out[4598] = ~layer1_out[2052] | layer1_out[2051];
    assign layer2_out[4599] = ~(layer1_out[6266] ^ layer1_out[6267]);
    assign layer2_out[4600] = layer1_out[3017];
    assign layer2_out[4601] = layer1_out[142] & layer1_out[143];
    assign layer2_out[4602] = 1'b1;
    assign layer2_out[4603] = layer1_out[5338] & layer1_out[5339];
    assign layer2_out[4604] = ~layer1_out[6411];
    assign layer2_out[4605] = ~(layer1_out[3937] ^ layer1_out[3938]);
    assign layer2_out[4606] = layer1_out[6832] | layer1_out[6833];
    assign layer2_out[4607] = layer1_out[226] | layer1_out[227];
    assign layer2_out[4608] = ~layer1_out[6944];
    assign layer2_out[4609] = layer1_out[7952];
    assign layer2_out[4610] = layer1_out[4584];
    assign layer2_out[4611] = layer1_out[1862];
    assign layer2_out[4612] = ~(layer1_out[642] & layer1_out[643]);
    assign layer2_out[4613] = layer1_out[4774] & layer1_out[4775];
    assign layer2_out[4614] = 1'b1;
    assign layer2_out[4615] = ~(layer1_out[3642] & layer1_out[3643]);
    assign layer2_out[4616] = ~layer1_out[7145];
    assign layer2_out[4617] = ~(layer1_out[5404] | layer1_out[5405]);
    assign layer2_out[4618] = ~(layer1_out[2250] & layer1_out[2251]);
    assign layer2_out[4619] = layer1_out[4968] & ~layer1_out[4969];
    assign layer2_out[4620] = 1'b1;
    assign layer2_out[4621] = ~layer1_out[7153];
    assign layer2_out[4622] = layer1_out[3790];
    assign layer2_out[4623] = ~layer1_out[3858];
    assign layer2_out[4624] = layer1_out[3185] & ~layer1_out[3186];
    assign layer2_out[4625] = ~layer1_out[2689];
    assign layer2_out[4626] = ~layer1_out[7009] | layer1_out[7010];
    assign layer2_out[4627] = layer1_out[3504] & ~layer1_out[3503];
    assign layer2_out[4628] = ~layer1_out[7918] | layer1_out[7917];
    assign layer2_out[4629] = ~(layer1_out[1332] & layer1_out[1333]);
    assign layer2_out[4630] = layer1_out[5348];
    assign layer2_out[4631] = ~layer1_out[1002];
    assign layer2_out[4632] = ~layer1_out[2076];
    assign layer2_out[4633] = layer1_out[1236];
    assign layer2_out[4634] = ~(layer1_out[5910] | layer1_out[5911]);
    assign layer2_out[4635] = layer1_out[2276] ^ layer1_out[2277];
    assign layer2_out[4636] = layer1_out[6082] | layer1_out[6083];
    assign layer2_out[4637] = layer1_out[6597];
    assign layer2_out[4638] = ~(layer1_out[5154] | layer1_out[5155]);
    assign layer2_out[4639] = layer1_out[1134];
    assign layer2_out[4640] = layer1_out[5242] & ~layer1_out[5241];
    assign layer2_out[4641] = layer1_out[4462];
    assign layer2_out[4642] = ~(layer1_out[2213] | layer1_out[2214]);
    assign layer2_out[4643] = ~layer1_out[3814];
    assign layer2_out[4644] = layer1_out[7813];
    assign layer2_out[4645] = layer1_out[7284];
    assign layer2_out[4646] = ~(layer1_out[1666] ^ layer1_out[1667]);
    assign layer2_out[4647] = 1'b0;
    assign layer2_out[4648] = layer1_out[5871];
    assign layer2_out[4649] = layer1_out[2904] & layer1_out[2905];
    assign layer2_out[4650] = layer1_out[3691] & ~layer1_out[3692];
    assign layer2_out[4651] = ~(layer1_out[825] ^ layer1_out[826]);
    assign layer2_out[4652] = layer1_out[887];
    assign layer2_out[4653] = 1'b1;
    assign layer2_out[4654] = layer1_out[5709] & ~layer1_out[5708];
    assign layer2_out[4655] = layer1_out[616] | layer1_out[617];
    assign layer2_out[4656] = ~(layer1_out[3828] | layer1_out[3829]);
    assign layer2_out[4657] = ~(layer1_out[5649] ^ layer1_out[5650]);
    assign layer2_out[4658] = ~layer1_out[4848] | layer1_out[4849];
    assign layer2_out[4659] = layer1_out[1929] ^ layer1_out[1930];
    assign layer2_out[4660] = layer1_out[3160];
    assign layer2_out[4661] = layer1_out[5095] & ~layer1_out[5094];
    assign layer2_out[4662] = ~layer1_out[4557];
    assign layer2_out[4663] = ~(layer1_out[4828] & layer1_out[4829]);
    assign layer2_out[4664] = ~layer1_out[7114];
    assign layer2_out[4665] = ~layer1_out[2504] | layer1_out[2503];
    assign layer2_out[4666] = layer1_out[2766];
    assign layer2_out[4667] = layer1_out[4383];
    assign layer2_out[4668] = ~layer1_out[1227];
    assign layer2_out[4669] = 1'b1;
    assign layer2_out[4670] = ~layer1_out[847];
    assign layer2_out[4671] = layer1_out[2135] ^ layer1_out[2136];
    assign layer2_out[4672] = ~(layer1_out[856] ^ layer1_out[857]);
    assign layer2_out[4673] = layer1_out[2611] | layer1_out[2612];
    assign layer2_out[4674] = ~(layer1_out[6979] | layer1_out[6980]);
    assign layer2_out[4675] = layer1_out[4147];
    assign layer2_out[4676] = ~(layer1_out[7441] & layer1_out[7442]);
    assign layer2_out[4677] = ~(layer1_out[3632] ^ layer1_out[3633]);
    assign layer2_out[4678] = layer1_out[5000] & layer1_out[5001];
    assign layer2_out[4679] = layer1_out[290];
    assign layer2_out[4680] = ~layer1_out[426];
    assign layer2_out[4681] = ~layer1_out[4752];
    assign layer2_out[4682] = 1'b1;
    assign layer2_out[4683] = layer1_out[2032];
    assign layer2_out[4684] = layer1_out[366];
    assign layer2_out[4685] = ~layer1_out[7482];
    assign layer2_out[4686] = layer1_out[3655] & layer1_out[3656];
    assign layer2_out[4687] = layer1_out[703];
    assign layer2_out[4688] = layer1_out[7856] & ~layer1_out[7855];
    assign layer2_out[4689] = ~(layer1_out[4592] & layer1_out[4593]);
    assign layer2_out[4690] = ~layer1_out[2857] | layer1_out[2856];
    assign layer2_out[4691] = ~(layer1_out[583] | layer1_out[584]);
    assign layer2_out[4692] = layer1_out[4836] & ~layer1_out[4835];
    assign layer2_out[4693] = ~layer1_out[1553];
    assign layer2_out[4694] = layer1_out[3640] & ~layer1_out[3641];
    assign layer2_out[4695] = ~(layer1_out[7315] & layer1_out[7316]);
    assign layer2_out[4696] = ~(layer1_out[6046] & layer1_out[6047]);
    assign layer2_out[4697] = layer1_out[787] | layer1_out[788];
    assign layer2_out[4698] = layer1_out[7503];
    assign layer2_out[4699] = layer1_out[3414] & layer1_out[3415];
    assign layer2_out[4700] = layer1_out[2608];
    assign layer2_out[4701] = layer1_out[4010] & ~layer1_out[4011];
    assign layer2_out[4702] = layer1_out[6220] | layer1_out[6221];
    assign layer2_out[4703] = ~layer1_out[2123] | layer1_out[2124];
    assign layer2_out[4704] = layer1_out[667] & layer1_out[668];
    assign layer2_out[4705] = layer1_out[6775];
    assign layer2_out[4706] = layer1_out[172] & ~layer1_out[173];
    assign layer2_out[4707] = layer1_out[507] & ~layer1_out[508];
    assign layer2_out[4708] = ~layer1_out[101] | layer1_out[100];
    assign layer2_out[4709] = ~layer1_out[4274];
    assign layer2_out[4710] = layer1_out[4783] & layer1_out[4784];
    assign layer2_out[4711] = layer1_out[3491];
    assign layer2_out[4712] = ~layer1_out[3108];
    assign layer2_out[4713] = ~layer1_out[1953];
    assign layer2_out[4714] = ~layer1_out[4933] | layer1_out[4934];
    assign layer2_out[4715] = ~layer1_out[2116];
    assign layer2_out[4716] = layer1_out[6089] & ~layer1_out[6090];
    assign layer2_out[4717] = ~(layer1_out[2458] | layer1_out[2459]);
    assign layer2_out[4718] = layer1_out[4914];
    assign layer2_out[4719] = ~(layer1_out[7529] | layer1_out[7530]);
    assign layer2_out[4720] = ~(layer1_out[1994] | layer1_out[1995]);
    assign layer2_out[4721] = ~layer1_out[2539];
    assign layer2_out[4722] = layer1_out[7662] & ~layer1_out[7661];
    assign layer2_out[4723] = layer1_out[6487];
    assign layer2_out[4724] = layer1_out[1736] & layer1_out[1737];
    assign layer2_out[4725] = layer1_out[722] & ~layer1_out[723];
    assign layer2_out[4726] = 1'b0;
    assign layer2_out[4727] = layer1_out[1372] & ~layer1_out[1371];
    assign layer2_out[4728] = layer1_out[4001] & layer1_out[4002];
    assign layer2_out[4729] = ~(layer1_out[5996] | layer1_out[5997]);
    assign layer2_out[4730] = layer1_out[5657] | layer1_out[5658];
    assign layer2_out[4731] = ~(layer1_out[2426] | layer1_out[2427]);
    assign layer2_out[4732] = 1'b0;
    assign layer2_out[4733] = ~(layer1_out[858] ^ layer1_out[859]);
    assign layer2_out[4734] = layer1_out[3160] & ~layer1_out[3159];
    assign layer2_out[4735] = ~(layer1_out[6243] | layer1_out[6244]);
    assign layer2_out[4736] = layer1_out[6469];
    assign layer2_out[4737] = layer1_out[2901];
    assign layer2_out[4738] = layer1_out[4366] | layer1_out[4367];
    assign layer2_out[4739] = ~layer1_out[4062];
    assign layer2_out[4740] = ~layer1_out[650] | layer1_out[649];
    assign layer2_out[4741] = layer1_out[2890] & layer1_out[2891];
    assign layer2_out[4742] = layer1_out[7833] ^ layer1_out[7834];
    assign layer2_out[4743] = layer1_out[7047] ^ layer1_out[7048];
    assign layer2_out[4744] = ~(layer1_out[4877] | layer1_out[4878]);
    assign layer2_out[4745] = layer1_out[6553];
    assign layer2_out[4746] = ~(layer1_out[4770] | layer1_out[4771]);
    assign layer2_out[4747] = ~layer1_out[6718];
    assign layer2_out[4748] = ~layer1_out[719];
    assign layer2_out[4749] = 1'b1;
    assign layer2_out[4750] = ~layer1_out[2298] | layer1_out[2297];
    assign layer2_out[4751] = layer1_out[7673] | layer1_out[7674];
    assign layer2_out[4752] = layer1_out[912];
    assign layer2_out[4753] = layer1_out[5157] ^ layer1_out[5158];
    assign layer2_out[4754] = layer1_out[3902] & ~layer1_out[3903];
    assign layer2_out[4755] = 1'b0;
    assign layer2_out[4756] = layer1_out[5341];
    assign layer2_out[4757] = layer1_out[4989];
    assign layer2_out[4758] = layer1_out[1303] | layer1_out[1304];
    assign layer2_out[4759] = ~(layer1_out[2995] | layer1_out[2996]);
    assign layer2_out[4760] = ~(layer1_out[6322] ^ layer1_out[6323]);
    assign layer2_out[4761] = ~layer1_out[972];
    assign layer2_out[4762] = ~(layer1_out[5495] | layer1_out[5496]);
    assign layer2_out[4763] = layer1_out[5423];
    assign layer2_out[4764] = ~layer1_out[3340];
    assign layer2_out[4765] = ~layer1_out[780] | layer1_out[781];
    assign layer2_out[4766] = ~layer1_out[3888] | layer1_out[3889];
    assign layer2_out[4767] = ~(layer1_out[4339] & layer1_out[4340]);
    assign layer2_out[4768] = layer1_out[4342];
    assign layer2_out[4769] = layer1_out[5476] & layer1_out[5477];
    assign layer2_out[4770] = ~(layer1_out[4868] & layer1_out[4869]);
    assign layer2_out[4771] = layer1_out[2266];
    assign layer2_out[4772] = layer1_out[5583] & ~layer1_out[5584];
    assign layer2_out[4773] = ~layer1_out[4376] | layer1_out[4377];
    assign layer2_out[4774] = layer1_out[1635] ^ layer1_out[1636];
    assign layer2_out[4775] = ~(layer1_out[3125] ^ layer1_out[3126]);
    assign layer2_out[4776] = ~layer1_out[2066] | layer1_out[2067];
    assign layer2_out[4777] = ~layer1_out[5701];
    assign layer2_out[4778] = ~(layer1_out[3995] | layer1_out[3996]);
    assign layer2_out[4779] = layer1_out[29];
    assign layer2_out[4780] = ~layer1_out[4029];
    assign layer2_out[4781] = ~layer1_out[5288];
    assign layer2_out[4782] = layer1_out[3107];
    assign layer2_out[4783] = ~layer1_out[5930];
    assign layer2_out[4784] = ~(layer1_out[109] & layer1_out[110]);
    assign layer2_out[4785] = ~layer1_out[2722] | layer1_out[2721];
    assign layer2_out[4786] = layer1_out[7621] | layer1_out[7622];
    assign layer2_out[4787] = layer1_out[4932] | layer1_out[4933];
    assign layer2_out[4788] = layer1_out[6385] & layer1_out[6386];
    assign layer2_out[4789] = layer1_out[5659] ^ layer1_out[5660];
    assign layer2_out[4790] = layer1_out[3863];
    assign layer2_out[4791] = ~(layer1_out[4150] & layer1_out[4151]);
    assign layer2_out[4792] = layer1_out[4785] & ~layer1_out[4784];
    assign layer2_out[4793] = ~layer1_out[906];
    assign layer2_out[4794] = layer1_out[7977] & layer1_out[7978];
    assign layer2_out[4795] = ~layer1_out[7948];
    assign layer2_out[4796] = ~(layer1_out[1533] & layer1_out[1534]);
    assign layer2_out[4797] = ~layer1_out[841];
    assign layer2_out[4798] = ~layer1_out[5812];
    assign layer2_out[4799] = layer1_out[6435];
    assign layer2_out[4800] = ~layer1_out[260] | layer1_out[259];
    assign layer2_out[4801] = ~layer1_out[20];
    assign layer2_out[4802] = ~(layer1_out[7400] & layer1_out[7401]);
    assign layer2_out[4803] = layer1_out[2728];
    assign layer2_out[4804] = ~layer1_out[5446];
    assign layer2_out[4805] = ~(layer1_out[2110] | layer1_out[2111]);
    assign layer2_out[4806] = layer1_out[314] & ~layer1_out[315];
    assign layer2_out[4807] = ~(layer1_out[3061] ^ layer1_out[3062]);
    assign layer2_out[4808] = ~layer1_out[6] | layer1_out[7];
    assign layer2_out[4809] = ~layer1_out[5706];
    assign layer2_out[4810] = ~layer1_out[733];
    assign layer2_out[4811] = ~layer1_out[6658];
    assign layer2_out[4812] = ~layer1_out[7216] | layer1_out[7215];
    assign layer2_out[4813] = ~layer1_out[6816] | layer1_out[6815];
    assign layer2_out[4814] = layer1_out[4564] ^ layer1_out[4565];
    assign layer2_out[4815] = ~layer1_out[2998] | layer1_out[2997];
    assign layer2_out[4816] = ~(layer1_out[1355] & layer1_out[1356]);
    assign layer2_out[4817] = layer1_out[6918] | layer1_out[6919];
    assign layer2_out[4818] = ~(layer1_out[5892] ^ layer1_out[5893]);
    assign layer2_out[4819] = 1'b1;
    assign layer2_out[4820] = ~(layer1_out[1908] | layer1_out[1909]);
    assign layer2_out[4821] = layer1_out[3480];
    assign layer2_out[4822] = ~layer1_out[1336];
    assign layer2_out[4823] = layer1_out[5183];
    assign layer2_out[4824] = layer1_out[1644] & ~layer1_out[1643];
    assign layer2_out[4825] = layer1_out[6280] & ~layer1_out[6281];
    assign layer2_out[4826] = ~layer1_out[248] | layer1_out[249];
    assign layer2_out[4827] = ~layer1_out[5470] | layer1_out[5469];
    assign layer2_out[4828] = ~layer1_out[919];
    assign layer2_out[4829] = layer1_out[1277] & layer1_out[1278];
    assign layer2_out[4830] = ~layer1_out[3563] | layer1_out[3562];
    assign layer2_out[4831] = layer1_out[1038];
    assign layer2_out[4832] = ~layer1_out[5864] | layer1_out[5863];
    assign layer2_out[4833] = ~layer1_out[1881] | layer1_out[1882];
    assign layer2_out[4834] = layer1_out[4882];
    assign layer2_out[4835] = layer1_out[2468] & ~layer1_out[2469];
    assign layer2_out[4836] = layer1_out[2052] | layer1_out[2053];
    assign layer2_out[4837] = ~(layer1_out[5757] | layer1_out[5758]);
    assign layer2_out[4838] = layer1_out[6790];
    assign layer2_out[4839] = layer1_out[161];
    assign layer2_out[4840] = layer1_out[4866] & layer1_out[4867];
    assign layer2_out[4841] = layer1_out[5904];
    assign layer2_out[4842] = ~layer1_out[5759] | layer1_out[5758];
    assign layer2_out[4843] = ~(layer1_out[6559] | layer1_out[6560]);
    assign layer2_out[4844] = ~(layer1_out[519] ^ layer1_out[520]);
    assign layer2_out[4845] = ~(layer1_out[2169] ^ layer1_out[2170]);
    assign layer2_out[4846] = layer1_out[3736] & ~layer1_out[3737];
    assign layer2_out[4847] = layer1_out[7665];
    assign layer2_out[4848] = ~layer1_out[5875] | layer1_out[5876];
    assign layer2_out[4849] = layer1_out[6531] & ~layer1_out[6532];
    assign layer2_out[4850] = layer1_out[6206] | layer1_out[6207];
    assign layer2_out[4851] = layer1_out[7588] & ~layer1_out[7587];
    assign layer2_out[4852] = layer1_out[6525];
    assign layer2_out[4853] = 1'b1;
    assign layer2_out[4854] = layer1_out[6702] | layer1_out[6703];
    assign layer2_out[4855] = ~(layer1_out[1668] | layer1_out[1669]);
    assign layer2_out[4856] = layer1_out[7763] & layer1_out[7764];
    assign layer2_out[4857] = ~(layer1_out[6614] & layer1_out[6615]);
    assign layer2_out[4858] = ~layer1_out[2461];
    assign layer2_out[4859] = 1'b1;
    assign layer2_out[4860] = ~layer1_out[5944];
    assign layer2_out[4861] = ~layer1_out[7539];
    assign layer2_out[4862] = 1'b1;
    assign layer2_out[4863] = layer1_out[3189] & ~layer1_out[3190];
    assign layer2_out[4864] = layer1_out[2210] ^ layer1_out[2211];
    assign layer2_out[4865] = ~(layer1_out[7819] & layer1_out[7820]);
    assign layer2_out[4866] = ~(layer1_out[5300] & layer1_out[5301]);
    assign layer2_out[4867] = layer1_out[7550];
    assign layer2_out[4868] = layer1_out[6622] ^ layer1_out[6623];
    assign layer2_out[4869] = layer1_out[2712] & layer1_out[2713];
    assign layer2_out[4870] = ~layer1_out[1111] | layer1_out[1110];
    assign layer2_out[4871] = ~layer1_out[1307] | layer1_out[1308];
    assign layer2_out[4872] = layer1_out[6496];
    assign layer2_out[4873] = ~layer1_out[4125] | layer1_out[4124];
    assign layer2_out[4874] = layer1_out[4658] & layer1_out[4659];
    assign layer2_out[4875] = layer1_out[7079];
    assign layer2_out[4876] = layer1_out[192] & ~layer1_out[191];
    assign layer2_out[4877] = layer1_out[3640] & ~layer1_out[3639];
    assign layer2_out[4878] = layer1_out[3119];
    assign layer2_out[4879] = layer1_out[3285];
    assign layer2_out[4880] = ~(layer1_out[5085] & layer1_out[5086]);
    assign layer2_out[4881] = layer1_out[2629];
    assign layer2_out[4882] = layer1_out[7256];
    assign layer2_out[4883] = layer1_out[531];
    assign layer2_out[4884] = layer1_out[3797] & layer1_out[3798];
    assign layer2_out[4885] = layer1_out[2736] & layer1_out[2737];
    assign layer2_out[4886] = layer1_out[2369];
    assign layer2_out[4887] = layer1_out[5442] | layer1_out[5443];
    assign layer2_out[4888] = ~layer1_out[1212] | layer1_out[1213];
    assign layer2_out[4889] = 1'b0;
    assign layer2_out[4890] = ~(layer1_out[4091] & layer1_out[4092]);
    assign layer2_out[4891] = layer1_out[984] | layer1_out[985];
    assign layer2_out[4892] = layer1_out[3890] ^ layer1_out[3891];
    assign layer2_out[4893] = ~layer1_out[2434];
    assign layer2_out[4894] = ~layer1_out[6067] | layer1_out[6066];
    assign layer2_out[4895] = 1'b1;
    assign layer2_out[4896] = ~layer1_out[228] | layer1_out[227];
    assign layer2_out[4897] = ~layer1_out[4934] | layer1_out[4935];
    assign layer2_out[4898] = layer1_out[1207] | layer1_out[1208];
    assign layer2_out[4899] = ~(layer1_out[5462] | layer1_out[5463]);
    assign layer2_out[4900] = layer1_out[5820] & ~layer1_out[5819];
    assign layer2_out[4901] = layer1_out[5696] ^ layer1_out[5697];
    assign layer2_out[4902] = ~(layer1_out[7810] | layer1_out[7811]);
    assign layer2_out[4903] = ~layer1_out[7596];
    assign layer2_out[4904] = layer1_out[3117];
    assign layer2_out[4905] = ~layer1_out[1201] | layer1_out[1202];
    assign layer2_out[4906] = ~(layer1_out[5045] & layer1_out[5046]);
    assign layer2_out[4907] = ~layer1_out[7137];
    assign layer2_out[4908] = ~(layer1_out[2025] ^ layer1_out[2026]);
    assign layer2_out[4909] = layer1_out[1272] & ~layer1_out[1271];
    assign layer2_out[4910] = layer1_out[4558] ^ layer1_out[4559];
    assign layer2_out[4911] = ~(layer1_out[7990] | layer1_out[7991]);
    assign layer2_out[4912] = layer1_out[6999] & ~layer1_out[7000];
    assign layer2_out[4913] = layer1_out[2430] & ~layer1_out[2431];
    assign layer2_out[4914] = 1'b1;
    assign layer2_out[4915] = 1'b0;
    assign layer2_out[4916] = layer1_out[2232];
    assign layer2_out[4917] = 1'b1;
    assign layer2_out[4918] = layer1_out[5812];
    assign layer2_out[4919] = ~layer1_out[5916];
    assign layer2_out[4920] = layer1_out[2089] | layer1_out[2090];
    assign layer2_out[4921] = layer1_out[221] & ~layer1_out[220];
    assign layer2_out[4922] = ~(layer1_out[5068] & layer1_out[5069]);
    assign layer2_out[4923] = ~layer1_out[3083];
    assign layer2_out[4924] = ~(layer1_out[5213] & layer1_out[5214]);
    assign layer2_out[4925] = ~layer1_out[4657] | layer1_out[4658];
    assign layer2_out[4926] = ~layer1_out[680] | layer1_out[679];
    assign layer2_out[4927] = layer1_out[5853];
    assign layer2_out[4928] = ~layer1_out[7590] | layer1_out[7589];
    assign layer2_out[4929] = layer1_out[3314] & layer1_out[3315];
    assign layer2_out[4930] = layer1_out[5230] | layer1_out[5231];
    assign layer2_out[4931] = ~layer1_out[5926];
    assign layer2_out[4932] = layer1_out[1985] | layer1_out[1986];
    assign layer2_out[4933] = layer1_out[7158];
    assign layer2_out[4934] = ~layer1_out[5598] | layer1_out[5597];
    assign layer2_out[4935] = ~layer1_out[3919] | layer1_out[3918];
    assign layer2_out[4936] = layer1_out[2287] & layer1_out[2288];
    assign layer2_out[4937] = ~layer1_out[1802];
    assign layer2_out[4938] = ~(layer1_out[7862] | layer1_out[7863]);
    assign layer2_out[4939] = layer1_out[7908] & layer1_out[7909];
    assign layer2_out[4940] = ~layer1_out[3238];
    assign layer2_out[4941] = ~layer1_out[7869];
    assign layer2_out[4942] = layer1_out[6899] | layer1_out[6900];
    assign layer2_out[4943] = ~layer1_out[7453];
    assign layer2_out[4944] = layer1_out[1019];
    assign layer2_out[4945] = ~(layer1_out[315] & layer1_out[316]);
    assign layer2_out[4946] = ~layer1_out[2950];
    assign layer2_out[4947] = ~layer1_out[4362] | layer1_out[4363];
    assign layer2_out[4948] = layer1_out[1969];
    assign layer2_out[4949] = layer1_out[6013] & ~layer1_out[6014];
    assign layer2_out[4950] = layer1_out[573];
    assign layer2_out[4951] = layer1_out[6189] & ~layer1_out[6190];
    assign layer2_out[4952] = ~layer1_out[2868];
    assign layer2_out[4953] = layer1_out[1964];
    assign layer2_out[4954] = layer1_out[3453] | layer1_out[3454];
    assign layer2_out[4955] = layer1_out[3472] & ~layer1_out[3473];
    assign layer2_out[4956] = ~layer1_out[978];
    assign layer2_out[4957] = layer1_out[5331];
    assign layer2_out[4958] = layer1_out[4610] ^ layer1_out[4611];
    assign layer2_out[4959] = layer1_out[4673] & ~layer1_out[4672];
    assign layer2_out[4960] = layer1_out[3680] & ~layer1_out[3681];
    assign layer2_out[4961] = layer1_out[4912] | layer1_out[4913];
    assign layer2_out[4962] = layer1_out[3576] & ~layer1_out[3575];
    assign layer2_out[4963] = ~layer1_out[118];
    assign layer2_out[4964] = ~layer1_out[273] | layer1_out[274];
    assign layer2_out[4965] = layer1_out[2139] | layer1_out[2140];
    assign layer2_out[4966] = layer1_out[4876] & layer1_out[4877];
    assign layer2_out[4967] = layer1_out[4099] & layer1_out[4100];
    assign layer2_out[4968] = layer1_out[2823] & layer1_out[2824];
    assign layer2_out[4969] = layer1_out[427];
    assign layer2_out[4970] = ~layer1_out[7170];
    assign layer2_out[4971] = ~layer1_out[4171] | layer1_out[4170];
    assign layer2_out[4972] = ~(layer1_out[1369] | layer1_out[1370]);
    assign layer2_out[4973] = layer1_out[3423] ^ layer1_out[3424];
    assign layer2_out[4974] = layer1_out[1725] & ~layer1_out[1726];
    assign layer2_out[4975] = ~layer1_out[4443] | layer1_out[4442];
    assign layer2_out[4976] = layer1_out[7877] & ~layer1_out[7876];
    assign layer2_out[4977] = layer1_out[6683] & ~layer1_out[6682];
    assign layer2_out[4978] = ~layer1_out[6451];
    assign layer2_out[4979] = layer1_out[2675] | layer1_out[2676];
    assign layer2_out[4980] = ~layer1_out[2837] | layer1_out[2838];
    assign layer2_out[4981] = layer1_out[1066];
    assign layer2_out[4982] = ~layer1_out[6190];
    assign layer2_out[4983] = layer1_out[7727];
    assign layer2_out[4984] = ~layer1_out[1263] | layer1_out[1262];
    assign layer2_out[4985] = ~layer1_out[1956] | layer1_out[1955];
    assign layer2_out[4986] = ~(layer1_out[1000] | layer1_out[1001]);
    assign layer2_out[4987] = ~(layer1_out[1598] & layer1_out[1599]);
    assign layer2_out[4988] = layer1_out[2951];
    assign layer2_out[4989] = 1'b1;
    assign layer2_out[4990] = ~(layer1_out[6843] & layer1_out[6844]);
    assign layer2_out[4991] = layer1_out[1782] & layer1_out[1783];
    assign layer2_out[4992] = layer1_out[7087] & ~layer1_out[7088];
    assign layer2_out[4993] = ~(layer1_out[6987] | layer1_out[6988]);
    assign layer2_out[4994] = layer1_out[5611] & layer1_out[5612];
    assign layer2_out[4995] = layer1_out[1830];
    assign layer2_out[4996] = ~layer1_out[1626];
    assign layer2_out[4997] = ~layer1_out[1681];
    assign layer2_out[4998] = layer1_out[4756] | layer1_out[4757];
    assign layer2_out[4999] = layer1_out[7426] & ~layer1_out[7427];
    assign layer2_out[5000] = ~(layer1_out[1063] | layer1_out[1064]);
    assign layer2_out[5001] = ~(layer1_out[3405] & layer1_out[3406]);
    assign layer2_out[5002] = layer1_out[5712];
    assign layer2_out[5003] = ~layer1_out[5284] | layer1_out[5285];
    assign layer2_out[5004] = layer1_out[7832] & layer1_out[7833];
    assign layer2_out[5005] = ~layer1_out[5101] | layer1_out[5102];
    assign layer2_out[5006] = layer1_out[1068] & ~layer1_out[1067];
    assign layer2_out[5007] = layer1_out[1304] | layer1_out[1305];
    assign layer2_out[5008] = layer1_out[4271] & ~layer1_out[4270];
    assign layer2_out[5009] = layer1_out[5312] & ~layer1_out[5311];
    assign layer2_out[5010] = ~(layer1_out[6779] & layer1_out[6780]);
    assign layer2_out[5011] = ~layer1_out[4573] | layer1_out[4574];
    assign layer2_out[5012] = layer1_out[3931] & ~layer1_out[3930];
    assign layer2_out[5013] = layer1_out[6304] & ~layer1_out[6305];
    assign layer2_out[5014] = layer1_out[3066];
    assign layer2_out[5015] = layer1_out[7028] & layer1_out[7029];
    assign layer2_out[5016] = layer1_out[4148] ^ layer1_out[4149];
    assign layer2_out[5017] = layer1_out[387] ^ layer1_out[388];
    assign layer2_out[5018] = ~(layer1_out[2420] | layer1_out[2421]);
    assign layer2_out[5019] = layer1_out[7348] & ~layer1_out[7349];
    assign layer2_out[5020] = ~layer1_out[1600];
    assign layer2_out[5021] = layer1_out[3336] | layer1_out[3337];
    assign layer2_out[5022] = layer1_out[5079];
    assign layer2_out[5023] = layer1_out[975] | layer1_out[976];
    assign layer2_out[5024] = ~layer1_out[2547] | layer1_out[2548];
    assign layer2_out[5025] = layer1_out[5774] ^ layer1_out[5775];
    assign layer2_out[5026] = layer1_out[6809];
    assign layer2_out[5027] = layer1_out[5707] & layer1_out[5708];
    assign layer2_out[5028] = ~layer1_out[151] | layer1_out[152];
    assign layer2_out[5029] = 1'b1;
    assign layer2_out[5030] = 1'b0;
    assign layer2_out[5031] = layer1_out[5465];
    assign layer2_out[5032] = ~layer1_out[2935];
    assign layer2_out[5033] = ~layer1_out[5650];
    assign layer2_out[5034] = ~layer1_out[6227] | layer1_out[6228];
    assign layer2_out[5035] = ~layer1_out[2130] | layer1_out[2131];
    assign layer2_out[5036] = ~layer1_out[534];
    assign layer2_out[5037] = layer1_out[4265] ^ layer1_out[4266];
    assign layer2_out[5038] = layer1_out[5511] & layer1_out[5512];
    assign layer2_out[5039] = ~(layer1_out[5718] & layer1_out[5719]);
    assign layer2_out[5040] = ~layer1_out[2228];
    assign layer2_out[5041] = 1'b1;
    assign layer2_out[5042] = ~layer1_out[1562];
    assign layer2_out[5043] = ~layer1_out[1660];
    assign layer2_out[5044] = 1'b1;
    assign layer2_out[5045] = ~layer1_out[266];
    assign layer2_out[5046] = 1'b1;
    assign layer2_out[5047] = layer1_out[7224] & ~layer1_out[7225];
    assign layer2_out[5048] = layer1_out[3461];
    assign layer2_out[5049] = layer1_out[3637] & ~layer1_out[3638];
    assign layer2_out[5050] = layer1_out[5074];
    assign layer2_out[5051] = ~(layer1_out[1440] | layer1_out[1441]);
    assign layer2_out[5052] = ~(layer1_out[5630] ^ layer1_out[5631]);
    assign layer2_out[5053] = layer1_out[5677] & ~layer1_out[5676];
    assign layer2_out[5054] = ~layer1_out[4819] | layer1_out[4818];
    assign layer2_out[5055] = ~(layer1_out[3034] | layer1_out[3035]);
    assign layer2_out[5056] = layer1_out[3492] & layer1_out[3493];
    assign layer2_out[5057] = ~layer1_out[3660] | layer1_out[3661];
    assign layer2_out[5058] = layer1_out[2939] | layer1_out[2940];
    assign layer2_out[5059] = layer1_out[445] & layer1_out[446];
    assign layer2_out[5060] = ~(layer1_out[3679] | layer1_out[3680]);
    assign layer2_out[5061] = ~layer1_out[2965];
    assign layer2_out[5062] = layer1_out[6201];
    assign layer2_out[5063] = ~(layer1_out[2158] & layer1_out[2159]);
    assign layer2_out[5064] = layer1_out[169];
    assign layer2_out[5065] = ~layer1_out[6059];
    assign layer2_out[5066] = ~layer1_out[3579];
    assign layer2_out[5067] = layer1_out[512] & ~layer1_out[511];
    assign layer2_out[5068] = layer1_out[5006] & ~layer1_out[5005];
    assign layer2_out[5069] = layer1_out[7848];
    assign layer2_out[5070] = ~layer1_out[7747];
    assign layer2_out[5071] = ~layer1_out[7947] | layer1_out[7946];
    assign layer2_out[5072] = layer1_out[3325];
    assign layer2_out[5073] = ~layer1_out[6991] | layer1_out[6990];
    assign layer2_out[5074] = ~(layer1_out[7692] ^ layer1_out[7693]);
    assign layer2_out[5075] = ~layer1_out[5023];
    assign layer2_out[5076] = 1'b1;
    assign layer2_out[5077] = layer1_out[443] & layer1_out[444];
    assign layer2_out[5078] = layer1_out[7523];
    assign layer2_out[5079] = ~layer1_out[5298];
    assign layer2_out[5080] = layer1_out[1892];
    assign layer2_out[5081] = ~layer1_out[2341];
    assign layer2_out[5082] = layer1_out[5350] & ~layer1_out[5349];
    assign layer2_out[5083] = ~layer1_out[597];
    assign layer2_out[5084] = ~(layer1_out[4792] & layer1_out[4793]);
    assign layer2_out[5085] = ~(layer1_out[3798] & layer1_out[3799]);
    assign layer2_out[5086] = layer1_out[1548] & layer1_out[1549];
    assign layer2_out[5087] = ~layer1_out[3369] | layer1_out[3370];
    assign layer2_out[5088] = layer1_out[4102] & layer1_out[4103];
    assign layer2_out[5089] = layer1_out[2593] & layer1_out[2594];
    assign layer2_out[5090] = layer1_out[357];
    assign layer2_out[5091] = layer1_out[5035] & ~layer1_out[5034];
    assign layer2_out[5092] = layer1_out[497] | layer1_out[498];
    assign layer2_out[5093] = ~layer1_out[7683];
    assign layer2_out[5094] = layer1_out[4838];
    assign layer2_out[5095] = ~(layer1_out[4453] & layer1_out[4454]);
    assign layer2_out[5096] = 1'b1;
    assign layer2_out[5097] = layer1_out[2983];
    assign layer2_out[5098] = layer1_out[3099] & ~layer1_out[3098];
    assign layer2_out[5099] = layer1_out[6321] ^ layer1_out[6322];
    assign layer2_out[5100] = ~layer1_out[5037] | layer1_out[5036];
    assign layer2_out[5101] = layer1_out[1443];
    assign layer2_out[5102] = layer1_out[705] & layer1_out[706];
    assign layer2_out[5103] = ~layer1_out[4193];
    assign layer2_out[5104] = layer1_out[6072] & layer1_out[6073];
    assign layer2_out[5105] = layer1_out[3555] & ~layer1_out[3554];
    assign layer2_out[5106] = ~(layer1_out[2068] | layer1_out[2069]);
    assign layer2_out[5107] = layer1_out[7706];
    assign layer2_out[5108] = ~layer1_out[5872];
    assign layer2_out[5109] = ~(layer1_out[5397] & layer1_out[5398]);
    assign layer2_out[5110] = layer1_out[4470] & layer1_out[4471];
    assign layer2_out[5111] = layer1_out[6643] | layer1_out[6644];
    assign layer2_out[5112] = ~layer1_out[7359];
    assign layer2_out[5113] = ~layer1_out[31] | layer1_out[30];
    assign layer2_out[5114] = ~layer1_out[7130];
    assign layer2_out[5115] = ~(layer1_out[2926] & layer1_out[2927]);
    assign layer2_out[5116] = ~layer1_out[7785];
    assign layer2_out[5117] = layer1_out[969] | layer1_out[970];
    assign layer2_out[5118] = layer1_out[2968] ^ layer1_out[2969];
    assign layer2_out[5119] = ~layer1_out[13] | layer1_out[14];
    assign layer2_out[5120] = ~(layer1_out[5193] | layer1_out[5194]);
    assign layer2_out[5121] = layer1_out[7066] & layer1_out[7067];
    assign layer2_out[5122] = ~layer1_out[5814];
    assign layer2_out[5123] = ~layer1_out[3080];
    assign layer2_out[5124] = layer1_out[2865] & ~layer1_out[2864];
    assign layer2_out[5125] = 1'b1;
    assign layer2_out[5126] = layer1_out[4675] ^ layer1_out[4676];
    assign layer2_out[5127] = ~layer1_out[2691];
    assign layer2_out[5128] = layer1_out[1591];
    assign layer2_out[5129] = 1'b0;
    assign layer2_out[5130] = layer1_out[926] & ~layer1_out[925];
    assign layer2_out[5131] = ~(layer1_out[3760] | layer1_out[3761]);
    assign layer2_out[5132] = ~(layer1_out[2119] | layer1_out[2120]);
    assign layer2_out[5133] = ~(layer1_out[3770] | layer1_out[3771]);
    assign layer2_out[5134] = ~layer1_out[2249] | layer1_out[2248];
    assign layer2_out[5135] = ~(layer1_out[5842] | layer1_out[5843]);
    assign layer2_out[5136] = ~(layer1_out[2940] ^ layer1_out[2941]);
    assign layer2_out[5137] = layer1_out[1654] & ~layer1_out[1655];
    assign layer2_out[5138] = layer1_out[1958] & layer1_out[1959];
    assign layer2_out[5139] = layer1_out[6145] ^ layer1_out[6146];
    assign layer2_out[5140] = ~layer1_out[4287];
    assign layer2_out[5141] = ~layer1_out[6887] | layer1_out[6886];
    assign layer2_out[5142] = ~layer1_out[4991];
    assign layer2_out[5143] = layer1_out[5040] | layer1_out[5041];
    assign layer2_out[5144] = ~layer1_out[1738] | layer1_out[1737];
    assign layer2_out[5145] = layer1_out[4355] & layer1_out[4356];
    assign layer2_out[5146] = layer1_out[6792] | layer1_out[6793];
    assign layer2_out[5147] = ~layer1_out[6589];
    assign layer2_out[5148] = layer1_out[3915] ^ layer1_out[3916];
    assign layer2_out[5149] = ~(layer1_out[7356] | layer1_out[7357]);
    assign layer2_out[5150] = 1'b1;
    assign layer2_out[5151] = ~(layer1_out[4255] ^ layer1_out[4256]);
    assign layer2_out[5152] = ~layer1_out[431] | layer1_out[430];
    assign layer2_out[5153] = layer1_out[1653];
    assign layer2_out[5154] = 1'b1;
    assign layer2_out[5155] = layer1_out[1544] & ~layer1_out[1543];
    assign layer2_out[5156] = ~layer1_out[5590] | layer1_out[5589];
    assign layer2_out[5157] = ~layer1_out[1580];
    assign layer2_out[5158] = layer1_out[4108] | layer1_out[4109];
    assign layer2_out[5159] = layer1_out[161] | layer1_out[162];
    assign layer2_out[5160] = ~layer1_out[2592];
    assign layer2_out[5161] = layer1_out[3558] & ~layer1_out[3559];
    assign layer2_out[5162] = layer1_out[3525];
    assign layer2_out[5163] = layer1_out[5755] & ~layer1_out[5754];
    assign layer2_out[5164] = layer1_out[2184];
    assign layer2_out[5165] = layer1_out[5127] & ~layer1_out[5128];
    assign layer2_out[5166] = layer1_out[6063] ^ layer1_out[6064];
    assign layer2_out[5167] = ~layer1_out[735] | layer1_out[734];
    assign layer2_out[5168] = ~layer1_out[7668];
    assign layer2_out[5169] = ~layer1_out[7800];
    assign layer2_out[5170] = layer1_out[648];
    assign layer2_out[5171] = layer1_out[3214] & ~layer1_out[3213];
    assign layer2_out[5172] = layer1_out[5816] & ~layer1_out[5815];
    assign layer2_out[5173] = ~layer1_out[662];
    assign layer2_out[5174] = layer1_out[2569] & ~layer1_out[2568];
    assign layer2_out[5175] = layer1_out[2359];
    assign layer2_out[5176] = layer1_out[4230];
    assign layer2_out[5177] = ~(layer1_out[4245] | layer1_out[4246]);
    assign layer2_out[5178] = ~layer1_out[744];
    assign layer2_out[5179] = ~(layer1_out[4326] | layer1_out[4327]);
    assign layer2_out[5180] = ~layer1_out[1224];
    assign layer2_out[5181] = ~layer1_out[6236] | layer1_out[6237];
    assign layer2_out[5182] = ~(layer1_out[3922] | layer1_out[3923]);
    assign layer2_out[5183] = layer1_out[2909] & ~layer1_out[2910];
    assign layer2_out[5184] = layer1_out[1142];
    assign layer2_out[5185] = ~layer1_out[4609];
    assign layer2_out[5186] = ~layer1_out[7510] | layer1_out[7511];
    assign layer2_out[5187] = 1'b0;
    assign layer2_out[5188] = layer1_out[7765];
    assign layer2_out[5189] = layer1_out[4426];
    assign layer2_out[5190] = layer1_out[1149] ^ layer1_out[1150];
    assign layer2_out[5191] = layer1_out[1452];
    assign layer2_out[5192] = layer1_out[1328] & ~layer1_out[1327];
    assign layer2_out[5193] = ~layer1_out[937] | layer1_out[936];
    assign layer2_out[5194] = ~layer1_out[1971];
    assign layer2_out[5195] = ~layer1_out[2064];
    assign layer2_out[5196] = ~layer1_out[975];
    assign layer2_out[5197] = ~layer1_out[4790] | layer1_out[4789];
    assign layer2_out[5198] = ~(layer1_out[6458] & layer1_out[6459]);
    assign layer2_out[5199] = ~(layer1_out[6265] ^ layer1_out[6266]);
    assign layer2_out[5200] = layer1_out[166];
    assign layer2_out[5201] = ~(layer1_out[1604] & layer1_out[1605]);
    assign layer2_out[5202] = layer1_out[7030];
    assign layer2_out[5203] = ~(layer1_out[2114] | layer1_out[2115]);
    assign layer2_out[5204] = ~layer1_out[5584];
    assign layer2_out[5205] = layer1_out[5185] | layer1_out[5186];
    assign layer2_out[5206] = ~layer1_out[6675];
    assign layer2_out[5207] = ~layer1_out[6024];
    assign layer2_out[5208] = layer1_out[2559] & ~layer1_out[2560];
    assign layer2_out[5209] = 1'b1;
    assign layer2_out[5210] = layer1_out[7556] & ~layer1_out[7555];
    assign layer2_out[5211] = ~layer1_out[4199];
    assign layer2_out[5212] = layer1_out[3773] & ~layer1_out[3772];
    assign layer2_out[5213] = ~layer1_out[3713] | layer1_out[3712];
    assign layer2_out[5214] = ~layer1_out[4598] | layer1_out[4597];
    assign layer2_out[5215] = 1'b1;
    assign layer2_out[5216] = layer1_out[3035] | layer1_out[3036];
    assign layer2_out[5217] = layer1_out[5845] & layer1_out[5846];
    assign layer2_out[5218] = layer1_out[3796];
    assign layer2_out[5219] = ~layer1_out[4859];
    assign layer2_out[5220] = ~layer1_out[4861];
    assign layer2_out[5221] = layer1_out[6781];
    assign layer2_out[5222] = ~(layer1_out[4025] ^ layer1_out[4026]);
    assign layer2_out[5223] = ~layer1_out[1] | layer1_out[2];
    assign layer2_out[5224] = ~(layer1_out[2976] | layer1_out[2977]);
    assign layer2_out[5225] = ~layer1_out[3059];
    assign layer2_out[5226] = layer1_out[6366];
    assign layer2_out[5227] = ~(layer1_out[5102] | layer1_out[5103]);
    assign layer2_out[5228] = ~layer1_out[1202] | layer1_out[1203];
    assign layer2_out[5229] = ~layer1_out[7178] | layer1_out[7177];
    assign layer2_out[5230] = layer1_out[282];
    assign layer2_out[5231] = layer1_out[4406] & layer1_out[4407];
    assign layer2_out[5232] = ~layer1_out[3779] | layer1_out[3778];
    assign layer2_out[5233] = ~layer1_out[575] | layer1_out[576];
    assign layer2_out[5234] = layer1_out[4957];
    assign layer2_out[5235] = layer1_out[4364];
    assign layer2_out[5236] = layer1_out[2785];
    assign layer2_out[5237] = layer1_out[3298] & ~layer1_out[3299];
    assign layer2_out[5238] = ~layer1_out[6302] | layer1_out[6303];
    assign layer2_out[5239] = ~layer1_out[4263];
    assign layer2_out[5240] = layer1_out[1325] ^ layer1_out[1326];
    assign layer2_out[5241] = layer1_out[7695];
    assign layer2_out[5242] = layer1_out[7714] ^ layer1_out[7715];
    assign layer2_out[5243] = layer1_out[3544] & layer1_out[3545];
    assign layer2_out[5244] = ~(layer1_out[4126] | layer1_out[4127]);
    assign layer2_out[5245] = ~layer1_out[5841];
    assign layer2_out[5246] = layer1_out[1296] & layer1_out[1297];
    assign layer2_out[5247] = ~(layer1_out[6621] & layer1_out[6622]);
    assign layer2_out[5248] = layer1_out[2372];
    assign layer2_out[5249] = ~(layer1_out[3880] | layer1_out[3881]);
    assign layer2_out[5250] = layer1_out[6697];
    assign layer2_out[5251] = ~layer1_out[1699];
    assign layer2_out[5252] = ~layer1_out[6316];
    assign layer2_out[5253] = layer1_out[93] ^ layer1_out[94];
    assign layer2_out[5254] = 1'b0;
    assign layer2_out[5255] = layer1_out[2500] & ~layer1_out[2499];
    assign layer2_out[5256] = ~layer1_out[1490];
    assign layer2_out[5257] = ~(layer1_out[180] | layer1_out[181]);
    assign layer2_out[5258] = layer1_out[309] & ~layer1_out[308];
    assign layer2_out[5259] = ~layer1_out[6518];
    assign layer2_out[5260] = layer1_out[127];
    assign layer2_out[5261] = ~(layer1_out[6381] | layer1_out[6382]);
    assign layer2_out[5262] = layer1_out[7878];
    assign layer2_out[5263] = 1'b1;
    assign layer2_out[5264] = ~layer1_out[775] | layer1_out[776];
    assign layer2_out[5265] = 1'b0;
    assign layer2_out[5266] = ~(layer1_out[7196] ^ layer1_out[7197]);
    assign layer2_out[5267] = ~(layer1_out[7581] & layer1_out[7582]);
    assign layer2_out[5268] = ~layer1_out[3462] | layer1_out[3463];
    assign layer2_out[5269] = ~layer1_out[5969] | layer1_out[5970];
    assign layer2_out[5270] = ~layer1_out[1425] | layer1_out[1424];
    assign layer2_out[5271] = layer1_out[2263] ^ layer1_out[2264];
    assign layer2_out[5272] = layer1_out[3008] & ~layer1_out[3009];
    assign layer2_out[5273] = layer1_out[818];
    assign layer2_out[5274] = layer1_out[358];
    assign layer2_out[5275] = layer1_out[6096] & ~layer1_out[6095];
    assign layer2_out[5276] = ~layer1_out[1934] | layer1_out[1933];
    assign layer2_out[5277] = ~layer1_out[700];
    assign layer2_out[5278] = layer1_out[1374];
    assign layer2_out[5279] = layer1_out[4526];
    assign layer2_out[5280] = layer1_out[2339];
    assign layer2_out[5281] = layer1_out[2369] | layer1_out[2370];
    assign layer2_out[5282] = layer1_out[5556] ^ layer1_out[5557];
    assign layer2_out[5283] = 1'b1;
    assign layer2_out[5284] = ~layer1_out[6153];
    assign layer2_out[5285] = ~layer1_out[5167] | layer1_out[5168];
    assign layer2_out[5286] = ~layer1_out[7265] | layer1_out[7264];
    assign layer2_out[5287] = ~layer1_out[3010];
    assign layer2_out[5288] = layer1_out[2504];
    assign layer2_out[5289] = ~layer1_out[2464] | layer1_out[2465];
    assign layer2_out[5290] = 1'b0;
    assign layer2_out[5291] = ~(layer1_out[6865] ^ layer1_out[6866]);
    assign layer2_out[5292] = ~layer1_out[6173] | layer1_out[6174];
    assign layer2_out[5293] = layer1_out[7361];
    assign layer2_out[5294] = layer1_out[2643] | layer1_out[2644];
    assign layer2_out[5295] = layer1_out[6653];
    assign layer2_out[5296] = layer1_out[4067];
    assign layer2_out[5297] = layer1_out[7268] | layer1_out[7269];
    assign layer2_out[5298] = layer1_out[92] & layer1_out[93];
    assign layer2_out[5299] = layer1_out[3091];
    assign layer2_out[5300] = ~layer1_out[188];
    assign layer2_out[5301] = ~(layer1_out[6742] & layer1_out[6743]);
    assign layer2_out[5302] = layer1_out[1811] & ~layer1_out[1810];
    assign layer2_out[5303] = layer1_out[1889];
    assign layer2_out[5304] = ~layer1_out[5952] | layer1_out[5953];
    assign layer2_out[5305] = ~(layer1_out[7945] | layer1_out[7946]);
    assign layer2_out[5306] = ~layer1_out[7691] | layer1_out[7690];
    assign layer2_out[5307] = ~(layer1_out[3758] & layer1_out[3759]);
    assign layer2_out[5308] = layer1_out[5880] | layer1_out[5881];
    assign layer2_out[5309] = layer1_out[6694];
    assign layer2_out[5310] = ~layer1_out[5734] | layer1_out[5735];
    assign layer2_out[5311] = ~layer1_out[5320];
    assign layer2_out[5312] = ~layer1_out[2871] | layer1_out[2872];
    assign layer2_out[5313] = ~layer1_out[6578];
    assign layer2_out[5314] = 1'b0;
    assign layer2_out[5315] = layer1_out[5192];
    assign layer2_out[5316] = layer1_out[7574] & ~layer1_out[7575];
    assign layer2_out[5317] = layer1_out[5689] & ~layer1_out[5690];
    assign layer2_out[5318] = layer1_out[1826] & layer1_out[1827];
    assign layer2_out[5319] = ~layer1_out[5787];
    assign layer2_out[5320] = layer1_out[3991] & layer1_out[3992];
    assign layer2_out[5321] = layer1_out[7899] & ~layer1_out[7900];
    assign layer2_out[5322] = layer1_out[6384] & ~layer1_out[6385];
    assign layer2_out[5323] = layer1_out[4747] ^ layer1_out[4748];
    assign layer2_out[5324] = layer1_out[1011] & ~layer1_out[1012];
    assign layer2_out[5325] = layer1_out[6370] & ~layer1_out[6369];
    assign layer2_out[5326] = ~layer1_out[1793];
    assign layer2_out[5327] = layer1_out[7392] & layer1_out[7393];
    assign layer2_out[5328] = ~layer1_out[4993] | layer1_out[4992];
    assign layer2_out[5329] = ~(layer1_out[7432] | layer1_out[7433]);
    assign layer2_out[5330] = ~layer1_out[3358];
    assign layer2_out[5331] = ~(layer1_out[7895] | layer1_out[7896]);
    assign layer2_out[5332] = ~layer1_out[5038];
    assign layer2_out[5333] = layer1_out[5244] & ~layer1_out[5245];
    assign layer2_out[5334] = layer1_out[6279] & ~layer1_out[6278];
    assign layer2_out[5335] = layer1_out[3718];
    assign layer2_out[5336] = layer1_out[1508] ^ layer1_out[1509];
    assign layer2_out[5337] = layer1_out[1447];
    assign layer2_out[5338] = layer1_out[1911] | layer1_out[1912];
    assign layer2_out[5339] = ~(layer1_out[3906] | layer1_out[3907]);
    assign layer2_out[5340] = ~layer1_out[2889] | layer1_out[2888];
    assign layer2_out[5341] = layer1_out[326];
    assign layer2_out[5342] = layer1_out[2992];
    assign layer2_out[5343] = ~(layer1_out[1684] | layer1_out[1685]);
    assign layer2_out[5344] = layer1_out[154] & ~layer1_out[155];
    assign layer2_out[5345] = ~layer1_out[1273];
    assign layer2_out[5346] = ~layer1_out[6080];
    assign layer2_out[5347] = layer1_out[3074] & ~layer1_out[3073];
    assign layer2_out[5348] = ~layer1_out[7617];
    assign layer2_out[5349] = layer1_out[5440] & ~layer1_out[5439];
    assign layer2_out[5350] = ~(layer1_out[401] | layer1_out[402]);
    assign layer2_out[5351] = ~layer1_out[1522];
    assign layer2_out[5352] = ~layer1_out[1849];
    assign layer2_out[5353] = ~layer1_out[5114] | layer1_out[5115];
    assign layer2_out[5354] = layer1_out[7125];
    assign layer2_out[5355] = ~layer1_out[1722];
    assign layer2_out[5356] = ~layer1_out[6172] | layer1_out[6173];
    assign layer2_out[5357] = ~layer1_out[7636];
    assign layer2_out[5358] = ~(layer1_out[1767] | layer1_out[1768]);
    assign layer2_out[5359] = ~(layer1_out[7543] & layer1_out[7544]);
    assign layer2_out[5360] = ~layer1_out[3624];
    assign layer2_out[5361] = layer1_out[2641] & ~layer1_out[2642];
    assign layer2_out[5362] = ~(layer1_out[6991] | layer1_out[6992]);
    assign layer2_out[5363] = layer1_out[4304] | layer1_out[4305];
    assign layer2_out[5364] = layer1_out[4801];
    assign layer2_out[5365] = ~layer1_out[7248] | layer1_out[7247];
    assign layer2_out[5366] = ~layer1_out[20] | layer1_out[19];
    assign layer2_out[5367] = ~layer1_out[3239];
    assign layer2_out[5368] = 1'b0;
    assign layer2_out[5369] = ~layer1_out[4677] | layer1_out[4678];
    assign layer2_out[5370] = layer1_out[3567] & layer1_out[3568];
    assign layer2_out[5371] = layer1_out[7597];
    assign layer2_out[5372] = ~layer1_out[2023];
    assign layer2_out[5373] = ~layer1_out[4967] | layer1_out[4966];
    assign layer2_out[5374] = layer1_out[6233] & ~layer1_out[6232];
    assign layer2_out[5375] = 1'b0;
    assign layer2_out[5376] = layer1_out[1647];
    assign layer2_out[5377] = layer1_out[3541] & ~layer1_out[3540];
    assign layer2_out[5378] = ~(layer1_out[7657] | layer1_out[7658]);
    assign layer2_out[5379] = ~layer1_out[2001] | layer1_out[2000];
    assign layer2_out[5380] = ~layer1_out[3470];
    assign layer2_out[5381] = layer1_out[1727] & layer1_out[1728];
    assign layer2_out[5382] = ~(layer1_out[7326] & layer1_out[7327]);
    assign layer2_out[5383] = ~layer1_out[782];
    assign layer2_out[5384] = layer1_out[2116];
    assign layer2_out[5385] = ~layer1_out[389] | layer1_out[388];
    assign layer2_out[5386] = ~layer1_out[7519];
    assign layer2_out[5387] = layer1_out[6552];
    assign layer2_out[5388] = ~layer1_out[7445];
    assign layer2_out[5389] = ~layer1_out[1321] | layer1_out[1322];
    assign layer2_out[5390] = ~layer1_out[1791] | layer1_out[1790];
    assign layer2_out[5391] = ~layer1_out[2489];
    assign layer2_out[5392] = ~(layer1_out[5081] ^ layer1_out[5082]);
    assign layer2_out[5393] = ~(layer1_out[5753] & layer1_out[5754]);
    assign layer2_out[5394] = ~layer1_out[2025];
    assign layer2_out[5395] = layer1_out[1021] & ~layer1_out[1022];
    assign layer2_out[5396] = layer1_out[5409] & layer1_out[5410];
    assign layer2_out[5397] = layer1_out[6699] & ~layer1_out[6700];
    assign layer2_out[5398] = ~layer1_out[7488];
    assign layer2_out[5399] = layer1_out[6629] & ~layer1_out[6628];
    assign layer2_out[5400] = layer1_out[7886] & layer1_out[7887];
    assign layer2_out[5401] = layer1_out[5473] | layer1_out[5474];
    assign layer2_out[5402] = layer1_out[804] ^ layer1_out[805];
    assign layer2_out[5403] = layer1_out[6621];
    assign layer2_out[5404] = ~layer1_out[6275] | layer1_out[6274];
    assign layer2_out[5405] = ~layer1_out[2044];
    assign layer2_out[5406] = ~layer1_out[6802] | layer1_out[6801];
    assign layer2_out[5407] = layer1_out[4451] ^ layer1_out[4452];
    assign layer2_out[5408] = ~layer1_out[1423] | layer1_out[1424];
    assign layer2_out[5409] = ~layer1_out[2245];
    assign layer2_out[5410] = ~(layer1_out[7915] | layer1_out[7916]);
    assign layer2_out[5411] = layer1_out[1384];
    assign layer2_out[5412] = ~layer1_out[3928];
    assign layer2_out[5413] = layer1_out[3909];
    assign layer2_out[5414] = layer1_out[895];
    assign layer2_out[5415] = layer1_out[1486];
    assign layer2_out[5416] = layer1_out[2370] & ~layer1_out[2371];
    assign layer2_out[5417] = layer1_out[7909];
    assign layer2_out[5418] = layer1_out[549];
    assign layer2_out[5419] = ~layer1_out[7716] | layer1_out[7717];
    assign layer2_out[5420] = layer1_out[2205] | layer1_out[2206];
    assign layer2_out[5421] = layer1_out[627];
    assign layer2_out[5422] = ~layer1_out[1096] | layer1_out[1097];
    assign layer2_out[5423] = layer1_out[4853] & ~layer1_out[4852];
    assign layer2_out[5424] = ~layer1_out[7564];
    assign layer2_out[5425] = layer1_out[5179] & layer1_out[5180];
    assign layer2_out[5426] = layer1_out[7126];
    assign layer2_out[5427] = ~layer1_out[2625];
    assign layer2_out[5428] = layer1_out[1136];
    assign layer2_out[5429] = layer1_out[5508] & ~layer1_out[5509];
    assign layer2_out[5430] = ~(layer1_out[6112] ^ layer1_out[6113]);
    assign layer2_out[5431] = 1'b1;
    assign layer2_out[5432] = ~(layer1_out[1105] & layer1_out[1106]);
    assign layer2_out[5433] = layer1_out[7104];
    assign layer2_out[5434] = ~layer1_out[7487];
    assign layer2_out[5435] = layer1_out[4365];
    assign layer2_out[5436] = layer1_out[4446];
    assign layer2_out[5437] = layer1_out[469] & layer1_out[470];
    assign layer2_out[5438] = layer1_out[455];
    assign layer2_out[5439] = ~layer1_out[2803];
    assign layer2_out[5440] = layer1_out[2984] & ~layer1_out[2983];
    assign layer2_out[5441] = ~layer1_out[746];
    assign layer2_out[5442] = layer1_out[1912] | layer1_out[1913];
    assign layer2_out[5443] = ~layer1_out[731];
    assign layer2_out[5444] = ~layer1_out[6948];
    assign layer2_out[5445] = layer1_out[3104];
    assign layer2_out[5446] = ~layer1_out[7784];
    assign layer2_out[5447] = ~layer1_out[5092];
    assign layer2_out[5448] = ~layer1_out[5294];
    assign layer2_out[5449] = layer1_out[1476] | layer1_out[1477];
    assign layer2_out[5450] = layer1_out[3255] ^ layer1_out[3256];
    assign layer2_out[5451] = layer1_out[6846] & ~layer1_out[6847];
    assign layer2_out[5452] = ~layer1_out[206] | layer1_out[207];
    assign layer2_out[5453] = layer1_out[2079] ^ layer1_out[2080];
    assign layer2_out[5454] = layer1_out[1131];
    assign layer2_out[5455] = layer1_out[891];
    assign layer2_out[5456] = layer1_out[769] | layer1_out[770];
    assign layer2_out[5457] = layer1_out[3420] & ~layer1_out[3421];
    assign layer2_out[5458] = ~(layer1_out[950] ^ layer1_out[951]);
    assign layer2_out[5459] = layer1_out[258];
    assign layer2_out[5460] = ~layer1_out[4104];
    assign layer2_out[5461] = ~layer1_out[3644] | layer1_out[3643];
    assign layer2_out[5462] = layer1_out[1400] | layer1_out[1401];
    assign layer2_out[5463] = layer1_out[6164] & layer1_out[6165];
    assign layer2_out[5464] = layer1_out[3883] ^ layer1_out[3884];
    assign layer2_out[5465] = layer1_out[5233];
    assign layer2_out[5466] = 1'b1;
    assign layer2_out[5467] = layer1_out[3935];
    assign layer2_out[5468] = ~layer1_out[1613] | layer1_out[1614];
    assign layer2_out[5469] = layer1_out[1663] & ~layer1_out[1662];
    assign layer2_out[5470] = layer1_out[7985];
    assign layer2_out[5471] = 1'b0;
    assign layer2_out[5472] = layer1_out[4604] & ~layer1_out[4603];
    assign layer2_out[5473] = layer1_out[4622];
    assign layer2_out[5474] = layer1_out[1203];
    assign layer2_out[5475] = ~layer1_out[4216];
    assign layer2_out[5476] = ~layer1_out[1903] | layer1_out[1902];
    assign layer2_out[5477] = layer1_out[3889];
    assign layer2_out[5478] = layer1_out[6778] & layer1_out[6779];
    assign layer2_out[5479] = ~layer1_out[6318];
    assign layer2_out[5480] = ~layer1_out[7539];
    assign layer2_out[5481] = layer1_out[7802] & ~layer1_out[7801];
    assign layer2_out[5482] = ~(layer1_out[3152] | layer1_out[3153]);
    assign layer2_out[5483] = ~layer1_out[2527] | layer1_out[2528];
    assign layer2_out[5484] = ~layer1_out[5441];
    assign layer2_out[5485] = ~(layer1_out[1346] | layer1_out[1347]);
    assign layer2_out[5486] = 1'b0;
    assign layer2_out[5487] = ~(layer1_out[2262] | layer1_out[2263]);
    assign layer2_out[5488] = 1'b0;
    assign layer2_out[5489] = layer1_out[2106];
    assign layer2_out[5490] = layer1_out[2618] & layer1_out[2619];
    assign layer2_out[5491] = layer1_out[3078] | layer1_out[3079];
    assign layer2_out[5492] = ~layer1_out[1868] | layer1_out[1869];
    assign layer2_out[5493] = layer1_out[4088];
    assign layer2_out[5494] = ~layer1_out[4730];
    assign layer2_out[5495] = ~(layer1_out[3732] | layer1_out[3733]);
    assign layer2_out[5496] = layer1_out[1605];
    assign layer2_out[5497] = ~layer1_out[7734] | layer1_out[7735];
    assign layer2_out[5498] = ~layer1_out[844];
    assign layer2_out[5499] = ~layer1_out[721];
    assign layer2_out[5500] = layer1_out[7018];
    assign layer2_out[5501] = ~layer1_out[1346];
    assign layer2_out[5502] = layer1_out[6619] | layer1_out[6620];
    assign layer2_out[5503] = layer1_out[4281] & ~layer1_out[4280];
    assign layer2_out[5504] = ~(layer1_out[792] & layer1_out[793]);
    assign layer2_out[5505] = ~layer1_out[2913];
    assign layer2_out[5506] = ~layer1_out[121];
    assign layer2_out[5507] = ~layer1_out[969];
    assign layer2_out[5508] = layer1_out[5899];
    assign layer2_out[5509] = layer1_out[1856] | layer1_out[1857];
    assign layer2_out[5510] = layer1_out[6739] & ~layer1_out[6738];
    assign layer2_out[5511] = layer1_out[7561];
    assign layer2_out[5512] = layer1_out[3267];
    assign layer2_out[5513] = layer1_out[395] & ~layer1_out[394];
    assign layer2_out[5514] = layer1_out[490] | layer1_out[491];
    assign layer2_out[5515] = ~layer1_out[5308];
    assign layer2_out[5516] = layer1_out[5016] | layer1_out[5017];
    assign layer2_out[5517] = layer1_out[6320] & ~layer1_out[6321];
    assign layer2_out[5518] = ~layer1_out[2160];
    assign layer2_out[5519] = layer1_out[7147];
    assign layer2_out[5520] = layer1_out[6644] | layer1_out[6645];
    assign layer2_out[5521] = layer1_out[1947] & ~layer1_out[1948];
    assign layer2_out[5522] = layer1_out[1218];
    assign layer2_out[5523] = ~(layer1_out[1864] | layer1_out[1865]);
    assign layer2_out[5524] = layer1_out[2243];
    assign layer2_out[5525] = layer1_out[3494] & ~layer1_out[3495];
    assign layer2_out[5526] = ~layer1_out[802] | layer1_out[801];
    assign layer2_out[5527] = ~layer1_out[7987] | layer1_out[7986];
    assign layer2_out[5528] = layer1_out[666];
    assign layer2_out[5529] = layer1_out[531] & ~layer1_out[530];
    assign layer2_out[5530] = ~layer1_out[7210];
    assign layer2_out[5531] = ~layer1_out[686];
    assign layer2_out[5532] = ~layer1_out[6701];
    assign layer2_out[5533] = layer1_out[2839] | layer1_out[2840];
    assign layer2_out[5534] = ~(layer1_out[6757] ^ layer1_out[6758]);
    assign layer2_out[5535] = ~(layer1_out[2396] & layer1_out[2397]);
    assign layer2_out[5536] = layer1_out[806];
    assign layer2_out[5537] = 1'b1;
    assign layer2_out[5538] = layer1_out[1126] ^ layer1_out[1127];
    assign layer2_out[5539] = layer1_out[4565] & ~layer1_out[4566];
    assign layer2_out[5540] = layer1_out[3308] | layer1_out[3309];
    assign layer2_out[5541] = 1'b0;
    assign layer2_out[5542] = ~layer1_out[2957] | layer1_out[2956];
    assign layer2_out[5543] = layer1_out[5993];
    assign layer2_out[5544] = ~(layer1_out[2582] | layer1_out[2583]);
    assign layer2_out[5545] = ~layer1_out[2409];
    assign layer2_out[5546] = layer1_out[6584] & layer1_out[6585];
    assign layer2_out[5547] = ~layer1_out[7161];
    assign layer2_out[5548] = layer1_out[6505] | layer1_out[6506];
    assign layer2_out[5549] = ~layer1_out[6648];
    assign layer2_out[5550] = layer1_out[258] | layer1_out[259];
    assign layer2_out[5551] = ~layer1_out[779];
    assign layer2_out[5552] = layer1_out[307] & ~layer1_out[308];
    assign layer2_out[5553] = ~layer1_out[7113];
    assign layer2_out[5554] = ~(layer1_out[6858] | layer1_out[6859]);
    assign layer2_out[5555] = layer1_out[2748] & ~layer1_out[2747];
    assign layer2_out[5556] = 1'b1;
    assign layer2_out[5557] = ~(layer1_out[4893] | layer1_out[4894]);
    assign layer2_out[5558] = ~layer1_out[384];
    assign layer2_out[5559] = layer1_out[2454];
    assign layer2_out[5560] = ~(layer1_out[6029] ^ layer1_out[6030]);
    assign layer2_out[5561] = ~layer1_out[1990] | layer1_out[1989];
    assign layer2_out[5562] = layer1_out[1328] & ~layer1_out[1329];
    assign layer2_out[5563] = layer1_out[5356];
    assign layer2_out[5564] = ~(layer1_out[6711] | layer1_out[6712]);
    assign layer2_out[5565] = ~layer1_out[3720];
    assign layer2_out[5566] = 1'b0;
    assign layer2_out[5567] = ~layer1_out[7808];
    assign layer2_out[5568] = layer1_out[1301] & ~layer1_out[1302];
    assign layer2_out[5569] = layer1_out[4416] & layer1_out[4417];
    assign layer2_out[5570] = ~(layer1_out[7610] | layer1_out[7611]);
    assign layer2_out[5571] = ~(layer1_out[1503] | layer1_out[1504]);
    assign layer2_out[5572] = layer1_out[7049] | layer1_out[7050];
    assign layer2_out[5573] = ~layer1_out[6396] | layer1_out[6395];
    assign layer2_out[5574] = layer1_out[2147];
    assign layer2_out[5575] = ~layer1_out[3612];
    assign layer2_out[5576] = layer1_out[819];
    assign layer2_out[5577] = ~layer1_out[5645];
    assign layer2_out[5578] = ~layer1_out[5398];
    assign layer2_out[5579] = layer1_out[454];
    assign layer2_out[5580] = 1'b1;
    assign layer2_out[5581] = ~(layer1_out[477] | layer1_out[478]);
    assign layer2_out[5582] = ~(layer1_out[3302] ^ layer1_out[3303]);
    assign layer2_out[5583] = ~layer1_out[6291];
    assign layer2_out[5584] = layer1_out[1603];
    assign layer2_out[5585] = layer1_out[3688];
    assign layer2_out[5586] = layer1_out[4141];
    assign layer2_out[5587] = ~layer1_out[6065] | layer1_out[6064];
    assign layer2_out[5588] = layer1_out[2820] & layer1_out[2821];
    assign layer2_out[5589] = ~layer1_out[1501];
    assign layer2_out[5590] = layer1_out[1787] & layer1_out[1788];
    assign layer2_out[5591] = layer1_out[2934] & ~layer1_out[2933];
    assign layer2_out[5592] = ~layer1_out[370];
    assign layer2_out[5593] = layer1_out[1020] & ~layer1_out[1021];
    assign layer2_out[5594] = layer1_out[3318];
    assign layer2_out[5595] = ~(layer1_out[7531] & layer1_out[7532]);
    assign layer2_out[5596] = layer1_out[6996];
    assign layer2_out[5597] = layer1_out[1284];
    assign layer2_out[5598] = layer1_out[1992] & ~layer1_out[1991];
    assign layer2_out[5599] = layer1_out[176] & ~layer1_out[175];
    assign layer2_out[5600] = ~layer1_out[2788] | layer1_out[2789];
    assign layer2_out[5601] = layer1_out[4507] & ~layer1_out[4506];
    assign layer2_out[5602] = layer1_out[4698];
    assign layer2_out[5603] = layer1_out[6031];
    assign layer2_out[5604] = layer1_out[3148] & ~layer1_out[3147];
    assign layer2_out[5605] = ~layer1_out[5971];
    assign layer2_out[5606] = layer1_out[2157] | layer1_out[2158];
    assign layer2_out[5607] = layer1_out[2081] | layer1_out[2082];
    assign layer2_out[5608] = layer1_out[7524] & ~layer1_out[7525];
    assign layer2_out[5609] = ~layer1_out[2514];
    assign layer2_out[5610] = layer1_out[3313] & layer1_out[3314];
    assign layer2_out[5611] = ~layer1_out[5476] | layer1_out[5475];
    assign layer2_out[5612] = ~layer1_out[4664] | layer1_out[4665];
    assign layer2_out[5613] = layer1_out[3348];
    assign layer2_out[5614] = ~layer1_out[7311] | layer1_out[7312];
    assign layer2_out[5615] = ~(layer1_out[632] ^ layer1_out[633]);
    assign layer2_out[5616] = layer1_out[1542];
    assign layer2_out[5617] = layer1_out[1220] & ~layer1_out[1219];
    assign layer2_out[5618] = layer1_out[328] & ~layer1_out[327];
    assign layer2_out[5619] = ~(layer1_out[245] | layer1_out[246]);
    assign layer2_out[5620] = ~(layer1_out[1939] & layer1_out[1940]);
    assign layer2_out[5621] = 1'b1;
    assign layer2_out[5622] = ~layer1_out[795];
    assign layer2_out[5623] = layer1_out[561] & ~layer1_out[560];
    assign layer2_out[5624] = layer1_out[2082] & layer1_out[2083];
    assign layer2_out[5625] = ~layer1_out[6027];
    assign layer2_out[5626] = layer1_out[5223] & ~layer1_out[5224];
    assign layer2_out[5627] = layer1_out[1915] ^ layer1_out[1916];
    assign layer2_out[5628] = layer1_out[6734] & ~layer1_out[6733];
    assign layer2_out[5629] = ~(layer1_out[1364] & layer1_out[1365]);
    assign layer2_out[5630] = ~(layer1_out[4962] ^ layer1_out[4963]);
    assign layer2_out[5631] = ~(layer1_out[5902] & layer1_out[5903]);
    assign layer2_out[5632] = layer1_out[7200] & layer1_out[7201];
    assign layer2_out[5633] = layer1_out[3301];
    assign layer2_out[5634] = ~(layer1_out[957] | layer1_out[958]);
    assign layer2_out[5635] = layer1_out[2650];
    assign layer2_out[5636] = layer1_out[5176] & ~layer1_out[5177];
    assign layer2_out[5637] = ~layer1_out[1556];
    assign layer2_out[5638] = layer1_out[3886] & layer1_out[3887];
    assign layer2_out[5639] = ~(layer1_out[977] & layer1_out[978]);
    assign layer2_out[5640] = 1'b0;
    assign layer2_out[5641] = ~layer1_out[5117];
    assign layer2_out[5642] = layer1_out[3636];
    assign layer2_out[5643] = ~layer1_out[3444] | layer1_out[3443];
    assign layer2_out[5644] = layer1_out[5058];
    assign layer2_out[5645] = ~layer1_out[5935] | layer1_out[5934];
    assign layer2_out[5646] = layer1_out[5017] & ~layer1_out[5018];
    assign layer2_out[5647] = ~layer1_out[4831];
    assign layer2_out[5648] = ~layer1_out[778] | layer1_out[777];
    assign layer2_out[5649] = ~(layer1_out[2541] ^ layer1_out[2542]);
    assign layer2_out[5650] = ~(layer1_out[652] & layer1_out[653]);
    assign layer2_out[5651] = ~layer1_out[2002];
    assign layer2_out[5652] = ~layer1_out[5742];
    assign layer2_out[5653] = ~layer1_out[5211] | layer1_out[5212];
    assign layer2_out[5654] = layer1_out[735] | layer1_out[736];
    assign layer2_out[5655] = layer1_out[3407] & ~layer1_out[3408];
    assign layer2_out[5656] = ~layer1_out[3346];
    assign layer2_out[5657] = ~layer1_out[940] | layer1_out[941];
    assign layer2_out[5658] = ~(layer1_out[5405] ^ layer1_out[5406]);
    assign layer2_out[5659] = layer1_out[5654] ^ layer1_out[5655];
    assign layer2_out[5660] = layer1_out[34];
    assign layer2_out[5661] = ~layer1_out[7669];
    assign layer2_out[5662] = ~(layer1_out[5077] ^ layer1_out[5078]);
    assign layer2_out[5663] = ~(layer1_out[2531] | layer1_out[2532]);
    assign layer2_out[5664] = layer1_out[4271] | layer1_out[4272];
    assign layer2_out[5665] = layer1_out[6784] & ~layer1_out[6783];
    assign layer2_out[5666] = layer1_out[4689] ^ layer1_out[4690];
    assign layer2_out[5667] = 1'b1;
    assign layer2_out[5668] = layer1_out[4737] | layer1_out[4738];
    assign layer2_out[5669] = layer1_out[5883];
    assign layer2_out[5670] = layer1_out[1747] & layer1_out[1748];
    assign layer2_out[5671] = ~layer1_out[6641];
    assign layer2_out[5672] = layer1_out[4344] & ~layer1_out[4345];
    assign layer2_out[5673] = layer1_out[4307] & ~layer1_out[4308];
    assign layer2_out[5674] = ~(layer1_out[1180] ^ layer1_out[1181]);
    assign layer2_out[5675] = ~(layer1_out[7323] | layer1_out[7324]);
    assign layer2_out[5676] = layer1_out[5054] | layer1_out[5055];
    assign layer2_out[5677] = ~layer1_out[4341] | layer1_out[4342];
    assign layer2_out[5678] = ~(layer1_out[7647] | layer1_out[7648]);
    assign layer2_out[5679] = ~layer1_out[4689] | layer1_out[4688];
    assign layer2_out[5680] = layer1_out[7754] & ~layer1_out[7753];
    assign layer2_out[5681] = layer1_out[3496] & ~layer1_out[3495];
    assign layer2_out[5682] = ~layer1_out[4301] | layer1_out[4302];
    assign layer2_out[5683] = ~layer1_out[23] | layer1_out[22];
    assign layer2_out[5684] = ~layer1_out[540] | layer1_out[541];
    assign layer2_out[5685] = ~layer1_out[5769];
    assign layer2_out[5686] = ~layer1_out[5692];
    assign layer2_out[5687] = ~layer1_out[7156];
    assign layer2_out[5688] = ~layer1_out[574];
    assign layer2_out[5689] = layer1_out[6835] ^ layer1_out[6836];
    assign layer2_out[5690] = ~layer1_out[4104];
    assign layer2_out[5691] = layer1_out[842] & ~layer1_out[843];
    assign layer2_out[5692] = ~(layer1_out[2239] & layer1_out[2240]);
    assign layer2_out[5693] = layer1_out[4958];
    assign layer2_out[5694] = layer1_out[994] & ~layer1_out[995];
    assign layer2_out[5695] = ~layer1_out[6389];
    assign layer2_out[5696] = ~layer1_out[224] | layer1_out[225];
    assign layer2_out[5697] = layer1_out[474] | layer1_out[475];
    assign layer2_out[5698] = layer1_out[4883];
    assign layer2_out[5699] = ~(layer1_out[6039] & layer1_out[6040]);
    assign layer2_out[5700] = ~layer1_out[6382];
    assign layer2_out[5701] = ~layer1_out[1244];
    assign layer2_out[5702] = layer1_out[4721] & ~layer1_out[4722];
    assign layer2_out[5703] = layer1_out[2748] & layer1_out[2749];
    assign layer2_out[5704] = ~(layer1_out[5295] | layer1_out[5296]);
    assign layer2_out[5705] = layer1_out[3050] & ~layer1_out[3049];
    assign layer2_out[5706] = layer1_out[146] & ~layer1_out[145];
    assign layer2_out[5707] = layer1_out[287] & layer1_out[288];
    assign layer2_out[5708] = layer1_out[2347] & layer1_out[2348];
    assign layer2_out[5709] = ~layer1_out[3621];
    assign layer2_out[5710] = ~layer1_out[3951];
    assign layer2_out[5711] = ~layer1_out[5148] | layer1_out[5149];
    assign layer2_out[5712] = layer1_out[118] ^ layer1_out[119];
    assign layer2_out[5713] = ~layer1_out[5198] | layer1_out[5199];
    assign layer2_out[5714] = ~layer1_out[3608] | layer1_out[3607];
    assign layer2_out[5715] = ~(layer1_out[2730] ^ layer1_out[2731]);
    assign layer2_out[5716] = layer1_out[691] & layer1_out[692];
    assign layer2_out[5717] = layer1_out[4086] & ~layer1_out[4085];
    assign layer2_out[5718] = layer1_out[3172] ^ layer1_out[3173];
    assign layer2_out[5719] = ~layer1_out[4306] | layer1_out[4307];
    assign layer2_out[5720] = layer1_out[1405];
    assign layer2_out[5721] = ~(layer1_out[5215] ^ layer1_out[5216]);
    assign layer2_out[5722] = layer1_out[6556];
    assign layer2_out[5723] = layer1_out[4562] & ~layer1_out[4563];
    assign layer2_out[5724] = layer1_out[3206] & ~layer1_out[3207];
    assign layer2_out[5725] = ~(layer1_out[300] & layer1_out[301]);
    assign layer2_out[5726] = ~layer1_out[3116] | layer1_out[3115];
    assign layer2_out[5727] = layer1_out[7628] | layer1_out[7629];
    assign layer2_out[5728] = layer1_out[3538] & ~layer1_out[3539];
    assign layer2_out[5729] = ~(layer1_out[2494] & layer1_out[2495]);
    assign layer2_out[5730] = ~layer1_out[1901];
    assign layer2_out[5731] = ~(layer1_out[2211] & layer1_out[2212]);
    assign layer2_out[5732] = 1'b0;
    assign layer2_out[5733] = layer1_out[5567] & ~layer1_out[5568];
    assign layer2_out[5734] = ~layer1_out[6479] | layer1_out[6478];
    assign layer2_out[5735] = ~layer1_out[5027];
    assign layer2_out[5736] = ~(layer1_out[6273] & layer1_out[6274]);
    assign layer2_out[5737] = 1'b0;
    assign layer2_out[5738] = layer1_out[2981] & ~layer1_out[2982];
    assign layer2_out[5739] = layer1_out[727] & layer1_out[728];
    assign layer2_out[5740] = layer1_out[5479] & layer1_out[5480];
    assign layer2_out[5741] = layer1_out[2771];
    assign layer2_out[5742] = ~(layer1_out[3577] | layer1_out[3578]);
    assign layer2_out[5743] = ~layer1_out[2024] | layer1_out[2023];
    assign layer2_out[5744] = ~(layer1_out[7646] | layer1_out[7647]);
    assign layer2_out[5745] = layer1_out[2467] & layer1_out[2468];
    assign layer2_out[5746] = ~layer1_out[4291];
    assign layer2_out[5747] = ~layer1_out[7895] | layer1_out[7894];
    assign layer2_out[5748] = ~layer1_out[4865] | layer1_out[4864];
    assign layer2_out[5749] = layer1_out[2970] & ~layer1_out[2971];
    assign layer2_out[5750] = layer1_out[3244] & layer1_out[3245];
    assign layer2_out[5751] = 1'b0;
    assign layer2_out[5752] = ~layer1_out[6271];
    assign layer2_out[5753] = layer1_out[4378];
    assign layer2_out[5754] = ~layer1_out[1381] | layer1_out[1382];
    assign layer2_out[5755] = layer1_out[5797] & ~layer1_out[5798];
    assign layer2_out[5756] = ~(layer1_out[1877] | layer1_out[1878]);
    assign layer2_out[5757] = ~layer1_out[6760];
    assign layer2_out[5758] = layer1_out[2818] & ~layer1_out[2819];
    assign layer2_out[5759] = layer1_out[450] & ~layer1_out[451];
    assign layer2_out[5760] = 1'b1;
    assign layer2_out[5761] = ~layer1_out[3988];
    assign layer2_out[5762] = ~(layer1_out[710] | layer1_out[711]);
    assign layer2_out[5763] = ~layer1_out[6114] | layer1_out[6113];
    assign layer2_out[5764] = 1'b0;
    assign layer2_out[5765] = ~layer1_out[5695] | layer1_out[5694];
    assign layer2_out[5766] = ~layer1_out[3223] | layer1_out[3224];
    assign layer2_out[5767] = ~layer1_out[5071];
    assign layer2_out[5768] = layer1_out[3757] & layer1_out[3758];
    assign layer2_out[5769] = ~layer1_out[1046];
    assign layer2_out[5770] = layer1_out[1379];
    assign layer2_out[5771] = ~(layer1_out[675] | layer1_out[676]);
    assign layer2_out[5772] = layer1_out[3908] & layer1_out[3909];
    assign layer2_out[5773] = ~layer1_out[932];
    assign layer2_out[5774] = layer1_out[7414] & ~layer1_out[7413];
    assign layer2_out[5775] = ~layer1_out[7093];
    assign layer2_out[5776] = ~layer1_out[6138];
    assign layer2_out[5777] = layer1_out[7333] & ~layer1_out[7334];
    assign layer2_out[5778] = ~layer1_out[1380];
    assign layer2_out[5779] = layer1_out[3241] & layer1_out[3242];
    assign layer2_out[5780] = layer1_out[2911] & ~layer1_out[2910];
    assign layer2_out[5781] = layer1_out[3057] & ~layer1_out[3058];
    assign layer2_out[5782] = ~layer1_out[1434];
    assign layer2_out[5783] = ~layer1_out[7565];
    assign layer2_out[5784] = layer1_out[2109] & ~layer1_out[2110];
    assign layer2_out[5785] = layer1_out[4907] ^ layer1_out[4908];
    assign layer2_out[5786] = layer1_out[4390] & ~layer1_out[4389];
    assign layer2_out[5787] = ~layer1_out[3664] | layer1_out[3663];
    assign layer2_out[5788] = layer1_out[2830];
    assign layer2_out[5789] = ~layer1_out[1855] | layer1_out[1856];
    assign layer2_out[5790] = layer1_out[2199] | layer1_out[2200];
    assign layer2_out[5791] = ~layer1_out[6967];
    assign layer2_out[5792] = ~layer1_out[6750];
    assign layer2_out[5793] = layer1_out[5175];
    assign layer2_out[5794] = ~layer1_out[5902] | layer1_out[5901];
    assign layer2_out[5795] = layer1_out[6670] & layer1_out[6671];
    assign layer2_out[5796] = ~layer1_out[1874] | layer1_out[1875];
    assign layer2_out[5797] = layer1_out[7641] & layer1_out[7642];
    assign layer2_out[5798] = ~layer1_out[2440];
    assign layer2_out[5799] = layer1_out[4897] & layer1_out[4898];
    assign layer2_out[5800] = layer1_out[1265];
    assign layer2_out[5801] = layer1_out[5356] & ~layer1_out[5355];
    assign layer2_out[5802] = layer1_out[2505];
    assign layer2_out[5803] = ~(layer1_out[2212] & layer1_out[2213]);
    assign layer2_out[5804] = ~layer1_out[7323];
    assign layer2_out[5805] = ~layer1_out[2572];
    assign layer2_out[5806] = ~layer1_out[2257] | layer1_out[2258];
    assign layer2_out[5807] = 1'b1;
    assign layer2_out[5808] = layer1_out[7085] ^ layer1_out[7086];
    assign layer2_out[5809] = ~layer1_out[2781] | layer1_out[2780];
    assign layer2_out[5810] = layer1_out[6551];
    assign layer2_out[5811] = layer1_out[2706] | layer1_out[2707];
    assign layer2_out[5812] = ~layer1_out[95] | layer1_out[96];
    assign layer2_out[5813] = 1'b1;
    assign layer2_out[5814] = layer1_out[7133] & ~layer1_out[7134];
    assign layer2_out[5815] = layer1_out[3235] | layer1_out[3236];
    assign layer2_out[5816] = ~layer1_out[6735];
    assign layer2_out[5817] = ~(layer1_out[3442] & layer1_out[3443]);
    assign layer2_out[5818] = layer1_out[6018] & ~layer1_out[6019];
    assign layer2_out[5819] = ~(layer1_out[2616] & layer1_out[2617]);
    assign layer2_out[5820] = ~layer1_out[821] | layer1_out[822];
    assign layer2_out[5821] = ~(layer1_out[1376] | layer1_out[1377]);
    assign layer2_out[5822] = layer1_out[428] & ~layer1_out[429];
    assign layer2_out[5823] = ~layer1_out[4810] | layer1_out[4811];
    assign layer2_out[5824] = ~layer1_out[833] | layer1_out[834];
    assign layer2_out[5825] = ~layer1_out[3773];
    assign layer2_out[5826] = layer1_out[6085] & layer1_out[6086];
    assign layer2_out[5827] = ~(layer1_out[3199] | layer1_out[3200]);
    assign layer2_out[5828] = ~layer1_out[2096];
    assign layer2_out[5829] = layer1_out[1531];
    assign layer2_out[5830] = layer1_out[951];
    assign layer2_out[5831] = layer1_out[2758] & ~layer1_out[2757];
    assign layer2_out[5832] = ~(layer1_out[5129] & layer1_out[5130]);
    assign layer2_out[5833] = layer1_out[1070] & layer1_out[1071];
    assign layer2_out[5834] = layer1_out[2333];
    assign layer2_out[5835] = layer1_out[7333];
    assign layer2_out[5836] = layer1_out[7762];
    assign layer2_out[5837] = layer1_out[1397] & layer1_out[1398];
    assign layer2_out[5838] = 1'b0;
    assign layer2_out[5839] = ~layer1_out[6219] | layer1_out[6218];
    assign layer2_out[5840] = layer1_out[4421];
    assign layer2_out[5841] = layer1_out[5331] | layer1_out[5332];
    assign layer2_out[5842] = layer1_out[7557];
    assign layer2_out[5843] = ~layer1_out[2351];
    assign layer2_out[5844] = layer1_out[3676];
    assign layer2_out[5845] = layer1_out[4681];
    assign layer2_out[5846] = layer1_out[7857];
    assign layer2_out[5847] = layer1_out[5256];
    assign layer2_out[5848] = layer1_out[5763] & ~layer1_out[5762];
    assign layer2_out[5849] = layer1_out[6506];
    assign layer2_out[5850] = ~layer1_out[7578];
    assign layer2_out[5851] = ~layer1_out[7341] | layer1_out[7342];
    assign layer2_out[5852] = ~layer1_out[899];
    assign layer2_out[5853] = ~layer1_out[3059];
    assign layer2_out[5854] = ~(layer1_out[3176] | layer1_out[3177]);
    assign layer2_out[5855] = layer1_out[4505];
    assign layer2_out[5856] = layer1_out[5639] ^ layer1_out[5640];
    assign layer2_out[5857] = layer1_out[1844] | layer1_out[1845];
    assign layer2_out[5858] = ~(layer1_out[2634] & layer1_out[2635]);
    assign layer2_out[5859] = layer1_out[5299] & layer1_out[5300];
    assign layer2_out[5860] = layer1_out[2259];
    assign layer2_out[5861] = layer1_out[1225];
    assign layer2_out[5862] = ~(layer1_out[771] & layer1_out[772]);
    assign layer2_out[5863] = ~(layer1_out[2638] | layer1_out[2639]);
    assign layer2_out[5864] = layer1_out[614];
    assign layer2_out[5865] = layer1_out[4606] & ~layer1_out[4605];
    assign layer2_out[5866] = layer1_out[5166] | layer1_out[5167];
    assign layer2_out[5867] = ~layer1_out[2610];
    assign layer2_out[5868] = layer1_out[1234] | layer1_out[1235];
    assign layer2_out[5869] = ~layer1_out[4372] | layer1_out[4373];
    assign layer2_out[5870] = layer1_out[3538] & ~layer1_out[3537];
    assign layer2_out[5871] = layer1_out[2787];
    assign layer2_out[5872] = ~layer1_out[4812];
    assign layer2_out[5873] = ~(layer1_out[6544] ^ layer1_out[6545]);
    assign layer2_out[5874] = ~(layer1_out[1403] | layer1_out[1404]);
    assign layer2_out[5875] = ~layer1_out[5160];
    assign layer2_out[5876] = layer1_out[7497];
    assign layer2_out[5877] = 1'b0;
    assign layer2_out[5878] = ~(layer1_out[5217] | layer1_out[5218]);
    assign layer2_out[5879] = layer1_out[7132] & ~layer1_out[7131];
    assign layer2_out[5880] = layer1_out[2311] & layer1_out[2312];
    assign layer2_out[5881] = layer1_out[1007] & ~layer1_out[1008];
    assign layer2_out[5882] = ~layer1_out[6696];
    assign layer2_out[5883] = layer1_out[7621];
    assign layer2_out[5884] = layer1_out[2943];
    assign layer2_out[5885] = ~layer1_out[1007];
    assign layer2_out[5886] = ~layer1_out[1144];
    assign layer2_out[5887] = ~layer1_out[2310] | layer1_out[2309];
    assign layer2_out[5888] = ~layer1_out[5582];
    assign layer2_out[5889] = ~layer1_out[945];
    assign layer2_out[5890] = layer1_out[7318];
    assign layer2_out[5891] = ~(layer1_out[7146] & layer1_out[7147]);
    assign layer2_out[5892] = layer1_out[3010];
    assign layer2_out[5893] = layer1_out[7015];
    assign layer2_out[5894] = 1'b0;
    assign layer2_out[5895] = ~layer1_out[1578];
    assign layer2_out[5896] = ~(layer1_out[375] & layer1_out[376]);
    assign layer2_out[5897] = ~layer1_out[4620];
    assign layer2_out[5898] = layer1_out[3935] & ~layer1_out[3936];
    assign layer2_out[5899] = 1'b1;
    assign layer2_out[5900] = ~(layer1_out[2320] | layer1_out[2321]);
    assign layer2_out[5901] = layer1_out[7454];
    assign layer2_out[5902] = layer1_out[4055] & layer1_out[4056];
    assign layer2_out[5903] = ~layer1_out[6155];
    assign layer2_out[5904] = layer1_out[3164] & layer1_out[3165];
    assign layer2_out[5905] = ~layer1_out[4818];
    assign layer2_out[5906] = ~layer1_out[4782] | layer1_out[4783];
    assign layer2_out[5907] = ~(layer1_out[1003] & layer1_out[1004]);
    assign layer2_out[5908] = layer1_out[5572] & ~layer1_out[5571];
    assign layer2_out[5909] = layer1_out[4825] ^ layer1_out[4826];
    assign layer2_out[5910] = layer1_out[5695] & layer1_out[5696];
    assign layer2_out[5911] = layer1_out[1034];
    assign layer2_out[5912] = 1'b1;
    assign layer2_out[5913] = layer1_out[4485] & layer1_out[4486];
    assign layer2_out[5914] = layer1_out[6003] & layer1_out[6004];
    assign layer2_out[5915] = layer1_out[5714] ^ layer1_out[5715];
    assign layer2_out[5916] = layer1_out[6127] & ~layer1_out[6128];
    assign layer2_out[5917] = ~layer1_out[3986];
    assign layer2_out[5918] = ~layer1_out[56];
    assign layer2_out[5919] = layer1_out[2528];
    assign layer2_out[5920] = 1'b0;
    assign layer2_out[5921] = layer1_out[4850] & ~layer1_out[4851];
    assign layer2_out[5922] = ~layer1_out[6863];
    assign layer2_out[5923] = layer1_out[3134] | layer1_out[3135];
    assign layer2_out[5924] = ~layer1_out[6650] | layer1_out[6651];
    assign layer2_out[5925] = layer1_out[679];
    assign layer2_out[5926] = ~(layer1_out[2269] ^ layer1_out[2270]);
    assign layer2_out[5927] = ~(layer1_out[3488] | layer1_out[3489]);
    assign layer2_out[5928] = layer1_out[1937];
    assign layer2_out[5929] = ~(layer1_out[0] ^ layer1_out[2]);
    assign layer2_out[5930] = layer1_out[2653] & ~layer1_out[2652];
    assign layer2_out[5931] = ~layer1_out[4368];
    assign layer2_out[5932] = ~layer1_out[4132] | layer1_out[4131];
    assign layer2_out[5933] = layer1_out[7034];
    assign layer2_out[5934] = ~layer1_out[1961] | layer1_out[1960];
    assign layer2_out[5935] = ~layer1_out[7848] | layer1_out[7847];
    assign layer2_out[5936] = ~layer1_out[365];
    assign layer2_out[5937] = ~layer1_out[5681];
    assign layer2_out[5938] = ~layer1_out[2892];
    assign layer2_out[5939] = ~layer1_out[6532];
    assign layer2_out[5940] = ~layer1_out[5889];
    assign layer2_out[5941] = ~layer1_out[4614];
    assign layer2_out[5942] = layer1_out[5030] & layer1_out[5031];
    assign layer2_out[5943] = ~(layer1_out[5453] | layer1_out[5454]);
    assign layer2_out[5944] = ~layer1_out[2383];
    assign layer2_out[5945] = layer1_out[786];
    assign layer2_out[5946] = ~(layer1_out[1821] | layer1_out[1822]);
    assign layer2_out[5947] = ~layer1_out[5623];
    assign layer2_out[5948] = layer1_out[1675];
    assign layer2_out[5949] = ~layer1_out[5436] | layer1_out[5437];
    assign layer2_out[5950] = layer1_out[2055] & ~layer1_out[2056];
    assign layer2_out[5951] = layer1_out[1294] | layer1_out[1295];
    assign layer2_out[5952] = layer1_out[2294];
    assign layer2_out[5953] = ~layer1_out[1367];
    assign layer2_out[5954] = ~layer1_out[4340] | layer1_out[4341];
    assign layer2_out[5955] = ~layer1_out[6522];
    assign layer2_out[5956] = ~layer1_out[1706] | layer1_out[1707];
    assign layer2_out[5957] = layer1_out[4080] & ~layer1_out[4081];
    assign layer2_out[5958] = ~layer1_out[709];
    assign layer2_out[5959] = ~(layer1_out[6200] | layer1_out[6201]);
    assign layer2_out[5960] = ~layer1_out[7832];
    assign layer2_out[5961] = ~layer1_out[3650] | layer1_out[3649];
    assign layer2_out[5962] = layer1_out[6852] & ~layer1_out[6853];
    assign layer2_out[5963] = layer1_out[392];
    assign layer2_out[5964] = layer1_out[4577];
    assign layer2_out[5965] = layer1_out[6737];
    assign layer2_out[5966] = ~layer1_out[6324];
    assign layer2_out[5967] = ~layer1_out[5589];
    assign layer2_out[5968] = ~layer1_out[7851];
    assign layer2_out[5969] = ~layer1_out[2153];
    assign layer2_out[5970] = 1'b1;
    assign layer2_out[5971] = 1'b0;
    assign layer2_out[5972] = ~layer1_out[5084] | layer1_out[5085];
    assign layer2_out[5973] = ~layer1_out[7662] | layer1_out[7663];
    assign layer2_out[5974] = ~layer1_out[2308] | layer1_out[2307];
    assign layer2_out[5975] = ~(layer1_out[1264] & layer1_out[1265]);
    assign layer2_out[5976] = ~(layer1_out[5109] ^ layer1_out[5110]);
    assign layer2_out[5977] = ~layer1_out[5514] | layer1_out[5515];
    assign layer2_out[5978] = layer1_out[3694];
    assign layer2_out[5979] = layer1_out[6666] & ~layer1_out[6665];
    assign layer2_out[5980] = layer1_out[1865];
    assign layer2_out[5981] = ~layer1_out[6150];
    assign layer2_out[5982] = layer1_out[5478];
    assign layer2_out[5983] = layer1_out[5015];
    assign layer2_out[5984] = ~layer1_out[7942];
    assign layer2_out[5985] = layer1_out[7091];
    assign layer2_out[5986] = layer1_out[7202] | layer1_out[7203];
    assign layer2_out[5987] = ~layer1_out[5645];
    assign layer2_out[5988] = ~(layer1_out[23] | layer1_out[24]);
    assign layer2_out[5989] = ~layer1_out[1819];
    assign layer2_out[5990] = layer1_out[2440];
    assign layer2_out[5991] = layer1_out[1688] ^ layer1_out[1689];
    assign layer2_out[5992] = layer1_out[4055];
    assign layer2_out[5993] = 1'b0;
    assign layer2_out[5994] = layer1_out[3271];
    assign layer2_out[5995] = layer1_out[284];
    assign layer2_out[5996] = ~(layer1_out[6921] | layer1_out[6922]);
    assign layer2_out[5997] = ~layer1_out[7281];
    assign layer2_out[5998] = ~layer1_out[5053] | layer1_out[5052];
    assign layer2_out[5999] = layer1_out[3600];
    assign layer2_out[6000] = layer1_out[7937] & ~layer1_out[7938];
    assign layer2_out[6001] = layer1_out[3269] & layer1_out[3270];
    assign layer2_out[6002] = layer1_out[5387];
    assign layer2_out[6003] = ~(layer1_out[1230] | layer1_out[1231]);
    assign layer2_out[6004] = layer1_out[5608];
    assign layer2_out[6005] = layer1_out[468] | layer1_out[469];
    assign layer2_out[6006] = ~layer1_out[1920];
    assign layer2_out[6007] = ~layer1_out[5633];
    assign layer2_out[6008] = layer1_out[2744];
    assign layer2_out[6009] = ~layer1_out[582];
    assign layer2_out[6010] = ~layer1_out[1859] | layer1_out[1860];
    assign layer2_out[6011] = layer1_out[3292] & ~layer1_out[3293];
    assign layer2_out[6012] = ~(layer1_out[2374] & layer1_out[2375]);
    assign layer2_out[6013] = layer1_out[5588];
    assign layer2_out[6014] = layer1_out[3835] | layer1_out[3836];
    assign layer2_out[6015] = layer1_out[1211] & ~layer1_out[1212];
    assign layer2_out[6016] = ~(layer1_out[1428] | layer1_out[1429]);
    assign layer2_out[6017] = ~(layer1_out[1132] & layer1_out[1133]);
    assign layer2_out[6018] = ~(layer1_out[6984] & layer1_out[6985]);
    assign layer2_out[6019] = ~layer1_out[4640];
    assign layer2_out[6020] = layer1_out[7343];
    assign layer2_out[6021] = layer1_out[2009];
    assign layer2_out[6022] = layer1_out[6684];
    assign layer2_out[6023] = layer1_out[6511];
    assign layer2_out[6024] = ~layer1_out[2410];
    assign layer2_out[6025] = ~layer1_out[2949] | layer1_out[2948];
    assign layer2_out[6026] = ~layer1_out[3713];
    assign layer2_out[6027] = ~layer1_out[2980] | layer1_out[2981];
    assign layer2_out[6028] = layer1_out[7438] & ~layer1_out[7439];
    assign layer2_out[6029] = ~layer1_out[7288];
    assign layer2_out[6030] = ~layer1_out[2948];
    assign layer2_out[6031] = ~layer1_out[2238];
    assign layer2_out[6032] = ~(layer1_out[127] | layer1_out[128]);
    assign layer2_out[6033] = 1'b1;
    assign layer2_out[6034] = layer1_out[3403];
    assign layer2_out[6035] = ~(layer1_out[6109] | layer1_out[6110]);
    assign layer2_out[6036] = layer1_out[2451] & ~layer1_out[2452];
    assign layer2_out[6037] = ~layer1_out[6580];
    assign layer2_out[6038] = ~layer1_out[2758];
    assign layer2_out[6039] = ~(layer1_out[3731] ^ layer1_out[3732]);
    assign layer2_out[6040] = layer1_out[5466] & ~layer1_out[5467];
    assign layer2_out[6041] = ~(layer1_out[3257] & layer1_out[3258]);
    assign layer2_out[6042] = layer1_out[255];
    assign layer2_out[6043] = 1'b1;
    assign layer2_out[6044] = ~layer1_out[4298];
    assign layer2_out[6045] = layer1_out[650] & ~layer1_out[651];
    assign layer2_out[6046] = layer1_out[7081] & ~layer1_out[7080];
    assign layer2_out[6047] = layer1_out[1722] & ~layer1_out[1723];
    assign layer2_out[6048] = ~layer1_out[4581] | layer1_out[4580];
    assign layer2_out[6049] = ~(layer1_out[4530] ^ layer1_out[4531]);
    assign layer2_out[6050] = ~(layer1_out[3352] ^ layer1_out[3353]);
    assign layer2_out[6051] = ~(layer1_out[3404] & layer1_out[3405]);
    assign layer2_out[6052] = ~(layer1_out[3341] & layer1_out[3342]);
    assign layer2_out[6053] = layer1_out[4974];
    assign layer2_out[6054] = layer1_out[1456];
    assign layer2_out[6055] = ~layer1_out[5521] | layer1_out[5522];
    assign layer2_out[6056] = layer1_out[2460];
    assign layer2_out[6057] = layer1_out[6345] & ~layer1_out[6346];
    assign layer2_out[6058] = layer1_out[4402];
    assign layer2_out[6059] = ~layer1_out[439] | layer1_out[438];
    assign layer2_out[6060] = ~(layer1_out[1498] & layer1_out[1499]);
    assign layer2_out[6061] = layer1_out[4548] | layer1_out[4549];
    assign layer2_out[6062] = ~(layer1_out[4480] ^ layer1_out[4481]);
    assign layer2_out[6063] = ~(layer1_out[5201] & layer1_out[5202]);
    assign layer2_out[6064] = ~layer1_out[6834];
    assign layer2_out[6065] = ~(layer1_out[6948] & layer1_out[6949]);
    assign layer2_out[6066] = layer1_out[6958] & layer1_out[6959];
    assign layer2_out[6067] = ~layer1_out[2041] | layer1_out[2042];
    assign layer2_out[6068] = ~layer1_out[5803];
    assign layer2_out[6069] = layer1_out[6287] ^ layer1_out[6288];
    assign layer2_out[6070] = layer1_out[705];
    assign layer2_out[6071] = ~(layer1_out[5565] & layer1_out[5566]);
    assign layer2_out[6072] = layer1_out[5136] & ~layer1_out[5135];
    assign layer2_out[6073] = ~layer1_out[7534];
    assign layer2_out[6074] = ~(layer1_out[1665] ^ layer1_out[1666]);
    assign layer2_out[6075] = layer1_out[4596] & ~layer1_out[4597];
    assign layer2_out[6076] = ~(layer1_out[268] & layer1_out[269]);
    assign layer2_out[6077] = layer1_out[2533] ^ layer1_out[2534];
    assign layer2_out[6078] = ~layer1_out[7020] | layer1_out[7019];
    assign layer2_out[6079] = ~layer1_out[4639] | layer1_out[4640];
    assign layer2_out[6080] = layer1_out[4917];
    assign layer2_out[6081] = layer1_out[1209] & ~layer1_out[1210];
    assign layer2_out[6082] = layer1_out[688] & ~layer1_out[687];
    assign layer2_out[6083] = layer1_out[6354] & layer1_out[6355];
    assign layer2_out[6084] = ~(layer1_out[3730] & layer1_out[3731]);
    assign layer2_out[6085] = layer1_out[4765] | layer1_out[4766];
    assign layer2_out[6086] = ~(layer1_out[2237] & layer1_out[2238]);
    assign layer2_out[6087] = 1'b0;
    assign layer2_out[6088] = ~(layer1_out[5907] ^ layer1_out[5908]);
    assign layer2_out[6089] = layer1_out[7754];
    assign layer2_out[6090] = layer1_out[4779] & ~layer1_out[4778];
    assign layer2_out[6091] = ~layer1_out[973] | layer1_out[974];
    assign layer2_out[6092] = ~(layer1_out[4786] ^ layer1_out[4787]);
    assign layer2_out[6093] = ~layer1_out[6203];
    assign layer2_out[6094] = ~(layer1_out[2606] | layer1_out[2607]);
    assign layer2_out[6095] = layer1_out[3905] | layer1_out[3906];
    assign layer2_out[6096] = ~layer1_out[7665];
    assign layer2_out[6097] = layer1_out[3042] & ~layer1_out[3043];
    assign layer2_out[6098] = layer1_out[2817];
    assign layer2_out[6099] = ~layer1_out[4886];
    assign layer2_out[6100] = layer1_out[361];
    assign layer2_out[6101] = layer1_out[2705];
    assign layer2_out[6102] = layer1_out[2564];
    assign layer2_out[6103] = ~layer1_out[4892] | layer1_out[4893];
    assign layer2_out[6104] = layer1_out[6752];
    assign layer2_out[6105] = layer1_out[210] | layer1_out[211];
    assign layer2_out[6106] = ~layer1_out[4392] | layer1_out[4393];
    assign layer2_out[6107] = ~layer1_out[4277];
    assign layer2_out[6108] = layer1_out[698] & ~layer1_out[697];
    assign layer2_out[6109] = ~layer1_out[2813] | layer1_out[2814];
    assign layer2_out[6110] = layer1_out[3505];
    assign layer2_out[6111] = layer1_out[1517] & layer1_out[1518];
    assign layer2_out[6112] = layer1_out[7608];
    assign layer2_out[6113] = ~(layer1_out[4320] | layer1_out[4321]);
    assign layer2_out[6114] = 1'b0;
    assign layer2_out[6115] = layer1_out[5337] & ~layer1_out[5336];
    assign layer2_out[6116] = 1'b0;
    assign layer2_out[6117] = layer1_out[1926];
    assign layer2_out[6118] = ~(layer1_out[378] | layer1_out[379]);
    assign layer2_out[6119] = layer1_out[4144];
    assign layer2_out[6120] = layer1_out[5427] & ~layer1_out[5426];
    assign layer2_out[6121] = layer1_out[5701] | layer1_out[5702];
    assign layer2_out[6122] = 1'b1;
    assign layer2_out[6123] = ~(layer1_out[6352] & layer1_out[6353]);
    assign layer2_out[6124] = ~(layer1_out[249] | layer1_out[250]);
    assign layer2_out[6125] = ~(layer1_out[5037] ^ layer1_out[5038]);
    assign layer2_out[6126] = layer1_out[2126] ^ layer1_out[2127];
    assign layer2_out[6127] = layer1_out[5080] ^ layer1_out[5081];
    assign layer2_out[6128] = layer1_out[556] & layer1_out[557];
    assign layer2_out[6129] = ~(layer1_out[5507] & layer1_out[5508]);
    assign layer2_out[6130] = ~(layer1_out[6497] & layer1_out[6498]);
    assign layer2_out[6131] = 1'b0;
    assign layer2_out[6132] = layer1_out[348];
    assign layer2_out[6133] = ~(layer1_out[5744] ^ layer1_out[5745]);
    assign layer2_out[6134] = layer1_out[3015];
    assign layer2_out[6135] = ~(layer1_out[3394] | layer1_out[3395]);
    assign layer2_out[6136] = layer1_out[523];
    assign layer2_out[6137] = layer1_out[5249];
    assign layer2_out[6138] = ~layer1_out[1819];
    assign layer2_out[6139] = layer1_out[3834] & ~layer1_out[3835];
    assign layer2_out[6140] = ~(layer1_out[848] & layer1_out[849]);
    assign layer2_out[6141] = layer1_out[6548] | layer1_out[6549];
    assign layer2_out[6142] = ~layer1_out[7995];
    assign layer2_out[6143] = layer1_out[1869];
    assign layer2_out[6144] = layer1_out[1246] & layer1_out[1247];
    assign layer2_out[6145] = 1'b1;
    assign layer2_out[6146] = layer1_out[3722] & layer1_out[3723];
    assign layer2_out[6147] = ~layer1_out[4381];
    assign layer2_out[6148] = ~layer1_out[1221] | layer1_out[1222];
    assign layer2_out[6149] = layer1_out[4670];
    assign layer2_out[6150] = ~layer1_out[2865];
    assign layer2_out[6151] = ~layer1_out[5827];
    assign layer2_out[6152] = 1'b0;
    assign layer2_out[6153] = ~layer1_out[6126] | layer1_out[6127];
    assign layer2_out[6154] = layer1_out[4924];
    assign layer2_out[6155] = layer1_out[878] & ~layer1_out[879];
    assign layer2_out[6156] = layer1_out[7592] ^ layer1_out[7593];
    assign layer2_out[6157] = layer1_out[5474] | layer1_out[5475];
    assign layer2_out[6158] = layer1_out[5662] & ~layer1_out[5661];
    assign layer2_out[6159] = ~layer1_out[6139];
    assign layer2_out[6160] = ~layer1_out[7871];
    assign layer2_out[6161] = layer1_out[7597];
    assign layer2_out[6162] = layer1_out[6876] & ~layer1_out[6877];
    assign layer2_out[6163] = ~(layer1_out[5329] | layer1_out[5330]);
    assign layer2_out[6164] = layer1_out[6488];
    assign layer2_out[6165] = ~layer1_out[4715] | layer1_out[4714];
    assign layer2_out[6166] = ~layer1_out[1547];
    assign layer2_out[6167] = layer1_out[3601] ^ layer1_out[3602];
    assign layer2_out[6168] = layer1_out[686];
    assign layer2_out[6169] = ~(layer1_out[5939] ^ layer1_out[5940]);
    assign layer2_out[6170] = 1'b1;
    assign layer2_out[6171] = layer1_out[3641] | layer1_out[3642];
    assign layer2_out[6172] = 1'b1;
    assign layer2_out[6173] = ~layer1_out[6584] | layer1_out[6583];
    assign layer2_out[6174] = ~layer1_out[265];
    assign layer2_out[6175] = ~layer1_out[2430];
    assign layer2_out[6176] = 1'b0;
    assign layer2_out[6177] = 1'b1;
    assign layer2_out[6178] = layer1_out[1554];
    assign layer2_out[6179] = layer1_out[4289] ^ layer1_out[4290];
    assign layer2_out[6180] = layer1_out[2626] & layer1_out[2627];
    assign layer2_out[6181] = ~layer1_out[3738];
    assign layer2_out[6182] = 1'b1;
    assign layer2_out[6183] = ~(layer1_out[2792] & layer1_out[2793]);
    assign layer2_out[6184] = layer1_out[6562] & ~layer1_out[6563];
    assign layer2_out[6185] = 1'b1;
    assign layer2_out[6186] = ~layer1_out[5924];
    assign layer2_out[6187] = layer1_out[5576] | layer1_out[5577];
    assign layer2_out[6188] = ~layer1_out[7026];
    assign layer2_out[6189] = layer1_out[6088];
    assign layer2_out[6190] = layer1_out[3910] & layer1_out[3911];
    assign layer2_out[6191] = ~(layer1_out[1081] ^ layer1_out[1082]);
    assign layer2_out[6192] = ~layer1_out[6340];
    assign layer2_out[6193] = layer1_out[5011];
    assign layer2_out[6194] = ~layer1_out[4686];
    assign layer2_out[6195] = layer1_out[7705] & ~layer1_out[7704];
    assign layer2_out[6196] = layer1_out[302] & ~layer1_out[301];
    assign layer2_out[6197] = ~layer1_out[664];
    assign layer2_out[6198] = ~(layer1_out[3970] | layer1_out[3971]);
    assign layer2_out[6199] = layer1_out[2692] | layer1_out[2693];
    assign layer2_out[6200] = layer1_out[6557];
    assign layer2_out[6201] = layer1_out[1441];
    assign layer2_out[6202] = layer1_out[265] & ~layer1_out[264];
    assign layer2_out[6203] = layer1_out[1248];
    assign layer2_out[6204] = layer1_out[277];
    assign layer2_out[6205] = ~layer1_out[3287];
    assign layer2_out[6206] = layer1_out[6617] & layer1_out[6618];
    assign layer2_out[6207] = layer1_out[965] & ~layer1_out[966];
    assign layer2_out[6208] = ~layer1_out[1618] | layer1_out[1619];
    assign layer2_out[6209] = ~layer1_out[2444] | layer1_out[2443];
    assign layer2_out[6210] = ~(layer1_out[3933] | layer1_out[3934]);
    assign layer2_out[6211] = layer1_out[7677];
    assign layer2_out[6212] = layer1_out[7305];
    assign layer2_out[6213] = ~layer1_out[505];
    assign layer2_out[6214] = layer1_out[285] & layer1_out[286];
    assign layer2_out[6215] = layer1_out[6509];
    assign layer2_out[6216] = layer1_out[4020];
    assign layer2_out[6217] = layer1_out[5549] & ~layer1_out[5550];
    assign layer2_out[6218] = layer1_out[2750];
    assign layer2_out[6219] = ~layer1_out[4461] | layer1_out[4462];
    assign layer2_out[6220] = ~layer1_out[536] | layer1_out[537];
    assign layer2_out[6221] = 1'b1;
    assign layer2_out[6222] = ~layer1_out[6672] | layer1_out[6673];
    assign layer2_out[6223] = ~layer1_out[1733] | layer1_out[1734];
    assign layer2_out[6224] = ~layer1_out[672];
    assign layer2_out[6225] = 1'b0;
    assign layer2_out[6226] = 1'b0;
    assign layer2_out[6227] = ~(layer1_out[2065] | layer1_out[2066]);
    assign layer2_out[6228] = layer1_out[3626];
    assign layer2_out[6229] = layer1_out[2165];
    assign layer2_out[6230] = ~layer1_out[2953];
    assign layer2_out[6231] = ~(layer1_out[5113] & layer1_out[5114]);
    assign layer2_out[6232] = layer1_out[231];
    assign layer2_out[6233] = ~(layer1_out[7971] ^ layer1_out[7972]);
    assign layer2_out[6234] = layer1_out[3286] & ~layer1_out[3287];
    assign layer2_out[6235] = layer1_out[4491];
    assign layer2_out[6236] = layer1_out[7837];
    assign layer2_out[6237] = layer1_out[4369] | layer1_out[4370];
    assign layer2_out[6238] = ~(layer1_out[3868] ^ layer1_out[3869]);
    assign layer2_out[6239] = ~(layer1_out[1009] | layer1_out[1010]);
    assign layer2_out[6240] = ~layer1_out[435];
    assign layer2_out[6241] = ~(layer1_out[2398] | layer1_out[2399]);
    assign layer2_out[6242] = layer1_out[6836] & layer1_out[6837];
    assign layer2_out[6243] = layer1_out[4862];
    assign layer2_out[6244] = ~layer1_out[5282] | layer1_out[5283];
    assign layer2_out[6245] = ~layer1_out[2236];
    assign layer2_out[6246] = ~(layer1_out[7314] | layer1_out[7315]);
    assign layer2_out[6247] = ~layer1_out[6175];
    assign layer2_out[6248] = layer1_out[2347];
    assign layer2_out[6249] = ~layer1_out[634];
    assign layer2_out[6250] = ~(layer1_out[5147] ^ layer1_out[5148]);
    assign layer2_out[6251] = layer1_out[1587];
    assign layer2_out[6252] = layer1_out[966];
    assign layer2_out[6253] = 1'b0;
    assign layer2_out[6254] = layer1_out[6578];
    assign layer2_out[6255] = layer1_out[288] & ~layer1_out[289];
    assign layer2_out[6256] = ~layer1_out[5228];
    assign layer2_out[6257] = layer1_out[4379];
    assign layer2_out[6258] = layer1_out[3167] & layer1_out[3168];
    assign layer2_out[6259] = ~(layer1_out[2753] ^ layer1_out[2754]);
    assign layer2_out[6260] = ~(layer1_out[2234] | layer1_out[2235]);
    assign layer2_out[6261] = ~layer1_out[6527];
    assign layer2_out[6262] = ~layer1_out[3451];
    assign layer2_out[6263] = layer1_out[6479] | layer1_out[6480];
    assign layer2_out[6264] = ~(layer1_out[657] & layer1_out[658]);
    assign layer2_out[6265] = ~(layer1_out[6770] | layer1_out[6771]);
    assign layer2_out[6266] = layer1_out[6985] & ~layer1_out[6986];
    assign layer2_out[6267] = ~layer1_out[4630] | layer1_out[4631];
    assign layer2_out[6268] = ~layer1_out[6727];
    assign layer2_out[6269] = layer1_out[636] & ~layer1_out[635];
    assign layer2_out[6270] = ~layer1_out[7700] | layer1_out[7699];
    assign layer2_out[6271] = layer1_out[6406] & ~layer1_out[6407];
    assign layer2_out[6272] = ~(layer1_out[2120] ^ layer1_out[2121]);
    assign layer2_out[6273] = layer1_out[2273] & ~layer1_out[2274];
    assign layer2_out[6274] = layer1_out[6409] & layer1_out[6410];
    assign layer2_out[6275] = layer1_out[6874] | layer1_out[6875];
    assign layer2_out[6276] = ~layer1_out[7157];
    assign layer2_out[6277] = ~layer1_out[1432];
    assign layer2_out[6278] = layer1_out[3441];
    assign layer2_out[6279] = ~(layer1_out[2281] & layer1_out[2282]);
    assign layer2_out[6280] = ~layer1_out[2240];
    assign layer2_out[6281] = ~layer1_out[1391];
    assign layer2_out[6282] = ~(layer1_out[5761] | layer1_out[5762]);
    assign layer2_out[6283] = layer1_out[7513];
    assign layer2_out[6284] = layer1_out[1487] & ~layer1_out[1488];
    assign layer2_out[6285] = 1'b1;
    assign layer2_out[6286] = layer1_out[1276];
    assign layer2_out[6287] = ~(layer1_out[1083] | layer1_out[1084]);
    assign layer2_out[6288] = ~(layer1_out[986] | layer1_out[987]);
    assign layer2_out[6289] = layer1_out[2895] & ~layer1_out[2896];
    assign layer2_out[6290] = layer1_out[2490] ^ layer1_out[2491];
    assign layer2_out[6291] = ~layer1_out[437];
    assign layer2_out[6292] = layer1_out[4070];
    assign layer2_out[6293] = layer1_out[90] & ~layer1_out[89];
    assign layer2_out[6294] = ~layer1_out[7777];
    assign layer2_out[6295] = ~layer1_out[5881];
    assign layer2_out[6296] = layer1_out[7671] & ~layer1_out[7670];
    assign layer2_out[6297] = layer1_out[196];
    assign layer2_out[6298] = layer1_out[1422] ^ layer1_out[1423];
    assign layer2_out[6299] = layer1_out[7579];
    assign layer2_out[6300] = layer1_out[6519] & layer1_out[6520];
    assign layer2_out[6301] = ~(layer1_out[2229] & layer1_out[2230]);
    assign layer2_out[6302] = 1'b1;
    assign layer2_out[6303] = layer1_out[4781] ^ layer1_out[4782];
    assign layer2_out[6304] = layer1_out[2144];
    assign layer2_out[6305] = layer1_out[600];
    assign layer2_out[6306] = layer1_out[2178] & layer1_out[2179];
    assign layer2_out[6307] = ~layer1_out[2991];
    assign layer2_out[6308] = ~layer1_out[1137] | layer1_out[1136];
    assign layer2_out[6309] = ~(layer1_out[6890] & layer1_out[6891]);
    assign layer2_out[6310] = layer1_out[1098] | layer1_out[1099];
    assign layer2_out[6311] = layer1_out[2138];
    assign layer2_out[6312] = ~layer1_out[6381];
    assign layer2_out[6313] = 1'b1;
    assign layer2_out[6314] = ~(layer1_out[7098] ^ layer1_out[7099]);
    assign layer2_out[6315] = layer1_out[471] & ~layer1_out[470];
    assign layer2_out[6316] = ~layer1_out[7500];
    assign layer2_out[6317] = ~layer1_out[53] | layer1_out[52];
    assign layer2_out[6318] = layer1_out[2501];
    assign layer2_out[6319] = layer1_out[4701];
    assign layer2_out[6320] = 1'b0;
    assign layer2_out[6321] = ~(layer1_out[119] ^ layer1_out[120]);
    assign layer2_out[6322] = layer1_out[2147] & ~layer1_out[2148];
    assign layer2_out[6323] = layer1_out[2006] & ~layer1_out[2005];
    assign layer2_out[6324] = ~(layer1_out[6373] & layer1_out[6374]);
    assign layer2_out[6325] = layer1_out[2418];
    assign layer2_out[6326] = layer1_out[5879] | layer1_out[5880];
    assign layer2_out[6327] = ~layer1_out[3125];
    assign layer2_out[6328] = layer1_out[6165] | layer1_out[6166];
    assign layer2_out[6329] = layer1_out[4163];
    assign layer2_out[6330] = ~layer1_out[3520];
    assign layer2_out[6331] = layer1_out[2842];
    assign layer2_out[6332] = layer1_out[7792] ^ layer1_out[7793];
    assign layer2_out[6333] = layer1_out[1056] & ~layer1_out[1055];
    assign layer2_out[6334] = layer1_out[4824] | layer1_out[4825];
    assign layer2_out[6335] = ~layer1_out[5834] | layer1_out[5833];
    assign layer2_out[6336] = ~layer1_out[4872] | layer1_out[4871];
    assign layer2_out[6337] = ~layer1_out[2090];
    assign layer2_out[6338] = layer1_out[222] ^ layer1_out[223];
    assign layer2_out[6339] = 1'b0;
    assign layer2_out[6340] = ~layer1_out[7397];
    assign layer2_out[6341] = layer1_out[4713] & ~layer1_out[4714];
    assign layer2_out[6342] = ~(layer1_out[6255] & layer1_out[6256]);
    assign layer2_out[6343] = ~layer1_out[1652];
    assign layer2_out[6344] = ~(layer1_out[1746] | layer1_out[1747]);
    assign layer2_out[6345] = layer1_out[4225];
    assign layer2_out[6346] = layer1_out[1673] & ~layer1_out[1672];
    assign layer2_out[6347] = layer1_out[1718] | layer1_out[1719];
    assign layer2_out[6348] = layer1_out[896] & layer1_out[897];
    assign layer2_out[6349] = layer1_out[783];
    assign layer2_out[6350] = ~layer1_out[914];
    assign layer2_out[6351] = 1'b1;
    assign layer2_out[6352] = layer1_out[3151] | layer1_out[3152];
    assign layer2_out[6353] = layer1_out[5618] & layer1_out[5619];
    assign layer2_out[6354] = layer1_out[3259] & ~layer1_out[3260];
    assign layer2_out[6355] = ~layer1_out[1994];
    assign layer2_out[6356] = layer1_out[5060] & ~layer1_out[5061];
    assign layer2_out[6357] = layer1_out[4871];
    assign layer2_out[6358] = ~layer1_out[2296] | layer1_out[2297];
    assign layer2_out[6359] = ~layer1_out[4058];
    assign layer2_out[6360] = layer1_out[1796] | layer1_out[1797];
    assign layer2_out[6361] = layer1_out[1861];
    assign layer2_out[6362] = ~layer1_out[2119];
    assign layer2_out[6363] = ~(layer1_out[6769] & layer1_out[6770]);
    assign layer2_out[6364] = layer1_out[4054] & ~layer1_out[4053];
    assign layer2_out[6365] = layer1_out[546];
    assign layer2_out[6366] = ~(layer1_out[7989] & layer1_out[7990]);
    assign layer2_out[6367] = layer1_out[3465];
    assign layer2_out[6368] = ~(layer1_out[7974] | layer1_out[7975]);
    assign layer2_out[6369] = layer1_out[5783];
    assign layer2_out[6370] = layer1_out[1041];
    assign layer2_out[6371] = ~(layer1_out[1245] & layer1_out[1246]);
    assign layer2_out[6372] = layer1_out[4789];
    assign layer2_out[6373] = layer1_out[7493] & ~layer1_out[7494];
    assign layer2_out[6374] = ~layer1_out[6624] | layer1_out[6625];
    assign layer2_out[6375] = ~layer1_out[7555] | layer1_out[7554];
    assign layer2_out[6376] = 1'b0;
    assign layer2_out[6377] = layer1_out[2914];
    assign layer2_out[6378] = layer1_out[407];
    assign layer2_out[6379] = ~(layer1_out[5229] & layer1_out[5230]);
    assign layer2_out[6380] = layer1_out[2009] & layer1_out[2010];
    assign layer2_out[6381] = 1'b1;
    assign layer2_out[6382] = layer1_out[2547] & ~layer1_out[2546];
    assign layer2_out[6383] = ~(layer1_out[496] & layer1_out[497]);
    assign layer2_out[6384] = layer1_out[1038] | layer1_out[1039];
    assign layer2_out[6385] = layer1_out[962] & layer1_out[963];
    assign layer2_out[6386] = layer1_out[3431] | layer1_out[3432];
    assign layer2_out[6387] = layer1_out[1072] & layer1_out[1073];
    assign layer2_out[6388] = layer1_out[6468];
    assign layer2_out[6389] = layer1_out[1578] & layer1_out[1579];
    assign layer2_out[6390] = ~layer1_out[2822];
    assign layer2_out[6391] = ~layer1_out[6387];
    assign layer2_out[6392] = ~(layer1_out[7953] ^ layer1_out[7954]);
    assign layer2_out[6393] = layer1_out[5452] & layer1_out[5453];
    assign layer2_out[6394] = ~layer1_out[5890] | layer1_out[5891];
    assign layer2_out[6395] = layer1_out[2087];
    assign layer2_out[6396] = layer1_out[7245] & layer1_out[7246];
    assign layer2_out[6397] = layer1_out[4802] | layer1_out[4803];
    assign layer2_out[6398] = layer1_out[6896] ^ layer1_out[6897];
    assign layer2_out[6399] = layer1_out[2172];
    assign layer2_out[6400] = ~(layer1_out[5381] | layer1_out[5382]);
    assign layer2_out[6401] = layer1_out[3594] & ~layer1_out[3593];
    assign layer2_out[6402] = ~layer1_out[7929] | layer1_out[7930];
    assign layer2_out[6403] = ~(layer1_out[4156] & layer1_out[4157]);
    assign layer2_out[6404] = layer1_out[1909] | layer1_out[1910];
    assign layer2_out[6405] = ~layer1_out[4265] | layer1_out[4264];
    assign layer2_out[6406] = ~layer1_out[3335] | layer1_out[3336];
    assign layer2_out[6407] = ~layer1_out[4519];
    assign layer2_out[6408] = layer1_out[6794];
    assign layer2_out[6409] = layer1_out[6744];
    assign layer2_out[6410] = ~layer1_out[6292];
    assign layer2_out[6411] = layer1_out[230];
    assign layer2_out[6412] = layer1_out[6741];
    assign layer2_out[6413] = ~(layer1_out[807] & layer1_out[808]);
    assign layer2_out[6414] = layer1_out[3748] | layer1_out[3749];
    assign layer2_out[6415] = ~(layer1_out[5400] & layer1_out[5401]);
    assign layer2_out[6416] = layer1_out[2566] & layer1_out[2567];
    assign layer2_out[6417] = 1'b0;
    assign layer2_out[6418] = layer1_out[200] & ~layer1_out[201];
    assign layer2_out[6419] = layer1_out[3385] & ~layer1_out[3384];
    assign layer2_out[6420] = ~layer1_out[1153] | layer1_out[1154];
    assign layer2_out[6421] = ~layer1_out[6823];
    assign layer2_out[6422] = layer1_out[6297] & ~layer1_out[6296];
    assign layer2_out[6423] = layer1_out[2380];
    assign layer2_out[6424] = ~layer1_out[7007];
    assign layer2_out[6425] = ~layer1_out[6707];
    assign layer2_out[6426] = layer1_out[128] ^ layer1_out[129];
    assign layer2_out[6427] = ~(layer1_out[7132] & layer1_out[7133]);
    assign layer2_out[6428] = layer1_out[4666] & ~layer1_out[4667];
    assign layer2_out[6429] = ~layer1_out[2387];
    assign layer2_out[6430] = ~layer1_out[84] | layer1_out[83];
    assign layer2_out[6431] = 1'b1;
    assign layer2_out[6432] = ~layer1_out[495];
    assign layer2_out[6433] = ~layer1_out[7106];
    assign layer2_out[6434] = ~(layer1_out[2679] ^ layer1_out[2680]);
    assign layer2_out[6435] = layer1_out[2433] ^ layer1_out[2434];
    assign layer2_out[6436] = layer1_out[3140] & ~layer1_out[3139];
    assign layer2_out[6437] = layer1_out[1765];
    assign layer2_out[6438] = layer1_out[7766];
    assign layer2_out[6439] = ~(layer1_out[7805] | layer1_out[7806]);
    assign layer2_out[6440] = layer1_out[5226] & ~layer1_out[5225];
    assign layer2_out[6441] = ~layer1_out[1888];
    assign layer2_out[6442] = layer1_out[2755];
    assign layer2_out[6443] = ~layer1_out[4046];
    assign layer2_out[6444] = ~layer1_out[7464] | layer1_out[7463];
    assign layer2_out[6445] = ~(layer1_out[1017] ^ layer1_out[1018]);
    assign layer2_out[6446] = layer1_out[5760] & layer1_out[5761];
    assign layer2_out[6447] = ~(layer1_out[2121] & layer1_out[2122]);
    assign layer2_out[6448] = ~layer1_out[7561];
    assign layer2_out[6449] = ~layer1_out[1210];
    assign layer2_out[6450] = ~layer1_out[464];
    assign layer2_out[6451] = ~(layer1_out[2219] | layer1_out[2220]);
    assign layer2_out[6452] = layer1_out[2741];
    assign layer2_out[6453] = layer1_out[7582];
    assign layer2_out[6454] = layer1_out[7188] & ~layer1_out[7189];
    assign layer2_out[6455] = 1'b1;
    assign layer2_out[6456] = ~layer1_out[624];
    assign layer2_out[6457] = layer1_out[858];
    assign layer2_out[6458] = ~layer1_out[3813];
    assign layer2_out[6459] = ~layer1_out[6277] | layer1_out[6276];
    assign layer2_out[6460] = layer1_out[7435] & layer1_out[7436];
    assign layer2_out[6461] = layer1_out[5145] ^ layer1_out[5146];
    assign layer2_out[6462] = layer1_out[5357] | layer1_out[5358];
    assign layer2_out[6463] = ~layer1_out[2573];
    assign layer2_out[6464] = ~layer1_out[3792] | layer1_out[3793];
    assign layer2_out[6465] = layer1_out[3572] | layer1_out[3573];
    assign layer2_out[6466] = ~layer1_out[4594];
    assign layer2_out[6467] = layer1_out[4624];
    assign layer2_out[6468] = ~(layer1_out[1088] & layer1_out[1089]);
    assign layer2_out[6469] = layer1_out[6494] & ~layer1_out[6493];
    assign layer2_out[6470] = layer1_out[6923];
    assign layer2_out[6471] = layer1_out[5945];
    assign layer2_out[6472] = layer1_out[5403] & ~layer1_out[5402];
    assign layer2_out[6473] = layer1_out[1466];
    assign layer2_out[6474] = layer1_out[2900] | layer1_out[2901];
    assign layer2_out[6475] = layer1_out[4040] | layer1_out[4041];
    assign layer2_out[6476] = layer1_out[3316] ^ layer1_out[3317];
    assign layer2_out[6477] = ~layer1_out[3583];
    assign layer2_out[6478] = ~layer1_out[270];
    assign layer2_out[6479] = ~layer1_out[2318] | layer1_out[2319];
    assign layer2_out[6480] = ~layer1_out[3775];
    assign layer2_out[6481] = ~layer1_out[4704];
    assign layer2_out[6482] = ~layer1_out[2867] | layer1_out[2866];
    assign layer2_out[6483] = ~layer1_out[2387];
    assign layer2_out[6484] = layer1_out[1703] & ~layer1_out[1704];
    assign layer2_out[6485] = layer1_out[5274] & ~layer1_out[5273];
    assign layer2_out[6486] = ~layer1_out[502];
    assign layer2_out[6487] = layer1_out[3658] & ~layer1_out[3657];
    assign layer2_out[6488] = ~layer1_out[3785] | layer1_out[3784];
    assign layer2_out[6489] = layer1_out[5123];
    assign layer2_out[6490] = ~layer1_out[3192] | layer1_out[3193];
    assign layer2_out[6491] = layer1_out[3068] ^ layer1_out[3069];
    assign layer2_out[6492] = layer1_out[6521] & ~layer1_out[6520];
    assign layer2_out[6493] = ~layer1_out[2561];
    assign layer2_out[6494] = ~layer1_out[4850] | layer1_out[4849];
    assign layer2_out[6495] = layer1_out[7213] | layer1_out[7214];
    assign layer2_out[6496] = ~(layer1_out[4005] & layer1_out[4006]);
    assign layer2_out[6497] = ~layer1_out[5507] | layer1_out[5506];
    assign layer2_out[6498] = ~layer1_out[5345];
    assign layer2_out[6499] = ~layer1_out[518];
    assign layer2_out[6500] = ~(layer1_out[140] ^ layer1_out[141]);
    assign layer2_out[6501] = layer1_out[6439];
    assign layer2_out[6502] = ~layer1_out[7824];
    assign layer2_out[6503] = layer1_out[5847];
    assign layer2_out[6504] = layer1_out[4335] & ~layer1_out[4336];
    assign layer2_out[6505] = layer1_out[69] & layer1_out[70];
    assign layer2_out[6506] = ~(layer1_out[887] & layer1_out[888]);
    assign layer2_out[6507] = ~layer1_out[5060] | layer1_out[5059];
    assign layer2_out[6508] = layer1_out[5570] | layer1_out[5571];
    assign layer2_out[6509] = ~layer1_out[1754] | layer1_out[1753];
    assign layer2_out[6510] = ~(layer1_out[317] | layer1_out[318]);
    assign layer2_out[6511] = layer1_out[5967] & ~layer1_out[5966];
    assign layer2_out[6512] = ~(layer1_out[3752] & layer1_out[3753]);
    assign layer2_out[6513] = ~layer1_out[6019] | layer1_out[6020];
    assign layer2_out[6514] = layer1_out[2153];
    assign layer2_out[6515] = ~layer1_out[6689];
    assign layer2_out[6516] = 1'b0;
    assign layer2_out[6517] = layer1_out[4232] ^ layer1_out[4233];
    assign layer2_out[6518] = ~(layer1_out[1165] ^ layer1_out[1166]);
    assign layer2_out[6519] = ~(layer1_out[1075] | layer1_out[1076]);
    assign layer2_out[6520] = layer1_out[7349];
    assign layer2_out[6521] = ~layer1_out[6683];
    assign layer2_out[6522] = ~layer1_out[1931];
    assign layer2_out[6523] = 1'b0;
    assign layer2_out[6524] = layer1_out[3416];
    assign layer2_out[6525] = ~layer1_out[2467];
    assign layer2_out[6526] = ~layer1_out[5542] | layer1_out[5541];
    assign layer2_out[6527] = layer1_out[700] & layer1_out[701];
    assign layer2_out[6528] = layer1_out[3788] & layer1_out[3789];
    assign layer2_out[6529] = layer1_out[5010] ^ layer1_out[5011];
    assign layer2_out[6530] = layer1_out[486];
    assign layer2_out[6531] = layer1_out[1907];
    assign layer2_out[6532] = layer1_out[6887] & ~layer1_out[6888];
    assign layer2_out[6533] = layer1_out[677];
    assign layer2_out[6534] = ~layer1_out[7470] | layer1_out[7469];
    assign layer2_out[6535] = layer1_out[267];
    assign layer2_out[6536] = ~(layer1_out[7035] | layer1_out[7036]);
    assign layer2_out[6537] = layer1_out[5471] & ~layer1_out[5472];
    assign layer2_out[6538] = ~layer1_out[796] | layer1_out[795];
    assign layer2_out[6539] = ~(layer1_out[7076] | layer1_out[7077]);
    assign layer2_out[6540] = ~layer1_out[7164] | layer1_out[7163];
    assign layer2_out[6541] = ~layer1_out[175] | layer1_out[174];
    assign layer2_out[6542] = layer1_out[6421] & ~layer1_out[6420];
    assign layer2_out[6543] = layer1_out[5170];
    assign layer2_out[6544] = layer1_out[6447];
    assign layer2_out[6545] = layer1_out[4725] | layer1_out[4726];
    assign layer2_out[6546] = layer1_out[2294];
    assign layer2_out[6547] = ~layer1_out[3484];
    assign layer2_out[6548] = ~(layer1_out[681] | layer1_out[682]);
    assign layer2_out[6549] = layer1_out[500] & ~layer1_out[501];
    assign layer2_out[6550] = layer1_out[2441] ^ layer1_out[2442];
    assign layer2_out[6551] = ~layer1_out[1674];
    assign layer2_out[6552] = ~layer1_out[7187];
    assign layer2_out[6553] = layer1_out[7389] & layer1_out[7390];
    assign layer2_out[6554] = ~layer1_out[7086];
    assign layer2_out[6555] = ~layer1_out[1735];
    assign layer2_out[6556] = layer1_out[2442];
    assign layer2_out[6557] = layer1_out[6981];
    assign layer2_out[6558] = layer1_out[6393];
    assign layer2_out[6559] = ~layer1_out[7890];
    assign layer2_out[6560] = layer1_out[495] ^ layer1_out[496];
    assign layer2_out[6561] = ~layer1_out[7344];
    assign layer2_out[6562] = ~(layer1_out[5945] | layer1_out[5946]);
    assign layer2_out[6563] = layer1_out[6075] | layer1_out[6076];
    assign layer2_out[6564] = ~(layer1_out[6241] | layer1_out[6242]);
    assign layer2_out[6565] = 1'b0;
    assign layer2_out[6566] = layer1_out[1755];
    assign layer2_out[6567] = layer1_out[7419] & ~layer1_out[7418];
    assign layer2_out[6568] = ~layer1_out[6474] | layer1_out[6475];
    assign layer2_out[6569] = layer1_out[6024];
    assign layer2_out[6570] = layer1_out[374] & ~layer1_out[373];
    assign layer2_out[6571] = layer1_out[4837] & layer1_out[4838];
    assign layer2_out[6572] = layer1_out[7375];
    assign layer2_out[6573] = layer1_out[4033] & layer1_out[4034];
    assign layer2_out[6574] = layer1_out[1893] | layer1_out[1894];
    assign layer2_out[6575] = layer1_out[7573];
    assign layer2_out[6576] = layer1_out[2807];
    assign layer2_out[6577] = layer1_out[7097];
    assign layer2_out[6578] = layer1_out[6133] & layer1_out[6134];
    assign layer2_out[6579] = ~(layer1_out[6375] | layer1_out[6376]);
    assign layer2_out[6580] = layer1_out[6379];
    assign layer2_out[6581] = ~layer1_out[5747] | layer1_out[5746];
    assign layer2_out[6582] = ~(layer1_out[7269] | layer1_out[7270]);
    assign layer2_out[6583] = layer1_out[1151];
    assign layer2_out[6584] = ~layer1_out[17] | layer1_out[18];
    assign layer2_out[6585] = layer1_out[71] | layer1_out[72];
    assign layer2_out[6586] = ~(layer1_out[3454] & layer1_out[3455]);
    assign layer2_out[6587] = ~(layer1_out[2133] ^ layer1_out[2134]);
    assign layer2_out[6588] = layer1_out[7141] & ~layer1_out[7140];
    assign layer2_out[6589] = ~layer1_out[4066];
    assign layer2_out[6590] = layer1_out[381];
    assign layer2_out[6591] = layer1_out[2096];
    assign layer2_out[6592] = ~(layer1_out[892] | layer1_out[893]);
    assign layer2_out[6593] = layer1_out[4458];
    assign layer2_out[6594] = layer1_out[107] | layer1_out[108];
    assign layer2_out[6595] = ~layer1_out[5484] | layer1_out[5485];
    assign layer2_out[6596] = ~layer1_out[3468];
    assign layer2_out[6597] = ~layer1_out[262];
    assign layer2_out[6598] = layer1_out[467];
    assign layer2_out[6599] = layer1_out[736];
    assign layer2_out[6600] = layer1_out[3520] & layer1_out[3521];
    assign layer2_out[6601] = ~(layer1_out[6091] | layer1_out[6092]);
    assign layer2_out[6602] = ~(layer1_out[551] ^ layer1_out[552]);
    assign layer2_out[6603] = ~(layer1_out[5100] & layer1_out[5101]);
    assign layer2_out[6604] = layer1_out[568] ^ layer1_out[569];
    assign layer2_out[6605] = layer1_out[6636] | layer1_out[6637];
    assign layer2_out[6606] = ~layer1_out[7654];
    assign layer2_out[6607] = ~(layer1_out[4250] & layer1_out[4251]);
    assign layer2_out[6608] = ~layer1_out[2074];
    assign layer2_out[6609] = layer1_out[2488] & ~layer1_out[2487];
    assign layer2_out[6610] = ~layer1_out[7708] | layer1_out[7709];
    assign layer2_out[6611] = ~(layer1_out[3446] & layer1_out[3447]);
    assign layer2_out[6612] = layer1_out[1741] & layer1_out[1742];
    assign layer2_out[6613] = ~(layer1_out[3201] ^ layer1_out[3202]);
    assign layer2_out[6614] = layer1_out[196];
    assign layer2_out[6615] = ~(layer1_out[4706] ^ layer1_out[4707]);
    assign layer2_out[6616] = ~layer1_out[6871];
    assign layer2_out[6617] = layer1_out[6636] & ~layer1_out[6635];
    assign layer2_out[6618] = ~(layer1_out[7295] | layer1_out[7296]);
    assign layer2_out[6619] = ~(layer1_out[6973] & layer1_out[6974]);
    assign layer2_out[6620] = ~(layer1_out[2569] | layer1_out[2570]);
    assign layer2_out[6621] = 1'b0;
    assign layer2_out[6622] = layer1_out[5323] & ~layer1_out[5322];
    assign layer2_out[6623] = ~layer1_out[5407];
    assign layer2_out[6624] = layer1_out[1017] & ~layer1_out[1016];
    assign layer2_out[6625] = ~layer1_out[1861];
    assign layer2_out[6626] = layer1_out[3113] & ~layer1_out[3112];
    assign layer2_out[6627] = ~layer1_out[5255] | layer1_out[5254];
    assign layer2_out[6628] = ~layer1_out[1331] | layer1_out[1330];
    assign layer2_out[6629] = ~layer1_out[6268] | layer1_out[6269];
    assign layer2_out[6630] = ~layer1_out[6048];
    assign layer2_out[6631] = layer1_out[2904];
    assign layer2_out[6632] = layer1_out[3787] ^ layer1_out[3788];
    assign layer2_out[6633] = ~layer1_out[2880];
    assign layer2_out[6634] = layer1_out[305];
    assign layer2_out[6635] = layer1_out[6716] ^ layer1_out[6717];
    assign layer2_out[6636] = ~(layer1_out[7602] ^ layer1_out[7603]);
    assign layer2_out[6637] = ~layer1_out[5702];
    assign layer2_out[6638] = layer1_out[1310];
    assign layer2_out[6639] = ~layer1_out[3018] | layer1_out[3017];
    assign layer2_out[6640] = layer1_out[5024];
    assign layer2_out[6641] = ~layer1_out[5794] | layer1_out[5793];
    assign layer2_out[6642] = layer1_out[2788];
    assign layer2_out[6643] = layer1_out[6942] | layer1_out[6943];
    assign layer2_out[6644] = ~layer1_out[7372];
    assign layer2_out[6645] = layer1_out[2127] & layer1_out[2128];
    assign layer2_out[6646] = 1'b0;
    assign layer2_out[6647] = ~(layer1_out[2057] | layer1_out[2058]);
    assign layer2_out[6648] = ~(layer1_out[7501] & layer1_out[7502]);
    assign layer2_out[6649] = layer1_out[7241] & layer1_out[7242];
    assign layer2_out[6650] = layer1_out[3205] & ~layer1_out[3206];
    assign layer2_out[6651] = layer1_out[6945];
    assign layer2_out[6652] = ~(layer1_out[2352] & layer1_out[2353]);
    assign layer2_out[6653] = ~layer1_out[3965];
    assign layer2_out[6654] = layer1_out[7991] | layer1_out[7992];
    assign layer2_out[6655] = ~layer1_out[7958];
    assign layer2_out[6656] = ~(layer1_out[2129] ^ layer1_out[2130]);
    assign layer2_out[6657] = ~(layer1_out[6831] & layer1_out[6832]);
    assign layer2_out[6658] = ~layer1_out[4195];
    assign layer2_out[6659] = layer1_out[6730] | layer1_out[6731];
    assign layer2_out[6660] = layer1_out[112];
    assign layer2_out[6661] = layer1_out[591];
    assign layer2_out[6662] = ~layer1_out[6782];
    assign layer2_out[6663] = ~layer1_out[7711];
    assign layer2_out[6664] = ~layer1_out[6818] | layer1_out[6817];
    assign layer2_out[6665] = ~(layer1_out[2617] ^ layer1_out[2618]);
    assign layer2_out[6666] = layer1_out[2404];
    assign layer2_out[6667] = layer1_out[6610] & ~layer1_out[6609];
    assign layer2_out[6668] = layer1_out[4646] | layer1_out[4647];
    assign layer2_out[6669] = ~layer1_out[1590] | layer1_out[1591];
    assign layer2_out[6670] = 1'b1;
    assign layer2_out[6671] = layer1_out[7590] & layer1_out[7591];
    assign layer2_out[6672] = layer1_out[7569] & layer1_out[7570];
    assign layer2_out[6673] = layer1_out[1145] & layer1_out[1146];
    assign layer2_out[6674] = layer1_out[4266] ^ layer1_out[4267];
    assign layer2_out[6675] = layer1_out[4078] & layer1_out[4079];
    assign layer2_out[6676] = layer1_out[90] & layer1_out[91];
    assign layer2_out[6677] = ~(layer1_out[7363] ^ layer1_out[7364]);
    assign layer2_out[6678] = ~layer1_out[3042];
    assign layer2_out[6679] = layer1_out[4328];
    assign layer2_out[6680] = ~(layer1_out[762] ^ layer1_out[763]);
    assign layer2_out[6681] = ~(layer1_out[332] ^ layer1_out[333]);
    assign layer2_out[6682] = layer1_out[5743] ^ layer1_out[5744];
    assign layer2_out[6683] = layer1_out[1014] & layer1_out[1015];
    assign layer2_out[6684] = ~layer1_out[3535];
    assign layer2_out[6685] = layer1_out[397];
    assign layer2_out[6686] = ~layer1_out[7119];
    assign layer2_out[6687] = layer1_out[7968];
    assign layer2_out[6688] = layer1_out[4653] | layer1_out[4654];
    assign layer2_out[6689] = ~(layer1_out[1723] & layer1_out[1724]);
    assign layer2_out[6690] = ~(layer1_out[4035] ^ layer1_out[4036]);
    assign layer2_out[6691] = layer1_out[7822];
    assign layer2_out[6692] = layer1_out[5415] | layer1_out[5416];
    assign layer2_out[6693] = layer1_out[4822];
    assign layer2_out[6694] = layer1_out[4736] & ~layer1_out[4735];
    assign layer2_out[6695] = ~layer1_out[5168] | layer1_out[5169];
    assign layer2_out[6696] = layer1_out[3914] & ~layer1_out[3913];
    assign layer2_out[6697] = layer1_out[6005] & ~layer1_out[6004];
    assign layer2_out[6698] = ~layer1_out[7492];
    assign layer2_out[6699] = layer1_out[963] ^ layer1_out[964];
    assign layer2_out[6700] = layer1_out[6163];
    assign layer2_out[6701] = ~(layer1_out[1532] & layer1_out[1533]);
    assign layer2_out[6702] = ~(layer1_out[3938] & layer1_out[3939]);
    assign layer2_out[6703] = ~layer1_out[5314];
    assign layer2_out[6704] = ~layer1_out[3716] | layer1_out[3717];
    assign layer2_out[6705] = ~layer1_out[1229] | layer1_out[1228];
    assign layer2_out[6706] = layer1_out[6070] | layer1_out[6071];
    assign layer2_out[6707] = layer1_out[2163];
    assign layer2_out[6708] = ~(layer1_out[5802] & layer1_out[5803]);
    assign layer2_out[6709] = layer1_out[7386] & layer1_out[7387];
    assign layer2_out[6710] = ~layer1_out[773] | layer1_out[772];
    assign layer2_out[6711] = ~(layer1_out[2908] ^ layer1_out[2909]);
    assign layer2_out[6712] = ~layer1_out[2156];
    assign layer2_out[6713] = layer1_out[5554];
    assign layer2_out[6714] = 1'b0;
    assign layer2_out[6715] = layer1_out[5478] | layer1_out[5479];
    assign layer2_out[6716] = layer1_out[291];
    assign layer2_out[6717] = layer1_out[1530];
    assign layer2_out[6718] = ~layer1_out[3551];
    assign layer2_out[6719] = layer1_out[1500];
    assign layer2_out[6720] = layer1_out[2760] & layer1_out[2761];
    assign layer2_out[6721] = layer1_out[5133];
    assign layer2_out[6722] = layer1_out[4382];
    assign layer2_out[6723] = layer1_out[2010] & ~layer1_out[2011];
    assign layer2_out[6724] = layer1_out[2392];
    assign layer2_out[6725] = ~(layer1_out[4200] | layer1_out[4201]);
    assign layer2_out[6726] = layer1_out[275];
    assign layer2_out[6727] = 1'b1;
    assign layer2_out[6728] = ~(layer1_out[5773] ^ layer1_out[5774]);
    assign layer2_out[6729] = 1'b1;
    assign layer2_out[6730] = ~layer1_out[1852];
    assign layer2_out[6731] = ~(layer1_out[7267] | layer1_out[7268]);
    assign layer2_out[6732] = ~layer1_out[632];
    assign layer2_out[6733] = layer1_out[5448] & ~layer1_out[5449];
    assign layer2_out[6734] = layer1_out[7099];
    assign layer2_out[6735] = layer1_out[6307] & layer1_out[6308];
    assign layer2_out[6736] = ~(layer1_out[4152] ^ layer1_out[4153]);
    assign layer2_out[6737] = ~layer1_out[595] | layer1_out[594];
    assign layer2_out[6738] = ~(layer1_out[5394] ^ layer1_out[5395]);
    assign layer2_out[6739] = layer1_out[5814] & ~layer1_out[5815];
    assign layer2_out[6740] = ~(layer1_out[7082] | layer1_out[7083]);
    assign layer2_out[6741] = layer1_out[1682];
    assign layer2_out[6742] = layer1_out[3417] & ~layer1_out[3418];
    assign layer2_out[6743] = ~layer1_out[6842];
    assign layer2_out[6744] = layer1_out[3984] | layer1_out[3985];
    assign layer2_out[6745] = layer1_out[4822] & ~layer1_out[4821];
    assign layer2_out[6746] = layer1_out[6010];
    assign layer2_out[6747] = layer1_out[7982];
    assign layer2_out[6748] = layer1_out[5209];
    assign layer2_out[6749] = ~layer1_out[4052] | layer1_out[4053];
    assign layer2_out[6750] = ~layer1_out[5144];
    assign layer2_out[6751] = layer1_out[3003];
    assign layer2_out[6752] = 1'b1;
    assign layer2_out[6753] = ~layer1_out[6561];
    assign layer2_out[6754] = 1'b1;
    assign layer2_out[6755] = layer1_out[5620];
    assign layer2_out[6756] = ~(layer1_out[4375] & layer1_out[4376]);
    assign layer2_out[6757] = layer1_out[2071];
    assign layer2_out[6758] = layer1_out[2184] & ~layer1_out[2183];
    assign layer2_out[6759] = ~layer1_out[3050] | layer1_out[3051];
    assign layer2_out[6760] = layer1_out[4205];
    assign layer2_out[6761] = layer1_out[2932] & layer1_out[2933];
    assign layer2_out[6762] = layer1_out[1446] & ~layer1_out[1447];
    assign layer2_out[6763] = ~layer1_out[6267] | layer1_out[6268];
    assign layer2_out[6764] = layer1_out[1656];
    assign layer2_out[6765] = ~layer1_out[6510] | layer1_out[6509];
    assign layer2_out[6766] = layer1_out[1535];
    assign layer2_out[6767] = ~layer1_out[4669];
    assign layer2_out[6768] = ~layer1_out[4023];
    assign layer2_out[6769] = layer1_out[6412] & layer1_out[6413];
    assign layer2_out[6770] = layer1_out[6502];
    assign layer2_out[6771] = ~(layer1_out[4727] & layer1_out[4728]);
    assign layer2_out[6772] = ~(layer1_out[4293] | layer1_out[4294]);
    assign layer2_out[6773] = layer1_out[1833] | layer1_out[1834];
    assign layer2_out[6774] = layer1_out[4300] & ~layer1_out[4301];
    assign layer2_out[6775] = layer1_out[5995];
    assign layer2_out[6776] = ~layer1_out[6299] | layer1_out[6298];
    assign layer2_out[6777] = layer1_out[4538];
    assign layer2_out[6778] = ~layer1_out[3393] | layer1_out[3392];
    assign layer2_out[6779] = ~(layer1_out[5451] ^ layer1_out[5452]);
    assign layer2_out[6780] = ~layer1_out[3434] | layer1_out[3433];
    assign layer2_out[6781] = ~layer1_out[7688] | layer1_out[7687];
    assign layer2_out[6782] = ~layer1_out[2723];
    assign layer2_out[6783] = layer1_out[5247] ^ layer1_out[5248];
    assign layer2_out[6784] = ~layer1_out[3870] | layer1_out[3871];
    assign layer2_out[6785] = layer1_out[7243] & ~layer1_out[7242];
    assign layer2_out[6786] = layer1_out[1351];
    assign layer2_out[6787] = layer1_out[3450];
    assign layer2_out[6788] = ~(layer1_out[6411] | layer1_out[6412]);
    assign layer2_out[6789] = ~(layer1_out[7535] | layer1_out[7536]);
    assign layer2_out[6790] = layer1_out[5724] | layer1_out[5725];
    assign layer2_out[6791] = layer1_out[7107] & layer1_out[7108];
    assign layer2_out[6792] = layer1_out[5365] & ~layer1_out[5364];
    assign layer2_out[6793] = ~layer1_out[7039];
    assign layer2_out[6794] = layer1_out[87] & ~layer1_out[86];
    assign layer2_out[6795] = layer1_out[3401] | layer1_out[3402];
    assign layer2_out[6796] = ~layer1_out[1972];
    assign layer2_out[6797] = ~layer1_out[2361] | layer1_out[2362];
    assign layer2_out[6798] = ~layer1_out[1575];
    assign layer2_out[6799] = ~layer1_out[7301];
    assign layer2_out[6800] = layer1_out[2767] | layer1_out[2768];
    assign layer2_out[6801] = layer1_out[2397] ^ layer1_out[2398];
    assign layer2_out[6802] = ~layer1_out[1980];
    assign layer2_out[6803] = layer1_out[4662];
    assign layer2_out[6804] = layer1_out[7355] | layer1_out[7356];
    assign layer2_out[6805] = ~layer1_out[3411] | layer1_out[3410];
    assign layer2_out[6806] = layer1_out[7789];
    assign layer2_out[6807] = ~(layer1_out[3705] & layer1_out[3706]);
    assign layer2_out[6808] = layer1_out[5740] | layer1_out[5741];
    assign layer2_out[6809] = layer1_out[7779] & ~layer1_out[7778];
    assign layer2_out[6810] = layer1_out[3974] | layer1_out[3975];
    assign layer2_out[6811] = layer1_out[2384] | layer1_out[2385];
    assign layer2_out[6812] = ~(layer1_out[3493] ^ layer1_out[3494]);
    assign layer2_out[6813] = layer1_out[3008];
    assign layer2_out[6814] = ~layer1_out[1538] | layer1_out[1539];
    assign layer2_out[6815] = layer1_out[828] & layer1_out[829];
    assign layer2_out[6816] = layer1_out[2451] & ~layer1_out[2450];
    assign layer2_out[6817] = ~layer1_out[6699] | layer1_out[6698];
    assign layer2_out[6818] = ~layer1_out[6171] | layer1_out[6170];
    assign layer2_out[6819] = 1'b0;
    assign layer2_out[6820] = ~layer1_out[2425];
    assign layer2_out[6821] = layer1_out[3948] & ~layer1_out[3947];
    assign layer2_out[6822] = ~layer1_out[5909] | layer1_out[5908];
    assign layer2_out[6823] = ~layer1_out[4581] | layer1_out[4582];
    assign layer2_out[6824] = ~(layer1_out[1996] & layer1_out[1997]);
    assign layer2_out[6825] = ~layer1_out[2131];
    assign layer2_out[6826] = layer1_out[1633];
    assign layer2_out[6827] = layer1_out[6309];
    assign layer2_out[6828] = ~layer1_out[58];
    assign layer2_out[6829] = 1'b1;
    assign layer2_out[6830] = ~layer1_out[190] | layer1_out[189];
    assign layer2_out[6831] = ~(layer1_out[2801] | layer1_out[2802]);
    assign layer2_out[6832] = layer1_out[7568] ^ layer1_out[7569];
    assign layer2_out[6833] = layer1_out[2794] & layer1_out[2795];
    assign layer2_out[6834] = layer1_out[4139];
    assign layer2_out[6835] = layer1_out[4834];
    assign layer2_out[6836] = layer1_out[1275] | layer1_out[1276];
    assign layer2_out[6837] = layer1_out[976] & ~layer1_out[977];
    assign layer2_out[6838] = ~layer1_out[1459];
    assign layer2_out[6839] = ~(layer1_out[2132] & layer1_out[2133]);
    assign layer2_out[6840] = layer1_out[3233];
    assign layer2_out[6841] = ~layer1_out[3932] | layer1_out[3931];
    assign layer2_out[6842] = ~layer1_out[1704];
    assign layer2_out[6843] = layer1_out[7844] & ~layer1_out[7845];
    assign layer2_out[6844] = ~layer1_out[7383];
    assign layer2_out[6845] = ~layer1_out[2069] | layer1_out[2070];
    assign layer2_out[6846] = layer1_out[3123] & layer1_out[3124];
    assign layer2_out[6847] = layer1_out[3695];
    assign layer2_out[6848] = layer1_out[7894];
    assign layer2_out[6849] = layer1_out[352];
    assign layer2_out[6850] = ~layer1_out[5382];
    assign layer2_out[6851] = layer1_out[2445] | layer1_out[2446];
    assign layer2_out[6852] = ~layer1_out[4829] | layer1_out[4830];
    assign layer2_out[6853] = ~(layer1_out[955] & layer1_out[956]);
    assign layer2_out[6854] = layer1_out[1975] | layer1_out[1976];
    assign layer2_out[6855] = layer1_out[4510] & ~layer1_out[4511];
    assign layer2_out[6856] = ~(layer1_out[3378] & layer1_out[3379]);
    assign layer2_out[6857] = layer1_out[1453] | layer1_out[1454];
    assign layer2_out[6858] = 1'b0;
    assign layer2_out[6859] = layer1_out[7784];
    assign layer2_out[6860] = ~layer1_out[5028] | layer1_out[5029];
    assign layer2_out[6861] = ~(layer1_out[2117] ^ layer1_out[2118]);
    assign layer2_out[6862] = layer1_out[6100];
    assign layer2_out[6863] = ~(layer1_out[6652] ^ layer1_out[6653]);
    assign layer2_out[6864] = ~layer1_out[2278] | layer1_out[2277];
    assign layer2_out[6865] = layer1_out[7913];
    assign layer2_out[6866] = layer1_out[5563] & ~layer1_out[5562];
    assign layer2_out[6867] = ~(layer1_out[2899] & layer1_out[2900]);
    assign layer2_out[6868] = layer1_out[749] & layer1_out[750];
    assign layer2_out[6869] = layer1_out[4759] ^ layer1_out[4760];
    assign layer2_out[6870] = layer1_out[7128] | layer1_out[7129];
    assign layer2_out[6871] = ~layer1_out[7296];
    assign layer2_out[6872] = ~layer1_out[5195];
    assign layer2_out[6873] = layer1_out[4800];
    assign layer2_out[6874] = ~layer1_out[7166] | layer1_out[7165];
    assign layer2_out[6875] = layer1_out[6975];
    assign layer2_out[6876] = ~layer1_out[3005];
    assign layer2_out[6877] = ~(layer1_out[3921] | layer1_out[3922]);
    assign layer2_out[6878] = ~layer1_out[5208] | layer1_out[5207];
    assign layer2_out[6879] = ~layer1_out[5595] | layer1_out[5596];
    assign layer2_out[6880] = ~layer1_out[3719];
    assign layer2_out[6881] = ~layer1_out[3291] | layer1_out[3290];
    assign layer2_out[6882] = layer1_out[3943];
    assign layer2_out[6883] = layer1_out[1166];
    assign layer2_out[6884] = ~(layer1_out[2456] & layer1_out[2457]);
    assign layer2_out[6885] = ~(layer1_out[2897] ^ layer1_out[2898]);
    assign layer2_out[6886] = layer1_out[1675] & ~layer1_out[1676];
    assign layer2_out[6887] = layer1_out[4532] | layer1_out[4533];
    assign layer2_out[6888] = ~layer1_out[2056];
    assign layer2_out[6889] = layer1_out[5328] & ~layer1_out[5327];
    assign layer2_out[6890] = layer1_out[263] | layer1_out[264];
    assign layer2_out[6891] = ~(layer1_out[290] ^ layer1_out[291]);
    assign layer2_out[6892] = layer1_out[1419];
    assign layer2_out[6893] = layer1_out[5560];
    assign layer2_out[6894] = layer1_out[6883];
    assign layer2_out[6895] = ~layer1_out[359];
    assign layer2_out[6896] = layer1_out[2217] ^ layer1_out[2218];
    assign layer2_out[6897] = ~layer1_out[2018];
    assign layer2_out[6898] = layer1_out[924] & ~layer1_out[925];
    assign layer2_out[6899] = layer1_out[898];
    assign layer2_out[6900] = layer1_out[4898];
    assign layer2_out[6901] = layer1_out[5982] & ~layer1_out[5983];
    assign layer2_out[6902] = layer1_out[7630];
    assign layer2_out[6903] = layer1_out[6147];
    assign layer2_out[6904] = layer1_out[3054];
    assign layer2_out[6905] = layer1_out[4612];
    assign layer2_out[6906] = layer1_out[6523] & layer1_out[6524];
    assign layer2_out[6907] = layer1_out[4260] & ~layer1_out[4261];
    assign layer2_out[6908] = layer1_out[1695] & ~layer1_out[1696];
    assign layer2_out[6909] = ~layer1_out[306] | layer1_out[307];
    assign layer2_out[6910] = layer1_out[670];
    assign layer2_out[6911] = layer1_out[4353];
    assign layer2_out[6912] = layer1_out[1515];
    assign layer2_out[6913] = ~layer1_out[7273] | layer1_out[7274];
    assign layer2_out[6914] = ~layer1_out[5275];
    assign layer2_out[6915] = layer1_out[2077] & layer1_out[2078];
    assign layer2_out[6916] = ~layer1_out[5278];
    assign layer2_out[6917] = layer1_out[3398] | layer1_out[3399];
    assign layer2_out[6918] = layer1_out[3356] & ~layer1_out[3357];
    assign layer2_out[6919] = layer1_out[5861] & ~layer1_out[5860];
    assign layer2_out[6920] = layer1_out[851] ^ layer1_out[852];
    assign layer2_out[6921] = ~layer1_out[338];
    assign layer2_out[6922] = layer1_out[6829];
    assign layer2_out[6923] = layer1_out[1800] & ~layer1_out[1801];
    assign layer2_out[6924] = ~(layer1_out[7254] | layer1_out[7255]);
    assign layer2_out[6925] = ~layer1_out[7835];
    assign layer2_out[6926] = layer1_out[6351] | layer1_out[6352];
    assign layer2_out[6927] = ~(layer1_out[6558] & layer1_out[6559]);
    assign layer2_out[6928] = ~(layer1_out[5517] ^ layer1_out[5518]);
    assign layer2_out[6929] = ~layer1_out[409] | layer1_out[408];
    assign layer2_out[6930] = ~layer1_out[6819] | layer1_out[6820];
    assign layer2_out[6931] = layer1_out[3440];
    assign layer2_out[6932] = ~layer1_out[2145];
    assign layer2_out[6933] = layer1_out[5413] & ~layer1_out[5414];
    assign layer2_out[6934] = layer1_out[3250] & layer1_out[3251];
    assign layer2_out[6935] = ~layer1_out[1798];
    assign layer2_out[6936] = layer1_out[6962];
    assign layer2_out[6937] = ~layer1_out[7526] | layer1_out[7527];
    assign layer2_out[6938] = ~layer1_out[6452];
    assign layer2_out[6939] = layer1_out[7724] & ~layer1_out[7723];
    assign layer2_out[6940] = ~layer1_out[2327];
    assign layer2_out[6941] = layer1_out[1484] ^ layer1_out[1485];
    assign layer2_out[6942] = ~layer1_out[6378];
    assign layer2_out[6943] = ~layer1_out[1043];
    assign layer2_out[6944] = ~layer1_out[5335];
    assign layer2_out[6945] = ~layer1_out[2791] | layer1_out[2790];
    assign layer2_out[6946] = ~layer1_out[3095];
    assign layer2_out[6947] = layer1_out[7838] & layer1_out[7839];
    assign layer2_out[6948] = layer1_out[5004];
    assign layer2_out[6949] = layer1_out[5383] & ~layer1_out[5384];
    assign layer2_out[6950] = layer1_out[637] & ~layer1_out[636];
    assign layer2_out[6951] = ~(layer1_out[4127] ^ layer1_out[4128]);
    assign layer2_out[6952] = ~(layer1_out[2600] ^ layer1_out[2601]);
    assign layer2_out[6953] = ~layer1_out[1138];
    assign layer2_out[6954] = ~layer1_out[774];
    assign layer2_out[6955] = ~(layer1_out[2314] & layer1_out[2315]);
    assign layer2_out[6956] = layer1_out[7044];
    assign layer2_out[6957] = 1'b1;
    assign layer2_out[6958] = layer1_out[4042];
    assign layer2_out[6959] = ~layer1_out[5090] | layer1_out[5091];
    assign layer2_out[6960] = ~layer1_out[3973] | layer1_out[3974];
    assign layer2_out[6961] = ~layer1_out[1788];
    assign layer2_out[6962] = ~layer1_out[2475];
    assign layer2_out[6963] = layer1_out[6100] ^ layer1_out[6101];
    assign layer2_out[6964] = ~layer1_out[6549];
    assign layer2_out[6965] = layer1_out[2553] & layer1_out[2554];
    assign layer2_out[6966] = layer1_out[7756] | layer1_out[7757];
    assign layer2_out[6967] = ~layer1_out[3726];
    assign layer2_out[6968] = ~layer1_out[1493];
    assign layer2_out[6969] = layer1_out[1559] & ~layer1_out[1558];
    assign layer2_out[6970] = layer1_out[3353] & ~layer1_out[3354];
    assign layer2_out[6971] = layer1_out[5529];
    assign layer2_out[6972] = ~layer1_out[2037];
    assign layer2_out[6973] = 1'b0;
    assign layer2_out[6974] = ~layer1_out[2011] | layer1_out[2012];
    assign layer2_out[6975] = ~(layer1_out[7905] & layer1_out[7906]);
    assign layer2_out[6976] = layer1_out[4599];
    assign layer2_out[6977] = ~(layer1_out[4171] ^ layer1_out[4172]);
    assign layer2_out[6978] = layer1_out[7307] & ~layer1_out[7308];
    assign layer2_out[6979] = layer1_out[6008];
    assign layer2_out[6980] = layer1_out[6913] & layer1_out[6914];
    assign layer2_out[6981] = layer1_out[1758] ^ layer1_out[1759];
    assign layer2_out[6982] = layer1_out[1445] & ~layer1_out[1446];
    assign layer2_out[6983] = ~(layer1_out[1290] | layer1_out[1291]);
    assign layer2_out[6984] = ~(layer1_out[2870] ^ layer1_out[2871]);
    assign layer2_out[6985] = layer1_out[1455] & layer1_out[1456];
    assign layer2_out[6986] = layer1_out[7117];
    assign layer2_out[6987] = layer1_out[3089];
    assign layer2_out[6988] = layer1_out[5958] | layer1_out[5959];
    assign layer2_out[6989] = ~layer1_out[4848];
    assign layer2_out[6990] = 1'b1;
    assign layer2_out[6991] = ~layer1_out[1207];
    assign layer2_out[6992] = ~(layer1_out[7626] & layer1_out[7627]);
    assign layer2_out[6993] = ~(layer1_out[6071] | layer1_out[6072]);
    assign layer2_out[6994] = ~layer1_out[7951];
    assign layer2_out[6995] = layer1_out[2083];
    assign layer2_out[6996] = layer1_out[323] ^ layer1_out[324];
    assign layer2_out[6997] = layer1_out[7262];
    assign layer2_out[6998] = ~(layer1_out[4212] ^ layer1_out[4213]);
    assign layer2_out[6999] = layer1_out[3406] ^ layer1_out[3407];
    assign layer2_out[7000] = ~(layer1_out[7056] | layer1_out[7057]);
    assign layer2_out[7001] = layer1_out[2292] & ~layer1_out[2293];
    assign layer2_out[7002] = ~layer1_out[5137];
    assign layer2_out[7003] = layer1_out[4130] | layer1_out[4131];
    assign layer2_out[7004] = layer1_out[1564] & ~layer1_out[1563];
    assign layer2_out[7005] = layer1_out[3726];
    assign layer2_out[7006] = ~layer1_out[1312] | layer1_out[1311];
    assign layer2_out[7007] = layer1_out[7758] & ~layer1_out[7759];
    assign layer2_out[7008] = layer1_out[2578] & layer1_out[2579];
    assign layer2_out[7009] = ~layer1_out[5418] | layer1_out[5419];
    assign layer2_out[7010] = ~layer1_out[4887];
    assign layer2_out[7011] = ~layer1_out[1958];
    assign layer2_out[7012] = layer1_out[1702] & ~layer1_out[1703];
    assign layer2_out[7013] = ~layer1_out[1067] | layer1_out[1066];
    assign layer2_out[7014] = layer1_out[1195];
    assign layer2_out[7015] = layer1_out[1193];
    assign layer2_out[7016] = ~layer1_out[2400];
    assign layer2_out[7017] = ~(layer1_out[2779] | layer1_out[2780]);
    assign layer2_out[7018] = ~layer1_out[1282] | layer1_out[1283];
    assign layer2_out[7019] = 1'b0;
    assign layer2_out[7020] = layer1_out[6346] & layer1_out[6347];
    assign layer2_out[7021] = layer1_out[3480];
    assign layer2_out[7022] = ~layer1_out[2575] | layer1_out[2574];
    assign layer2_out[7023] = layer1_out[1836] | layer1_out[1837];
    assign layer2_out[7024] = layer1_out[1771] & ~layer1_out[1772];
    assign layer2_out[7025] = layer1_out[2864];
    assign layer2_out[7026] = ~(layer1_out[4663] & layer1_out[4664]);
    assign layer2_out[7027] = ~layer1_out[1332];
    assign layer2_out[7028] = ~layer1_out[6366];
    assign layer2_out[7029] = layer1_out[2683];
    assign layer2_out[7030] = ~layer1_out[1777] | layer1_out[1778];
    assign layer2_out[7031] = ~layer1_out[303] | layer1_out[302];
    assign layer2_out[7032] = ~(layer1_out[5558] & layer1_out[5559]);
    assign layer2_out[7033] = layer1_out[7371] & layer1_out[7372];
    assign layer2_out[7034] = layer1_out[4994] ^ layer1_out[4995];
    assign layer2_out[7035] = ~layer1_out[4499];
    assign layer2_out[7036] = ~layer1_out[796];
    assign layer2_out[7037] = ~layer1_out[3226] | layer1_out[3225];
    assign layer2_out[7038] = ~(layer1_out[7343] ^ layer1_out[7344]);
    assign layer2_out[7039] = layer1_out[6995] | layer1_out[6996];
    assign layer2_out[7040] = ~layer1_out[4384];
    assign layer2_out[7041] = layer1_out[5631];
    assign layer2_out[7042] = ~layer1_out[5699] | layer1_out[5698];
    assign layer2_out[7043] = layer1_out[5403] | layer1_out[5404];
    assign layer2_out[7044] = ~layer1_out[1138] | layer1_out[1137];
    assign layer2_out[7045] = ~layer1_out[6528];
    assign layer2_out[7046] = ~layer1_out[6314] | layer1_out[6313];
    assign layer2_out[7047] = ~layer1_out[682] | layer1_out[683];
    assign layer2_out[7048] = layer1_out[3924];
    assign layer2_out[7049] = ~layer1_out[1216] | layer1_out[1217];
    assign layer2_out[7050] = layer1_out[3804] & ~layer1_out[3803];
    assign layer2_out[7051] = ~(layer1_out[1752] | layer1_out[1753]);
    assign layer2_out[7052] = ~layer1_out[4396];
    assign layer2_out[7053] = layer1_out[7176] | layer1_out[7177];
    assign layer2_out[7054] = layer1_out[684] & ~layer1_out[683];
    assign layer2_out[7055] = ~(layer1_out[617] | layer1_out[618]);
    assign layer2_out[7056] = ~layer1_out[6867];
    assign layer2_out[7057] = ~layer1_out[5498];
    assign layer2_out[7058] = ~layer1_out[197] | layer1_out[198];
    assign layer2_out[7059] = layer1_out[73] & ~layer1_out[74];
    assign layer2_out[7060] = layer1_out[6314];
    assign layer2_out[7061] = 1'b0;
    assign layer2_out[7062] = 1'b0;
    assign layer2_out[7063] = ~(layer1_out[2421] | layer1_out[2422]);
    assign layer2_out[7064] = 1'b0;
    assign layer2_out[7065] = layer1_out[1528] | layer1_out[1529];
    assign layer2_out[7066] = layer1_out[4487];
    assign layer2_out[7067] = ~layer1_out[2322];
    assign layer2_out[7068] = layer1_out[3249] | layer1_out[3250];
    assign layer2_out[7069] = ~layer1_out[6677];
    assign layer2_out[7070] = layer1_out[5286];
    assign layer2_out[7071] = layer1_out[620];
    assign layer2_out[7072] = ~(layer1_out[5862] ^ layer1_out[5863]);
    assign layer2_out[7073] = ~(layer1_out[6565] & layer1_out[6566]);
    assign layer2_out[7074] = ~(layer1_out[1118] | layer1_out[1119]);
    assign layer2_out[7075] = ~layer1_out[2336];
    assign layer2_out[7076] = ~layer1_out[4881] | layer1_out[4880];
    assign layer2_out[7077] = ~(layer1_out[5682] | layer1_out[5683]);
    assign layer2_out[7078] = ~layer1_out[4652];
    assign layer2_out[7079] = ~layer1_out[6169] | layer1_out[6170];
    assign layer2_out[7080] = ~layer1_out[178];
    assign layer2_out[7081] = layer1_out[7547] & ~layer1_out[7548];
    assign layer2_out[7082] = 1'b1;
    assign layer2_out[7083] = layer1_out[873];
    assign layer2_out[7084] = ~(layer1_out[5895] | layer1_out[5896]);
    assign layer2_out[7085] = ~(layer1_out[3215] ^ layer1_out[3216]);
    assign layer2_out[7086] = ~layer1_out[2482];
    assign layer2_out[7087] = ~(layer1_out[7452] | layer1_out[7453]);
    assign layer2_out[7088] = ~layer1_out[6935] | layer1_out[6934];
    assign layer2_out[7089] = layer1_out[1144];
    assign layer2_out[7090] = ~layer1_out[4134] | layer1_out[4135];
    assign layer2_out[7091] = layer1_out[3161] | layer1_out[3162];
    assign layer2_out[7092] = ~layer1_out[5362];
    assign layer2_out[7093] = 1'b0;
    assign layer2_out[7094] = 1'b0;
    assign layer2_out[7095] = layer1_out[7215];
    assign layer2_out[7096] = ~(layer1_out[6602] & layer1_out[6603]);
    assign layer2_out[7097] = layer1_out[335];
    assign layer2_out[7098] = ~layer1_out[3742];
    assign layer2_out[7099] = ~layer1_out[923];
    assign layer2_out[7100] = ~layer1_out[5345] | layer1_out[5344];
    assign layer2_out[7101] = ~(layer1_out[3136] ^ layer1_out[3137]);
    assign layer2_out[7102] = ~(layer1_out[7297] & layer1_out[7298]);
    assign layer2_out[7103] = ~layer1_out[4444] | layer1_out[4445];
    assign layer2_out[7104] = ~layer1_out[5333];
    assign layer2_out[7105] = layer1_out[2984] & ~layer1_out[2985];
    assign layer2_out[7106] = ~(layer1_out[7057] | layer1_out[7058]);
    assign layer2_out[7107] = 1'b1;
    assign layer2_out[7108] = ~(layer1_out[6917] ^ layer1_out[6918]);
    assign layer2_out[7109] = ~layer1_out[7958];
    assign layer2_out[7110] = ~layer1_out[414];
    assign layer2_out[7111] = ~(layer1_out[4172] | layer1_out[4173]);
    assign layer2_out[7112] = ~(layer1_out[7666] & layer1_out[7667]);
    assign layer2_out[7113] = layer1_out[4232] & ~layer1_out[4231];
    assign layer2_out[7114] = ~(layer1_out[3476] & layer1_out[3477]);
    assign layer2_out[7115] = ~(layer1_out[6902] | layer1_out[6903]);
    assign layer2_out[7116] = ~layer1_out[4249] | layer1_out[4248];
    assign layer2_out[7117] = layer1_out[3291] | layer1_out[3292];
    assign layer2_out[7118] = ~(layer1_out[1173] | layer1_out[1174]);
    assign layer2_out[7119] = ~layer1_out[6829] | layer1_out[6830];
    assign layer2_out[7120] = layer1_out[2449] & ~layer1_out[2450];
    assign layer2_out[7121] = ~layer1_out[4547] | layer1_out[4546];
    assign layer2_out[7122] = 1'b1;
    assign layer2_out[7123] = layer1_out[3159] & ~layer1_out[3158];
    assign layer2_out[7124] = ~layer1_out[2936];
    assign layer2_out[7125] = ~layer1_out[5417];
    assign layer2_out[7126] = ~(layer1_out[7892] | layer1_out[7893]);
    assign layer2_out[7127] = ~layer1_out[7096];
    assign layer2_out[7128] = ~layer1_out[2196] | layer1_out[2195];
    assign layer2_out[7129] = ~(layer1_out[4209] & layer1_out[4210]);
    assign layer2_out[7130] = ~(layer1_out[4607] | layer1_out[4608]);
    assign layer2_out[7131] = layer1_out[5104] ^ layer1_out[5105];
    assign layer2_out[7132] = ~layer1_out[39];
    assign layer2_out[7133] = ~layer1_out[5222];
    assign layer2_out[7134] = layer1_out[247];
    assign layer2_out[7135] = layer1_out[1324] & layer1_out[1325];
    assign layer2_out[7136] = layer1_out[6701] & ~layer1_out[6702];
    assign layer2_out[7137] = layer1_out[7700];
    assign layer2_out[7138] = ~layer1_out[422];
    assign layer2_out[7139] = ~layer1_out[3707] | layer1_out[3708];
    assign layer2_out[7140] = ~layer1_out[2428];
    assign layer2_out[7141] = ~(layer1_out[7903] ^ layer1_out[7904]);
    assign layer2_out[7142] = layer1_out[1161];
    assign layer2_out[7143] = layer1_out[6335] | layer1_out[6336];
    assign layer2_out[7144] = layer1_out[4123] & layer1_out[4124];
    assign layer2_out[7145] = layer1_out[2778];
    assign layer2_out[7146] = ~layer1_out[836];
    assign layer2_out[7147] = ~layer1_out[7543] | layer1_out[7542];
    assign layer2_out[7148] = layer1_out[1233] & layer1_out[1234];
    assign layer2_out[7149] = layer1_out[1726] & layer1_out[1727];
    assign layer2_out[7150] = layer1_out[5566] ^ layer1_out[5567];
    assign layer2_out[7151] = 1'b1;
    assign layer2_out[7152] = ~layer1_out[2774] | layer1_out[2775];
    assign layer2_out[7153] = layer1_out[5122] & layer1_out[5123];
    assign layer2_out[7154] = ~(layer1_out[7724] | layer1_out[7725]);
    assign layer2_out[7155] = ~(layer1_out[7618] ^ layer1_out[7619]);
    assign layer2_out[7156] = ~(layer1_out[4183] | layer1_out[4184]);
    assign layer2_out[7157] = ~(layer1_out[5638] | layer1_out[5639]);
    assign layer2_out[7158] = layer1_out[615];
    assign layer2_out[7159] = layer1_out[7196];
    assign layer2_out[7160] = layer1_out[4345] & layer1_out[4346];
    assign layer2_out[7161] = layer1_out[4764];
    assign layer2_out[7162] = layer1_out[4322] & ~layer1_out[4323];
    assign layer2_out[7163] = layer1_out[7512] & layer1_out[7513];
    assign layer2_out[7164] = ~layer1_out[3331] | layer1_out[3330];
    assign layer2_out[7165] = layer1_out[6372] & layer1_out[6373];
    assign layer2_out[7166] = ~layer1_out[7102] | layer1_out[7101];
    assign layer2_out[7167] = ~layer1_out[1213] | layer1_out[1214];
    assign layer2_out[7168] = 1'b1;
    assign layer2_out[7169] = ~layer1_out[2859];
    assign layer2_out[7170] = layer1_out[4132] & layer1_out[4133];
    assign layer2_out[7171] = layer1_out[4555] ^ layer1_out[4556];
    assign layer2_out[7172] = ~layer1_out[5106];
    assign layer2_out[7173] = layer1_out[689];
    assign layer2_out[7174] = layer1_out[7088] & ~layer1_out[7089];
    assign layer2_out[7175] = layer1_out[5042] & layer1_out[5043];
    assign layer2_out[7176] = layer1_out[7033];
    assign layer2_out[7177] = layer1_out[1086];
    assign layer2_out[7178] = ~layer1_out[1478];
    assign layer2_out[7179] = layer1_out[6640] | layer1_out[6641];
    assign layer2_out[7180] = layer1_out[3028];
    assign layer2_out[7181] = layer1_out[5427] & layer1_out[5428];
    assign layer2_out[7182] = ~(layer1_out[7636] & layer1_out[7637]);
    assign layer2_out[7183] = ~layer1_out[304] | layer1_out[303];
    assign layer2_out[7184] = layer1_out[5746];
    assign layer2_out[7185] = ~(layer1_out[6012] | layer1_out[6013]);
    assign layer2_out[7186] = ~(layer1_out[2084] | layer1_out[2085]);
    assign layer2_out[7187] = 1'b0;
    assign layer2_out[7188] = ~layer1_out[7199];
    assign layer2_out[7189] = layer1_out[3857] & layer1_out[3858];
    assign layer2_out[7190] = ~layer1_out[3324];
    assign layer2_out[7191] = ~layer1_out[4690] | layer1_out[4691];
    assign layer2_out[7192] = ~layer1_out[6697] | layer1_out[6698];
    assign layer2_out[7193] = ~layer1_out[7193];
    assign layer2_out[7194] = layer1_out[3556] & ~layer1_out[3555];
    assign layer2_out[7195] = ~(layer1_out[5663] | layer1_out[5664]);
    assign layer2_out[7196] = ~layer1_out[103] | layer1_out[104];
    assign layer2_out[7197] = layer1_out[3155] | layer1_out[3156];
    assign layer2_out[7198] = layer1_out[1832];
    assign layer2_out[7199] = 1'b1;
    assign layer2_out[7200] = layer1_out[4728];
    assign layer2_out[7201] = layer1_out[1108] & ~layer1_out[1107];
    assign layer2_out[7202] = ~layer1_out[2516];
    assign layer2_out[7203] = ~layer1_out[1099] | layer1_out[1100];
    assign layer2_out[7204] = layer1_out[1054];
    assign layer2_out[7205] = ~(layer1_out[3144] | layer1_out[3145]);
    assign layer2_out[7206] = ~layer1_out[453];
    assign layer2_out[7207] = ~layer1_out[7744];
    assign layer2_out[7208] = ~(layer1_out[5738] ^ layer1_out[5739]);
    assign layer2_out[7209] = layer1_out[6188];
    assign layer2_out[7210] = layer1_out[3869] | layer1_out[3870];
    assign layer2_out[7211] = layer1_out[1269];
    assign layer2_out[7212] = ~layer1_out[2415] | layer1_out[2416];
    assign layer2_out[7213] = layer1_out[3263] & layer1_out[3264];
    assign layer2_out[7214] = ~layer1_out[7385] | layer1_out[7384];
    assign layer2_out[7215] = ~(layer1_out[5851] & layer1_out[5852]);
    assign layer2_out[7216] = ~(layer1_out[6764] | layer1_out[6765]);
    assign layer2_out[7217] = layer1_out[3811] & layer1_out[3812];
    assign layer2_out[7218] = layer1_out[4419] & ~layer1_out[4420];
    assign layer2_out[7219] = layer1_out[6263];
    assign layer2_out[7220] = ~layer1_out[2886] | layer1_out[2885];
    assign layer2_out[7221] = layer1_out[7941];
    assign layer2_out[7222] = layer1_out[3793] ^ layer1_out[3794];
    assign layer2_out[7223] = layer1_out[144] | layer1_out[145];
    assign layer2_out[7224] = ~layer1_out[3461];
    assign layer2_out[7225] = ~(layer1_out[7668] | layer1_out[7669]);
    assign layer2_out[7226] = ~(layer1_out[7606] ^ layer1_out[7607]);
    assign layer2_out[7227] = layer1_out[6333];
    assign layer2_out[7228] = layer1_out[2714] & layer1_out[2715];
    assign layer2_out[7229] = ~layer1_out[7759] | layer1_out[7760];
    assign layer2_out[7230] = ~layer1_out[3567] | layer1_out[3566];
    assign layer2_out[7231] = layer1_out[5074];
    assign layer2_out[7232] = 1'b1;
    assign layer2_out[7233] = layer1_out[1750] & ~layer1_out[1749];
    assign layer2_out[7234] = 1'b1;
    assign layer2_out[7235] = layer1_out[2190] ^ layer1_out[2191];
    assign layer2_out[7236] = layer1_out[5006];
    assign layer2_out[7237] = ~(layer1_out[7423] | layer1_out[7424]);
    assign layer2_out[7238] = layer1_out[1241] | layer1_out[1242];
    assign layer2_out[7239] = layer1_out[6045];
    assign layer2_out[7240] = ~layer1_out[3297];
    assign layer2_out[7241] = layer1_out[7559] & ~layer1_out[7560];
    assign layer2_out[7242] = layer1_out[3305];
    assign layer2_out[7243] = ~layer1_out[7360];
    assign layer2_out[7244] = ~(layer1_out[4428] & layer1_out[4429]);
    assign layer2_out[7245] = layer1_out[7227];
    assign layer2_out[7246] = layer1_out[1967] & ~layer1_out[1968];
    assign layer2_out[7247] = ~layer1_out[1428];
    assign layer2_out[7248] = 1'b1;
    assign layer2_out[7249] = layer1_out[2532] & ~layer1_out[2533];
    assign layer2_out[7250] = ~(layer1_out[2570] ^ layer1_out[2571]);
    assign layer2_out[7251] = ~layer1_out[5486];
    assign layer2_out[7252] = ~(layer1_out[6119] & layer1_out[6120]);
    assign layer2_out[7253] = ~(layer1_out[6014] | layer1_out[6015]);
    assign layer2_out[7254] = layer1_out[1164] & ~layer1_out[1163];
    assign layer2_out[7255] = ~(layer1_out[1623] & layer1_out[1624]);
    assign layer2_out[7256] = ~layer1_out[7143] | layer1_out[7142];
    assign layer2_out[7257] = ~layer1_out[3818] | layer1_out[3817];
    assign layer2_out[7258] = ~layer1_out[1479];
    assign layer2_out[7259] = layer1_out[2298];
    assign layer2_out[7260] = ~layer1_out[4083];
    assign layer2_out[7261] = layer1_out[939] & ~layer1_out[940];
    assign layer2_out[7262] = layer1_out[5424] | layer1_out[5425];
    assign layer2_out[7263] = ~(layer1_out[7046] | layer1_out[7047]);
    assign layer2_out[7264] = ~layer1_out[7805];
    assign layer2_out[7265] = ~layer1_out[4323];
    assign layer2_out[7266] = layer1_out[364] & ~layer1_out[363];
    assign layer2_out[7267] = ~(layer1_out[1486] ^ layer1_out[1487]);
    assign layer2_out[7268] = layer1_out[1857] & layer1_out[1858];
    assign layer2_out[7269] = layer1_out[6195];
    assign layer2_out[7270] = ~layer1_out[7943];
    assign layer2_out[7271] = ~layer1_out[3528];
    assign layer2_out[7272] = ~(layer1_out[5732] ^ layer1_out[5733]);
    assign layer2_out[7273] = ~layer1_out[4311] | layer1_out[4310];
    assign layer2_out[7274] = ~layer1_out[6797];
    assign layer2_out[7275] = ~layer1_out[5781];
    assign layer2_out[7276] = ~layer1_out[1879] | layer1_out[1880];
    assign layer2_out[7277] = ~layer1_out[3179];
    assign layer2_out[7278] = layer1_out[7584];
    assign layer2_out[7279] = layer1_out[7738] & ~layer1_out[7737];
    assign layer2_out[7280] = layer1_out[7781] ^ layer1_out[7782];
    assign layer2_out[7281] = ~(layer1_out[7793] ^ layer1_out[7794]);
    assign layer2_out[7282] = layer1_out[2898] & layer1_out[2899];
    assign layer2_out[7283] = layer1_out[6669] & ~layer1_out[6668];
    assign layer2_out[7284] = ~layer1_out[1498];
    assign layer2_out[7285] = layer1_out[658] | layer1_out[659];
    assign layer2_out[7286] = ~(layer1_out[3114] ^ layer1_out[3115]);
    assign layer2_out[7287] = ~(layer1_out[7548] & layer1_out[7549]);
    assign layer2_out[7288] = layer1_out[7594] & layer1_out[7595];
    assign layer2_out[7289] = ~layer1_out[3836] | layer1_out[3837];
    assign layer2_out[7290] = layer1_out[1694] & layer1_out[1695];
    assign layer2_out[7291] = layer1_out[4846];
    assign layer2_out[7292] = ~(layer1_out[1824] | layer1_out[1825]);
    assign layer2_out[7293] = ~layer1_out[180];
    assign layer2_out[7294] = ~layer1_out[6330];
    assign layer2_out[7295] = ~layer1_out[6337] | layer1_out[6338];
    assign layer2_out[7296] = ~layer1_out[3856];
    assign layer2_out[7297] = layer1_out[7172] & layer1_out[7173];
    assign layer2_out[7298] = ~layer1_out[37] | layer1_out[38];
    assign layer2_out[7299] = ~layer1_out[3983] | layer1_out[3984];
    assign layer2_out[7300] = ~(layer1_out[337] & layer1_out[338]);
    assign layer2_out[7301] = ~(layer1_out[2344] | layer1_out[2345]);
    assign layer2_out[7302] = layer1_out[1388];
    assign layer2_out[7303] = ~layer1_out[2394] | layer1_out[2393];
    assign layer2_out[7304] = ~(layer1_out[7340] ^ layer1_out[7341]);
    assign layer2_out[7305] = layer1_out[7866];
    assign layer2_out[7306] = layer1_out[6857] & ~layer1_out[6858];
    assign layer2_out[7307] = layer1_out[7979];
    assign layer2_out[7308] = layer1_out[6547] & ~layer1_out[6548];
    assign layer2_out[7309] = layer1_out[493] ^ layer1_out[494];
    assign layer2_out[7310] = layer1_out[6608] & ~layer1_out[6607];
    assign layer2_out[7311] = layer1_out[163];
    assign layer2_out[7312] = layer1_out[4980] & ~layer1_out[4979];
    assign layer2_out[7313] = ~(layer1_out[3542] | layer1_out[3543]);
    assign layer2_out[7314] = layer1_out[879] | layer1_out[880];
    assign layer2_out[7315] = 1'b1;
    assign layer2_out[7316] = layer1_out[6535] & ~layer1_out[6534];
    assign layer2_out[7317] = ~layer1_out[7562];
    assign layer2_out[7318] = ~layer1_out[6498];
    assign layer2_out[7319] = ~layer1_out[5885];
    assign layer2_out[7320] = layer1_out[78] & layer1_out[79];
    assign layer2_out[7321] = layer1_out[4204];
    assign layer2_out[7322] = layer1_out[3926] ^ layer1_out[3927];
    assign layer2_out[7323] = layer1_out[7586] ^ layer1_out[7587];
    assign layer2_out[7324] = ~layer1_out[1189] | layer1_out[1190];
    assign layer2_out[7325] = layer1_out[4371] & ~layer1_out[4372];
    assign layer2_out[7326] = ~layer1_out[5954];
    assign layer2_out[7327] = 1'b1;
    assign layer2_out[7328] = ~layer1_out[4185] | layer1_out[4184];
    assign layer2_out[7329] = ~(layer1_out[7465] | layer1_out[7466]);
    assign layer2_out[7330] = layer1_out[5266] & ~layer1_out[5265];
    assign layer2_out[7331] = layer1_out[4772] & ~layer1_out[4771];
    assign layer2_out[7332] = layer1_out[619];
    assign layer2_out[7333] = ~layer1_out[4208];
    assign layer2_out[7334] = layer1_out[4807] & ~layer1_out[4806];
    assign layer2_out[7335] = layer1_out[5143] ^ layer1_out[5144];
    assign layer2_out[7336] = ~layer1_out[6184];
    assign layer2_out[7337] = layer1_out[5069];
    assign layer2_out[7338] = layer1_out[4179] & ~layer1_out[4180];
    assign layer2_out[7339] = ~(layer1_out[2742] | layer1_out[2743]);
    assign layer2_out[7340] = layer1_out[2243] & ~layer1_out[2244];
    assign layer2_out[7341] = ~layer1_out[1045] | layer1_out[1046];
    assign layer2_out[7342] = layer1_out[7384];
    assign layer2_out[7343] = layer1_out[723];
    assign layer2_out[7344] = ~(layer1_out[835] & layer1_out[836]);
    assign layer2_out[7345] = layer1_out[1310] | layer1_out[1311];
    assign layer2_out[7346] = layer1_out[7763];
    assign layer2_out[7347] = layer1_out[7516];
    assign layer2_out[7348] = ~layer1_out[5764] | layer1_out[5765];
    assign layer2_out[7349] = layer1_out[368] | layer1_out[369];
    assign layer2_out[7350] = layer1_out[634] & ~layer1_out[635];
    assign layer2_out[7351] = layer1_out[893] ^ layer1_out[894];
    assign layer2_out[7352] = ~layer1_out[3189] | layer1_out[3188];
    assign layer2_out[7353] = ~(layer1_out[3385] & layer1_out[3386]);
    assign layer2_out[7354] = layer1_out[5494] & layer1_out[5495];
    assign layer2_out[7355] = ~(layer1_out[5263] ^ layer1_out[5264]);
    assign layer2_out[7356] = ~layer1_out[3997];
    assign layer2_out[7357] = layer1_out[7218];
    assign layer2_out[7358] = layer1_out[3819];
    assign layer2_out[7359] = ~layer1_out[215];
    assign layer2_out[7360] = ~layer1_out[2343] | layer1_out[2342];
    assign layer2_out[7361] = layer1_out[6393] & layer1_out[6394];
    assign layer2_out[7362] = ~layer1_out[4613];
    assign layer2_out[7363] = layer1_out[2332] & ~layer1_out[2333];
    assign layer2_out[7364] = ~layer1_out[4629];
    assign layer2_out[7365] = layer1_out[6671] & layer1_out[6672];
    assign layer2_out[7366] = ~layer1_out[5392] | layer1_out[5393];
    assign layer2_out[7367] = layer1_out[4347];
    assign layer2_out[7368] = layer1_out[3672];
    assign layer2_out[7369] = ~layer1_out[4155];
    assign layer2_out[7370] = layer1_out[7676];
    assign layer2_out[7371] = layer1_out[2060] & ~layer1_out[2061];
    assign layer2_out[7372] = layer1_out[7968];
    assign layer2_out[7373] = ~layer1_out[6357];
    assign layer2_out[7374] = ~layer1_out[6659] | layer1_out[6660];
    assign layer2_out[7375] = 1'b1;
    assign layer2_out[7376] = layer1_out[2046] ^ layer1_out[2047];
    assign layer2_out[7377] = ~layer1_out[5748];
    assign layer2_out[7378] = ~layer1_out[4824];
    assign layer2_out[7379] = layer1_out[4910];
    assign layer2_out[7380] = ~layer1_out[2764];
    assign layer2_out[7381] = ~layer1_out[1999];
    assign layer2_out[7382] = ~layer1_out[4638] | layer1_out[4637];
    assign layer2_out[7383] = ~layer1_out[613];
    assign layer2_out[7384] = ~layer1_out[6767] | layer1_out[6766];
    assign layer2_out[7385] = layer1_out[121] & ~layer1_out[120];
    assign layer2_out[7386] = ~layer1_out[3382] | layer1_out[3383];
    assign layer2_out[7387] = ~(layer1_out[4939] & layer1_out[4940]);
    assign layer2_out[7388] = ~layer1_out[4764] | layer1_out[4765];
    assign layer2_out[7389] = ~(layer1_out[7210] & layer1_out[7211]);
    assign layer2_out[7390] = layer1_out[7788];
    assign layer2_out[7391] = ~(layer1_out[3786] & layer1_out[3787]);
    assign layer2_out[7392] = ~layer1_out[2640] | layer1_out[2639];
    assign layer2_out[7393] = ~layer1_out[7095] | layer1_out[7094];
    assign layer2_out[7394] = ~(layer1_out[2085] | layer1_out[2086]);
    assign layer2_out[7395] = ~layer1_out[3690] | layer1_out[3689];
    assign layer2_out[7396] = layer1_out[1734] & layer1_out[1735];
    assign layer2_out[7397] = layer1_out[1743] | layer1_out[1744];
    assign layer2_out[7398] = layer1_out[3190];
    assign layer2_out[7399] = 1'b1;
    assign layer2_out[7400] = ~layer1_out[702];
    assign layer2_out[7401] = layer1_out[7751] & ~layer1_out[7752];
    assign layer2_out[7402] = ~layer1_out[7001] | layer1_out[7000];
    assign layer2_out[7403] = ~layer1_out[3842];
    assign layer2_out[7404] = ~(layer1_out[2815] | layer1_out[2816]);
    assign layer2_out[7405] = layer1_out[111];
    assign layer2_out[7406] = ~layer1_out[3150] | layer1_out[3149];
    assign layer2_out[7407] = ~layer1_out[1785];
    assign layer2_out[7408] = ~(layer1_out[2847] & layer1_out[2848]);
    assign layer2_out[7409] = layer1_out[1116] | layer1_out[1117];
    assign layer2_out[7410] = ~(layer1_out[3305] & layer1_out[3306]);
    assign layer2_out[7411] = layer1_out[2725] & layer1_out[2726];
    assign layer2_out[7412] = layer1_out[3282];
    assign layer2_out[7413] = ~layer1_out[1031];
    assign layer2_out[7414] = ~layer1_out[667] | layer1_out[666];
    assign layer2_out[7415] = layer1_out[3925];
    assign layer2_out[7416] = ~(layer1_out[7865] ^ layer1_out[7866]);
    assign layer2_out[7417] = layer1_out[6502] | layer1_out[6503];
    assign layer2_out[7418] = layer1_out[1056] & ~layer1_out[1057];
    assign layer2_out[7419] = ~layer1_out[2332] | layer1_out[2331];
    assign layer2_out[7420] = layer1_out[1254];
    assign layer2_out[7421] = ~layer1_out[294] | layer1_out[295];
    assign layer2_out[7422] = layer1_out[7703] & layer1_out[7704];
    assign layer2_out[7423] = layer1_out[2634];
    assign layer2_out[7424] = ~layer1_out[6990];
    assign layer2_out[7425] = 1'b1;
    assign layer2_out[7426] = layer1_out[7864];
    assign layer2_out[7427] = layer1_out[6241];
    assign layer2_out[7428] = ~(layer1_out[6184] & layer1_out[6185]);
    assign layer2_out[7429] = ~layer1_out[4035];
    assign layer2_out[7430] = layer1_out[3377] & ~layer1_out[3378];
    assign layer2_out[7431] = ~layer1_out[3901];
    assign layer2_out[7432] = layer1_out[7815] | layer1_out[7816];
    assign layer2_out[7433] = ~layer1_out[4251];
    assign layer2_out[7434] = ~layer1_out[1709];
    assign layer2_out[7435] = ~layer1_out[4935];
    assign layer2_out[7436] = 1'b1;
    assign layer2_out[7437] = layer1_out[2073];
    assign layer2_out[7438] = layer1_out[238] & ~layer1_out[237];
    assign layer2_out[7439] = layer1_out[2029] & layer1_out[2030];
    assign layer2_out[7440] = ~layer1_out[2861];
    assign layer2_out[7441] = ~(layer1_out[7091] ^ layer1_out[7092]);
    assign layer2_out[7442] = layer1_out[2835] ^ layer1_out[2836];
    assign layer2_out[7443] = layer1_out[3822] & ~layer1_out[3823];
    assign layer2_out[7444] = 1'b1;
    assign layer2_out[7445] = layer1_out[3864] | layer1_out[3865];
    assign layer2_out[7446] = layer1_out[6248] & ~layer1_out[6247];
    assign layer2_out[7447] = layer1_out[4481] ^ layer1_out[4482];
    assign layer2_out[7448] = ~(layer1_out[5097] & layer1_out[5098]);
    assign layer2_out[7449] = ~(layer1_out[3781] & layer1_out[3782]);
    assign layer2_out[7450] = ~(layer1_out[761] | layer1_out[762]);
    assign layer2_out[7451] = layer1_out[7963];
    assign layer2_out[7452] = ~(layer1_out[1751] ^ layer1_out[1752]);
    assign layer2_out[7453] = layer1_out[6611] ^ layer1_out[6612];
    assign layer2_out[7454] = ~(layer1_out[2588] | layer1_out[2589]);
    assign layer2_out[7455] = layer1_out[3075] & ~layer1_out[3076];
    assign layer2_out[7456] = 1'b1;
    assign layer2_out[7457] = layer1_out[2067];
    assign layer2_out[7458] = ~(layer1_out[2437] ^ layer1_out[2438]);
    assign layer2_out[7459] = ~layer1_out[6558] | layer1_out[6557];
    assign layer2_out[7460] = ~layer1_out[5121] | layer1_out[5122];
    assign layer2_out[7461] = ~layer1_out[6551];
    assign layer2_out[7462] = ~layer1_out[7575] | layer1_out[7576];
    assign layer2_out[7463] = layer1_out[6712];
    assign layer2_out[7464] = layer1_out[4841];
    assign layer2_out[7465] = ~layer1_out[910];
    assign layer2_out[7466] = layer1_out[6432];
    assign layer2_out[7467] = ~(layer1_out[7174] ^ layer1_out[7175]);
    assign layer2_out[7468] = ~layer1_out[7854] | layer1_out[7853];
    assign layer2_out[7469] = ~(layer1_out[1652] & layer1_out[1653]);
    assign layer2_out[7470] = ~layer1_out[5875] | layer1_out[5874];
    assign layer2_out[7471] = layer1_out[48] & ~layer1_out[47];
    assign layer2_out[7472] = ~layer1_out[4567];
    assign layer2_out[7473] = layer1_out[6658] & ~layer1_out[6659];
    assign layer2_out[7474] = ~layer1_out[7381];
    assign layer2_out[7475] = layer1_out[684];
    assign layer2_out[7476] = layer1_out[7680];
    assign layer2_out[7477] = ~layer1_out[2539];
    assign layer2_out[7478] = 1'b0;
    assign layer2_out[7479] = layer1_out[6778];
    assign layer2_out[7480] = 1'b0;
    assign layer2_out[7481] = layer1_out[1292] ^ layer1_out[1293];
    assign layer2_out[7482] = ~layer1_out[4517];
    assign layer2_out[7483] = ~layer1_out[6294] | layer1_out[6293];
    assign layer2_out[7484] = layer1_out[3815];
    assign layer2_out[7485] = 1'b0;
    assign layer2_out[7486] = ~layer1_out[812];
    assign layer2_out[7487] = layer1_out[6444];
    assign layer2_out[7488] = ~(layer1_out[1521] | layer1_out[1522]);
    assign layer2_out[7489] = layer1_out[5976] & layer1_out[5977];
    assign layer2_out[7490] = ~(layer1_out[57] & layer1_out[58]);
    assign layer2_out[7491] = layer1_out[538] & layer1_out[539];
    assign layer2_out[7492] = layer1_out[5819];
    assign layer2_out[7493] = ~(layer1_out[2805] & layer1_out[2806]);
    assign layer2_out[7494] = layer1_out[5270];
    assign layer2_out[7495] = layer1_out[5313];
    assign layer2_out[7496] = ~layer1_out[1259] | layer1_out[1258];
    assign layer2_out[7497] = ~layer1_out[3228];
    assign layer2_out[7498] = ~layer1_out[319];
    assign layer2_out[7499] = ~(layer1_out[4423] | layer1_out[4424]);
    assign layer2_out[7500] = ~layer1_out[6144];
    assign layer2_out[7501] = ~layer1_out[2092] | layer1_out[2093];
    assign layer2_out[7502] = layer1_out[492] | layer1_out[493];
    assign layer2_out[7503] = ~layer1_out[3163];
    assign layer2_out[7504] = ~layer1_out[1794] | layer1_out[1795];
    assign layer2_out[7505] = 1'b0;
    assign layer2_out[7506] = layer1_out[6533] | layer1_out[6534];
    assign layer2_out[7507] = ~layer1_out[6217];
    assign layer2_out[7508] = layer1_out[4956] | layer1_out[4957];
    assign layer2_out[7509] = ~layer1_out[2760] | layer1_out[2759];
    assign layer2_out[7510] = layer1_out[7154] | layer1_out[7155];
    assign layer2_out[7511] = ~layer1_out[1576] | layer1_out[1575];
    assign layer2_out[7512] = ~(layer1_out[4540] | layer1_out[4541]);
    assign layer2_out[7513] = layer1_out[2235] & layer1_out[2236];
    assign layer2_out[7514] = ~layer1_out[3653] | layer1_out[3654];
    assign layer2_out[7515] = layer1_out[6485];
    assign layer2_out[7516] = layer1_out[2555] | layer1_out[2556];
    assign layer2_out[7517] = layer1_out[1028] & ~layer1_out[1029];
    assign layer2_out[7518] = layer1_out[767] ^ layer1_out[768];
    assign layer2_out[7519] = ~(layer1_out[5713] | layer1_out[5714]);
    assign layer2_out[7520] = layer1_out[3911] | layer1_out[3912];
    assign layer2_out[7521] = layer1_out[6357] & ~layer1_out[6358];
    assign layer2_out[7522] = ~(layer1_out[6083] & layer1_out[6084]);
    assign layer2_out[7523] = ~layer1_out[1280] | layer1_out[1279];
    assign layer2_out[7524] = layer1_out[373] & ~layer1_out[372];
    assign layer2_out[7525] = ~layer1_out[874];
    assign layer2_out[7526] = layer1_out[690];
    assign layer2_out[7527] = layer1_out[3297] & layer1_out[3298];
    assign layer2_out[7528] = ~layer1_out[4418];
    assign layer2_out[7529] = ~(layer1_out[411] | layer1_out[412]);
    assign layer2_out[7530] = layer1_out[4984] & layer1_out[4985];
    assign layer2_out[7531] = ~(layer1_out[4780] | layer1_out[4781]);
    assign layer2_out[7532] = ~layer1_out[2773];
    assign layer2_out[7533] = ~layer1_out[7768];
    assign layer2_out[7534] = ~layer1_out[1087];
    assign layer2_out[7535] = ~(layer1_out[7482] | layer1_out[7483]);
    assign layer2_out[7536] = layer1_out[4654] ^ layer1_out[4655];
    assign layer2_out[7537] = 1'b0;
    assign layer2_out[7538] = ~(layer1_out[6904] & layer1_out[6905]);
    assign layer2_out[7539] = ~(layer1_out[1995] & layer1_out[1996]);
    assign layer2_out[7540] = layer1_out[3753];
    assign layer2_out[7541] = layer1_out[105];
    assign layer2_out[7542] = layer1_out[6885] & layer1_out[6886];
    assign layer2_out[7543] = ~layer1_out[6162];
    assign layer2_out[7544] = ~(layer1_out[7772] ^ layer1_out[7773]);
    assign layer2_out[7545] = ~layer1_out[3789] | layer1_out[3790];
    assign layer2_out[7546] = layer1_out[2104] & layer1_out[2105];
    assign layer2_out[7547] = ~layer1_out[4005];
    assign layer2_out[7548] = ~(layer1_out[637] & layer1_out[638]);
    assign layer2_out[7549] = layer1_out[7617] & ~layer1_out[7616];
    assign layer2_out[7550] = ~(layer1_out[5673] & layer1_out[5674]);
    assign layer2_out[7551] = layer1_out[6042];
    assign layer2_out[7552] = ~(layer1_out[3600] & layer1_out[3601]);
    assign layer2_out[7553] = ~(layer1_out[7741] | layer1_out[7742]);
    assign layer2_out[7554] = layer1_out[2850] & ~layer1_out[2849];
    assign layer2_out[7555] = layer1_out[1820] & ~layer1_out[1821];
    assign layer2_out[7556] = ~layer1_out[672];
    assign layer2_out[7557] = ~layer1_out[6211] | layer1_out[6212];
    assign layer2_out[7558] = layer1_out[3745] & layer1_out[3746];
    assign layer2_out[7559] = layer1_out[7231];
    assign layer2_out[7560] = ~layer1_out[7780] | layer1_out[7781];
    assign layer2_out[7561] = ~layer1_out[1293] | layer1_out[1294];
    assign layer2_out[7562] = ~layer1_out[888];
    assign layer2_out[7563] = ~layer1_out[1577] | layer1_out[1576];
    assign layer2_out[7564] = layer1_out[1480] ^ layer1_out[1481];
    assign layer2_out[7565] = ~layer1_out[7709] | layer1_out[7710];
    assign layer2_out[7566] = ~layer1_out[5022];
    assign layer2_out[7567] = ~(layer1_out[7189] | layer1_out[7190]);
    assign layer2_out[7568] = layer1_out[6631] & layer1_out[6632];
    assign layer2_out[7569] = layer1_out[1799] & layer1_out[1800];
    assign layer2_out[7570] = ~(layer1_out[2810] | layer1_out[2811]);
    assign layer2_out[7571] = 1'b0;
    assign layer2_out[7572] = layer1_out[6568] & ~layer1_out[6569];
    assign layer2_out[7573] = layer1_out[2234];
    assign layer2_out[7574] = ~layer1_out[370] | layer1_out[369];
    assign layer2_out[7575] = layer1_out[4029];
    assign layer2_out[7576] = layer1_out[6144];
    assign layer2_out[7577] = ~layer1_out[915] | layer1_out[916];
    assign layer2_out[7578] = layer1_out[6627];
    assign layer2_out[7579] = ~(layer1_out[4474] & layer1_out[4475]);
    assign layer2_out[7580] = ~layer1_out[44];
    assign layer2_out[7581] = layer1_out[13];
    assign layer2_out[7582] = ~layer1_out[7611] | layer1_out[7612];
    assign layer2_out[7583] = layer1_out[7235] ^ layer1_out[7236];
    assign layer2_out[7584] = layer1_out[352] & ~layer1_out[351];
    assign layer2_out[7585] = ~layer1_out[42];
    assign layer2_out[7586] = ~layer1_out[244] | layer1_out[245];
    assign layer2_out[7587] = ~layer1_out[627] | layer1_out[626];
    assign layer2_out[7588] = ~layer1_out[4326];
    assign layer2_out[7589] = ~(layer1_out[5828] ^ layer1_out[5829]);
    assign layer2_out[7590] = ~layer1_out[1496] | layer1_out[1497];
    assign layer2_out[7591] = layer1_out[5859] & ~layer1_out[5858];
    assign layer2_out[7592] = ~(layer1_out[1627] | layer1_out[1628]);
    assign layer2_out[7593] = layer1_out[6133];
    assign layer2_out[7594] = ~layer1_out[2579] | layer1_out[2580];
    assign layer2_out[7595] = layer1_out[6193] | layer1_out[6194];
    assign layer2_out[7596] = ~layer1_out[5337] | layer1_out[5338];
    assign layer2_out[7597] = layer1_out[3329] | layer1_out[3330];
    assign layer2_out[7598] = layer1_out[4313] & ~layer1_out[4312];
    assign layer2_out[7599] = ~layer1_out[5339];
    assign layer2_out[7600] = ~layer1_out[2241] | layer1_out[2242];
    assign layer2_out[7601] = ~(layer1_out[3989] & layer1_out[3990]);
    assign layer2_out[7602] = layer1_out[7940];
    assign layer2_out[7603] = layer1_out[928];
    assign layer2_out[7604] = ~layer1_out[6791] | layer1_out[6792];
    assign layer2_out[7605] = 1'b1;
    assign layer2_out[7606] = ~layer1_out[1984];
    assign layer2_out[7607] = layer1_out[3597];
    assign layer2_out[7608] = layer1_out[3534] & layer1_out[3535];
    assign layer2_out[7609] = ~layer1_out[476];
    assign layer2_out[7610] = ~layer1_out[6688] | layer1_out[6689];
    assign layer2_out[7611] = layer1_out[2520] | layer1_out[2521];
    assign layer2_out[7612] = ~layer1_out[608];
    assign layer2_out[7613] = layer1_out[4009] & layer1_out[4010];
    assign layer2_out[7614] = ~layer1_out[7550];
    assign layer2_out[7615] = ~layer1_out[2432] | layer1_out[2431];
    assign layer2_out[7616] = layer1_out[1419];
    assign layer2_out[7617] = layer1_out[7922] | layer1_out[7923];
    assign layer2_out[7618] = ~layer1_out[3767];
    assign layer2_out[7619] = ~(layer1_out[5538] ^ layer1_out[5539]);
    assign layer2_out[7620] = layer1_out[1593] ^ layer1_out[1594];
    assign layer2_out[7621] = ~(layer1_out[1395] & layer1_out[1396]);
    assign layer2_out[7622] = ~layer1_out[4528];
    assign layer2_out[7623] = layer1_out[4651] & layer1_out[4652];
    assign layer2_out[7624] = ~layer1_out[7234] | layer1_out[7233];
    assign layer2_out[7625] = ~layer1_out[79];
    assign layer2_out[7626] = ~layer1_out[2557] | layer1_out[2558];
    assign layer2_out[7627] = ~(layer1_out[7415] & layer1_out[7416]);
    assign layer2_out[7628] = ~layer1_out[1524] | layer1_out[1525];
    assign layer2_out[7629] = layer1_out[6888] ^ layer1_out[6889];
    assign layer2_out[7630] = layer1_out[5444] & ~layer1_out[5443];
    assign layer2_out[7631] = ~(layer1_out[725] | layer1_out[726]);
    assign layer2_out[7632] = layer1_out[527] | layer1_out[528];
    assign layer2_out[7633] = layer1_out[3603] | layer1_out[3604];
    assign layer2_out[7634] = ~(layer1_out[6076] | layer1_out[6077]);
    assign layer2_out[7635] = ~(layer1_out[6138] | layer1_out[6139]);
    assign layer2_out[7636] = ~(layer1_out[4805] & layer1_out[4806]);
    assign layer2_out[7637] = layer1_out[1807];
    assign layer2_out[7638] = ~layer1_out[2197] | layer1_out[2198];
    assign layer2_out[7639] = 1'b0;
    assign layer2_out[7640] = ~(layer1_out[7026] & layer1_out[7027]);
    assign layer2_out[7641] = 1'b1;
    assign layer2_out[7642] = layer1_out[4463] & ~layer1_out[4464];
    assign layer2_out[7643] = ~layer1_out[2613] | layer1_out[2612];
    assign layer2_out[7644] = ~layer1_out[3348];
    assign layer2_out[7645] = layer1_out[2853] & ~layer1_out[2854];
    assign layer2_out[7646] = ~layer1_out[7960];
    assign layer2_out[7647] = layer1_out[3432] ^ layer1_out[3433];
    assign layer2_out[7648] = 1'b0;
    assign layer2_out[7649] = layer1_out[7619] & layer1_out[7620];
    assign layer2_out[7650] = 1'b0;
    assign layer2_out[7651] = layer1_out[399] & ~layer1_out[400];
    assign layer2_out[7652] = layer1_out[5688] & ~layer1_out[5689];
    assign layer2_out[7653] = layer1_out[7471];
    assign layer2_out[7654] = layer1_out[4164] & ~layer1_out[4163];
    assign layer2_out[7655] = ~(layer1_out[7100] | layer1_out[7101]);
    assign layer2_out[7656] = layer1_out[203];
    assign layer2_out[7657] = layer1_out[2280];
    assign layer2_out[7658] = layer1_out[5677] & ~layer1_out[5678];
    assign layer2_out[7659] = layer1_out[4744] & ~layer1_out[4743];
    assign layer2_out[7660] = layer1_out[3645];
    assign layer2_out[7661] = ~(layer1_out[5425] | layer1_out[5426]);
    assign layer2_out[7662] = layer1_out[785];
    assign layer2_out[7663] = layer1_out[920] ^ layer1_out[921];
    assign layer2_out[7664] = ~layer1_out[3032];
    assign layer2_out[7665] = ~layer1_out[7957];
    assign layer2_out[7666] = ~(layer1_out[7461] ^ layer1_out[7462]);
    assign layer2_out[7667] = ~layer1_out[7330];
    assign layer2_out[7668] = layer1_out[5960] & ~layer1_out[5959];
    assign layer2_out[7669] = layer1_out[7236];
    assign layer2_out[7670] = ~layer1_out[3808];
    assign layer2_out[7671] = ~layer1_out[3976] | layer1_out[3975];
    assign layer2_out[7672] = ~(layer1_out[321] | layer1_out[322]);
    assign layer2_out[7673] = layer1_out[1586] ^ layer1_out[1587];
    assign layer2_out[7674] = layer1_out[6760];
    assign layer2_out[7675] = ~layer1_out[7519];
    assign layer2_out[7676] = layer1_out[983] | layer1_out[984];
    assign layer2_out[7677] = ~layer1_out[2094];
    assign layer2_out[7678] = layer1_out[7729];
    assign layer2_out[7679] = layer1_out[1959];
    assign layer2_out[7680] = ~layer1_out[6417] | layer1_out[6418];
    assign layer2_out[7681] = layer1_out[4050] | layer1_out[4051];
    assign layer2_out[7682] = layer1_out[4249] & layer1_out[4250];
    assign layer2_out[7683] = ~layer1_out[7467] | layer1_out[7466];
    assign layer2_out[7684] = layer1_out[1804];
    assign layer2_out[7685] = ~layer1_out[2551];
    assign layer2_out[7686] = layer1_out[2576] & ~layer1_out[2575];
    assign layer2_out[7687] = ~(layer1_out[6961] & layer1_out[6962]);
    assign layer2_out[7688] = ~layer1_out[164];
    assign layer2_out[7689] = layer1_out[1123] & layer1_out[1124];
    assign layer2_out[7690] = ~(layer1_out[6005] ^ layer1_out[6006]);
    assign layer2_out[7691] = layer1_out[3475];
    assign layer2_out[7692] = layer1_out[322];
    assign layer2_out[7693] = 1'b1;
    assign layer2_out[7694] = ~(layer1_out[6141] | layer1_out[6142]);
    assign layer2_out[7695] = ~(layer1_out[2498] & layer1_out[2499]);
    assign layer2_out[7696] = ~(layer1_out[6239] & layer1_out[6240]);
    assign layer2_out[7697] = ~(layer1_out[6821] & layer1_out[6822]);
    assign layer2_out[7698] = ~(layer1_out[4560] | layer1_out[4561]);
    assign layer2_out[7699] = layer1_out[2017] & layer1_out[2018];
    assign layer2_out[7700] = ~layer1_out[823];
    assign layer2_out[7701] = ~layer1_out[6465] | layer1_out[6466];
    assign layer2_out[7702] = layer1_out[967] ^ layer1_out[968];
    assign layer2_out[7703] = ~(layer1_out[1488] | layer1_out[1489]);
    assign layer2_out[7704] = layer1_out[7565];
    assign layer2_out[7705] = layer1_out[4891];
    assign layer2_out[7706] = layer1_out[6454] ^ layer1_out[6455];
    assign layer2_out[7707] = layer1_out[3389] & layer1_out[3390];
    assign layer2_out[7708] = layer1_out[2519];
    assign layer2_out[7709] = layer1_out[6146] | layer1_out[6147];
    assign layer2_out[7710] = ~layer1_out[6009];
    assign layer2_out[7711] = ~layer1_out[3852] | layer1_out[3851];
    assign layer2_out[7712] = layer1_out[3004];
    assign layer2_out[7713] = ~layer1_out[1180];
    assign layer2_out[7714] = ~layer1_out[2882];
    assign layer2_out[7715] = ~layer1_out[2226] | layer1_out[2227];
    assign layer2_out[7716] = ~(layer1_out[7631] & layer1_out[7632]);
    assign layer2_out[7717] = ~layer1_out[885] | layer1_out[884];
    assign layer2_out[7718] = layer1_out[6074] & ~layer1_out[6073];
    assign layer2_out[7719] = ~layer1_out[3138];
    assign layer2_out[7720] = ~(layer1_out[2649] & layer1_out[2650]);
    assign layer2_out[7721] = ~layer1_out[7828];
    assign layer2_out[7722] = ~layer1_out[4452];
    assign layer2_out[7723] = ~layer1_out[5109];
    assign layer2_out[7724] = ~layer1_out[4517] | layer1_out[4518];
    assign layer2_out[7725] = layer1_out[1728] & ~layer1_out[1729];
    assign layer2_out[7726] = ~layer1_out[5942];
    assign layer2_out[7727] = ~layer1_out[4167];
    assign layer2_out[7728] = layer1_out[2846] & layer1_out[2847];
    assign layer2_out[7729] = layer1_out[3393];
    assign layer2_out[7730] = layer1_out[922];
    assign layer2_out[7731] = ~layer1_out[5147] | layer1_out[5146];
    assign layer2_out[7732] = layer1_out[2337] & ~layer1_out[2338];
    assign layer2_out[7733] = layer1_out[1416] & ~layer1_out[1417];
    assign layer2_out[7734] = layer1_out[4776] & layer1_out[4777];
    assign layer2_out[7735] = layer1_out[3360];
    assign layer2_out[7736] = ~layer1_out[3893];
    assign layer2_out[7737] = ~layer1_out[7082] | layer1_out[7081];
    assign layer2_out[7738] = ~(layer1_out[6390] & layer1_out[6391]);
    assign layer2_out[7739] = layer1_out[4531];
    assign layer2_out[7740] = ~(layer1_out[6292] | layer1_out[6293]);
    assign layer2_out[7741] = ~layer1_out[2201] | layer1_out[2200];
    assign layer2_out[7742] = ~layer1_out[81];
    assign layer2_out[7743] = ~layer1_out[4929];
    assign layer2_out[7744] = layer1_out[6766] & ~layer1_out[6765];
    assign layer2_out[7745] = layer1_out[3007] & ~layer1_out[3006];
    assign layer2_out[7746] = ~layer1_out[2101];
    assign layer2_out[7747] = layer1_out[1319];
    assign layer2_out[7748] = layer1_out[2139] & ~layer1_out[2138];
    assign layer2_out[7749] = layer1_out[1357] | layer1_out[1358];
    assign layer2_out[7750] = layer1_out[1082] ^ layer1_out[1083];
    assign layer2_out[7751] = ~layer1_out[2314];
    assign layer2_out[7752] = layer1_out[1664];
    assign layer2_out[7753] = ~(layer1_out[7944] & layer1_out[7945]);
    assign layer2_out[7754] = ~layer1_out[2417] | layer1_out[2416];
    assign layer2_out[7755] = ~layer1_out[3863] | layer1_out[3864];
    assign layer2_out[7756] = ~layer1_out[4306];
    assign layer2_out[7757] = ~layer1_out[6107];
    assign layer2_out[7758] = ~(layer1_out[7702] ^ layer1_out[7703]);
    assign layer2_out[7759] = layer1_out[6687] & ~layer1_out[6686];
    assign layer2_out[7760] = layer1_out[2166] | layer1_out[2167];
    assign layer2_out[7761] = ~(layer1_out[855] & layer1_out[856]);
    assign layer2_out[7762] = layer1_out[1198];
    assign layer2_out[7763] = layer1_out[812];
    assign layer2_out[7764] = layer1_out[1320];
    assign layer2_out[7765] = layer1_out[3025] | layer1_out[3026];
    assign layer2_out[7766] = ~(layer1_out[797] & layer1_out[798]);
    assign layer2_out[7767] = 1'b0;
    assign layer2_out[7768] = layer1_out[3597] ^ layer1_out[3598];
    assign layer2_out[7769] = layer1_out[2664] & layer1_out[2665];
    assign layer2_out[7770] = 1'b0;
    assign layer2_out[7771] = ~(layer1_out[4450] & layer1_out[4451]);
    assign layer2_out[7772] = ~layer1_out[535];
    assign layer2_out[7773] = layer1_out[1589] & ~layer1_out[1588];
    assign layer2_out[7774] = ~layer1_out[1373];
    assign layer2_out[7775] = ~layer1_out[3856];
    assign layer2_out[7776] = layer1_out[4946] & ~layer1_out[4945];
    assign layer2_out[7777] = ~layer1_out[1075];
    assign layer2_out[7778] = 1'b1;
    assign layer2_out[7779] = layer1_out[418] & ~layer1_out[419];
    assign layer2_out[7780] = layer1_out[515] & layer1_out[516];
    assign layer2_out[7781] = 1'b0;
    assign layer2_out[7782] = ~(layer1_out[5067] | layer1_out[5068]);
    assign layer2_out[7783] = ~layer1_out[2155];
    assign layer2_out[7784] = layer1_out[6601] ^ layer1_out[6602];
    assign layer2_out[7785] = 1'b1;
    assign layer2_out[7786] = layer1_out[3861] & ~layer1_out[3860];
    assign layer2_out[7787] = 1'b0;
    assign layer2_out[7788] = layer1_out[901] | layer1_out[902];
    assign layer2_out[7789] = ~layer1_out[3467];
    assign layer2_out[7790] = ~layer1_out[7209] | layer1_out[7208];
    assign layer2_out[7791] = layer1_out[5988];
    assign layer2_out[7792] = layer1_out[3912] & layer1_out[3913];
    assign layer2_out[7793] = layer1_out[6442] & ~layer1_out[6441];
    assign layer2_out[7794] = layer1_out[3812] & ~layer1_out[3813];
    assign layer2_out[7795] = ~(layer1_out[5433] & layer1_out[5434]);
    assign layer2_out[7796] = ~layer1_out[3606];
    assign layer2_out[7797] = ~layer1_out[1158];
    assign layer2_out[7798] = layer1_out[3948];
    assign layer2_out[7799] = layer1_out[2064];
    assign layer2_out[7800] = ~layer1_out[7448] | layer1_out[7449];
    assign layer2_out[7801] = layer1_out[2202] & ~layer1_out[2201];
    assign layer2_out[7802] = layer1_out[5504];
    assign layer2_out[7803] = layer1_out[3933] & ~layer1_out[3932];
    assign layer2_out[7804] = ~layer1_out[7752];
    assign layer2_out[7805] = ~layer1_out[6461];
    assign layer2_out[7806] = ~layer1_out[3762] | layer1_out[3761];
    assign layer2_out[7807] = layer1_out[3299] & layer1_out[3300];
    assign layer2_out[7808] = layer1_out[1972] | layer1_out[1973];
    assign layer2_out[7809] = layer1_out[5290] & layer1_out[5291];
    assign layer2_out[7810] = layer1_out[4350];
    assign layer2_out[7811] = layer1_out[2244] & layer1_out[2245];
    assign layer2_out[7812] = ~layer1_out[561] | layer1_out[562];
    assign layer2_out[7813] = layer1_out[3202];
    assign layer2_out[7814] = layer1_out[5894] & layer1_out[5895];
    assign layer2_out[7815] = ~(layer1_out[1181] & layer1_out[1182]);
    assign layer2_out[7816] = ~layer1_out[3545];
    assign layer2_out[7817] = layer1_out[506] & layer1_out[507];
    assign layer2_out[7818] = 1'b1;
    assign layer2_out[7819] = ~layer1_out[4284] | layer1_out[4283];
    assign layer2_out[7820] = layer1_out[4645];
    assign layer2_out[7821] = ~layer1_out[423] | layer1_out[424];
    assign layer2_out[7822] = ~(layer1_out[5772] ^ layer1_out[5773]);
    assign layer2_out[7823] = ~layer1_out[640];
    assign layer2_out[7824] = layer1_out[3222] | layer1_out[3223];
    assign layer2_out[7825] = ~(layer1_out[7599] & layer1_out[7600]);
    assign layer2_out[7826] = layer1_out[7240] & ~layer1_out[7241];
    assign layer2_out[7827] = ~layer1_out[4507] | layer1_out[4508];
    assign layer2_out[7828] = ~layer1_out[5348];
    assign layer2_out[7829] = ~layer1_out[6647];
    assign layer2_out[7830] = layer1_out[4976] & ~layer1_out[4977];
    assign layer2_out[7831] = layer1_out[4821] & ~layer1_out[4820];
    assign layer2_out[7832] = 1'b0;
    assign layer2_out[7833] = ~(layer1_out[589] ^ layer1_out[590]);
    assign layer2_out[7834] = ~layer1_out[2457];
    assign layer2_out[7835] = ~layer1_out[66];
    assign layer2_out[7836] = layer1_out[1792] & ~layer1_out[1791];
    assign layer2_out[7837] = layer1_out[4435] & ~layer1_out[4436];
    assign layer2_out[7838] = ~layer1_out[7779] | layer1_out[7780];
    assign layer2_out[7839] = ~(layer1_out[4003] | layer1_out[4004]);
    assign layer2_out[7840] = ~layer1_out[6812];
    assign layer2_out[7841] = layer1_out[2452] ^ layer1_out[2453];
    assign layer2_out[7842] = ~(layer1_out[7414] | layer1_out[7415]);
    assign layer2_out[7843] = ~(layer1_out[2972] | layer1_out[2973]);
    assign layer2_out[7844] = layer1_out[6720];
    assign layer2_out[7845] = ~(layer1_out[1696] ^ layer1_out[1697]);
    assign layer2_out[7846] = layer1_out[7495] | layer1_out[7496];
    assign layer2_out[7847] = ~(layer1_out[1815] | layer1_out[1816]);
    assign layer2_out[7848] = layer1_out[2630] & ~layer1_out[2629];
    assign layer2_out[7849] = layer1_out[6325] & ~layer1_out[6326];
    assign layer2_out[7850] = layer1_out[6992] | layer1_out[6993];
    assign layer2_out[7851] = layer1_out[1158];
    assign layer2_out[7852] = ~(layer1_out[6233] & layer1_out[6234]);
    assign layer2_out[7853] = layer1_out[5652] & layer1_out[5653];
    assign layer2_out[7854] = ~(layer1_out[7239] | layer1_out[7240]);
    assign layer2_out[7855] = layer1_out[7247];
    assign layer2_out[7856] = layer1_out[3087] & layer1_out[3088];
    assign layer2_out[7857] = ~(layer1_out[4136] | layer1_out[4137]);
    assign layer2_out[7858] = ~layer1_out[1061];
    assign layer2_out[7859] = layer1_out[5030];
    assign layer2_out[7860] = layer1_out[6762] & ~layer1_out[6763];
    assign layer2_out[7861] = layer1_out[5660] & layer1_out[5661];
    assign layer2_out[7862] = layer1_out[1992] & ~layer1_out[1993];
    assign layer2_out[7863] = layer1_out[2168];
    assign layer2_out[7864] = layer1_out[5128];
    assign layer2_out[7865] = ~(layer1_out[3003] ^ layer1_out[3004]);
    assign layer2_out[7866] = ~layer1_out[6628];
    assign layer2_out[7867] = layer1_out[1171];
    assign layer2_out[7868] = ~layer1_out[6527];
    assign layer2_out[7869] = layer1_out[5371];
    assign layer2_out[7870] = layer1_out[399];
    assign layer2_out[7871] = layer1_out[5968] & ~layer1_out[5969];
    assign layer2_out[7872] = ~layer1_out[7390] | layer1_out[7391];
    assign layer2_out[7873] = layer1_out[6333] & ~layer1_out[6332];
    assign layer2_out[7874] = layer1_out[6826] & layer1_out[6827];
    assign layer2_out[7875] = layer1_out[4202] | layer1_out[4203];
    assign layer2_out[7876] = layer1_out[3992] ^ layer1_out[3993];
    assign layer2_out[7877] = ~(layer1_out[603] & layer1_out[604]);
    assign layer2_out[7878] = layer1_out[571] & ~layer1_out[570];
    assign layer2_out[7879] = ~layer1_out[6471] | layer1_out[6472];
    assign layer2_out[7880] = layer1_out[1322];
    assign layer2_out[7881] = ~layer1_out[3364];
    assign layer2_out[7882] = ~layer1_out[4377] | layer1_out[4378];
    assign layer2_out[7883] = ~layer1_out[4247] | layer1_out[4246];
    assign layer2_out[7884] = ~layer1_out[5585];
    assign layer2_out[7885] = ~(layer1_out[788] & layer1_out[789]);
    assign layer2_out[7886] = layer1_out[88] & ~layer1_out[89];
    assign layer2_out[7887] = layer1_out[7544] | layer1_out[7545];
    assign layer2_out[7888] = ~(layer1_out[6433] ^ layer1_out[6434]);
    assign layer2_out[7889] = ~(layer1_out[3697] | layer1_out[3698]);
    assign layer2_out[7890] = layer1_out[3902];
    assign layer2_out[7891] = layer1_out[3046];
    assign layer2_out[7892] = ~layer1_out[4027];
    assign layer2_out[7893] = 1'b0;
    assign layer2_out[7894] = layer1_out[1152];
    assign layer2_out[7895] = layer1_out[2521] & ~layer1_out[2522];
    assign layer2_out[7896] = layer1_out[876] & ~layer1_out[875];
    assign layer2_out[7897] = layer1_out[1636] & layer1_out[1637];
    assign layer2_out[7898] = ~(layer1_out[2669] & layer1_out[2670]);
    assign layer2_out[7899] = layer1_out[2562] ^ layer1_out[2563];
    assign layer2_out[7900] = layer1_out[1716] & layer1_out[1717];
    assign layer2_out[7901] = layer1_out[3602] & layer1_out[3603];
    assign layer2_out[7902] = 1'b1;
    assign layer2_out[7903] = layer1_out[2517] ^ layer1_out[2518];
    assign layer2_out[7904] = ~(layer1_out[2621] | layer1_out[2622]);
    assign layer2_out[7905] = ~layer1_out[1614] | layer1_out[1615];
    assign layer2_out[7906] = layer1_out[5829] | layer1_out[5830];
    assign layer2_out[7907] = ~layer1_out[3673];
    assign layer2_out[7908] = layer1_out[5258] | layer1_out[5259];
    assign layer2_out[7909] = 1'b0;
    assign layer2_out[7910] = layer1_out[7973];
    assign layer2_out[7911] = ~(layer1_out[1468] | layer1_out[1469]);
    assign layer2_out[7912] = layer1_out[4673] ^ layer1_out[4674];
    assign layer2_out[7913] = ~(layer1_out[809] | layer1_out[810]);
    assign layer2_out[7914] = layer1_out[6163] & ~layer1_out[6164];
    assign layer2_out[7915] = layer1_out[7858] | layer1_out[7859];
    assign layer2_out[7916] = layer1_out[3077];
    assign layer2_out[7917] = ~(layer1_out[602] | layer1_out[603]);
    assign layer2_out[7918] = ~layer1_out[1573];
    assign layer2_out[7919] = ~(layer1_out[712] | layer1_out[713]);
    assign layer2_out[7920] = layer1_out[6571] & ~layer1_out[6572];
    assign layer2_out[7921] = layer1_out[5821] | layer1_out[5822];
    assign layer2_out[7922] = ~layer1_out[5134];
    assign layer2_out[7923] = layer1_out[5605] ^ layer1_out[5606];
    assign layer2_out[7924] = ~layer1_out[5750] | layer1_out[5751];
    assign layer2_out[7925] = ~(layer1_out[384] ^ layer1_out[385]);
    assign layer2_out[7926] = ~(layer1_out[5850] | layer1_out[5851]);
    assign layer2_out[7927] = ~layer1_out[4696];
    assign layer2_out[7928] = ~layer1_out[1366] | layer1_out[1365];
    assign layer2_out[7929] = layer1_out[6489] & layer1_out[6490];
    assign layer2_out[7930] = layer1_out[3617];
    assign layer2_out[7931] = ~layer1_out[2017] | layer1_out[2016];
    assign layer2_out[7932] = layer1_out[4927] & ~layer1_out[4926];
    assign layer2_out[7933] = layer1_out[5903];
    assign layer2_out[7934] = ~(layer1_out[2216] | layer1_out[2217]);
    assign layer2_out[7935] = layer1_out[3246] | layer1_out[3247];
    assign layer2_out[7936] = layer1_out[5019];
    assign layer2_out[7937] = ~layer1_out[3510];
    assign layer2_out[7938] = ~layer1_out[5862] | layer1_out[5861];
    assign layer2_out[7939] = layer1_out[655] | layer1_out[656];
    assign layer2_out[7940] = 1'b0;
    assign layer2_out[7941] = ~layer1_out[2496];
    assign layer2_out[7942] = layer1_out[727];
    assign layer2_out[7943] = ~layer1_out[4731];
    assign layer2_out[7944] = ~layer1_out[3178];
    assign layer2_out[7945] = ~(layer1_out[2955] & layer1_out[2956]);
    assign layer2_out[7946] = layer1_out[1427];
    assign layer2_out[7947] = ~layer1_out[1139];
    assign layer2_out[7948] = ~(layer1_out[4101] | layer1_out[4102]);
    assign layer2_out[7949] = ~layer1_out[7322];
    assign layer2_out[7950] = ~layer1_out[6131];
    assign layer2_out[7951] = layer1_out[4762];
    assign layer2_out[7952] = layer1_out[7924] & ~layer1_out[7925];
    assign layer2_out[7953] = layer1_out[6355] & layer1_out[6356];
    assign layer2_out[7954] = layer1_out[4017];
    assign layer2_out[7955] = ~layer1_out[3447];
    assign layer2_out[7956] = layer1_out[6397] ^ layer1_out[6398];
    assign layer2_out[7957] = ~layer1_out[5302];
    assign layer2_out[7958] = ~(layer1_out[4367] & layer1_out[4368]);
    assign layer2_out[7959] = ~(layer1_out[4627] ^ layer1_out[4628]);
    assign layer2_out[7960] = ~(layer1_out[5808] & layer1_out[5809]);
    assign layer2_out[7961] = 1'b1;
    assign layer2_out[7962] = ~layer1_out[5540];
    assign layer2_out[7963] = layer1_out[6172];
    assign layer2_out[7964] = layer1_out[3735] ^ layer1_out[3736];
    assign layer2_out[7965] = 1'b1;
    assign layer2_out[7966] = ~layer1_out[461] | layer1_out[460];
    assign layer2_out[7967] = ~layer1_out[300];
    assign layer2_out[7968] = ~layer1_out[3629] | layer1_out[3628];
    assign layer2_out[7969] = ~layer1_out[3766] | layer1_out[3767];
    assign layer2_out[7970] = ~(layer1_out[187] & layer1_out[188]);
    assign layer2_out[7971] = ~layer1_out[508];
    assign layer2_out[7972] = ~layer1_out[7265] | layer1_out[7266];
    assign layer2_out[7973] = ~layer1_out[2246];
    assign layer2_out[7974] = layer1_out[5253] & ~layer1_out[5252];
    assign layer2_out[7975] = ~(layer1_out[4334] & layer1_out[4335]);
    assign layer2_out[7976] = layer1_out[40];
    assign layer2_out[7977] = layer1_out[3820] & ~layer1_out[3819];
    assign layer2_out[7978] = ~(layer1_out[2225] & layer1_out[2226]);
    assign layer2_out[7979] = 1'b0;
    assign layer2_out[7980] = layer1_out[3693] | layer1_out[3694];
    assign layer2_out[7981] = ~(layer1_out[4937] ^ layer1_out[4938]);
    assign layer2_out[7982] = ~layer1_out[5980] | layer1_out[5981];
    assign layer2_out[7983] = layer1_out[6261];
    assign layer2_out[7984] = ~(layer1_out[3371] | layer1_out[3372]);
    assign layer2_out[7985] = layer1_out[949] & layer1_out[950];
    assign layer2_out[7986] = layer1_out[7148] | layer1_out[7149];
    assign layer2_out[7987] = layer1_out[6250];
    assign layer2_out[7988] = ~(layer1_out[2432] | layer1_out[2433]);
    assign layer2_out[7989] = layer1_out[5721] & ~layer1_out[5722];
    assign layer2_out[7990] = ~layer1_out[532];
    assign layer2_out[7991] = ~(layer1_out[3565] ^ layer1_out[3566]);
    assign layer2_out[7992] = 1'b0;
    assign layer2_out[7993] = ~layer1_out[1030];
    assign layer2_out[7994] = layer1_out[4960];
    assign layer2_out[7995] = layer1_out[7139] & ~layer1_out[7140];
    assign layer2_out[7996] = layer1_out[3437] | layer1_out[3438];
    assign layer2_out[7997] = layer1_out[595];
    assign layer2_out[7998] = ~(layer1_out[7900] & layer1_out[7901]);
    assign layer2_out[7999] = layer1_out[6221];
    assign layer3_out[0] = ~layer2_out[6022] | layer2_out[6021];
    assign layer3_out[1] = ~(layer2_out[6132] & layer2_out[6133]);
    assign layer3_out[2] = ~layer2_out[6080] | layer2_out[6081];
    assign layer3_out[3] = ~(layer2_out[271] ^ layer2_out[272]);
    assign layer3_out[4] = ~layer2_out[5951];
    assign layer3_out[5] = ~layer2_out[3519];
    assign layer3_out[6] = ~layer2_out[2936];
    assign layer3_out[7] = ~layer2_out[1664];
    assign layer3_out[8] = layer2_out[7286];
    assign layer3_out[9] = ~layer2_out[6222];
    assign layer3_out[10] = 1'b0;
    assign layer3_out[11] = ~(layer2_out[4722] | layer2_out[4723]);
    assign layer3_out[12] = 1'b0;
    assign layer3_out[13] = layer2_out[6346] & layer2_out[6347];
    assign layer3_out[14] = layer2_out[3338];
    assign layer3_out[15] = layer2_out[3842] & ~layer2_out[3841];
    assign layer3_out[16] = ~layer2_out[2908];
    assign layer3_out[17] = ~(layer2_out[4853] ^ layer2_out[4854]);
    assign layer3_out[18] = layer2_out[5117] | layer2_out[5118];
    assign layer3_out[19] = ~layer2_out[1645];
    assign layer3_out[20] = ~layer2_out[1234];
    assign layer3_out[21] = ~layer2_out[2549];
    assign layer3_out[22] = layer2_out[6650];
    assign layer3_out[23] = layer2_out[2418];
    assign layer3_out[24] = ~layer2_out[4258];
    assign layer3_out[25] = ~layer2_out[882] | layer2_out[881];
    assign layer3_out[26] = ~(layer2_out[6094] | layer2_out[6095]);
    assign layer3_out[27] = ~(layer2_out[5491] ^ layer2_out[5492]);
    assign layer3_out[28] = layer2_out[627];
    assign layer3_out[29] = ~layer2_out[513];
    assign layer3_out[30] = ~layer2_out[1669];
    assign layer3_out[31] = ~layer2_out[4118] | layer2_out[4117];
    assign layer3_out[32] = 1'b1;
    assign layer3_out[33] = layer2_out[1782];
    assign layer3_out[34] = layer2_out[4356];
    assign layer3_out[35] = ~(layer2_out[2975] | layer2_out[2976]);
    assign layer3_out[36] = ~(layer2_out[3356] | layer2_out[3357]);
    assign layer3_out[37] = ~layer2_out[7562];
    assign layer3_out[38] = ~layer2_out[1913] | layer2_out[1914];
    assign layer3_out[39] = ~layer2_out[6436];
    assign layer3_out[40] = ~layer2_out[5704] | layer2_out[5705];
    assign layer3_out[41] = layer2_out[2460];
    assign layer3_out[42] = ~(layer2_out[3937] | layer2_out[3938]);
    assign layer3_out[43] = layer2_out[139] | layer2_out[140];
    assign layer3_out[44] = 1'b0;
    assign layer3_out[45] = ~layer2_out[7135];
    assign layer3_out[46] = layer2_out[6887];
    assign layer3_out[47] = layer2_out[3135];
    assign layer3_out[48] = layer2_out[2295];
    assign layer3_out[49] = ~layer2_out[7322];
    assign layer3_out[50] = ~layer2_out[2403];
    assign layer3_out[51] = ~layer2_out[6462];
    assign layer3_out[52] = ~(layer2_out[4148] & layer2_out[4149]);
    assign layer3_out[53] = ~layer2_out[3508];
    assign layer3_out[54] = layer2_out[1355] ^ layer2_out[1356];
    assign layer3_out[55] = layer2_out[77];
    assign layer3_out[56] = layer2_out[1467];
    assign layer3_out[57] = ~layer2_out[6879];
    assign layer3_out[58] = ~layer2_out[6529];
    assign layer3_out[59] = layer2_out[774] & ~layer2_out[773];
    assign layer3_out[60] = layer2_out[3408];
    assign layer3_out[61] = ~layer2_out[2767] | layer2_out[2768];
    assign layer3_out[62] = 1'b1;
    assign layer3_out[63] = ~layer2_out[3592] | layer2_out[3591];
    assign layer3_out[64] = layer2_out[4488] ^ layer2_out[4489];
    assign layer3_out[65] = ~(layer2_out[3687] ^ layer2_out[3688]);
    assign layer3_out[66] = ~layer2_out[517];
    assign layer3_out[67] = layer2_out[138];
    assign layer3_out[68] = ~(layer2_out[3572] ^ layer2_out[3573]);
    assign layer3_out[69] = ~(layer2_out[4650] ^ layer2_out[4651]);
    assign layer3_out[70] = layer2_out[4317];
    assign layer3_out[71] = 1'b0;
    assign layer3_out[72] = layer2_out[7461];
    assign layer3_out[73] = layer2_out[5417];
    assign layer3_out[74] = layer2_out[3310] & ~layer2_out[3311];
    assign layer3_out[75] = layer2_out[5061] ^ layer2_out[5062];
    assign layer3_out[76] = layer2_out[2448] & layer2_out[2449];
    assign layer3_out[77] = ~(layer2_out[4352] & layer2_out[4353]);
    assign layer3_out[78] = layer2_out[1975];
    assign layer3_out[79] = layer2_out[194] & ~layer2_out[195];
    assign layer3_out[80] = layer2_out[6216];
    assign layer3_out[81] = ~(layer2_out[7205] | layer2_out[7206]);
    assign layer3_out[82] = layer2_out[19];
    assign layer3_out[83] = ~layer2_out[6190];
    assign layer3_out[84] = ~layer2_out[682];
    assign layer3_out[85] = layer2_out[575] & ~layer2_out[576];
    assign layer3_out[86] = ~layer2_out[1836] | layer2_out[1837];
    assign layer3_out[87] = ~layer2_out[7037] | layer2_out[7038];
    assign layer3_out[88] = ~(layer2_out[849] ^ layer2_out[850]);
    assign layer3_out[89] = ~layer2_out[1632];
    assign layer3_out[90] = ~(layer2_out[3366] & layer2_out[3367]);
    assign layer3_out[91] = ~layer2_out[1643];
    assign layer3_out[92] = ~layer2_out[1966];
    assign layer3_out[93] = layer2_out[1085] & ~layer2_out[1086];
    assign layer3_out[94] = layer2_out[6924] ^ layer2_out[6925];
    assign layer3_out[95] = ~layer2_out[2788];
    assign layer3_out[96] = layer2_out[5580] & layer2_out[5581];
    assign layer3_out[97] = ~layer2_out[4998] | layer2_out[4997];
    assign layer3_out[98] = layer2_out[5610] ^ layer2_out[5611];
    assign layer3_out[99] = ~layer2_out[7590] | layer2_out[7589];
    assign layer3_out[100] = layer2_out[5527];
    assign layer3_out[101] = layer2_out[5248];
    assign layer3_out[102] = layer2_out[537];
    assign layer3_out[103] = ~layer2_out[3685];
    assign layer3_out[104] = layer2_out[538] & layer2_out[539];
    assign layer3_out[105] = layer2_out[2638];
    assign layer3_out[106] = ~layer2_out[3707];
    assign layer3_out[107] = layer2_out[2606];
    assign layer3_out[108] = layer2_out[3073] ^ layer2_out[3074];
    assign layer3_out[109] = ~layer2_out[2504];
    assign layer3_out[110] = ~(layer2_out[1980] & layer2_out[1981]);
    assign layer3_out[111] = layer2_out[5180];
    assign layer3_out[112] = layer2_out[2701];
    assign layer3_out[113] = layer2_out[3264];
    assign layer3_out[114] = layer2_out[6418];
    assign layer3_out[115] = layer2_out[6220] & ~layer2_out[6219];
    assign layer3_out[116] = ~(layer2_out[6116] ^ layer2_out[6117]);
    assign layer3_out[117] = layer2_out[5300] & layer2_out[5301];
    assign layer3_out[118] = layer2_out[2839] | layer2_out[2840];
    assign layer3_out[119] = ~(layer2_out[5656] & layer2_out[5657]);
    assign layer3_out[120] = layer2_out[6777];
    assign layer3_out[121] = ~(layer2_out[7703] | layer2_out[7704]);
    assign layer3_out[122] = ~layer2_out[6837];
    assign layer3_out[123] = layer2_out[977] & layer2_out[978];
    assign layer3_out[124] = ~layer2_out[1215];
    assign layer3_out[125] = ~(layer2_out[4593] ^ layer2_out[4594]);
    assign layer3_out[126] = ~layer2_out[7336];
    assign layer3_out[127] = ~layer2_out[7497];
    assign layer3_out[128] = ~(layer2_out[7799] | layer2_out[7800]);
    assign layer3_out[129] = ~layer2_out[3317];
    assign layer3_out[130] = ~layer2_out[5945] | layer2_out[5946];
    assign layer3_out[131] = layer2_out[7686] | layer2_out[7687];
    assign layer3_out[132] = ~(layer2_out[6817] & layer2_out[6818]);
    assign layer3_out[133] = layer2_out[4282] & ~layer2_out[4283];
    assign layer3_out[134] = layer2_out[7963];
    assign layer3_out[135] = ~(layer2_out[7185] & layer2_out[7186]);
    assign layer3_out[136] = layer2_out[6051];
    assign layer3_out[137] = ~layer2_out[604] | layer2_out[603];
    assign layer3_out[138] = layer2_out[6779] & ~layer2_out[6778];
    assign layer3_out[139] = layer2_out[7476];
    assign layer3_out[140] = layer2_out[989] | layer2_out[990];
    assign layer3_out[141] = layer2_out[2891];
    assign layer3_out[142] = layer2_out[4835];
    assign layer3_out[143] = 1'b0;
    assign layer3_out[144] = ~layer2_out[7233];
    assign layer3_out[145] = layer2_out[7910] | layer2_out[7911];
    assign layer3_out[146] = layer2_out[5258];
    assign layer3_out[147] = layer2_out[6474] & ~layer2_out[6473];
    assign layer3_out[148] = ~layer2_out[6860];
    assign layer3_out[149] = layer2_out[7482] & ~layer2_out[7481];
    assign layer3_out[150] = ~(layer2_out[2879] & layer2_out[2880]);
    assign layer3_out[151] = ~(layer2_out[402] ^ layer2_out[403]);
    assign layer3_out[152] = ~layer2_out[2323] | layer2_out[2324];
    assign layer3_out[153] = ~layer2_out[775] | layer2_out[774];
    assign layer3_out[154] = ~layer2_out[5591] | layer2_out[5590];
    assign layer3_out[155] = ~(layer2_out[1772] | layer2_out[1773]);
    assign layer3_out[156] = layer2_out[335] & layer2_out[336];
    assign layer3_out[157] = layer2_out[2192] ^ layer2_out[2193];
    assign layer3_out[158] = ~(layer2_out[5048] ^ layer2_out[5049]);
    assign layer3_out[159] = ~(layer2_out[1323] ^ layer2_out[1324]);
    assign layer3_out[160] = ~(layer2_out[1739] | layer2_out[1740]);
    assign layer3_out[161] = layer2_out[1013] & ~layer2_out[1012];
    assign layer3_out[162] = layer2_out[6862] & ~layer2_out[6863];
    assign layer3_out[163] = layer2_out[5447];
    assign layer3_out[164] = layer2_out[6096];
    assign layer3_out[165] = ~(layer2_out[3601] | layer2_out[3602]);
    assign layer3_out[166] = ~(layer2_out[1517] ^ layer2_out[1518]);
    assign layer3_out[167] = layer2_out[3512] & ~layer2_out[3513];
    assign layer3_out[168] = layer2_out[4145] ^ layer2_out[4146];
    assign layer3_out[169] = layer2_out[700];
    assign layer3_out[170] = ~layer2_out[4173];
    assign layer3_out[171] = ~layer2_out[4391];
    assign layer3_out[172] = layer2_out[7979] & ~layer2_out[7980];
    assign layer3_out[173] = layer2_out[4010];
    assign layer3_out[174] = layer2_out[1122] & ~layer2_out[1121];
    assign layer3_out[175] = layer2_out[3219] & ~layer2_out[3220];
    assign layer3_out[176] = ~(layer2_out[1372] | layer2_out[1373]);
    assign layer3_out[177] = ~layer2_out[7649];
    assign layer3_out[178] = ~layer2_out[1522];
    assign layer3_out[179] = ~layer2_out[4012];
    assign layer3_out[180] = ~layer2_out[4141];
    assign layer3_out[181] = layer2_out[1495];
    assign layer3_out[182] = ~(layer2_out[2334] ^ layer2_out[2335]);
    assign layer3_out[183] = layer2_out[3339];
    assign layer3_out[184] = layer2_out[5812];
    assign layer3_out[185] = layer2_out[623] | layer2_out[624];
    assign layer3_out[186] = ~layer2_out[2094];
    assign layer3_out[187] = layer2_out[2905] & layer2_out[2906];
    assign layer3_out[188] = ~layer2_out[1716];
    assign layer3_out[189] = ~(layer2_out[3568] ^ layer2_out[3569]);
    assign layer3_out[190] = ~(layer2_out[1303] & layer2_out[1304]);
    assign layer3_out[191] = layer2_out[2440];
    assign layer3_out[192] = layer2_out[373];
    assign layer3_out[193] = ~layer2_out[3883];
    assign layer3_out[194] = layer2_out[88] & layer2_out[89];
    assign layer3_out[195] = layer2_out[2964] ^ layer2_out[2965];
    assign layer3_out[196] = layer2_out[46] & ~layer2_out[47];
    assign layer3_out[197] = layer2_out[5777];
    assign layer3_out[198] = 1'b0;
    assign layer3_out[199] = layer2_out[5201] & ~layer2_out[5200];
    assign layer3_out[200] = layer2_out[5811] ^ layer2_out[5812];
    assign layer3_out[201] = ~layer2_out[4528] | layer2_out[4529];
    assign layer3_out[202] = layer2_out[1201];
    assign layer3_out[203] = ~layer2_out[5567];
    assign layer3_out[204] = layer2_out[7810] | layer2_out[7811];
    assign layer3_out[205] = layer2_out[6197];
    assign layer3_out[206] = layer2_out[2058] & ~layer2_out[2057];
    assign layer3_out[207] = layer2_out[2998];
    assign layer3_out[208] = ~(layer2_out[7778] ^ layer2_out[7779]);
    assign layer3_out[209] = ~layer2_out[2864];
    assign layer3_out[210] = layer2_out[1389];
    assign layer3_out[211] = ~(layer2_out[893] & layer2_out[894]);
    assign layer3_out[212] = layer2_out[5964];
    assign layer3_out[213] = 1'b1;
    assign layer3_out[214] = layer2_out[7117] & ~layer2_out[7118];
    assign layer3_out[215] = ~layer2_out[4110] | layer2_out[4111];
    assign layer3_out[216] = layer2_out[1794] | layer2_out[1795];
    assign layer3_out[217] = layer2_out[2755];
    assign layer3_out[218] = layer2_out[1491];
    assign layer3_out[219] = layer2_out[1317];
    assign layer3_out[220] = ~layer2_out[5024] | layer2_out[5025];
    assign layer3_out[221] = ~layer2_out[740] | layer2_out[739];
    assign layer3_out[222] = ~(layer2_out[1741] ^ layer2_out[1742]);
    assign layer3_out[223] = layer2_out[3787] | layer2_out[3788];
    assign layer3_out[224] = layer2_out[4962];
    assign layer3_out[225] = layer2_out[4267] & ~layer2_out[4266];
    assign layer3_out[226] = layer2_out[7391];
    assign layer3_out[227] = ~(layer2_out[1242] ^ layer2_out[1243]);
    assign layer3_out[228] = layer2_out[6520];
    assign layer3_out[229] = layer2_out[3799] & ~layer2_out[3798];
    assign layer3_out[230] = ~layer2_out[6557];
    assign layer3_out[231] = ~layer2_out[4653] | layer2_out[4652];
    assign layer3_out[232] = ~layer2_out[1997];
    assign layer3_out[233] = layer2_out[154];
    assign layer3_out[234] = ~layer2_out[2314] | layer2_out[2315];
    assign layer3_out[235] = ~(layer2_out[1796] | layer2_out[1797]);
    assign layer3_out[236] = ~layer2_out[6252];
    assign layer3_out[237] = ~(layer2_out[4700] & layer2_out[4701]);
    assign layer3_out[238] = ~layer2_out[7859];
    assign layer3_out[239] = layer2_out[7130];
    assign layer3_out[240] = layer2_out[291] ^ layer2_out[292];
    assign layer3_out[241] = layer2_out[4246] & ~layer2_out[4245];
    assign layer3_out[242] = ~layer2_out[5179];
    assign layer3_out[243] = ~layer2_out[5585] | layer2_out[5584];
    assign layer3_out[244] = layer2_out[6815] & ~layer2_out[6816];
    assign layer3_out[245] = ~layer2_out[1247];
    assign layer3_out[246] = layer2_out[7030] & layer2_out[7031];
    assign layer3_out[247] = ~layer2_out[6699];
    assign layer3_out[248] = ~layer2_out[4584];
    assign layer3_out[249] = ~layer2_out[2899];
    assign layer3_out[250] = ~(layer2_out[810] ^ layer2_out[811]);
    assign layer3_out[251] = ~layer2_out[2713];
    assign layer3_out[252] = ~(layer2_out[350] & layer2_out[351]);
    assign layer3_out[253] = layer2_out[6037] & ~layer2_out[6038];
    assign layer3_out[254] = 1'b0;
    assign layer3_out[255] = layer2_out[2287] ^ layer2_out[2288];
    assign layer3_out[256] = layer2_out[7605] ^ layer2_out[7606];
    assign layer3_out[257] = layer2_out[6372] & layer2_out[6373];
    assign layer3_out[258] = layer2_out[3877] & ~layer2_out[3878];
    assign layer3_out[259] = ~layer2_out[4761] | layer2_out[4762];
    assign layer3_out[260] = layer2_out[1481] | layer2_out[1482];
    assign layer3_out[261] = layer2_out[2038] ^ layer2_out[2039];
    assign layer3_out[262] = layer2_out[1308];
    assign layer3_out[263] = layer2_out[2013] & ~layer2_out[2012];
    assign layer3_out[264] = layer2_out[1932] | layer2_out[1933];
    assign layer3_out[265] = ~(layer2_out[5543] ^ layer2_out[5544]);
    assign layer3_out[266] = layer2_out[2277] ^ layer2_out[2278];
    assign layer3_out[267] = ~(layer2_out[343] | layer2_out[344]);
    assign layer3_out[268] = ~layer2_out[1322] | layer2_out[1321];
    assign layer3_out[269] = ~layer2_out[3667];
    assign layer3_out[270] = layer2_out[4207] | layer2_out[4208];
    assign layer3_out[271] = layer2_out[861];
    assign layer3_out[272] = ~layer2_out[7798] | layer2_out[7799];
    assign layer3_out[273] = layer2_out[6304];
    assign layer3_out[274] = ~layer2_out[1087];
    assign layer3_out[275] = layer2_out[7143];
    assign layer3_out[276] = ~layer2_out[5463];
    assign layer3_out[277] = layer2_out[1875];
    assign layer3_out[278] = layer2_out[6092];
    assign layer3_out[279] = ~(layer2_out[7668] & layer2_out[7669]);
    assign layer3_out[280] = ~layer2_out[5037];
    assign layer3_out[281] = layer2_out[5400];
    assign layer3_out[282] = layer2_out[3057];
    assign layer3_out[283] = layer2_out[3079];
    assign layer3_out[284] = ~layer2_out[4780];
    assign layer3_out[285] = ~(layer2_out[368] ^ layer2_out[369]);
    assign layer3_out[286] = layer2_out[5643] & layer2_out[5644];
    assign layer3_out[287] = layer2_out[5908] | layer2_out[5909];
    assign layer3_out[288] = ~(layer2_out[6311] ^ layer2_out[6312]);
    assign layer3_out[289] = layer2_out[5874] ^ layer2_out[5875];
    assign layer3_out[290] = ~layer2_out[4650] | layer2_out[4649];
    assign layer3_out[291] = layer2_out[3050] & ~layer2_out[3049];
    assign layer3_out[292] = layer2_out[1302] & layer2_out[1303];
    assign layer3_out[293] = layer2_out[7701] & layer2_out[7702];
    assign layer3_out[294] = layer2_out[3768] & layer2_out[3769];
    assign layer3_out[295] = 1'b0;
    assign layer3_out[296] = 1'b0;
    assign layer3_out[297] = ~layer2_out[803];
    assign layer3_out[298] = ~layer2_out[4586];
    assign layer3_out[299] = layer2_out[3597] | layer2_out[3598];
    assign layer3_out[300] = layer2_out[2044] | layer2_out[2045];
    assign layer3_out[301] = layer2_out[2392] & ~layer2_out[2393];
    assign layer3_out[302] = ~layer2_out[7385];
    assign layer3_out[303] = ~layer2_out[2960];
    assign layer3_out[304] = ~(layer2_out[441] | layer2_out[442]);
    assign layer3_out[305] = layer2_out[6743];
    assign layer3_out[306] = layer2_out[7486] & ~layer2_out[7485];
    assign layer3_out[307] = layer2_out[1805] ^ layer2_out[1806];
    assign layer3_out[308] = ~layer2_out[6511] | layer2_out[6510];
    assign layer3_out[309] = layer2_out[2022] | layer2_out[2023];
    assign layer3_out[310] = layer2_out[2189] ^ layer2_out[2190];
    assign layer3_out[311] = layer2_out[6111] & ~layer2_out[6112];
    assign layer3_out[312] = ~(layer2_out[6] | layer2_out[7]);
    assign layer3_out[313] = layer2_out[2733] & ~layer2_out[2734];
    assign layer3_out[314] = ~layer2_out[1819];
    assign layer3_out[315] = ~layer2_out[2332] | layer2_out[2331];
    assign layer3_out[316] = layer2_out[357];
    assign layer3_out[317] = ~(layer2_out[5947] & layer2_out[5948]);
    assign layer3_out[318] = ~(layer2_out[3973] & layer2_out[3974]);
    assign layer3_out[319] = 1'b0;
    assign layer3_out[320] = layer2_out[2664];
    assign layer3_out[321] = ~layer2_out[3134];
    assign layer3_out[322] = layer2_out[6508] & ~layer2_out[6507];
    assign layer3_out[323] = ~layer2_out[6198] | layer2_out[6199];
    assign layer3_out[324] = layer2_out[3785];
    assign layer3_out[325] = ~layer2_out[7075];
    assign layer3_out[326] = layer2_out[2093] ^ layer2_out[2094];
    assign layer3_out[327] = layer2_out[4536];
    assign layer3_out[328] = layer2_out[5477];
    assign layer3_out[329] = layer2_out[7616] ^ layer2_out[7617];
    assign layer3_out[330] = layer2_out[55];
    assign layer3_out[331] = layer2_out[4350] & ~layer2_out[4349];
    assign layer3_out[332] = layer2_out[4431];
    assign layer3_out[333] = layer2_out[7038] & layer2_out[7039];
    assign layer3_out[334] = ~layer2_out[6477];
    assign layer3_out[335] = ~layer2_out[6452] | layer2_out[6451];
    assign layer3_out[336] = layer2_out[6949];
    assign layer3_out[337] = layer2_out[1501];
    assign layer3_out[338] = ~layer2_out[1800] | layer2_out[1799];
    assign layer3_out[339] = ~(layer2_out[2854] ^ layer2_out[2855]);
    assign layer3_out[340] = layer2_out[1472] | layer2_out[1473];
    assign layer3_out[341] = layer2_out[3747];
    assign layer3_out[342] = layer2_out[2077] | layer2_out[2078];
    assign layer3_out[343] = ~(layer2_out[7224] & layer2_out[7225]);
    assign layer3_out[344] = ~(layer2_out[4458] ^ layer2_out[4459]);
    assign layer3_out[345] = layer2_out[6614];
    assign layer3_out[346] = ~(layer2_out[5444] & layer2_out[5445]);
    assign layer3_out[347] = ~layer2_out[5060];
    assign layer3_out[348] = ~layer2_out[7529] | layer2_out[7528];
    assign layer3_out[349] = ~layer2_out[5046] | layer2_out[5047];
    assign layer3_out[350] = layer2_out[4269];
    assign layer3_out[351] = 1'b0;
    assign layer3_out[352] = layer2_out[2967];
    assign layer3_out[353] = ~layer2_out[2923];
    assign layer3_out[354] = ~layer2_out[6403];
    assign layer3_out[355] = ~layer2_out[4771];
    assign layer3_out[356] = layer2_out[971] & ~layer2_out[972];
    assign layer3_out[357] = ~(layer2_out[5762] | layer2_out[5763]);
    assign layer3_out[358] = ~layer2_out[255];
    assign layer3_out[359] = 1'b0;
    assign layer3_out[360] = ~layer2_out[4466];
    assign layer3_out[361] = layer2_out[3031] ^ layer2_out[3032];
    assign layer3_out[362] = layer2_out[4179] | layer2_out[4180];
    assign layer3_out[363] = ~layer2_out[6880];
    assign layer3_out[364] = layer2_out[905] | layer2_out[906];
    assign layer3_out[365] = ~layer2_out[7209];
    assign layer3_out[366] = ~layer2_out[1557];
    assign layer3_out[367] = ~(layer2_out[2580] & layer2_out[2581]);
    assign layer3_out[368] = 1'b0;
    assign layer3_out[369] = layer2_out[5901] & layer2_out[5902];
    assign layer3_out[370] = ~(layer2_out[4874] | layer2_out[4875]);
    assign layer3_out[371] = layer2_out[4594] ^ layer2_out[4595];
    assign layer3_out[372] = layer2_out[4685];
    assign layer3_out[373] = ~layer2_out[5007] | layer2_out[5008];
    assign layer3_out[374] = ~(layer2_out[6337] | layer2_out[6338]);
    assign layer3_out[375] = ~(layer2_out[5054] & layer2_out[5055]);
    assign layer3_out[376] = layer2_out[5053] & layer2_out[5054];
    assign layer3_out[377] = ~(layer2_out[5174] & layer2_out[5175]);
    assign layer3_out[378] = ~(layer2_out[3454] & layer2_out[3455]);
    assign layer3_out[379] = ~layer2_out[4955];
    assign layer3_out[380] = layer2_out[2512];
    assign layer3_out[381] = layer2_out[5317];
    assign layer3_out[382] = layer2_out[497] & ~layer2_out[496];
    assign layer3_out[383] = ~layer2_out[7702] | layer2_out[7703];
    assign layer3_out[384] = ~layer2_out[230] | layer2_out[231];
    assign layer3_out[385] = ~layer2_out[7030];
    assign layer3_out[386] = layer2_out[2073] | layer2_out[2074];
    assign layer3_out[387] = layer2_out[5810] & layer2_out[5811];
    assign layer3_out[388] = layer2_out[5829];
    assign layer3_out[389] = layer2_out[4192] | layer2_out[4193];
    assign layer3_out[390] = 1'b0;
    assign layer3_out[391] = layer2_out[4804];
    assign layer3_out[392] = 1'b0;
    assign layer3_out[393] = ~layer2_out[4104];
    assign layer3_out[394] = ~(layer2_out[5940] & layer2_out[5941]);
    assign layer3_out[395] = layer2_out[3156] & ~layer2_out[3155];
    assign layer3_out[396] = ~layer2_out[5302];
    assign layer3_out[397] = ~(layer2_out[3224] ^ layer2_out[3225]);
    assign layer3_out[398] = layer2_out[4238];
    assign layer3_out[399] = ~layer2_out[2368];
    assign layer3_out[400] = ~layer2_out[4967] | layer2_out[4966];
    assign layer3_out[401] = ~layer2_out[6658] | layer2_out[6659];
    assign layer3_out[402] = layer2_out[5268] & ~layer2_out[5269];
    assign layer3_out[403] = layer2_out[208];
    assign layer3_out[404] = ~(layer2_out[2438] & layer2_out[2439]);
    assign layer3_out[405] = layer2_out[2516] | layer2_out[2517];
    assign layer3_out[406] = ~layer2_out[2207];
    assign layer3_out[407] = layer2_out[4672] | layer2_out[4673];
    assign layer3_out[408] = ~(layer2_out[1593] ^ layer2_out[1594]);
    assign layer3_out[409] = ~layer2_out[1648] | layer2_out[1649];
    assign layer3_out[410] = layer2_out[6144];
    assign layer3_out[411] = layer2_out[7006];
    assign layer3_out[412] = ~layer2_out[1786];
    assign layer3_out[413] = layer2_out[7338] | layer2_out[7339];
    assign layer3_out[414] = layer2_out[3480] ^ layer2_out[3481];
    assign layer3_out[415] = layer2_out[5326];
    assign layer3_out[416] = ~layer2_out[1627] | layer2_out[1628];
    assign layer3_out[417] = layer2_out[2848];
    assign layer3_out[418] = ~layer2_out[2483];
    assign layer3_out[419] = ~(layer2_out[7794] & layer2_out[7795]);
    assign layer3_out[420] = layer2_out[2155] | layer2_out[2156];
    assign layer3_out[421] = ~(layer2_out[1340] ^ layer2_out[1341]);
    assign layer3_out[422] = ~layer2_out[6824] | layer2_out[6825];
    assign layer3_out[423] = ~(layer2_out[4842] & layer2_out[4843]);
    assign layer3_out[424] = ~(layer2_out[2868] | layer2_out[2869]);
    assign layer3_out[425] = ~(layer2_out[1945] | layer2_out[1946]);
    assign layer3_out[426] = ~layer2_out[1912];
    assign layer3_out[427] = layer2_out[5108];
    assign layer3_out[428] = ~layer2_out[7258];
    assign layer3_out[429] = ~layer2_out[2385] | layer2_out[2386];
    assign layer3_out[430] = ~(layer2_out[4319] & layer2_out[4320]);
    assign layer3_out[431] = layer2_out[6912];
    assign layer3_out[432] = ~layer2_out[5531] | layer2_out[5532];
    assign layer3_out[433] = ~layer2_out[4612];
    assign layer3_out[434] = ~layer2_out[5206];
    assign layer3_out[435] = ~layer2_out[3254];
    assign layer3_out[436] = layer2_out[5655] & ~layer2_out[5654];
    assign layer3_out[437] = layer2_out[6716] ^ layer2_out[6717];
    assign layer3_out[438] = ~(layer2_out[723] | layer2_out[724]);
    assign layer3_out[439] = ~(layer2_out[5855] ^ layer2_out[5856]);
    assign layer3_out[440] = layer2_out[7394] | layer2_out[7395];
    assign layer3_out[441] = 1'b0;
    assign layer3_out[442] = ~layer2_out[623];
    assign layer3_out[443] = layer2_out[3957] & layer2_out[3958];
    assign layer3_out[444] = ~layer2_out[7999];
    assign layer3_out[445] = ~layer2_out[4022];
    assign layer3_out[446] = ~(layer2_out[1300] ^ layer2_out[1301]);
    assign layer3_out[447] = layer2_out[3731] & ~layer2_out[3732];
    assign layer3_out[448] = ~(layer2_out[7204] | layer2_out[7205]);
    assign layer3_out[449] = ~(layer2_out[2191] & layer2_out[2192]);
    assign layer3_out[450] = ~layer2_out[7833];
    assign layer3_out[451] = layer2_out[3869] & ~layer2_out[3868];
    assign layer3_out[452] = ~layer2_out[6571];
    assign layer3_out[453] = ~(layer2_out[1132] & layer2_out[1133]);
    assign layer3_out[454] = ~layer2_out[4048];
    assign layer3_out[455] = layer2_out[1052];
    assign layer3_out[456] = layer2_out[2696];
    assign layer3_out[457] = layer2_out[6545] | layer2_out[6546];
    assign layer3_out[458] = ~layer2_out[2553] | layer2_out[2552];
    assign layer3_out[459] = layer2_out[6734] ^ layer2_out[6735];
    assign layer3_out[460] = ~layer2_out[4051] | layer2_out[4052];
    assign layer3_out[461] = ~layer2_out[5860] | layer2_out[5859];
    assign layer3_out[462] = ~(layer2_out[4689] & layer2_out[4690]);
    assign layer3_out[463] = layer2_out[4894];
    assign layer3_out[464] = layer2_out[390] & ~layer2_out[389];
    assign layer3_out[465] = ~(layer2_out[2429] & layer2_out[2430]);
    assign layer3_out[466] = layer2_out[1368] | layer2_out[1369];
    assign layer3_out[467] = ~(layer2_out[3759] & layer2_out[3760]);
    assign layer3_out[468] = ~layer2_out[1378];
    assign layer3_out[469] = ~layer2_out[7649];
    assign layer3_out[470] = layer2_out[5387] & layer2_out[5388];
    assign layer3_out[471] = ~(layer2_out[3341] ^ layer2_out[3342]);
    assign layer3_out[472] = layer2_out[6452] ^ layer2_out[6453];
    assign layer3_out[473] = ~layer2_out[1614] | layer2_out[1615];
    assign layer3_out[474] = layer2_out[5089] | layer2_out[5090];
    assign layer3_out[475] = layer2_out[6543];
    assign layer3_out[476] = layer2_out[21];
    assign layer3_out[477] = ~layer2_out[686];
    assign layer3_out[478] = ~layer2_out[6107] | layer2_out[6106];
    assign layer3_out[479] = ~layer2_out[4338] | layer2_out[4337];
    assign layer3_out[480] = layer2_out[6169] & ~layer2_out[6170];
    assign layer3_out[481] = layer2_out[4002] & ~layer2_out[4001];
    assign layer3_out[482] = layer2_out[2436];
    assign layer3_out[483] = layer2_out[1259] | layer2_out[1260];
    assign layer3_out[484] = layer2_out[3288] ^ layer2_out[3289];
    assign layer3_out[485] = layer2_out[6453] & ~layer2_out[6454];
    assign layer3_out[486] = ~layer2_out[3456];
    assign layer3_out[487] = layer2_out[4472];
    assign layer3_out[488] = layer2_out[6215];
    assign layer3_out[489] = layer2_out[4528] & ~layer2_out[4527];
    assign layer3_out[490] = layer2_out[4845];
    assign layer3_out[491] = layer2_out[2359] | layer2_out[2360];
    assign layer3_out[492] = layer2_out[7084] & ~layer2_out[7083];
    assign layer3_out[493] = layer2_out[6338];
    assign layer3_out[494] = layer2_out[578];
    assign layer3_out[495] = ~layer2_out[7245];
    assign layer3_out[496] = ~layer2_out[7919] | layer2_out[7918];
    assign layer3_out[497] = ~layer2_out[4433];
    assign layer3_out[498] = layer2_out[2843];
    assign layer3_out[499] = ~(layer2_out[7846] & layer2_out[7847]);
    assign layer3_out[500] = ~layer2_out[206];
    assign layer3_out[501] = ~layer2_out[763] | layer2_out[762];
    assign layer3_out[502] = ~layer2_out[5075];
    assign layer3_out[503] = ~layer2_out[5264];
    assign layer3_out[504] = layer2_out[2938];
    assign layer3_out[505] = layer2_out[7068] & layer2_out[7069];
    assign layer3_out[506] = layer2_out[4797] | layer2_out[4798];
    assign layer3_out[507] = layer2_out[354];
    assign layer3_out[508] = layer2_out[742] & ~layer2_out[743];
    assign layer3_out[509] = layer2_out[6684];
    assign layer3_out[510] = layer2_out[6096];
    assign layer3_out[511] = layer2_out[1091] & ~layer2_out[1092];
    assign layer3_out[512] = ~layer2_out[2866];
    assign layer3_out[513] = ~(layer2_out[2585] ^ layer2_out[2586]);
    assign layer3_out[514] = ~(layer2_out[7370] | layer2_out[7371]);
    assign layer3_out[515] = ~(layer2_out[6568] & layer2_out[6569]);
    assign layer3_out[516] = ~layer2_out[463];
    assign layer3_out[517] = ~layer2_out[1275] | layer2_out[1274];
    assign layer3_out[518] = ~(layer2_out[7410] | layer2_out[7411]);
    assign layer3_out[519] = layer2_out[3052];
    assign layer3_out[520] = layer2_out[3084] & ~layer2_out[3085];
    assign layer3_out[521] = ~layer2_out[1459];
    assign layer3_out[522] = layer2_out[4063] | layer2_out[4064];
    assign layer3_out[523] = ~layer2_out[979];
    assign layer3_out[524] = ~layer2_out[2080];
    assign layer3_out[525] = layer2_out[1630] ^ layer2_out[1631];
    assign layer3_out[526] = layer2_out[3005];
    assign layer3_out[527] = layer2_out[6489] | layer2_out[6490];
    assign layer3_out[528] = layer2_out[5050];
    assign layer3_out[529] = layer2_out[7319] ^ layer2_out[7320];
    assign layer3_out[530] = ~layer2_out[3364];
    assign layer3_out[531] = layer2_out[1480] ^ layer2_out[1481];
    assign layer3_out[532] = ~layer2_out[7769];
    assign layer3_out[533] = ~layer2_out[4715];
    assign layer3_out[534] = ~layer2_out[3072] | layer2_out[3073];
    assign layer3_out[535] = ~layer2_out[2642];
    assign layer3_out[536] = layer2_out[7034] ^ layer2_out[7035];
    assign layer3_out[537] = layer2_out[7086] | layer2_out[7087];
    assign layer3_out[538] = ~(layer2_out[6027] & layer2_out[6028]);
    assign layer3_out[539] = layer2_out[4729];
    assign layer3_out[540] = layer2_out[2428];
    assign layer3_out[541] = ~layer2_out[5634] | layer2_out[5633];
    assign layer3_out[542] = layer2_out[3297] ^ layer2_out[3298];
    assign layer3_out[543] = 1'b0;
    assign layer3_out[544] = 1'b1;
    assign layer3_out[545] = layer2_out[416];
    assign layer3_out[546] = ~layer2_out[4683] | layer2_out[4684];
    assign layer3_out[547] = ~layer2_out[6293];
    assign layer3_out[548] = ~(layer2_out[1004] & layer2_out[1005]);
    assign layer3_out[549] = layer2_out[6815];
    assign layer3_out[550] = layer2_out[1931];
    assign layer3_out[551] = layer2_out[2914];
    assign layer3_out[552] = ~(layer2_out[2956] & layer2_out[2957]);
    assign layer3_out[553] = ~(layer2_out[3985] ^ layer2_out[3986]);
    assign layer3_out[554] = layer2_out[5802] & ~layer2_out[5801];
    assign layer3_out[555] = ~layer2_out[2611] | layer2_out[2612];
    assign layer3_out[556] = ~layer2_out[3672];
    assign layer3_out[557] = ~(layer2_out[6282] | layer2_out[6283]);
    assign layer3_out[558] = ~layer2_out[4513];
    assign layer3_out[559] = ~(layer2_out[698] ^ layer2_out[699]);
    assign layer3_out[560] = ~(layer2_out[7218] & layer2_out[7219]);
    assign layer3_out[561] = ~layer2_out[2101] | layer2_out[2102];
    assign layer3_out[562] = layer2_out[2674];
    assign layer3_out[563] = ~(layer2_out[3952] | layer2_out[3953]);
    assign layer3_out[564] = layer2_out[2673];
    assign layer3_out[565] = ~layer2_out[6828];
    assign layer3_out[566] = ~layer2_out[478];
    assign layer3_out[567] = ~layer2_out[2985] | layer2_out[2984];
    assign layer3_out[568] = ~layer2_out[7656];
    assign layer3_out[569] = 1'b1;
    assign layer3_out[570] = layer2_out[5297];
    assign layer3_out[571] = ~layer2_out[2149];
    assign layer3_out[572] = layer2_out[3143];
    assign layer3_out[573] = layer2_out[3549] & layer2_out[3550];
    assign layer3_out[574] = layer2_out[7539] ^ layer2_out[7540];
    assign layer3_out[575] = ~(layer2_out[4195] | layer2_out[4196]);
    assign layer3_out[576] = layer2_out[471] & ~layer2_out[472];
    assign layer3_out[577] = ~(layer2_out[6927] ^ layer2_out[6928]);
    assign layer3_out[578] = ~layer2_out[6998];
    assign layer3_out[579] = layer2_out[6602];
    assign layer3_out[580] = layer2_out[363];
    assign layer3_out[581] = layer2_out[2289] & ~layer2_out[2290];
    assign layer3_out[582] = ~layer2_out[2240];
    assign layer3_out[583] = ~layer2_out[5930];
    assign layer3_out[584] = ~(layer2_out[1553] & layer2_out[1554]);
    assign layer3_out[585] = layer2_out[2912];
    assign layer3_out[586] = layer2_out[7694];
    assign layer3_out[587] = layer2_out[5349] & ~layer2_out[5348];
    assign layer3_out[588] = ~layer2_out[6935] | layer2_out[6936];
    assign layer3_out[589] = layer2_out[6652] & ~layer2_out[6651];
    assign layer3_out[590] = layer2_out[6341] ^ layer2_out[6342];
    assign layer3_out[591] = layer2_out[3919] | layer2_out[3920];
    assign layer3_out[592] = layer2_out[5529];
    assign layer3_out[593] = ~(layer2_out[1896] | layer2_out[1897]);
    assign layer3_out[594] = layer2_out[3837] & ~layer2_out[3838];
    assign layer3_out[595] = ~layer2_out[5245] | layer2_out[5246];
    assign layer3_out[596] = ~layer2_out[2508] | layer2_out[2509];
    assign layer3_out[597] = ~layer2_out[7585] | layer2_out[7586];
    assign layer3_out[598] = ~(layer2_out[5344] | layer2_out[5345]);
    assign layer3_out[599] = ~(layer2_out[5226] | layer2_out[5227]);
    assign layer3_out[600] = ~(layer2_out[3865] | layer2_out[3866]);
    assign layer3_out[601] = ~(layer2_out[6503] & layer2_out[6504]);
    assign layer3_out[602] = layer2_out[2301];
    assign layer3_out[603] = ~layer2_out[3555];
    assign layer3_out[604] = layer2_out[5602] ^ layer2_out[5603];
    assign layer3_out[605] = layer2_out[7833] | layer2_out[7834];
    assign layer3_out[606] = layer2_out[276] | layer2_out[277];
    assign layer3_out[607] = layer2_out[1442] | layer2_out[1443];
    assign layer3_out[608] = ~layer2_out[1692] | layer2_out[1693];
    assign layer3_out[609] = ~(layer2_out[2800] ^ layer2_out[2801]);
    assign layer3_out[610] = layer2_out[6269];
    assign layer3_out[611] = layer2_out[3698];
    assign layer3_out[612] = ~layer2_out[4766] | layer2_out[4767];
    assign layer3_out[613] = layer2_out[1554];
    assign layer3_out[614] = ~(layer2_out[2142] ^ layer2_out[2143]);
    assign layer3_out[615] = layer2_out[7562];
    assign layer3_out[616] = layer2_out[6845] ^ layer2_out[6846];
    assign layer3_out[617] = ~(layer2_out[4703] | layer2_out[4704]);
    assign layer3_out[618] = layer2_out[7894] & ~layer2_out[7895];
    assign layer3_out[619] = layer2_out[295] ^ layer2_out[296];
    assign layer3_out[620] = ~layer2_out[3847];
    assign layer3_out[621] = ~layer2_out[7257] | layer2_out[7256];
    assign layer3_out[622] = ~layer2_out[1215] | layer2_out[1214];
    assign layer3_out[623] = ~layer2_out[592];
    assign layer3_out[624] = layer2_out[4628] & ~layer2_out[4627];
    assign layer3_out[625] = ~(layer2_out[929] ^ layer2_out[930]);
    assign layer3_out[626] = layer2_out[3133] ^ layer2_out[3134];
    assign layer3_out[627] = layer2_out[5814] & ~layer2_out[5815];
    assign layer3_out[628] = layer2_out[4693] ^ layer2_out[4694];
    assign layer3_out[629] = layer2_out[3571] | layer2_out[3572];
    assign layer3_out[630] = layer2_out[1229] ^ layer2_out[1230];
    assign layer3_out[631] = ~layer2_out[1516];
    assign layer3_out[632] = 1'b0;
    assign layer3_out[633] = layer2_out[3528] | layer2_out[3529];
    assign layer3_out[634] = ~layer2_out[7347] | layer2_out[7346];
    assign layer3_out[635] = ~(layer2_out[5379] & layer2_out[5380]);
    assign layer3_out[636] = ~layer2_out[3281];
    assign layer3_out[637] = ~layer2_out[4578] | layer2_out[4577];
    assign layer3_out[638] = layer2_out[5278] & layer2_out[5279];
    assign layer3_out[639] = layer2_out[3563] & ~layer2_out[3564];
    assign layer3_out[640] = layer2_out[7628];
    assign layer3_out[641] = ~layer2_out[6956] | layer2_out[6955];
    assign layer3_out[642] = layer2_out[3249];
    assign layer3_out[643] = layer2_out[2615];
    assign layer3_out[644] = layer2_out[1705];
    assign layer3_out[645] = ~layer2_out[2331];
    assign layer3_out[646] = ~layer2_out[6813];
    assign layer3_out[647] = layer2_out[6895];
    assign layer3_out[648] = layer2_out[326];
    assign layer3_out[649] = ~layer2_out[5970];
    assign layer3_out[650] = ~layer2_out[2164];
    assign layer3_out[651] = layer2_out[2756] | layer2_out[2757];
    assign layer3_out[652] = layer2_out[1166];
    assign layer3_out[653] = ~layer2_out[3022] | layer2_out[3023];
    assign layer3_out[654] = layer2_out[7398] & layer2_out[7399];
    assign layer3_out[655] = ~(layer2_out[4746] ^ layer2_out[4747]);
    assign layer3_out[656] = layer2_out[3925] & ~layer2_out[3926];
    assign layer3_out[657] = ~layer2_out[2337];
    assign layer3_out[658] = ~layer2_out[533];
    assign layer3_out[659] = layer2_out[5647] & ~layer2_out[5646];
    assign layer3_out[660] = layer2_out[6766] & ~layer2_out[6767];
    assign layer3_out[661] = layer2_out[4338];
    assign layer3_out[662] = layer2_out[2578] & ~layer2_out[2577];
    assign layer3_out[663] = ~layer2_out[6519];
    assign layer3_out[664] = ~(layer2_out[7624] & layer2_out[7625]);
    assign layer3_out[665] = layer2_out[7556] & ~layer2_out[7557];
    assign layer3_out[666] = ~(layer2_out[6891] ^ layer2_out[6892]);
    assign layer3_out[667] = layer2_out[3450];
    assign layer3_out[668] = ~(layer2_out[3857] & layer2_out[3858]);
    assign layer3_out[669] = ~(layer2_out[7425] & layer2_out[7426]);
    assign layer3_out[670] = ~layer2_out[1862];
    assign layer3_out[671] = layer2_out[7770];
    assign layer3_out[672] = layer2_out[4170] & ~layer2_out[4169];
    assign layer3_out[673] = layer2_out[5981] ^ layer2_out[5982];
    assign layer3_out[674] = ~layer2_out[4973] | layer2_out[4974];
    assign layer3_out[675] = ~layer2_out[4290] | layer2_out[4291];
    assign layer3_out[676] = ~(layer2_out[6257] ^ layer2_out[6258]);
    assign layer3_out[677] = ~(layer2_out[1575] | layer2_out[1576]);
    assign layer3_out[678] = ~layer2_out[32];
    assign layer3_out[679] = layer2_out[6475] & layer2_out[6476];
    assign layer3_out[680] = ~layer2_out[1375] | layer2_out[1376];
    assign layer3_out[681] = layer2_out[4325];
    assign layer3_out[682] = layer2_out[6358];
    assign layer3_out[683] = ~layer2_out[4622];
    assign layer3_out[684] = ~(layer2_out[4448] | layer2_out[4449]);
    assign layer3_out[685] = ~layer2_out[5680] | layer2_out[5681];
    assign layer3_out[686] = layer2_out[7134];
    assign layer3_out[687] = layer2_out[5882] & ~layer2_out[5881];
    assign layer3_out[688] = ~layer2_out[2881];
    assign layer3_out[689] = layer2_out[4085] & layer2_out[4086];
    assign layer3_out[690] = ~(layer2_out[4113] & layer2_out[4114]);
    assign layer3_out[691] = layer2_out[1541];
    assign layer3_out[692] = ~(layer2_out[5582] & layer2_out[5583]);
    assign layer3_out[693] = ~layer2_out[4906];
    assign layer3_out[694] = ~layer2_out[3333];
    assign layer3_out[695] = layer2_out[6439] | layer2_out[6440];
    assign layer3_out[696] = ~layer2_out[4462];
    assign layer3_out[697] = ~(layer2_out[2603] & layer2_out[2604]);
    assign layer3_out[698] = ~layer2_out[7246];
    assign layer3_out[699] = layer2_out[4635];
    assign layer3_out[700] = layer2_out[6560] & ~layer2_out[6559];
    assign layer3_out[701] = ~(layer2_out[6878] & layer2_out[6879]);
    assign layer3_out[702] = 1'b0;
    assign layer3_out[703] = ~layer2_out[3439] | layer2_out[3438];
    assign layer3_out[704] = layer2_out[7744];
    assign layer3_out[705] = layer2_out[1353];
    assign layer3_out[706] = layer2_out[1470] ^ layer2_out[1471];
    assign layer3_out[707] = ~layer2_out[4191];
    assign layer3_out[708] = layer2_out[48] | layer2_out[49];
    assign layer3_out[709] = layer2_out[2661] & ~layer2_out[2662];
    assign layer3_out[710] = layer2_out[3490] & ~layer2_out[3491];
    assign layer3_out[711] = layer2_out[37] & ~layer2_out[36];
    assign layer3_out[712] = layer2_out[2597];
    assign layer3_out[713] = ~(layer2_out[4847] & layer2_out[4848]);
    assign layer3_out[714] = layer2_out[5868] | layer2_out[5869];
    assign layer3_out[715] = layer2_out[269] & ~layer2_out[270];
    assign layer3_out[716] = ~layer2_out[7518] | layer2_out[7517];
    assign layer3_out[717] = layer2_out[1762] & ~layer2_out[1763];
    assign layer3_out[718] = ~layer2_out[2458] | layer2_out[2459];
    assign layer3_out[719] = layer2_out[3070];
    assign layer3_out[720] = ~layer2_out[4052];
    assign layer3_out[721] = ~(layer2_out[6893] | layer2_out[6894]);
    assign layer3_out[722] = ~layer2_out[491];
    assign layer3_out[723] = layer2_out[4486] & layer2_out[4487];
    assign layer3_out[724] = layer2_out[6656];
    assign layer3_out[725] = ~(layer2_out[855] & layer2_out[856]);
    assign layer3_out[726] = ~layer2_out[6859];
    assign layer3_out[727] = layer2_out[7265] | layer2_out[7266];
    assign layer3_out[728] = layer2_out[3962] ^ layer2_out[3963];
    assign layer3_out[729] = layer2_out[4531] ^ layer2_out[4532];
    assign layer3_out[730] = layer2_out[3630];
    assign layer3_out[731] = 1'b1;
    assign layer3_out[732] = layer2_out[7867] & layer2_out[7868];
    assign layer3_out[733] = layer2_out[1123];
    assign layer3_out[734] = layer2_out[17];
    assign layer3_out[735] = ~layer2_out[4249] | layer2_out[4250];
    assign layer3_out[736] = layer2_out[3661];
    assign layer3_out[737] = ~layer2_out[4227] | layer2_out[4226];
    assign layer3_out[738] = layer2_out[3018] & layer2_out[3019];
    assign layer3_out[739] = ~layer2_out[1487];
    assign layer3_out[740] = ~layer2_out[415];
    assign layer3_out[741] = 1'b1;
    assign layer3_out[742] = ~(layer2_out[7254] ^ layer2_out[7255]);
    assign layer3_out[743] = ~layer2_out[1366];
    assign layer3_out[744] = layer2_out[2515] | layer2_out[2516];
    assign layer3_out[745] = layer2_out[4348] & ~layer2_out[4349];
    assign layer3_out[746] = layer2_out[3169] & ~layer2_out[3168];
    assign layer3_out[747] = layer2_out[4412] | layer2_out[4413];
    assign layer3_out[748] = layer2_out[3629];
    assign layer3_out[749] = ~(layer2_out[7469] ^ layer2_out[7470]);
    assign layer3_out[750] = 1'b1;
    assign layer3_out[751] = ~layer2_out[4801];
    assign layer3_out[752] = ~(layer2_out[4026] ^ layer2_out[4027]);
    assign layer3_out[753] = layer2_out[7838] & ~layer2_out[7839];
    assign layer3_out[754] = ~layer2_out[7368];
    assign layer3_out[755] = ~layer2_out[822] | layer2_out[821];
    assign layer3_out[756] = ~layer2_out[5285];
    assign layer3_out[757] = ~(layer2_out[6306] & layer2_out[6307]);
    assign layer3_out[758] = ~layer2_out[5978];
    assign layer3_out[759] = ~layer2_out[4406];
    assign layer3_out[760] = layer2_out[6283] | layer2_out[6284];
    assign layer3_out[761] = ~layer2_out[517];
    assign layer3_out[762] = ~layer2_out[995] | layer2_out[994];
    assign layer3_out[763] = layer2_out[3255] & layer2_out[3256];
    assign layer3_out[764] = layer2_out[1879];
    assign layer3_out[765] = ~layer2_out[359] | layer2_out[358];
    assign layer3_out[766] = ~layer2_out[3115] | layer2_out[3114];
    assign layer3_out[767] = ~layer2_out[134] | layer2_out[135];
    assign layer3_out[768] = layer2_out[332] | layer2_out[333];
    assign layer3_out[769] = layer2_out[4516];
    assign layer3_out[770] = ~(layer2_out[3369] & layer2_out[3370]);
    assign layer3_out[771] = layer2_out[5616];
    assign layer3_out[772] = layer2_out[545];
    assign layer3_out[773] = ~layer2_out[458] | layer2_out[459];
    assign layer3_out[774] = ~layer2_out[7546];
    assign layer3_out[775] = layer2_out[7147];
    assign layer3_out[776] = ~layer2_out[2542] | layer2_out[2543];
    assign layer3_out[777] = layer2_out[2566];
    assign layer3_out[778] = ~layer2_out[5352];
    assign layer3_out[779] = layer2_out[5500] ^ layer2_out[5501];
    assign layer3_out[780] = layer2_out[5641];
    assign layer3_out[781] = ~layer2_out[3260];
    assign layer3_out[782] = layer2_out[4386] & ~layer2_out[4385];
    assign layer3_out[783] = layer2_out[1694] ^ layer2_out[1695];
    assign layer3_out[784] = ~(layer2_out[1447] & layer2_out[1448]);
    assign layer3_out[785] = layer2_out[2689] | layer2_out[2690];
    assign layer3_out[786] = ~layer2_out[5781] | layer2_out[5782];
    assign layer3_out[787] = ~layer2_out[2952];
    assign layer3_out[788] = ~layer2_out[5322];
    assign layer3_out[789] = ~(layer2_out[3477] ^ layer2_out[3478]);
    assign layer3_out[790] = ~layer2_out[3182];
    assign layer3_out[791] = 1'b0;
    assign layer3_out[792] = ~layer2_out[1124];
    assign layer3_out[793] = layer2_out[5741] & ~layer2_out[5742];
    assign layer3_out[794] = ~layer2_out[1288];
    assign layer3_out[795] = ~layer2_out[2344];
    assign layer3_out[796] = layer2_out[308] ^ layer2_out[309];
    assign layer3_out[797] = 1'b0;
    assign layer3_out[798] = ~(layer2_out[2861] & layer2_out[2862]);
    assign layer3_out[799] = layer2_out[2681] | layer2_out[2682];
    assign layer3_out[800] = layer2_out[1778];
    assign layer3_out[801] = ~layer2_out[5915];
    assign layer3_out[802] = ~layer2_out[6230];
    assign layer3_out[803] = ~layer2_out[4657];
    assign layer3_out[804] = ~layer2_out[493];
    assign layer3_out[805] = ~layer2_out[6885];
    assign layer3_out[806] = ~layer2_out[5087];
    assign layer3_out[807] = layer2_out[6200] & layer2_out[6201];
    assign layer3_out[808] = layer2_out[3662];
    assign layer3_out[809] = layer2_out[1475] | layer2_out[1476];
    assign layer3_out[810] = layer2_out[2730];
    assign layer3_out[811] = ~(layer2_out[5120] | layer2_out[5121]);
    assign layer3_out[812] = layer2_out[4898] ^ layer2_out[4899];
    assign layer3_out[813] = layer2_out[3068];
    assign layer3_out[814] = ~(layer2_out[3911] & layer2_out[3912]);
    assign layer3_out[815] = layer2_out[2812];
    assign layer3_out[816] = layer2_out[5388];
    assign layer3_out[817] = ~layer2_out[436];
    assign layer3_out[818] = ~(layer2_out[6309] & layer2_out[6310]);
    assign layer3_out[819] = ~layer2_out[7553];
    assign layer3_out[820] = ~(layer2_out[2836] & layer2_out[2837]);
    assign layer3_out[821] = ~layer2_out[6927];
    assign layer3_out[822] = layer2_out[7342] & layer2_out[7343];
    assign layer3_out[823] = 1'b1;
    assign layer3_out[824] = ~layer2_out[7945];
    assign layer3_out[825] = ~(layer2_out[3354] | layer2_out[3355]);
    assign layer3_out[826] = layer2_out[3632] ^ layer2_out[3633];
    assign layer3_out[827] = ~layer2_out[854];
    assign layer3_out[828] = layer2_out[3373];
    assign layer3_out[829] = layer2_out[7274] & ~layer2_out[7273];
    assign layer3_out[830] = ~layer2_out[3167] | layer2_out[3168];
    assign layer3_out[831] = layer2_out[651] ^ layer2_out[652];
    assign layer3_out[832] = ~layer2_out[6869];
    assign layer3_out[833] = layer2_out[481] ^ layer2_out[482];
    assign layer3_out[834] = ~layer2_out[6693];
    assign layer3_out[835] = ~layer2_out[485];
    assign layer3_out[836] = ~layer2_out[7098];
    assign layer3_out[837] = layer2_out[2165] ^ layer2_out[2166];
    assign layer3_out[838] = ~layer2_out[1669];
    assign layer3_out[839] = layer2_out[3538] & ~layer2_out[3539];
    assign layer3_out[840] = layer2_out[2963];
    assign layer3_out[841] = layer2_out[1983];
    assign layer3_out[842] = layer2_out[2222] & ~layer2_out[2223];
    assign layer3_out[843] = ~layer2_out[6810];
    assign layer3_out[844] = layer2_out[1506] | layer2_out[1507];
    assign layer3_out[845] = ~(layer2_out[3928] & layer2_out[3929]);
    assign layer3_out[846] = ~(layer2_out[3963] & layer2_out[3964]);
    assign layer3_out[847] = layer2_out[5316] & ~layer2_out[5317];
    assign layer3_out[848] = layer2_out[635] | layer2_out[636];
    assign layer3_out[849] = layer2_out[7840] ^ layer2_out[7841];
    assign layer3_out[850] = ~layer2_out[697] | layer2_out[698];
    assign layer3_out[851] = layer2_out[5284];
    assign layer3_out[852] = ~layer2_out[6209] | layer2_out[6210];
    assign layer3_out[853] = ~layer2_out[7407];
    assign layer3_out[854] = layer2_out[4493] & layer2_out[4494];
    assign layer3_out[855] = layer2_out[5833];
    assign layer3_out[856] = layer2_out[7449] & ~layer2_out[7450];
    assign layer3_out[857] = ~(layer2_out[5734] & layer2_out[5735]);
    assign layer3_out[858] = layer2_out[6006];
    assign layer3_out[859] = ~layer2_out[652] | layer2_out[653];
    assign layer3_out[860] = ~(layer2_out[1431] ^ layer2_out[1432]);
    assign layer3_out[861] = ~(layer2_out[5792] ^ layer2_out[5793]);
    assign layer3_out[862] = layer2_out[4029] & ~layer2_out[4028];
    assign layer3_out[863] = layer2_out[1026];
    assign layer3_out[864] = ~layer2_out[7306] | layer2_out[7305];
    assign layer3_out[865] = ~layer2_out[4426];
    assign layer3_out[866] = layer2_out[99];
    assign layer3_out[867] = layer2_out[6675];
    assign layer3_out[868] = ~layer2_out[2986];
    assign layer3_out[869] = layer2_out[6847];
    assign layer3_out[870] = ~layer2_out[5026];
    assign layer3_out[871] = ~layer2_out[4171];
    assign layer3_out[872] = 1'b1;
    assign layer3_out[873] = layer2_out[2919] | layer2_out[2920];
    assign layer3_out[874] = ~layer2_out[7102] | layer2_out[7103];
    assign layer3_out[875] = layer2_out[4157];
    assign layer3_out[876] = ~(layer2_out[2099] ^ layer2_out[2100]);
    assign layer3_out[877] = layer2_out[2240] ^ layer2_out[2241];
    assign layer3_out[878] = layer2_out[2539] & ~layer2_out[2538];
    assign layer3_out[879] = layer2_out[4155] & ~layer2_out[4156];
    assign layer3_out[880] = layer2_out[1691] & layer2_out[1692];
    assign layer3_out[881] = layer2_out[5262];
    assign layer3_out[882] = ~(layer2_out[50] ^ layer2_out[51]);
    assign layer3_out[883] = layer2_out[2993] ^ layer2_out[2994];
    assign layer3_out[884] = ~layer2_out[2617];
    assign layer3_out[885] = layer2_out[4829] & layer2_out[4830];
    assign layer3_out[886] = layer2_out[7916] ^ layer2_out[7917];
    assign layer3_out[887] = ~layer2_out[3551];
    assign layer3_out[888] = ~layer2_out[3453] | layer2_out[3454];
    assign layer3_out[889] = ~layer2_out[1407];
    assign layer3_out[890] = ~(layer2_out[2128] ^ layer2_out[2129]);
    assign layer3_out[891] = layer2_out[4219] & layer2_out[4220];
    assign layer3_out[892] = ~(layer2_out[131] & layer2_out[132]);
    assign layer3_out[893] = ~layer2_out[4599] | layer2_out[4600];
    assign layer3_out[894] = ~layer2_out[6744];
    assign layer3_out[895] = ~layer2_out[5102] | layer2_out[5101];
    assign layer3_out[896] = layer2_out[3456];
    assign layer3_out[897] = layer2_out[5558] | layer2_out[5559];
    assign layer3_out[898] = layer2_out[1716];
    assign layer3_out[899] = ~layer2_out[3142];
    assign layer3_out[900] = layer2_out[3876] ^ layer2_out[3877];
    assign layer3_out[901] = layer2_out[2853] & ~layer2_out[2854];
    assign layer3_out[902] = layer2_out[3205] ^ layer2_out[3206];
    assign layer3_out[903] = ~layer2_out[2059];
    assign layer3_out[904] = ~(layer2_out[2903] ^ layer2_out[2904]);
    assign layer3_out[905] = layer2_out[3229] & ~layer2_out[3230];
    assign layer3_out[906] = ~(layer2_out[2434] & layer2_out[2435]);
    assign layer3_out[907] = layer2_out[3231] & layer2_out[3232];
    assign layer3_out[908] = layer2_out[6028] & layer2_out[6029];
    assign layer3_out[909] = ~(layer2_out[3698] ^ layer2_out[3699]);
    assign layer3_out[910] = layer2_out[6783];
    assign layer3_out[911] = layer2_out[4707];
    assign layer3_out[912] = ~layer2_out[5886];
    assign layer3_out[913] = layer2_out[7482];
    assign layer3_out[914] = ~(layer2_out[5328] & layer2_out[5329]);
    assign layer3_out[915] = layer2_out[7477] & ~layer2_out[7478];
    assign layer3_out[916] = layer2_out[1376];
    assign layer3_out[917] = ~layer2_out[3676];
    assign layer3_out[918] = ~(layer2_out[1146] | layer2_out[1147]);
    assign layer3_out[919] = ~(layer2_out[3484] ^ layer2_out[3485]);
    assign layer3_out[920] = ~layer2_out[4659];
    assign layer3_out[921] = layer2_out[7181] | layer2_out[7182];
    assign layer3_out[922] = 1'b0;
    assign layer3_out[923] = layer2_out[6548] & ~layer2_out[6547];
    assign layer3_out[924] = layer2_out[764] ^ layer2_out[765];
    assign layer3_out[925] = layer2_out[4641] | layer2_out[4642];
    assign layer3_out[926] = ~(layer2_out[2416] ^ layer2_out[2417]);
    assign layer3_out[927] = ~layer2_out[2611];
    assign layer3_out[928] = 1'b0;
    assign layer3_out[929] = ~(layer2_out[7920] & layer2_out[7921]);
    assign layer3_out[930] = ~layer2_out[7850] | layer2_out[7851];
    assign layer3_out[931] = layer2_out[171] & ~layer2_out[172];
    assign layer3_out[932] = ~layer2_out[4867];
    assign layer3_out[933] = ~layer2_out[3431] | layer2_out[3432];
    assign layer3_out[934] = layer2_out[3831] & ~layer2_out[3830];
    assign layer3_out[935] = 1'b0;
    assign layer3_out[936] = ~layer2_out[7021];
    assign layer3_out[937] = layer2_out[1635] & ~layer2_out[1636];
    assign layer3_out[938] = layer2_out[4806] & layer2_out[4807];
    assign layer3_out[939] = layer2_out[2345] ^ layer2_out[2346];
    assign layer3_out[940] = ~(layer2_out[2489] ^ layer2_out[2490]);
    assign layer3_out[941] = ~layer2_out[5659];
    assign layer3_out[942] = layer2_out[3573] ^ layer2_out[3574];
    assign layer3_out[943] = layer2_out[5334];
    assign layer3_out[944] = ~layer2_out[5744] | layer2_out[5745];
    assign layer3_out[945] = ~(layer2_out[2415] & layer2_out[2416]);
    assign layer3_out[946] = ~(layer2_out[5461] ^ layer2_out[5462]);
    assign layer3_out[947] = layer2_out[1909] | layer2_out[1910];
    assign layer3_out[948] = layer2_out[3091] ^ layer2_out[3092];
    assign layer3_out[949] = layer2_out[5390];
    assign layer3_out[950] = ~layer2_out[6165] | layer2_out[6164];
    assign layer3_out[951] = ~layer2_out[6807] | layer2_out[6806];
    assign layer3_out[952] = layer2_out[689] & layer2_out[690];
    assign layer3_out[953] = ~(layer2_out[7048] ^ layer2_out[7049]);
    assign layer3_out[954] = ~(layer2_out[344] ^ layer2_out[345]);
    assign layer3_out[955] = layer2_out[7972];
    assign layer3_out[956] = ~(layer2_out[7318] & layer2_out[7319]);
    assign layer3_out[957] = ~layer2_out[901];
    assign layer3_out[958] = layer2_out[3546] | layer2_out[3547];
    assign layer3_out[959] = layer2_out[4675] & layer2_out[4676];
    assign layer3_out[960] = ~(layer2_out[1284] | layer2_out[1285]);
    assign layer3_out[961] = ~(layer2_out[5528] & layer2_out[5529]);
    assign layer3_out[962] = layer2_out[4746];
    assign layer3_out[963] = ~layer2_out[7421];
    assign layer3_out[964] = layer2_out[5989] & layer2_out[5990];
    assign layer3_out[965] = layer2_out[3908];
    assign layer3_out[966] = layer2_out[5240] ^ layer2_out[5241];
    assign layer3_out[967] = layer2_out[4558] & layer2_out[4559];
    assign layer3_out[968] = ~(layer2_out[6995] ^ layer2_out[6996]);
    assign layer3_out[969] = ~layer2_out[421];
    assign layer3_out[970] = ~(layer2_out[5652] | layer2_out[5653]);
    assign layer3_out[971] = layer2_out[4371] & layer2_out[4372];
    assign layer3_out[972] = layer2_out[4218] & ~layer2_out[4219];
    assign layer3_out[973] = layer2_out[4793];
    assign layer3_out[974] = layer2_out[3152] & ~layer2_out[3151];
    assign layer3_out[975] = layer2_out[4459] & layer2_out[4460];
    assign layer3_out[976] = layer2_out[3116] ^ layer2_out[3117];
    assign layer3_out[977] = layer2_out[4383];
    assign layer3_out[978] = layer2_out[574] & layer2_out[575];
    assign layer3_out[979] = layer2_out[3478];
    assign layer3_out[980] = layer2_out[4227];
    assign layer3_out[981] = ~layer2_out[7235];
    assign layer3_out[982] = ~(layer2_out[3547] & layer2_out[3548]);
    assign layer3_out[983] = ~(layer2_out[4377] ^ layer2_out[4378]);
    assign layer3_out[984] = layer2_out[1279] | layer2_out[1280];
    assign layer3_out[985] = ~layer2_out[7821] | layer2_out[7822];
    assign layer3_out[986] = layer2_out[6068];
    assign layer3_out[987] = layer2_out[5852];
    assign layer3_out[988] = ~layer2_out[841];
    assign layer3_out[989] = ~layer2_out[5233];
    assign layer3_out[990] = ~layer2_out[6888] | layer2_out[6889];
    assign layer3_out[991] = ~layer2_out[3645] | layer2_out[3646];
    assign layer3_out[992] = layer2_out[5204] ^ layer2_out[5205];
    assign layer3_out[993] = layer2_out[4049] & ~layer2_out[4050];
    assign layer3_out[994] = layer2_out[1416];
    assign layer3_out[995] = layer2_out[2590] | layer2_out[2591];
    assign layer3_out[996] = ~layer2_out[2302];
    assign layer3_out[997] = layer2_out[5961] | layer2_out[5962];
    assign layer3_out[998] = 1'b0;
    assign layer3_out[999] = ~layer2_out[3691];
    assign layer3_out[1000] = ~layer2_out[2857];
    assign layer3_out[1001] = layer2_out[1319];
    assign layer3_out[1002] = ~layer2_out[617] | layer2_out[618];
    assign layer3_out[1003] = layer2_out[7439] | layer2_out[7440];
    assign layer3_out[1004] = ~layer2_out[3674] | layer2_out[3673];
    assign layer3_out[1005] = ~layer2_out[6353];
    assign layer3_out[1006] = layer2_out[3332] & ~layer2_out[3333];
    assign layer3_out[1007] = ~layer2_out[5182] | layer2_out[5183];
    assign layer3_out[1008] = ~layer2_out[757];
    assign layer3_out[1009] = layer2_out[4358] & ~layer2_out[4359];
    assign layer3_out[1010] = layer2_out[3981];
    assign layer3_out[1011] = layer2_out[5791] & ~layer2_out[5792];
    assign layer3_out[1012] = 1'b1;
    assign layer3_out[1013] = layer2_out[4045];
    assign layer3_out[1014] = ~layer2_out[4122];
    assign layer3_out[1015] = layer2_out[547];
    assign layer3_out[1016] = ~layer2_out[6944] | layer2_out[6943];
    assign layer3_out[1017] = ~(layer2_out[2703] & layer2_out[2704]);
    assign layer3_out[1018] = layer2_out[1898];
    assign layer3_out[1019] = layer2_out[3828];
    assign layer3_out[1020] = layer2_out[1362] ^ layer2_out[1363];
    assign layer3_out[1021] = ~(layer2_out[7418] | layer2_out[7419]);
    assign layer3_out[1022] = ~layer2_out[7869] | layer2_out[7870];
    assign layer3_out[1023] = layer2_out[6532] & ~layer2_out[6533];
    assign layer3_out[1024] = ~layer2_out[4599];
    assign layer3_out[1025] = layer2_out[4747] & layer2_out[4748];
    assign layer3_out[1026] = ~(layer2_out[3422] ^ layer2_out[3423]);
    assign layer3_out[1027] = layer2_out[2795] & ~layer2_out[2794];
    assign layer3_out[1028] = ~(layer2_out[5706] | layer2_out[5707]);
    assign layer3_out[1029] = layer2_out[6681] | layer2_out[6682];
    assign layer3_out[1030] = layer2_out[6420];
    assign layer3_out[1031] = layer2_out[2851];
    assign layer3_out[1032] = ~layer2_out[352] | layer2_out[353];
    assign layer3_out[1033] = layer2_out[3580];
    assign layer3_out[1034] = ~(layer2_out[4024] | layer2_out[4025]);
    assign layer3_out[1035] = 1'b1;
    assign layer3_out[1036] = ~layer2_out[3226];
    assign layer3_out[1037] = layer2_out[2550];
    assign layer3_out[1038] = ~layer2_out[5202];
    assign layer3_out[1039] = layer2_out[598];
    assign layer3_out[1040] = ~layer2_out[4137];
    assign layer3_out[1041] = ~layer2_out[6125] | layer2_out[6126];
    assign layer3_out[1042] = layer2_out[3576];
    assign layer3_out[1043] = layer2_out[4751] & layer2_out[4752];
    assign layer3_out[1044] = layer2_out[7340] & layer2_out[7341];
    assign layer3_out[1045] = layer2_out[70] ^ layer2_out[71];
    assign layer3_out[1046] = 1'b1;
    assign layer3_out[1047] = 1'b1;
    assign layer3_out[1048] = layer2_out[2426];
    assign layer3_out[1049] = layer2_out[3875];
    assign layer3_out[1050] = ~layer2_out[114];
    assign layer3_out[1051] = ~layer2_out[6398] | layer2_out[6397];
    assign layer3_out[1052] = layer2_out[3693] ^ layer2_out[3694];
    assign layer3_out[1053] = ~layer2_out[5205] | layer2_out[5206];
    assign layer3_out[1054] = layer2_out[1174];
    assign layer3_out[1055] = layer2_out[4379];
    assign layer3_out[1056] = ~layer2_out[3940];
    assign layer3_out[1057] = ~layer2_out[3873];
    assign layer3_out[1058] = ~layer2_out[3899];
    assign layer3_out[1059] = layer2_out[5904] | layer2_out[5905];
    assign layer3_out[1060] = ~(layer2_out[493] ^ layer2_out[494]);
    assign layer3_out[1061] = layer2_out[6408];
    assign layer3_out[1062] = ~(layer2_out[5959] | layer2_out[5960]);
    assign layer3_out[1063] = layer2_out[399];
    assign layer3_out[1064] = ~layer2_out[5183] | layer2_out[5184];
    assign layer3_out[1065] = layer2_out[6298];
    assign layer3_out[1066] = ~layer2_out[1078] | layer2_out[1077];
    assign layer3_out[1067] = layer2_out[1564] & layer2_out[1565];
    assign layer3_out[1068] = layer2_out[4168] & layer2_out[4169];
    assign layer3_out[1069] = layer2_out[1960] & layer2_out[1961];
    assign layer3_out[1070] = ~layer2_out[5172];
    assign layer3_out[1071] = layer2_out[1837] ^ layer2_out[1838];
    assign layer3_out[1072] = layer2_out[1017];
    assign layer3_out[1073] = layer2_out[357] & layer2_out[358];
    assign layer3_out[1074] = layer2_out[2173];
    assign layer3_out[1075] = ~layer2_out[302];
    assign layer3_out[1076] = layer2_out[398] | layer2_out[399];
    assign layer3_out[1077] = ~layer2_out[2300];
    assign layer3_out[1078] = ~(layer2_out[7191] & layer2_out[7192]);
    assign layer3_out[1079] = layer2_out[6202] & ~layer2_out[6203];
    assign layer3_out[1080] = ~(layer2_out[1804] ^ layer2_out[1805]);
    assign layer3_out[1081] = layer2_out[794] & ~layer2_out[793];
    assign layer3_out[1082] = ~layer2_out[4223];
    assign layer3_out[1083] = layer2_out[4079];
    assign layer3_out[1084] = layer2_out[1073];
    assign layer3_out[1085] = layer2_out[5893];
    assign layer3_out[1086] = ~(layer2_out[7213] & layer2_out[7214]);
    assign layer3_out[1087] = ~(layer2_out[2688] ^ layer2_out[2689]);
    assign layer3_out[1088] = ~layer2_out[4455] | layer2_out[4454];
    assign layer3_out[1089] = layer2_out[1906] & ~layer2_out[1907];
    assign layer3_out[1090] = ~layer2_out[5408] | layer2_out[5409];
    assign layer3_out[1091] = layer2_out[6920] & ~layer2_out[6919];
    assign layer3_out[1092] = layer2_out[5397] & layer2_out[5398];
    assign layer3_out[1093] = layer2_out[1764] & ~layer2_out[1763];
    assign layer3_out[1094] = layer2_out[4938];
    assign layer3_out[1095] = ~layer2_out[1184];
    assign layer3_out[1096] = layer2_out[787] & ~layer2_out[786];
    assign layer3_out[1097] = layer2_out[5346];
    assign layer3_out[1098] = ~layer2_out[3805];
    assign layer3_out[1099] = layer2_out[7777];
    assign layer3_out[1100] = ~layer2_out[570];
    assign layer3_out[1101] = layer2_out[4216];
    assign layer3_out[1102] = layer2_out[6414];
    assign layer3_out[1103] = layer2_out[3551];
    assign layer3_out[1104] = ~layer2_out[1353] | layer2_out[1354];
    assign layer3_out[1105] = 1'b1;
    assign layer3_out[1106] = ~(layer2_out[6792] ^ layer2_out[6793]);
    assign layer3_out[1107] = ~layer2_out[4910];
    assign layer3_out[1108] = ~layer2_out[3695];
    assign layer3_out[1109] = ~layer2_out[6270] | layer2_out[6271];
    assign layer3_out[1110] = layer2_out[4820];
    assign layer3_out[1111] = layer2_out[1172] & layer2_out[1173];
    assign layer3_out[1112] = layer2_out[7314];
    assign layer3_out[1113] = layer2_out[5728];
    assign layer3_out[1114] = ~layer2_out[3139];
    assign layer3_out[1115] = layer2_out[2847];
    assign layer3_out[1116] = ~layer2_out[6362] | layer2_out[6361];
    assign layer3_out[1117] = ~(layer2_out[3574] & layer2_out[3575]);
    assign layer3_out[1118] = ~(layer2_out[222] | layer2_out[223]);
    assign layer3_out[1119] = ~(layer2_out[5644] ^ layer2_out[5645]);
    assign layer3_out[1120] = layer2_out[2965] & ~layer2_out[2966];
    assign layer3_out[1121] = ~layer2_out[5224];
    assign layer3_out[1122] = ~layer2_out[6960] | layer2_out[6961];
    assign layer3_out[1123] = ~layer2_out[449] | layer2_out[448];
    assign layer3_out[1124] = layer2_out[3070];
    assign layer3_out[1125] = 1'b1;
    assign layer3_out[1126] = ~(layer2_out[5771] | layer2_out[5772]);
    assign layer3_out[1127] = layer2_out[4285] ^ layer2_out[4286];
    assign layer3_out[1128] = ~layer2_out[7721] | layer2_out[7722];
    assign layer3_out[1129] = layer2_out[5832] & ~layer2_out[5833];
    assign layer3_out[1130] = ~layer2_out[4486] | layer2_out[4485];
    assign layer3_out[1131] = layer2_out[2322] | layer2_out[2323];
    assign layer3_out[1132] = ~layer2_out[5309] | layer2_out[5310];
    assign layer3_out[1133] = ~(layer2_out[2228] & layer2_out[2229]);
    assign layer3_out[1134] = layer2_out[6073] & ~layer2_out[6072];
    assign layer3_out[1135] = ~layer2_out[1940];
    assign layer3_out[1136] = ~(layer2_out[5823] & layer2_out[5824]);
    assign layer3_out[1137] = layer2_out[3177] ^ layer2_out[3178];
    assign layer3_out[1138] = ~(layer2_out[6385] ^ layer2_out[6386]);
    assign layer3_out[1139] = layer2_out[1888] & layer2_out[1889];
    assign layer3_out[1140] = layer2_out[6131] | layer2_out[6132];
    assign layer3_out[1141] = layer2_out[7350] | layer2_out[7351];
    assign layer3_out[1142] = layer2_out[1507] & ~layer2_out[1508];
    assign layer3_out[1143] = layer2_out[1114] | layer2_out[1115];
    assign layer3_out[1144] = layer2_out[602];
    assign layer3_out[1145] = 1'b1;
    assign layer3_out[1146] = layer2_out[2172] ^ layer2_out[2173];
    assign layer3_out[1147] = ~(layer2_out[1291] ^ layer2_out[1292]);
    assign layer3_out[1148] = layer2_out[3038];
    assign layer3_out[1149] = ~layer2_out[1262];
    assign layer3_out[1150] = layer2_out[7493] ^ layer2_out[7494];
    assign layer3_out[1151] = layer2_out[4782] & ~layer2_out[4781];
    assign layer3_out[1152] = ~layer2_out[6411];
    assign layer3_out[1153] = ~(layer2_out[374] ^ layer2_out[375]);
    assign layer3_out[1154] = ~(layer2_out[3105] & layer2_out[3106]);
    assign layer3_out[1155] = layer2_out[3365] ^ layer2_out[3366];
    assign layer3_out[1156] = layer2_out[1725];
    assign layer3_out[1157] = ~layer2_out[2118] | layer2_out[2119];
    assign layer3_out[1158] = ~(layer2_out[7098] | layer2_out[7099]);
    assign layer3_out[1159] = ~layer2_out[3543];
    assign layer3_out[1160] = layer2_out[4974] & layer2_out[4975];
    assign layer3_out[1161] = ~layer2_out[1648];
    assign layer3_out[1162] = ~(layer2_out[7042] & layer2_out[7043]);
    assign layer3_out[1163] = ~(layer2_out[5650] & layer2_out[5651]);
    assign layer3_out[1164] = 1'b1;
    assign layer3_out[1165] = ~(layer2_out[5159] & layer2_out[5160]);
    assign layer3_out[1166] = ~(layer2_out[3075] & layer2_out[3076]);
    assign layer3_out[1167] = layer2_out[6635];
    assign layer3_out[1168] = ~layer2_out[7872] | layer2_out[7873];
    assign layer3_out[1169] = ~layer2_out[1159];
    assign layer3_out[1170] = layer2_out[2641];
    assign layer3_out[1171] = ~layer2_out[7622];
    assign layer3_out[1172] = ~(layer2_out[3074] | layer2_out[3075]);
    assign layer3_out[1173] = layer2_out[5770];
    assign layer3_out[1174] = layer2_out[7941];
    assign layer3_out[1175] = ~layer2_out[5147];
    assign layer3_out[1176] = ~layer2_out[5372];
    assign layer3_out[1177] = layer2_out[1359] & ~layer2_out[1360];
    assign layer3_out[1178] = layer2_out[7965] & layer2_out[7966];
    assign layer3_out[1179] = layer2_out[4784] & layer2_out[4785];
    assign layer3_out[1180] = layer2_out[1818];
    assign layer3_out[1181] = ~layer2_out[3670];
    assign layer3_out[1182] = layer2_out[4244];
    assign layer3_out[1183] = layer2_out[566] | layer2_out[567];
    assign layer3_out[1184] = layer2_out[1607];
    assign layer3_out[1185] = ~layer2_out[4824];
    assign layer3_out[1186] = ~layer2_out[2346] | layer2_out[2347];
    assign layer3_out[1187] = ~layer2_out[6978] | layer2_out[6979];
    assign layer3_out[1188] = layer2_out[385] & ~layer2_out[384];
    assign layer3_out[1189] = layer2_out[3340] & layer2_out[3341];
    assign layer3_out[1190] = layer2_out[7237] & layer2_out[7238];
    assign layer3_out[1191] = 1'b1;
    assign layer3_out[1192] = ~layer2_out[6558] | layer2_out[6559];
    assign layer3_out[1193] = ~layer2_out[3277];
    assign layer3_out[1194] = 1'b0;
    assign layer3_out[1195] = ~(layer2_out[1809] & layer2_out[1810]);
    assign layer3_out[1196] = ~layer2_out[3108];
    assign layer3_out[1197] = ~(layer2_out[927] ^ layer2_out[928]);
    assign layer3_out[1198] = layer2_out[6883] & layer2_out[6884];
    assign layer3_out[1199] = layer2_out[5907] & ~layer2_out[5906];
    assign layer3_out[1200] = layer2_out[3977];
    assign layer3_out[1201] = ~layer2_out[6163];
    assign layer3_out[1202] = layer2_out[7626] & ~layer2_out[7625];
    assign layer3_out[1203] = layer2_out[361] & layer2_out[362];
    assign layer3_out[1204] = layer2_out[7320] | layer2_out[7321];
    assign layer3_out[1205] = layer2_out[6141];
    assign layer3_out[1206] = ~(layer2_out[6336] | layer2_out[6337]);
    assign layer3_out[1207] = ~(layer2_out[3892] ^ layer2_out[3893]);
    assign layer3_out[1208] = layer2_out[4998] & layer2_out[4999];
    assign layer3_out[1209] = ~layer2_out[658];
    assign layer3_out[1210] = layer2_out[703] ^ layer2_out[704];
    assign layer3_out[1211] = layer2_out[4282] & ~layer2_out[4281];
    assign layer3_out[1212] = ~(layer2_out[4805] ^ layer2_out[4806]);
    assign layer3_out[1213] = layer2_out[7363];
    assign layer3_out[1214] = ~layer2_out[5069] | layer2_out[5070];
    assign layer3_out[1215] = layer2_out[2064] ^ layer2_out[2065];
    assign layer3_out[1216] = layer2_out[2217] | layer2_out[2218];
    assign layer3_out[1217] = layer2_out[2742];
    assign layer3_out[1218] = ~layer2_out[288] | layer2_out[289];
    assign layer3_out[1219] = ~layer2_out[2007] | layer2_out[2006];
    assign layer3_out[1220] = ~layer2_out[5409];
    assign layer3_out[1221] = ~layer2_out[707];
    assign layer3_out[1222] = layer2_out[74] & layer2_out[75];
    assign layer3_out[1223] = layer2_out[3926];
    assign layer3_out[1224] = layer2_out[6888];
    assign layer3_out[1225] = layer2_out[429] & ~layer2_out[430];
    assign layer3_out[1226] = layer2_out[1595];
    assign layer3_out[1227] = layer2_out[5898];
    assign layer3_out[1228] = layer2_out[7772];
    assign layer3_out[1229] = layer2_out[298];
    assign layer3_out[1230] = ~layer2_out[4297];
    assign layer3_out[1231] = ~(layer2_out[3183] ^ layer2_out[3184]);
    assign layer3_out[1232] = layer2_out[4104] & layer2_out[4105];
    assign layer3_out[1233] = layer2_out[901] & ~layer2_out[902];
    assign layer3_out[1234] = ~(layer2_out[3913] | layer2_out[3914]);
    assign layer3_out[1235] = layer2_out[856] ^ layer2_out[857];
    assign layer3_out[1236] = ~layer2_out[3174];
    assign layer3_out[1237] = layer2_out[3029] & ~layer2_out[3028];
    assign layer3_out[1238] = 1'b1;
    assign layer3_out[1239] = layer2_out[6605] ^ layer2_out[6606];
    assign layer3_out[1240] = 1'b0;
    assign layer3_out[1241] = ~(layer2_out[5597] ^ layer2_out[5598]);
    assign layer3_out[1242] = layer2_out[3791] & ~layer2_out[3792];
    assign layer3_out[1243] = layer2_out[3102];
    assign layer3_out[1244] = ~(layer2_out[1220] & layer2_out[1221]);
    assign layer3_out[1245] = layer2_out[5275];
    assign layer3_out[1246] = layer2_out[4108];
    assign layer3_out[1247] = ~layer2_out[1012];
    assign layer3_out[1248] = ~(layer2_out[6974] & layer2_out[6975]);
    assign layer3_out[1249] = layer2_out[2466] ^ layer2_out[2467];
    assign layer3_out[1250] = layer2_out[4507] & layer2_out[4508];
    assign layer3_out[1251] = layer2_out[2338] ^ layer2_out[2339];
    assign layer3_out[1252] = layer2_out[263];
    assign layer3_out[1253] = layer2_out[5495];
    assign layer3_out[1254] = layer2_out[4546] & ~layer2_out[4547];
    assign layer3_out[1255] = layer2_out[4308];
    assign layer3_out[1256] = layer2_out[1088] & layer2_out[1089];
    assign layer3_out[1257] = layer2_out[1394];
    assign layer3_out[1258] = ~layer2_out[3835];
    assign layer3_out[1259] = layer2_out[1225] | layer2_out[1226];
    assign layer3_out[1260] = ~layer2_out[2589];
    assign layer3_out[1261] = layer2_out[3426];
    assign layer3_out[1262] = layer2_out[7660];
    assign layer3_out[1263] = ~layer2_out[2265];
    assign layer3_out[1264] = layer2_out[3697] & ~layer2_out[3696];
    assign layer3_out[1265] = ~layer2_out[3664];
    assign layer3_out[1266] = layer2_out[2726] & ~layer2_out[2727];
    assign layer3_out[1267] = ~(layer2_out[4734] | layer2_out[4735]);
    assign layer3_out[1268] = ~(layer2_out[7550] & layer2_out[7551]);
    assign layer3_out[1269] = layer2_out[5396] & ~layer2_out[5395];
    assign layer3_out[1270] = 1'b0;
    assign layer3_out[1271] = layer2_out[4010] & layer2_out[4011];
    assign layer3_out[1272] = ~layer2_out[863];
    assign layer3_out[1273] = layer2_out[4455] & ~layer2_out[4456];
    assign layer3_out[1274] = ~(layer2_out[3727] ^ layer2_out[3728]);
    assign layer3_out[1275] = layer2_out[44] & ~layer2_out[43];
    assign layer3_out[1276] = layer2_out[1167] ^ layer2_out[1168];
    assign layer3_out[1277] = ~layer2_out[2762];
    assign layer3_out[1278] = ~(layer2_out[1050] & layer2_out[1051]);
    assign layer3_out[1279] = layer2_out[4628] & layer2_out[4629];
    assign layer3_out[1280] = ~layer2_out[7903];
    assign layer3_out[1281] = layer2_out[495] ^ layer2_out[496];
    assign layer3_out[1282] = layer2_out[187];
    assign layer3_out[1283] = layer2_out[3887] | layer2_out[3888];
    assign layer3_out[1284] = layer2_out[3460] & layer2_out[3461];
    assign layer3_out[1285] = ~layer2_out[2605] | layer2_out[2606];
    assign layer3_out[1286] = ~(layer2_out[2735] & layer2_out[2736]);
    assign layer3_out[1287] = layer2_out[4499] | layer2_out[4500];
    assign layer3_out[1288] = layer2_out[431] | layer2_out[432];
    assign layer3_out[1289] = ~layer2_out[6384];
    assign layer3_out[1290] = ~layer2_out[4999];
    assign layer3_out[1291] = layer2_out[655] | layer2_out[656];
    assign layer3_out[1292] = layer2_out[4640] ^ layer2_out[4641];
    assign layer3_out[1293] = ~(layer2_out[5667] ^ layer2_out[5668]);
    assign layer3_out[1294] = layer2_out[4334] & layer2_out[4335];
    assign layer3_out[1295] = layer2_out[591] & ~layer2_out[592];
    assign layer3_out[1296] = ~(layer2_out[6581] | layer2_out[6582]);
    assign layer3_out[1297] = layer2_out[3534];
    assign layer3_out[1298] = ~layer2_out[1502] | layer2_out[1501];
    assign layer3_out[1299] = ~(layer2_out[1953] | layer2_out[1954]);
    assign layer3_out[1300] = ~layer2_out[7442];
    assign layer3_out[1301] = layer2_out[695];
    assign layer3_out[1302] = ~(layer2_out[2558] & layer2_out[2559]);
    assign layer3_out[1303] = layer2_out[4882];
    assign layer3_out[1304] = ~(layer2_out[1756] | layer2_out[1757]);
    assign layer3_out[1305] = layer2_out[7080];
    assign layer3_out[1306] = layer2_out[4230] & ~layer2_out[4229];
    assign layer3_out[1307] = ~layer2_out[4646];
    assign layer3_out[1308] = ~(layer2_out[4318] ^ layer2_out[4319]);
    assign layer3_out[1309] = ~layer2_out[1167];
    assign layer3_out[1310] = ~layer2_out[6181];
    assign layer3_out[1311] = ~layer2_out[1757];
    assign layer3_out[1312] = ~(layer2_out[1590] ^ layer2_out[1591]);
    assign layer3_out[1313] = ~layer2_out[3506];
    assign layer3_out[1314] = layer2_out[2218] ^ layer2_out[2219];
    assign layer3_out[1315] = layer2_out[3043] & ~layer2_out[3042];
    assign layer3_out[1316] = ~(layer2_out[4309] ^ layer2_out[4310]);
    assign layer3_out[1317] = ~(layer2_out[5932] & layer2_out[5933]);
    assign layer3_out[1318] = layer2_out[6681];
    assign layer3_out[1319] = layer2_out[5207] ^ layer2_out[5208];
    assign layer3_out[1320] = layer2_out[2113];
    assign layer3_out[1321] = ~layer2_out[5944];
    assign layer3_out[1322] = layer2_out[5084] ^ layer2_out[5085];
    assign layer3_out[1323] = layer2_out[2706];
    assign layer3_out[1324] = ~layer2_out[7831];
    assign layer3_out[1325] = layer2_out[3751];
    assign layer3_out[1326] = layer2_out[7326] & ~layer2_out[7327];
    assign layer3_out[1327] = ~layer2_out[3241];
    assign layer3_out[1328] = ~layer2_out[3995];
    assign layer3_out[1329] = ~layer2_out[2242] | layer2_out[2241];
    assign layer3_out[1330] = layer2_out[5449] | layer2_out[5450];
    assign layer3_out[1331] = ~(layer2_out[3443] & layer2_out[3444]);
    assign layer3_out[1332] = layer2_out[6937] ^ layer2_out[6938];
    assign layer3_out[1333] = layer2_out[3262];
    assign layer3_out[1334] = ~layer2_out[5213];
    assign layer3_out[1335] = layer2_out[759];
    assign layer3_out[1336] = layer2_out[293] & ~layer2_out[294];
    assign layer3_out[1337] = layer2_out[2870] & ~layer2_out[2869];
    assign layer3_out[1338] = ~layer2_out[4013] | layer2_out[4012];
    assign layer3_out[1339] = ~layer2_out[4479];
    assign layer3_out[1340] = layer2_out[3751];
    assign layer3_out[1341] = 1'b0;
    assign layer3_out[1342] = ~layer2_out[3238] | layer2_out[3237];
    assign layer3_out[1343] = layer2_out[4202];
    assign layer3_out[1344] = ~layer2_out[5796] | layer2_out[5795];
    assign layer3_out[1345] = ~layer2_out[6285] | layer2_out[6286];
    assign layer3_out[1346] = ~layer2_out[4079] | layer2_out[4080];
    assign layer3_out[1347] = ~layer2_out[7542];
    assign layer3_out[1348] = layer2_out[6799];
    assign layer3_out[1349] = layer2_out[6657] & layer2_out[6658];
    assign layer3_out[1350] = ~(layer2_out[1487] ^ layer2_out[1488]);
    assign layer3_out[1351] = layer2_out[1614];
    assign layer3_out[1352] = layer2_out[2341] | layer2_out[2342];
    assign layer3_out[1353] = layer2_out[6113] ^ layer2_out[6114];
    assign layer3_out[1354] = layer2_out[5973] & layer2_out[5974];
    assign layer3_out[1355] = layer2_out[6352];
    assign layer3_out[1356] = layer2_out[3948] & ~layer2_out[3949];
    assign layer3_out[1357] = layer2_out[641];
    assign layer3_out[1358] = layer2_out[6721] & ~layer2_out[6722];
    assign layer3_out[1359] = layer2_out[1030] & layer2_out[1031];
    assign layer3_out[1360] = ~layer2_out[5166];
    assign layer3_out[1361] = ~layer2_out[2807] | layer2_out[2806];
    assign layer3_out[1362] = layer2_out[6909] ^ layer2_out[6910];
    assign layer3_out[1363] = ~(layer2_out[5960] & layer2_out[5961]);
    assign layer3_out[1364] = ~layer2_out[2277] | layer2_out[2276];
    assign layer3_out[1365] = layer2_out[428] & layer2_out[429];
    assign layer3_out[1366] = layer2_out[6999] | layer2_out[7000];
    assign layer3_out[1367] = ~layer2_out[5487];
    assign layer3_out[1368] = ~layer2_out[4202] | layer2_out[4201];
    assign layer3_out[1369] = ~(layer2_out[3201] | layer2_out[3202]);
    assign layer3_out[1370] = ~layer2_out[6384];
    assign layer3_out[1371] = ~layer2_out[1273];
    assign layer3_out[1372] = ~layer2_out[3453];
    assign layer3_out[1373] = ~layer2_out[5845];
    assign layer3_out[1374] = layer2_out[5770] & ~layer2_out[5771];
    assign layer3_out[1375] = ~layer2_out[4317];
    assign layer3_out[1376] = ~(layer2_out[887] ^ layer2_out[888]);
    assign layer3_out[1377] = ~layer2_out[3982];
    assign layer3_out[1378] = ~layer2_out[933];
    assign layer3_out[1379] = ~layer2_out[5969];
    assign layer3_out[1380] = ~(layer2_out[1492] & layer2_out[1493]);
    assign layer3_out[1381] = layer2_out[976];
    assign layer3_out[1382] = layer2_out[5921] & ~layer2_out[5922];
    assign layer3_out[1383] = layer2_out[903];
    assign layer3_out[1384] = layer2_out[186] & ~layer2_out[185];
    assign layer3_out[1385] = ~layer2_out[4417];
    assign layer3_out[1386] = ~layer2_out[5882];
    assign layer3_out[1387] = ~(layer2_out[100] | layer2_out[101]);
    assign layer3_out[1388] = layer2_out[1744] ^ layer2_out[1745];
    assign layer3_out[1389] = ~layer2_out[1575];
    assign layer3_out[1390] = layer2_out[4846];
    assign layer3_out[1391] = ~(layer2_out[4276] & layer2_out[4277]);
    assign layer3_out[1392] = ~layer2_out[3000];
    assign layer3_out[1393] = layer2_out[7409];
    assign layer3_out[1394] = layer2_out[4390];
    assign layer3_out[1395] = layer2_out[5253];
    assign layer3_out[1396] = ~layer2_out[2419];
    assign layer3_out[1397] = layer2_out[7148] & ~layer2_out[7147];
    assign layer3_out[1398] = layer2_out[4905] & layer2_out[4906];
    assign layer3_out[1399] = 1'b1;
    assign layer3_out[1400] = layer2_out[3623] & ~layer2_out[3622];
    assign layer3_out[1401] = layer2_out[7779] & ~layer2_out[7780];
    assign layer3_out[1402] = layer2_out[2643] & layer2_out[2644];
    assign layer3_out[1403] = layer2_out[7231];
    assign layer3_out[1404] = ~layer2_out[1403];
    assign layer3_out[1405] = layer2_out[285] & layer2_out[286];
    assign layer3_out[1406] = layer2_out[1094] | layer2_out[1095];
    assign layer3_out[1407] = layer2_out[5150] & ~layer2_out[5151];
    assign layer3_out[1408] = ~layer2_out[4870];
    assign layer3_out[1409] = ~layer2_out[4332];
    assign layer3_out[1410] = layer2_out[7615] & layer2_out[7616];
    assign layer3_out[1411] = ~layer2_out[6638];
    assign layer3_out[1412] = ~layer2_out[3198];
    assign layer3_out[1413] = layer2_out[1072];
    assign layer3_out[1414] = ~layer2_out[5572];
    assign layer3_out[1415] = ~(layer2_out[1200] ^ layer2_out[1201]);
    assign layer3_out[1416] = 1'b1;
    assign layer3_out[1417] = layer2_out[6808];
    assign layer3_out[1418] = layer2_out[2422] & ~layer2_out[2423];
    assign layer3_out[1419] = ~(layer2_out[2638] & layer2_out[2639]);
    assign layer3_out[1420] = layer2_out[588] & ~layer2_out[589];
    assign layer3_out[1421] = layer2_out[5292] & layer2_out[5293];
    assign layer3_out[1422] = layer2_out[979];
    assign layer3_out[1423] = 1'b0;
    assign layer3_out[1424] = layer2_out[6841] & ~layer2_out[6842];
    assign layer3_out[1425] = layer2_out[964] & ~layer2_out[963];
    assign layer3_out[1426] = ~(layer2_out[1620] & layer2_out[1621]);
    assign layer3_out[1427] = layer2_out[5142];
    assign layer3_out[1428] = layer2_out[6939];
    assign layer3_out[1429] = layer2_out[1406] ^ layer2_out[1407];
    assign layer3_out[1430] = ~(layer2_out[2909] | layer2_out[2910]);
    assign layer3_out[1431] = ~(layer2_out[6165] ^ layer2_out[6166]);
    assign layer3_out[1432] = layer2_out[5938];
    assign layer3_out[1433] = layer2_out[145] & ~layer2_out[146];
    assign layer3_out[1434] = layer2_out[6454];
    assign layer3_out[1435] = ~layer2_out[1799];
    assign layer3_out[1436] = layer2_out[1866];
    assign layer3_out[1437] = layer2_out[3350] & ~layer2_out[3351];
    assign layer3_out[1438] = layer2_out[822];
    assign layer3_out[1439] = layer2_out[3889] | layer2_out[3890];
    assign layer3_out[1440] = ~layer2_out[3458] | layer2_out[3457];
    assign layer3_out[1441] = ~layer2_out[7951];
    assign layer3_out[1442] = 1'b1;
    assign layer3_out[1443] = ~(layer2_out[6556] ^ layer2_out[6557]);
    assign layer3_out[1444] = layer2_out[1469];
    assign layer3_out[1445] = ~layer2_out[567] | layer2_out[568];
    assign layer3_out[1446] = layer2_out[3915] & layer2_out[3916];
    assign layer3_out[1447] = ~layer2_out[1512];
    assign layer3_out[1448] = layer2_out[923] & ~layer2_out[922];
    assign layer3_out[1449] = layer2_out[4231];
    assign layer3_out[1450] = ~layer2_out[2817] | layer2_out[2818];
    assign layer3_out[1451] = layer2_out[811] & ~layer2_out[812];
    assign layer3_out[1452] = layer2_out[2236];
    assign layer3_out[1453] = layer2_out[2112] ^ layer2_out[2113];
    assign layer3_out[1454] = layer2_out[328];
    assign layer3_out[1455] = ~layer2_out[7291] | layer2_out[7292];
    assign layer3_out[1456] = layer2_out[6181] & ~layer2_out[6182];
    assign layer3_out[1457] = layer2_out[6850];
    assign layer3_out[1458] = ~layer2_out[3581];
    assign layer3_out[1459] = layer2_out[5401];
    assign layer3_out[1460] = layer2_out[5596];
    assign layer3_out[1461] = ~(layer2_out[6994] & layer2_out[6995]);
    assign layer3_out[1462] = layer2_out[6678] ^ layer2_out[6679];
    assign layer3_out[1463] = ~(layer2_out[7238] | layer2_out[7239]);
    assign layer3_out[1464] = layer2_out[471];
    assign layer3_out[1465] = ~(layer2_out[1110] | layer2_out[1111]);
    assign layer3_out[1466] = ~layer2_out[2048];
    assign layer3_out[1467] = ~(layer2_out[6638] ^ layer2_out[6639]);
    assign layer3_out[1468] = ~layer2_out[2433] | layer2_out[2434];
    assign layer3_out[1469] = layer2_out[2260] & ~layer2_out[2259];
    assign layer3_out[1470] = layer2_out[7709];
    assign layer3_out[1471] = ~layer2_out[1322];
    assign layer3_out[1472] = layer2_out[6628] & ~layer2_out[6629];
    assign layer3_out[1473] = ~(layer2_out[5436] | layer2_out[5437]);
    assign layer3_out[1474] = layer2_out[750] & ~layer2_out[749];
    assign layer3_out[1475] = layer2_out[409];
    assign layer3_out[1476] = layer2_out[3318] & ~layer2_out[3319];
    assign layer3_out[1477] = ~(layer2_out[7563] & layer2_out[7564]);
    assign layer3_out[1478] = ~(layer2_out[6931] ^ layer2_out[6932]);
    assign layer3_out[1479] = ~layer2_out[6233];
    assign layer3_out[1480] = layer2_out[2170] | layer2_out[2171];
    assign layer3_out[1481] = layer2_out[125];
    assign layer3_out[1482] = ~layer2_out[5924];
    assign layer3_out[1483] = ~(layer2_out[3708] & layer2_out[3709]);
    assign layer3_out[1484] = layer2_out[61] & ~layer2_out[60];
    assign layer3_out[1485] = ~layer2_out[105];
    assign layer3_out[1486] = layer2_out[875] & ~layer2_out[876];
    assign layer3_out[1487] = ~layer2_out[5553] | layer2_out[5552];
    assign layer3_out[1488] = ~(layer2_out[1112] | layer2_out[1113]);
    assign layer3_out[1489] = layer2_out[2584];
    assign layer3_out[1490] = ~layer2_out[337];
    assign layer3_out[1491] = layer2_out[1531] ^ layer2_out[1532];
    assign layer3_out[1492] = layer2_out[2595];
    assign layer3_out[1493] = ~(layer2_out[1439] & layer2_out[1440]);
    assign layer3_out[1494] = layer2_out[1349] & layer2_out[1350];
    assign layer3_out[1495] = ~layer2_out[1006];
    assign layer3_out[1496] = ~(layer2_out[6717] & layer2_out[6718]);
    assign layer3_out[1497] = ~layer2_out[1629];
    assign layer3_out[1498] = 1'b0;
    assign layer3_out[1499] = ~layer2_out[3380];
    assign layer3_out[1500] = ~(layer2_out[5927] | layer2_out[5928]);
    assign layer3_out[1501] = layer2_out[7537] & ~layer2_out[7538];
    assign layer3_out[1502] = ~(layer2_out[5228] ^ layer2_out[5229]);
    assign layer3_out[1503] = layer2_out[1940];
    assign layer3_out[1504] = ~(layer2_out[833] | layer2_out[834]);
    assign layer3_out[1505] = layer2_out[2574];
    assign layer3_out[1506] = ~layer2_out[798];
    assign layer3_out[1507] = ~(layer2_out[7307] & layer2_out[7308]);
    assign layer3_out[1508] = layer2_out[1886] | layer2_out[1887];
    assign layer3_out[1509] = layer2_out[1151];
    assign layer3_out[1510] = layer2_out[2527];
    assign layer3_out[1511] = layer2_out[521] & layer2_out[522];
    assign layer3_out[1512] = layer2_out[5769] & ~layer2_out[5768];
    assign layer3_out[1513] = ~(layer2_out[675] & layer2_out[676]);
    assign layer3_out[1514] = ~layer2_out[3219];
    assign layer3_out[1515] = layer2_out[1466];
    assign layer3_out[1516] = layer2_out[1697];
    assign layer3_out[1517] = ~(layer2_out[3159] & layer2_out[3160]);
    assign layer3_out[1518] = ~layer2_out[5765];
    assign layer3_out[1519] = layer2_out[5989];
    assign layer3_out[1520] = ~(layer2_out[4444] ^ layer2_out[4445]);
    assign layer3_out[1521] = ~layer2_out[2306];
    assign layer3_out[1522] = layer2_out[5123] & ~layer2_out[5122];
    assign layer3_out[1523] = ~layer2_out[5526] | layer2_out[5525];
    assign layer3_out[1524] = ~layer2_out[1650] | layer2_out[1651];
    assign layer3_out[1525] = layer2_out[2889];
    assign layer3_out[1526] = layer2_out[7746];
    assign layer3_out[1527] = layer2_out[2882] & layer2_out[2883];
    assign layer3_out[1528] = ~(layer2_out[3638] & layer2_out[3639]);
    assign layer3_out[1529] = layer2_out[4552] & ~layer2_out[4553];
    assign layer3_out[1530] = layer2_out[1925] ^ layer2_out[1926];
    assign layer3_out[1531] = ~(layer2_out[6764] ^ layer2_out[6765]);
    assign layer3_out[1532] = ~layer2_out[1406];
    assign layer3_out[1533] = 1'b0;
    assign layer3_out[1534] = ~layer2_out[5118];
    assign layer3_out[1535] = ~(layer2_out[5123] ^ layer2_out[5124]);
    assign layer3_out[1536] = layer2_out[5707] | layer2_out[5708];
    assign layer3_out[1537] = layer2_out[2510] & layer2_out[2511];
    assign layer3_out[1538] = ~(layer2_out[4121] | layer2_out[4122]);
    assign layer3_out[1539] = layer2_out[510] & ~layer2_out[509];
    assign layer3_out[1540] = ~layer2_out[1025];
    assign layer3_out[1541] = ~(layer2_out[5414] | layer2_out[5415]);
    assign layer3_out[1542] = layer2_out[3522];
    assign layer3_out[1543] = layer2_out[6379] & ~layer2_out[6378];
    assign layer3_out[1544] = layer2_out[1142] & ~layer2_out[1141];
    assign layer3_out[1545] = layer2_out[7345] & layer2_out[7346];
    assign layer3_out[1546] = layer2_out[3473];
    assign layer3_out[1547] = layer2_out[208];
    assign layer3_out[1548] = layer2_out[3827] | layer2_out[3828];
    assign layer3_out[1549] = ~(layer2_out[7194] & layer2_out[7195]);
    assign layer3_out[1550] = ~layer2_out[2576];
    assign layer3_out[1551] = ~layer2_out[4890];
    assign layer3_out[1552] = layer2_out[7281] & layer2_out[7282];
    assign layer3_out[1553] = ~(layer2_out[2162] ^ layer2_out[2163]);
    assign layer3_out[1554] = ~layer2_out[3287];
    assign layer3_out[1555] = layer2_out[3611] | layer2_out[3612];
    assign layer3_out[1556] = layer2_out[6710];
    assign layer3_out[1557] = layer2_out[5434] | layer2_out[5435];
    assign layer3_out[1558] = ~layer2_out[7220];
    assign layer3_out[1559] = ~(layer2_out[5809] & layer2_out[5810]);
    assign layer3_out[1560] = layer2_out[5799] & ~layer2_out[5798];
    assign layer3_out[1561] = ~(layer2_out[4510] & layer2_out[4511]);
    assign layer3_out[1562] = ~(layer2_out[2994] | layer2_out[2995]);
    assign layer3_out[1563] = ~(layer2_out[7889] ^ layer2_out[7890]);
    assign layer3_out[1564] = layer2_out[2322];
    assign layer3_out[1565] = ~layer2_out[1791] | layer2_out[1790];
    assign layer3_out[1566] = layer2_out[1312] & ~layer2_out[1313];
    assign layer3_out[1567] = ~layer2_out[544] | layer2_out[543];
    assign layer3_out[1568] = ~layer2_out[3655] | layer2_out[3656];
    assign layer3_out[1569] = layer2_out[4194];
    assign layer3_out[1570] = layer2_out[7534] | layer2_out[7535];
    assign layer3_out[1571] = layer2_out[2259];
    assign layer3_out[1572] = ~layer2_out[2672];
    assign layer3_out[1573] = layer2_out[5931] ^ layer2_out[5932];
    assign layer3_out[1574] = layer2_out[527] ^ layer2_out[528];
    assign layer3_out[1575] = ~layer2_out[3522];
    assign layer3_out[1576] = ~(layer2_out[5203] & layer2_out[5204]);
    assign layer3_out[1577] = layer2_out[1916];
    assign layer3_out[1578] = layer2_out[1081] ^ layer2_out[1082];
    assign layer3_out[1579] = ~layer2_out[1223] | layer2_out[1222];
    assign layer3_out[1580] = 1'b0;
    assign layer3_out[1581] = layer2_out[5391];
    assign layer3_out[1582] = ~(layer2_out[5538] & layer2_out[5539]);
    assign layer3_out[1583] = layer2_out[903] | layer2_out[904];
    assign layer3_out[1584] = layer2_out[1047];
    assign layer3_out[1585] = layer2_out[7311] | layer2_out[7312];
    assign layer3_out[1586] = ~layer2_out[4402];
    assign layer3_out[1587] = ~layer2_out[1657];
    assign layer3_out[1588] = ~layer2_out[6013];
    assign layer3_out[1589] = layer2_out[6471] ^ layer2_out[6472];
    assign layer3_out[1590] = ~layer2_out[1687];
    assign layer3_out[1591] = ~layer2_out[1624] | layer2_out[1625];
    assign layer3_out[1592] = layer2_out[6812];
    assign layer3_out[1593] = layer2_out[3012] & ~layer2_out[3013];
    assign layer3_out[1594] = 1'b0;
    assign layer3_out[1595] = layer2_out[3384] & ~layer2_out[3385];
    assign layer3_out[1596] = layer2_out[2759] ^ layer2_out[2760];
    assign layer3_out[1597] = layer2_out[6329];
    assign layer3_out[1598] = layer2_out[5997] & ~layer2_out[5996];
    assign layer3_out[1599] = ~(layer2_out[6201] & layer2_out[6202]);
    assign layer3_out[1600] = ~layer2_out[1232];
    assign layer3_out[1601] = ~(layer2_out[1289] ^ layer2_out[1290]);
    assign layer3_out[1602] = layer2_out[5306];
    assign layer3_out[1603] = layer2_out[5603] | layer2_out[5604];
    assign layer3_out[1604] = layer2_out[3080];
    assign layer3_out[1605] = layer2_out[4175];
    assign layer3_out[1606] = layer2_out[5715] ^ layer2_out[5716];
    assign layer3_out[1607] = ~layer2_out[342];
    assign layer3_out[1608] = layer2_out[7788];
    assign layer3_out[1609] = ~(layer2_out[5299] | layer2_out[5300]);
    assign layer3_out[1610] = ~layer2_out[7422] | layer2_out[7421];
    assign layer3_out[1611] = layer2_out[1143] & ~layer2_out[1142];
    assign layer3_out[1612] = ~layer2_out[2119];
    assign layer3_out[1613] = layer2_out[6512] & ~layer2_out[6513];
    assign layer3_out[1614] = ~layer2_out[7930];
    assign layer3_out[1615] = layer2_out[7411] ^ layer2_out[7412];
    assign layer3_out[1616] = ~(layer2_out[734] & layer2_out[735]);
    assign layer3_out[1617] = layer2_out[2997] ^ layer2_out[2998];
    assign layer3_out[1618] = ~layer2_out[6207];
    assign layer3_out[1619] = layer2_out[7449] & ~layer2_out[7448];
    assign layer3_out[1620] = layer2_out[6218] & ~layer2_out[6219];
    assign layer3_out[1621] = layer2_out[1459] & ~layer2_out[1458];
    assign layer3_out[1622] = ~layer2_out[7003];
    assign layer3_out[1623] = ~layer2_out[791];
    assign layer3_out[1624] = layer2_out[2939];
    assign layer3_out[1625] = ~layer2_out[6049];
    assign layer3_out[1626] = layer2_out[5396] | layer2_out[5397];
    assign layer3_out[1627] = ~(layer2_out[1461] & layer2_out[1462]);
    assign layer3_out[1628] = ~(layer2_out[4657] & layer2_out[4658]);
    assign layer3_out[1629] = layer2_out[2665];
    assign layer3_out[1630] = 1'b0;
    assign layer3_out[1631] = ~layer2_out[380];
    assign layer3_out[1632] = layer2_out[3403];
    assign layer3_out[1633] = layer2_out[2317];
    assign layer3_out[1634] = layer2_out[6868] ^ layer2_out[6869];
    assign layer3_out[1635] = ~layer2_out[5020] | layer2_out[5021];
    assign layer3_out[1636] = layer2_out[2014];
    assign layer3_out[1637] = ~layer2_out[3223] | layer2_out[3224];
    assign layer3_out[1638] = layer2_out[5337] & layer2_out[5338];
    assign layer3_out[1639] = layer2_out[5062] & layer2_out[5063];
    assign layer3_out[1640] = layer2_out[1478];
    assign layer3_out[1641] = ~layer2_out[3058];
    assign layer3_out[1642] = ~(layer2_out[6526] & layer2_out[6527]);
    assign layer3_out[1643] = ~(layer2_out[307] | layer2_out[308]);
    assign layer3_out[1644] = layer2_out[3743];
    assign layer3_out[1645] = layer2_out[2134];
    assign layer3_out[1646] = ~(layer2_out[6229] ^ layer2_out[6230]);
    assign layer3_out[1647] = ~layer2_out[4592];
    assign layer3_out[1648] = ~layer2_out[6288];
    assign layer3_out[1649] = layer2_out[6154] ^ layer2_out[6155];
    assign layer3_out[1650] = ~layer2_out[840];
    assign layer3_out[1651] = layer2_out[7848] & ~layer2_out[7849];
    assign layer3_out[1652] = layer2_out[4083];
    assign layer3_out[1653] = ~layer2_out[5890];
    assign layer3_out[1654] = ~(layer2_out[4426] & layer2_out[4427]);
    assign layer3_out[1655] = layer2_out[1638] | layer2_out[1639];
    assign layer3_out[1656] = layer2_out[1711];
    assign layer3_out[1657] = layer2_out[973] | layer2_out[974];
    assign layer3_out[1658] = ~layer2_out[203];
    assign layer3_out[1659] = ~(layer2_out[7503] & layer2_out[7504]);
    assign layer3_out[1660] = layer2_out[6480] | layer2_out[6481];
    assign layer3_out[1661] = layer2_out[951] & ~layer2_out[950];
    assign layer3_out[1662] = layer2_out[800] & ~layer2_out[801];
    assign layer3_out[1663] = layer2_out[4932];
    assign layer3_out[1664] = ~layer2_out[608];
    assign layer3_out[1665] = ~(layer2_out[7724] | layer2_out[7725]);
    assign layer3_out[1666] = layer2_out[4005];
    assign layer3_out[1667] = ~layer2_out[7619] | layer2_out[7618];
    assign layer3_out[1668] = ~layer2_out[3095];
    assign layer3_out[1669] = layer2_out[287];
    assign layer3_out[1670] = layer2_out[6254];
    assign layer3_out[1671] = ~layer2_out[1784];
    assign layer3_out[1672] = ~(layer2_out[4364] ^ layer2_out[4365]);
    assign layer3_out[1673] = layer2_out[173] & ~layer2_out[174];
    assign layer3_out[1674] = layer2_out[5280];
    assign layer3_out[1675] = ~(layer2_out[6019] & layer2_out[6020]);
    assign layer3_out[1676] = layer2_out[1929] ^ layer2_out[1930];
    assign layer3_out[1677] = 1'b0;
    assign layer3_out[1678] = ~(layer2_out[2219] & layer2_out[2220]);
    assign layer3_out[1679] = layer2_out[3227];
    assign layer3_out[1680] = ~(layer2_out[5599] ^ layer2_out[5600]);
    assign layer3_out[1681] = layer2_out[1883];
    assign layer3_out[1682] = ~(layer2_out[3900] ^ layer2_out[3901]);
    assign layer3_out[1683] = 1'b1;
    assign layer3_out[1684] = ~layer2_out[1707];
    assign layer3_out[1685] = ~(layer2_out[473] | layer2_out[474]);
    assign layer3_out[1686] = layer2_out[3539] & ~layer2_out[3540];
    assign layer3_out[1687] = layer2_out[7152] & ~layer2_out[7151];
    assign layer3_out[1688] = ~layer2_out[5679];
    assign layer3_out[1689] = layer2_out[672];
    assign layer3_out[1690] = layer2_out[2725] & layer2_out[2726];
    assign layer3_out[1691] = ~layer2_out[3037] | layer2_out[3038];
    assign layer3_out[1692] = ~layer2_out[6992];
    assign layer3_out[1693] = layer2_out[1037] & ~layer2_out[1038];
    assign layer3_out[1694] = layer2_out[1009];
    assign layer3_out[1695] = layer2_out[4304];
    assign layer3_out[1696] = layer2_out[7121];
    assign layer3_out[1697] = ~layer2_out[66];
    assign layer3_out[1698] = layer2_out[361];
    assign layer3_out[1699] = ~(layer2_out[4160] | layer2_out[4161]);
    assign layer3_out[1700] = ~layer2_out[5751] | layer2_out[5750];
    assign layer3_out[1701] = layer2_out[2698] & ~layer2_out[2697];
    assign layer3_out[1702] = layer2_out[7888];
    assign layer3_out[1703] = ~layer2_out[5170];
    assign layer3_out[1704] = layer2_out[4926];
    assign layer3_out[1705] = layer2_out[939] & layer2_out[940];
    assign layer3_out[1706] = ~layer2_out[2826];
    assign layer3_out[1707] = layer2_out[3709] & layer2_out[3710];
    assign layer3_out[1708] = layer2_out[1314] & ~layer2_out[1313];
    assign layer3_out[1709] = layer2_out[2036] & ~layer2_out[2035];
    assign layer3_out[1710] = layer2_out[585] & layer2_out[586];
    assign layer3_out[1711] = ~(layer2_out[5246] & layer2_out[5247]);
    assign layer3_out[1712] = layer2_out[4114];
    assign layer3_out[1713] = ~layer2_out[3015];
    assign layer3_out[1714] = ~(layer2_out[6723] | layer2_out[6724]);
    assign layer3_out[1715] = layer2_out[2353] | layer2_out[2354];
    assign layer3_out[1716] = ~layer2_out[3616] | layer2_out[3615];
    assign layer3_out[1717] = layer2_out[3738] & ~layer2_out[3739];
    assign layer3_out[1718] = ~(layer2_out[7818] | layer2_out[7819]);
    assign layer3_out[1719] = ~(layer2_out[7472] | layer2_out[7473]);
    assign layer3_out[1720] = layer2_out[1770] & ~layer2_out[1769];
    assign layer3_out[1721] = ~layer2_out[1567];
    assign layer3_out[1722] = ~layer2_out[4222];
    assign layer3_out[1723] = layer2_out[1496] | layer2_out[1497];
    assign layer3_out[1724] = ~layer2_out[1841] | layer2_out[1842];
    assign layer3_out[1725] = layer2_out[330] | layer2_out[331];
    assign layer3_out[1726] = ~layer2_out[701];
    assign layer3_out[1727] = layer2_out[2720] & layer2_out[2721];
    assign layer3_out[1728] = layer2_out[3501];
    assign layer3_out[1729] = layer2_out[3312] & layer2_out[3313];
    assign layer3_out[1730] = ~layer2_out[2122] | layer2_out[2123];
    assign layer3_out[1731] = layer2_out[1276];
    assign layer3_out[1732] = ~(layer2_out[3486] ^ layer2_out[3487]);
    assign layer3_out[1733] = layer2_out[845] ^ layer2_out[846];
    assign layer3_out[1734] = ~layer2_out[3561] | layer2_out[3562];
    assign layer3_out[1735] = layer2_out[77] | layer2_out[78];
    assign layer3_out[1736] = layer2_out[7076];
    assign layer3_out[1737] = ~layer2_out[6281];
    assign layer3_out[1738] = layer2_out[3479] & ~layer2_out[3480];
    assign layer3_out[1739] = layer2_out[604] & layer2_out[605];
    assign layer3_out[1740] = ~(layer2_out[5330] & layer2_out[5331]);
    assign layer3_out[1741] = ~layer2_out[6991];
    assign layer3_out[1742] = layer2_out[4788];
    assign layer3_out[1743] = ~layer2_out[7632] | layer2_out[7631];
    assign layer3_out[1744] = layer2_out[1003] & ~layer2_out[1002];
    assign layer3_out[1745] = layer2_out[2097] & ~layer2_out[2096];
    assign layer3_out[1746] = layer2_out[5313];
    assign layer3_out[1747] = ~layer2_out[4006];
    assign layer3_out[1748] = layer2_out[2474] & layer2_out[2475];
    assign layer3_out[1749] = ~(layer2_out[5655] ^ layer2_out[5656]);
    assign layer3_out[1750] = ~layer2_out[2845];
    assign layer3_out[1751] = ~layer2_out[4178];
    assign layer3_out[1752] = ~layer2_out[6444] | layer2_out[6443];
    assign layer3_out[1753] = ~(layer2_out[2382] | layer2_out[2383]);
    assign layer3_out[1754] = ~(layer2_out[2626] ^ layer2_out[2627]);
    assign layer3_out[1755] = layer2_out[563] | layer2_out[564];
    assign layer3_out[1756] = layer2_out[6969] & ~layer2_out[6970];
    assign layer3_out[1757] = layer2_out[3990];
    assign layer3_out[1758] = layer2_out[4463];
    assign layer3_out[1759] = layer2_out[7830] ^ layer2_out[7831];
    assign layer3_out[1760] = ~layer2_out[2248];
    assign layer3_out[1761] = layer2_out[3169] & ~layer2_out[3170];
    assign layer3_out[1762] = ~(layer2_out[1702] ^ layer2_out[1703]);
    assign layer3_out[1763] = layer2_out[3691];
    assign layer3_out[1764] = ~layer2_out[7160] | layer2_out[7159];
    assign layer3_out[1765] = layer2_out[2509] & layer2_out[2510];
    assign layer3_out[1766] = ~layer2_out[3544] | layer2_out[3543];
    assign layer3_out[1767] = ~(layer2_out[7223] | layer2_out[7224]);
    assign layer3_out[1768] = 1'b0;
    assign layer3_out[1769] = layer2_out[1009];
    assign layer3_out[1770] = layer2_out[3586];
    assign layer3_out[1771] = layer2_out[5133] & ~layer2_out[5132];
    assign layer3_out[1772] = ~(layer2_out[3578] | layer2_out[3579]);
    assign layer3_out[1773] = ~layer2_out[5896];
    assign layer3_out[1774] = ~(layer2_out[5281] & layer2_out[5282]);
    assign layer3_out[1775] = layer2_out[6266];
    assign layer3_out[1776] = layer2_out[4636];
    assign layer3_out[1777] = 1'b0;
    assign layer3_out[1778] = layer2_out[7678] & ~layer2_out[7679];
    assign layer3_out[1779] = layer2_out[3041];
    assign layer3_out[1780] = ~layer2_out[3325];
    assign layer3_out[1781] = ~layer2_out[4714];
    assign layer3_out[1782] = layer2_out[2031];
    assign layer3_out[1783] = ~layer2_out[7329];
    assign layer3_out[1784] = layer2_out[1171] ^ layer2_out[1172];
    assign layer3_out[1785] = layer2_out[1092] & ~layer2_out[1093];
    assign layer3_out[1786] = layer2_out[920] | layer2_out[921];
    assign layer3_out[1787] = ~(layer2_out[4450] ^ layer2_out[4451]);
    assign layer3_out[1788] = ~layer2_out[1129];
    assign layer3_out[1789] = ~layer2_out[848];
    assign layer3_out[1790] = ~layer2_out[5594] | layer2_out[5595];
    assign layer3_out[1791] = layer2_out[7705];
    assign layer3_out[1792] = ~(layer2_out[7696] & layer2_out[7697]);
    assign layer3_out[1793] = ~(layer2_out[2414] & layer2_out[2415]);
    assign layer3_out[1794] = ~(layer2_out[2913] ^ layer2_out[2914]);
    assign layer3_out[1795] = layer2_out[1927];
    assign layer3_out[1796] = ~layer2_out[5913];
    assign layer3_out[1797] = ~(layer2_out[2954] | layer2_out[2955]);
    assign layer3_out[1798] = layer2_out[5417] ^ layer2_out[5418];
    assign layer3_out[1799] = layer2_out[7063];
    assign layer3_out[1800] = layer2_out[7764];
    assign layer3_out[1801] = ~layer2_out[7734] | layer2_out[7733];
    assign layer3_out[1802] = ~layer2_out[4231];
    assign layer3_out[1803] = layer2_out[5059];
    assign layer3_out[1804] = layer2_out[1762];
    assign layer3_out[1805] = ~layer2_out[2935];
    assign layer3_out[1806] = layer2_out[6259] | layer2_out[6260];
    assign layer3_out[1807] = layer2_out[7372] & ~layer2_out[7373];
    assign layer3_out[1808] = ~layer2_out[69];
    assign layer3_out[1809] = layer2_out[7728] | layer2_out[7729];
    assign layer3_out[1810] = ~(layer2_out[1600] ^ layer2_out[1601]);
    assign layer3_out[1811] = layer2_out[1910] ^ layer2_out[1911];
    assign layer3_out[1812] = layer2_out[6059];
    assign layer3_out[1813] = layer2_out[1855] & layer2_out[1856];
    assign layer3_out[1814] = ~(layer2_out[1249] & layer2_out[1250]);
    assign layer3_out[1815] = layer2_out[7756];
    assign layer3_out[1816] = layer2_out[2492];
    assign layer3_out[1817] = layer2_out[4843] ^ layer2_out[4844];
    assign layer3_out[1818] = ~layer2_out[229] | layer2_out[228];
    assign layer3_out[1819] = ~(layer2_out[394] & layer2_out[395]);
    assign layer3_out[1820] = ~layer2_out[7643];
    assign layer3_out[1821] = layer2_out[5497] & ~layer2_out[5496];
    assign layer3_out[1822] = ~layer2_out[3406] | layer2_out[3405];
    assign layer3_out[1823] = ~layer2_out[4358];
    assign layer3_out[1824] = ~layer2_out[7173];
    assign layer3_out[1825] = layer2_out[3719];
    assign layer3_out[1826] = ~(layer2_out[6673] ^ layer2_out[6674]);
    assign layer3_out[1827] = ~layer2_out[3277];
    assign layer3_out[1828] = layer2_out[2493];
    assign layer3_out[1829] = ~layer2_out[1942];
    assign layer3_out[1830] = ~layer2_out[982];
    assign layer3_out[1831] = 1'b1;
    assign layer3_out[1832] = ~layer2_out[3013] | layer2_out[3014];
    assign layer3_out[1833] = ~(layer2_out[7949] | layer2_out[7950]);
    assign layer3_out[1834] = layer2_out[5096];
    assign layer3_out[1835] = layer2_out[2809] & ~layer2_out[2810];
    assign layer3_out[1836] = layer2_out[5052] & layer2_out[5053];
    assign layer3_out[1837] = layer2_out[6684];
    assign layer3_out[1838] = ~layer2_out[830] | layer2_out[831];
    assign layer3_out[1839] = layer2_out[7479] & ~layer2_out[7478];
    assign layer3_out[1840] = ~layer2_out[2829];
    assign layer3_out[1841] = ~layer2_out[1661];
    assign layer3_out[1842] = ~(layer2_out[1866] & layer2_out[1867]);
    assign layer3_out[1843] = layer2_out[2315];
    assign layer3_out[1844] = ~(layer2_out[3196] ^ layer2_out[3197]);
    assign layer3_out[1845] = layer2_out[250];
    assign layer3_out[1846] = layer2_out[7820] | layer2_out[7821];
    assign layer3_out[1847] = layer2_out[226] ^ layer2_out[227];
    assign layer3_out[1848] = layer2_out[6753];
    assign layer3_out[1849] = layer2_out[1642] & layer2_out[1643];
    assign layer3_out[1850] = ~layer2_out[1262];
    assign layer3_out[1851] = layer2_out[467] & ~layer2_out[466];
    assign layer3_out[1852] = layer2_out[2653];
    assign layer3_out[1853] = ~layer2_out[1676];
    assign layer3_out[1854] = layer2_out[5641] & ~layer2_out[5642];
    assign layer3_out[1855] = ~layer2_out[7432];
    assign layer3_out[1856] = layer2_out[5170];
    assign layer3_out[1857] = 1'b1;
    assign layer3_out[1858] = ~layer2_out[1629];
    assign layer3_out[1859] = ~layer2_out[7435];
    assign layer3_out[1860] = layer2_out[2319] | layer2_out[2320];
    assign layer3_out[1861] = ~layer2_out[2465];
    assign layer3_out[1862] = layer2_out[4336] ^ layer2_out[4337];
    assign layer3_out[1863] = layer2_out[7736];
    assign layer3_out[1864] = ~(layer2_out[7597] ^ layer2_out[7598]);
    assign layer3_out[1865] = ~(layer2_out[2307] & layer2_out[2308]);
    assign layer3_out[1866] = layer2_out[6567];
    assign layer3_out[1867] = layer2_out[2407];
    assign layer3_out[1868] = ~layer2_out[7727] | layer2_out[7726];
    assign layer3_out[1869] = layer2_out[6511] & ~layer2_out[6512];
    assign layer3_out[1870] = 1'b1;
    assign layer3_out[1871] = ~layer2_out[3649] | layer2_out[3650];
    assign layer3_out[1872] = layer2_out[4716];
    assign layer3_out[1873] = layer2_out[6556];
    assign layer3_out[1874] = layer2_out[3979] & ~layer2_out[3980];
    assign layer3_out[1875] = ~layer2_out[1720] | layer2_out[1721];
    assign layer3_out[1876] = layer2_out[6956] & ~layer2_out[6957];
    assign layer3_out[1877] = ~layer2_out[6677] | layer2_out[6678];
    assign layer3_out[1878] = layer2_out[224] & layer2_out[225];
    assign layer3_out[1879] = layer2_out[4696] & layer2_out[4697];
    assign layer3_out[1880] = ~(layer2_out[7444] ^ layer2_out[7445]);
    assign layer3_out[1881] = ~layer2_out[4945] | layer2_out[4944];
    assign layer3_out[1882] = layer2_out[22];
    assign layer3_out[1883] = layer2_out[5411];
    assign layer3_out[1884] = ~layer2_out[2111];
    assign layer3_out[1885] = ~layer2_out[4439] | layer2_out[4438];
    assign layer3_out[1886] = ~layer2_out[6736];
    assign layer3_out[1887] = layer2_out[4789];
    assign layer3_out[1888] = layer2_out[0];
    assign layer3_out[1889] = layer2_out[5414];
    assign layer3_out[1890] = ~layer2_out[1230];
    assign layer3_out[1891] = layer2_out[4792];
    assign layer3_out[1892] = layer2_out[1825];
    assign layer3_out[1893] = layer2_out[108];
    assign layer3_out[1894] = ~(layer2_out[3404] | layer2_out[3405]);
    assign layer3_out[1895] = layer2_out[4147] & ~layer2_out[4146];
    assign layer3_out[1896] = layer2_out[5266];
    assign layer3_out[1897] = layer2_out[8] & ~layer2_out[9];
    assign layer3_out[1898] = ~layer2_out[7372];
    assign layer3_out[1899] = layer2_out[3239] | layer2_out[3240];
    assign layer3_out[1900] = layer2_out[1950] & layer2_out[1951];
    assign layer3_out[1901] = ~layer2_out[7538];
    assign layer3_out[1902] = ~(layer2_out[7751] | layer2_out[7752]);
    assign layer3_out[1903] = 1'b1;
    assign layer3_out[1904] = layer2_out[6946] ^ layer2_out[6947];
    assign layer3_out[1905] = layer2_out[3967];
    assign layer3_out[1906] = ~(layer2_out[1211] | layer2_out[1212]);
    assign layer3_out[1907] = ~layer2_out[5196];
    assign layer3_out[1908] = ~(layer2_out[782] ^ layer2_out[783]);
    assign layer3_out[1909] = layer2_out[5907];
    assign layer3_out[1910] = ~layer2_out[7772];
    assign layer3_out[1911] = layer2_out[1700] ^ layer2_out[1701];
    assign layer3_out[1912] = ~layer2_out[1663];
    assign layer3_out[1913] = layer2_out[5171] ^ layer2_out[5172];
    assign layer3_out[1914] = ~layer2_out[917] | layer2_out[918];
    assign layer3_out[1915] = ~(layer2_out[2499] ^ layer2_out[2500]);
    assign layer3_out[1916] = ~(layer2_out[2212] ^ layer2_out[2213]);
    assign layer3_out[1917] = ~(layer2_out[3080] | layer2_out[3081]);
    assign layer3_out[1918] = layer2_out[1410];
    assign layer3_out[1919] = layer2_out[2745];
    assign layer3_out[1920] = layer2_out[816] & ~layer2_out[815];
    assign layer3_out[1921] = layer2_out[6158] | layer2_out[6159];
    assign layer3_out[1922] = ~layer2_out[2791];
    assign layer3_out[1923] = ~(layer2_out[921] | layer2_out[922]);
    assign layer3_out[1924] = ~layer2_out[4769] | layer2_out[4770];
    assign layer3_out[1925] = layer2_out[3313] & layer2_out[3314];
    assign layer3_out[1926] = layer2_out[7220] ^ layer2_out[7221];
    assign layer3_out[1927] = layer2_out[4046] & ~layer2_out[4047];
    assign layer3_out[1928] = ~(layer2_out[3451] ^ layer2_out[3452]);
    assign layer3_out[1929] = ~layer2_out[3006];
    assign layer3_out[1930] = ~layer2_out[2896] | layer2_out[2897];
    assign layer3_out[1931] = 1'b1;
    assign layer3_out[1932] = 1'b0;
    assign layer3_out[1933] = ~layer2_out[3229] | layer2_out[3228];
    assign layer3_out[1934] = ~layer2_out[3409];
    assign layer3_out[1935] = layer2_out[1179];
    assign layer3_out[1936] = layer2_out[1493] ^ layer2_out[1494];
    assign layer3_out[1937] = 1'b0;
    assign layer3_out[1938] = ~(layer2_out[5355] & layer2_out[5356]);
    assign layer3_out[1939] = layer2_out[2688];
    assign layer3_out[1940] = ~layer2_out[6191] | layer2_out[6192];
    assign layer3_out[1941] = ~layer2_out[6748];
    assign layer3_out[1942] = ~layer2_out[5092];
    assign layer3_out[1943] = ~(layer2_out[7253] ^ layer2_out[7254]);
    assign layer3_out[1944] = layer2_out[72] & ~layer2_out[71];
    assign layer3_out[1945] = layer2_out[2765] & layer2_out[2766];
    assign layer3_out[1946] = ~layer2_out[7711] | layer2_out[7710];
    assign layer3_out[1947] = layer2_out[7520];
    assign layer3_out[1948] = layer2_out[3164] & layer2_out[3165];
    assign layer3_out[1949] = ~(layer2_out[2477] | layer2_out[2478]);
    assign layer3_out[1950] = layer2_out[7897] & layer2_out[7898];
    assign layer3_out[1951] = ~(layer2_out[7039] & layer2_out[7040]);
    assign layer3_out[1952] = ~layer2_out[579];
    assign layer3_out[1953] = layer2_out[7276] & layer2_out[7277];
    assign layer3_out[1954] = layer2_out[2941];
    assign layer3_out[1955] = ~layer2_out[3059] | layer2_out[3058];
    assign layer3_out[1956] = layer2_out[4543];
    assign layer3_out[1957] = layer2_out[3749] ^ layer2_out[3750];
    assign layer3_out[1958] = layer2_out[6493];
    assign layer3_out[1959] = ~layer2_out[695];
    assign layer3_out[1960] = layer2_out[7155] & ~layer2_out[7154];
    assign layer3_out[1961] = ~layer2_out[6725];
    assign layer3_out[1962] = layer2_out[563] & ~layer2_out[562];
    assign layer3_out[1963] = layer2_out[6234];
    assign layer3_out[1964] = layer2_out[1188] & layer2_out[1189];
    assign layer3_out[1965] = layer2_out[1619] | layer2_out[1620];
    assign layer3_out[1966] = layer2_out[4557];
    assign layer3_out[1967] = ~(layer2_out[7927] ^ layer2_out[7928]);
    assign layer3_out[1968] = layer2_out[6973] | layer2_out[6974];
    assign layer3_out[1969] = layer2_out[5394] ^ layer2_out[5395];
    assign layer3_out[1970] = layer2_out[2376];
    assign layer3_out[1971] = ~layer2_out[3439] | layer2_out[3440];
    assign layer3_out[1972] = layer2_out[5475] | layer2_out[5476];
    assign layer3_out[1973] = ~layer2_out[3435];
    assign layer3_out[1974] = ~(layer2_out[6404] | layer2_out[6405]);
    assign layer3_out[1975] = layer2_out[1044] & ~layer2_out[1043];
    assign layer3_out[1976] = ~layer2_out[5472];
    assign layer3_out[1977] = ~(layer2_out[1558] | layer2_out[1559]);
    assign layer3_out[1978] = layer2_out[3448];
    assign layer3_out[1979] = layer2_out[5136] & layer2_out[5137];
    assign layer3_out[1980] = ~layer2_out[4331];
    assign layer3_out[1981] = layer2_out[6466];
    assign layer3_out[1982] = ~layer2_out[7532];
    assign layer3_out[1983] = layer2_out[3752];
    assign layer3_out[1984] = layer2_out[3515];
    assign layer3_out[1985] = layer2_out[5031];
    assign layer3_out[1986] = ~layer2_out[461] | layer2_out[462];
    assign layer3_out[1987] = layer2_out[2321];
    assign layer3_out[1988] = ~(layer2_out[1678] | layer2_out[1679]);
    assign layer3_out[1989] = ~layer2_out[4977] | layer2_out[4978];
    assign layer3_out[1990] = layer2_out[4287] | layer2_out[4288];
    assign layer3_out[1991] = layer2_out[890];
    assign layer3_out[1992] = layer2_out[4498];
    assign layer3_out[1993] = layer2_out[3355];
    assign layer3_out[1994] = ~(layer2_out[1443] ^ layer2_out[1444]);
    assign layer3_out[1995] = ~layer2_out[1811];
    assign layer3_out[1996] = ~layer2_out[2402];
    assign layer3_out[1997] = layer2_out[3265] ^ layer2_out[3266];
    assign layer3_out[1998] = ~(layer2_out[6670] & layer2_out[6671]);
    assign layer3_out[1999] = layer2_out[6788];
    assign layer3_out[2000] = layer2_out[4830] & layer2_out[4831];
    assign layer3_out[2001] = layer2_out[5208] & layer2_out[5209];
    assign layer3_out[2002] = layer2_out[3470] & ~layer2_out[3469];
    assign layer3_out[2003] = ~layer2_out[2860] | layer2_out[2861];
    assign layer3_out[2004] = layer2_out[1413];
    assign layer3_out[2005] = ~(layer2_out[3822] & layer2_out[3823]);
    assign layer3_out[2006] = ~layer2_out[2621];
    assign layer3_out[2007] = layer2_out[376] | layer2_out[377];
    assign layer3_out[2008] = layer2_out[2026] & ~layer2_out[2025];
    assign layer3_out[2009] = ~layer2_out[6199];
    assign layer3_out[2010] = layer2_out[5107] & layer2_out[5108];
    assign layer3_out[2011] = ~layer2_out[6686] | layer2_out[6687];
    assign layer3_out[2012] = ~layer2_out[1946] | layer2_out[1947];
    assign layer3_out[2013] = layer2_out[1091] & ~layer2_out[1090];
    assign layer3_out[2014] = 1'b1;
    assign layer3_out[2015] = ~layer2_out[3271] | layer2_out[3270];
    assign layer3_out[2016] = layer2_out[673] | layer2_out[674];
    assign layer3_out[2017] = ~(layer2_out[2832] | layer2_out[2833]);
    assign layer3_out[2018] = layer2_out[5290] ^ layer2_out[5291];
    assign layer3_out[2019] = ~layer2_out[5872];
    assign layer3_out[2020] = layer2_out[3130] & ~layer2_out[3131];
    assign layer3_out[2021] = layer2_out[4275];
    assign layer3_out[2022] = ~layer2_out[3413];
    assign layer3_out[2023] = layer2_out[1126] & layer2_out[1127];
    assign layer3_out[2024] = layer2_out[1498];
    assign layer3_out[2025] = ~(layer2_out[993] ^ layer2_out[994]);
    assign layer3_out[2026] = layer2_out[910];
    assign layer3_out[2027] = ~layer2_out[606];
    assign layer3_out[2028] = layer2_out[3166];
    assign layer3_out[2029] = ~layer2_out[7964];
    assign layer3_out[2030] = layer2_out[7600] & ~layer2_out[7601];
    assign layer3_out[2031] = layer2_out[5216];
    assign layer3_out[2032] = ~layer2_out[4579];
    assign layer3_out[2033] = ~(layer2_out[3700] & layer2_out[3701]);
    assign layer3_out[2034] = ~(layer2_out[6043] & layer2_out[6044]);
    assign layer3_out[2035] = layer2_out[3678] | layer2_out[3679];
    assign layer3_out[2036] = ~(layer2_out[3338] & layer2_out[3339]);
    assign layer3_out[2037] = ~layer2_out[483];
    assign layer3_out[2038] = ~layer2_out[2257] | layer2_out[2256];
    assign layer3_out[2039] = layer2_out[1299];
    assign layer3_out[2040] = layer2_out[6124] & ~layer2_out[6125];
    assign layer3_out[2041] = ~layer2_out[3999] | layer2_out[4000];
    assign layer3_out[2042] = ~layer2_out[1737];
    assign layer3_out[2043] = layer2_out[6279] | layer2_out[6280];
    assign layer3_out[2044] = ~layer2_out[7514] | layer2_out[7513];
    assign layer3_out[2045] = ~layer2_out[4088] | layer2_out[4089];
    assign layer3_out[2046] = ~layer2_out[3402] | layer2_out[3401];
    assign layer3_out[2047] = ~(layer2_out[4852] & layer2_out[4853]);
    assign layer3_out[2048] = layer2_out[433] & ~layer2_out[434];
    assign layer3_out[2049] = ~layer2_out[3252] | layer2_out[3253];
    assign layer3_out[2050] = ~layer2_out[5355];
    assign layer3_out[2051] = layer2_out[7418] & ~layer2_out[7417];
    assign layer3_out[2052] = layer2_out[2324] | layer2_out[2325];
    assign layer3_out[2053] = layer2_out[4633] ^ layer2_out[4634];
    assign layer3_out[2054] = layer2_out[646];
    assign layer3_out[2055] = ~(layer2_out[1251] & layer2_out[1252]);
    assign layer3_out[2056] = ~(layer2_out[738] ^ layer2_out[739]);
    assign layer3_out[2057] = ~layer2_out[2293];
    assign layer3_out[2058] = layer2_out[2375] ^ layer2_out[2376];
    assign layer3_out[2059] = ~layer2_out[7116] | layer2_out[7115];
    assign layer3_out[2060] = ~layer2_out[2723];
    assign layer3_out[2061] = ~layer2_out[3077];
    assign layer3_out[2062] = ~(layer2_out[6114] & layer2_out[6115]);
    assign layer3_out[2063] = layer2_out[5502];
    assign layer3_out[2064] = layer2_out[3803] & ~layer2_out[3802];
    assign layer3_out[2065] = layer2_out[365] & layer2_out[366];
    assign layer3_out[2066] = layer2_out[39];
    assign layer3_out[2067] = layer2_out[4091];
    assign layer3_out[2068] = layer2_out[7253];
    assign layer3_out[2069] = layer2_out[3774] & ~layer2_out[3773];
    assign layer3_out[2070] = ~(layer2_out[650] & layer2_out[651]);
    assign layer3_out[2071] = layer2_out[539] | layer2_out[540];
    assign layer3_out[2072] = layer2_out[2457] & ~layer2_out[2458];
    assign layer3_out[2073] = ~(layer2_out[3878] | layer2_out[3879]);
    assign layer3_out[2074] = layer2_out[3126] ^ layer2_out[3127];
    assign layer3_out[2075] = ~(layer2_out[1186] & layer2_out[1187]);
    assign layer3_out[2076] = layer2_out[1081];
    assign layer3_out[2077] = ~(layer2_out[7464] | layer2_out[7465]);
    assign layer3_out[2078] = ~layer2_out[258];
    assign layer3_out[2079] = layer2_out[7535] | layer2_out[7536];
    assign layer3_out[2080] = layer2_out[2006];
    assign layer3_out[2081] = ~(layer2_out[4721] | layer2_out[4722]);
    assign layer3_out[2082] = layer2_out[548] | layer2_out[549];
    assign layer3_out[2083] = layer2_out[2842];
    assign layer3_out[2084] = layer2_out[1952];
    assign layer3_out[2085] = layer2_out[234] & ~layer2_out[235];
    assign layer3_out[2086] = ~layer2_out[4679] | layer2_out[4680];
    assign layer3_out[2087] = ~(layer2_out[195] ^ layer2_out[196]);
    assign layer3_out[2088] = ~(layer2_out[6803] & layer2_out[6804]);
    assign layer3_out[2089] = layer2_out[2803] & ~layer2_out[2802];
    assign layer3_out[2090] = layer2_out[662];
    assign layer3_out[2091] = ~layer2_out[3988];
    assign layer3_out[2092] = ~layer2_out[6703];
    assign layer3_out[2093] = layer2_out[2410] & layer2_out[2411];
    assign layer3_out[2094] = ~(layer2_out[4964] & layer2_out[4965]);
    assign layer3_out[2095] = layer2_out[2066] & ~layer2_out[2067];
    assign layer3_out[2096] = layer2_out[1402] | layer2_out[1403];
    assign layer3_out[2097] = ~layer2_out[5846];
    assign layer3_out[2098] = layer2_out[4581];
    assign layer3_out[2099] = ~layer2_out[7293] | layer2_out[7292];
    assign layer3_out[2100] = ~layer2_out[2147];
    assign layer3_out[2101] = layer2_out[6996] ^ layer2_out[6997];
    assign layer3_out[2102] = ~(layer2_out[4347] ^ layer2_out[4348]);
    assign layer3_out[2103] = 1'b1;
    assign layer3_out[2104] = layer2_out[5796] | layer2_out[5797];
    assign layer3_out[2105] = ~(layer2_out[4838] & layer2_out[4839]);
    assign layer3_out[2106] = ~(layer2_out[3081] ^ layer2_out[3082]);
    assign layer3_out[2107] = ~(layer2_out[397] & layer2_out[398]);
    assign layer3_out[2108] = layer2_out[825] & ~layer2_out[826];
    assign layer3_out[2109] = ~layer2_out[6321] | layer2_out[6322];
    assign layer3_out[2110] = ~layer2_out[1726];
    assign layer3_out[2111] = ~layer2_out[5104];
    assign layer3_out[2112] = 1'b1;
    assign layer3_out[2113] = layer2_out[7516];
    assign layer3_out[2114] = ~layer2_out[7783];
    assign layer3_out[2115] = layer2_out[3383] | layer2_out[3384];
    assign layer3_out[2116] = ~(layer2_out[3046] & layer2_out[3047]);
    assign layer3_out[2117] = layer2_out[5263] & ~layer2_out[5264];
    assign layer3_out[2118] = ~(layer2_out[532] | layer2_out[533]);
    assign layer3_out[2119] = ~layer2_out[4580];
    assign layer3_out[2120] = ~layer2_out[1482];
    assign layer3_out[2121] = ~layer2_out[6834] | layer2_out[6833];
    assign layer3_out[2122] = layer2_out[6590] ^ layer2_out[6591];
    assign layer3_out[2123] = ~layer2_out[7041];
    assign layer3_out[2124] = layer2_out[5986] & ~layer2_out[5987];
    assign layer3_out[2125] = 1'b1;
    assign layer3_out[2126] = layer2_out[1884];
    assign layer3_out[2127] = ~layer2_out[7886] | layer2_out[7887];
    assign layer3_out[2128] = layer2_out[7216] ^ layer2_out[7217];
    assign layer3_out[2129] = layer2_out[7970];
    assign layer3_out[2130] = layer2_out[2814] & ~layer2_out[2813];
    assign layer3_out[2131] = ~layer2_out[1591];
    assign layer3_out[2132] = ~layer2_out[6550];
    assign layer3_out[2133] = 1'b1;
    assign layer3_out[2134] = layer2_out[1484] ^ layer2_out[1485];
    assign layer3_out[2135] = ~layer2_out[4074];
    assign layer3_out[2136] = ~layer2_out[570] | layer2_out[569];
    assign layer3_out[2137] = ~layer2_out[3374];
    assign layer3_out[2138] = layer2_out[110] & ~layer2_out[111];
    assign layer3_out[2139] = ~layer2_out[6274];
    assign layer3_out[2140] = ~(layer2_out[5619] & layer2_out[5620]);
    assign layer3_out[2141] = ~layer2_out[3258];
    assign layer3_out[2142] = layer2_out[4434] ^ layer2_out[4435];
    assign layer3_out[2143] = ~layer2_out[1281] | layer2_out[1282];
    assign layer3_out[2144] = ~layer2_out[7083] | layer2_out[7082];
    assign layer3_out[2145] = layer2_out[5406] & ~layer2_out[5407];
    assign layer3_out[2146] = ~layer2_out[1580] | layer2_out[1579];
    assign layer3_out[2147] = layer2_out[5408] & ~layer2_out[5407];
    assign layer3_out[2148] = ~layer2_out[1381];
    assign layer3_out[2149] = layer2_out[1125] & ~layer2_out[1126];
    assign layer3_out[2150] = layer2_out[7883] ^ layer2_out[7884];
    assign layer3_out[2151] = ~layer2_out[355] | layer2_out[356];
    assign layer3_out[2152] = ~layer2_out[2811];
    assign layer3_out[2153] = ~layer2_out[4032] | layer2_out[4031];
    assign layer3_out[2154] = ~(layer2_out[2769] | layer2_out[2770]);
    assign layer3_out[2155] = layer2_out[3098] | layer2_out[3099];
    assign layer3_out[2156] = layer2_out[6977];
    assign layer3_out[2157] = 1'b1;
    assign layer3_out[2158] = layer2_out[836];
    assign layer3_out[2159] = layer2_out[5455] & ~layer2_out[5456];
    assign layer3_out[2160] = ~(layer2_out[4212] ^ layer2_out[4213]);
    assign layer3_out[2161] = ~(layer2_out[7849] | layer2_out[7850]);
    assign layer3_out[2162] = layer2_out[7808];
    assign layer3_out[2163] = layer2_out[613];
    assign layer3_out[2164] = ~(layer2_out[219] ^ layer2_out[220]);
    assign layer3_out[2165] = layer2_out[3017];
    assign layer3_out[2166] = layer2_out[221];
    assign layer3_out[2167] = layer2_out[7884];
    assign layer3_out[2168] = layer2_out[6150] & ~layer2_out[6149];
    assign layer3_out[2169] = ~(layer2_out[676] ^ layer2_out[677]);
    assign layer3_out[2170] = layer2_out[1451] & ~layer2_out[1452];
    assign layer3_out[2171] = ~(layer2_out[6497] ^ layer2_out[6498]);
    assign layer3_out[2172] = layer2_out[7807];
    assign layer3_out[2173] = layer2_out[3716] & ~layer2_out[3715];
    assign layer3_out[2174] = layer2_out[7176] | layer2_out[7177];
    assign layer3_out[2175] = ~layer2_out[1155];
    assign layer3_out[2176] = layer2_out[4588] | layer2_out[4589];
    assign layer3_out[2177] = layer2_out[2171] & ~layer2_out[2172];
    assign layer3_out[2178] = layer2_out[3780] & ~layer2_out[3779];
    assign layer3_out[2179] = layer2_out[3391] & ~layer2_out[3392];
    assign layer3_out[2180] = ~(layer2_out[4222] ^ layer2_out[4223]);
    assign layer3_out[2181] = layer2_out[657] & layer2_out[658];
    assign layer3_out[2182] = ~(layer2_out[5506] | layer2_out[5507]);
    assign layer3_out[2183] = layer2_out[1609];
    assign layer3_out[2184] = layer2_out[657];
    assign layer3_out[2185] = ~(layer2_out[3721] ^ layer2_out[3722]);
    assign layer3_out[2186] = ~(layer2_out[149] | layer2_out[150]);
    assign layer3_out[2187] = layer2_out[3415];
    assign layer3_out[2188] = ~(layer2_out[45] ^ layer2_out[46]);
    assign layer3_out[2189] = ~layer2_out[735] | layer2_out[736];
    assign layer3_out[2190] = ~layer2_out[799] | layer2_out[800];
    assign layer3_out[2191] = ~layer2_out[1488];
    assign layer3_out[2192] = layer2_out[5939] | layer2_out[5940];
    assign layer3_out[2193] = layer2_out[1980] & ~layer2_out[1979];
    assign layer3_out[2194] = layer2_out[3411] | layer2_out[3412];
    assign layer3_out[2195] = ~(layer2_out[718] | layer2_out[719]);
    assign layer3_out[2196] = ~(layer2_out[201] | layer2_out[202]);
    assign layer3_out[2197] = layer2_out[3251];
    assign layer3_out[2198] = ~layer2_out[6578];
    assign layer3_out[2199] = layer2_out[2827] | layer2_out[2828];
    assign layer3_out[2200] = layer2_out[4691];
    assign layer3_out[2201] = ~layer2_out[3793] | layer2_out[3794];
    assign layer3_out[2202] = layer2_out[2821] & ~layer2_out[2820];
    assign layer3_out[2203] = layer2_out[5464] & layer2_out[5465];
    assign layer3_out[2204] = layer2_out[22] & layer2_out[23];
    assign layer3_out[2205] = ~(layer2_out[3762] ^ layer2_out[3763]);
    assign layer3_out[2206] = ~layer2_out[5936];
    assign layer3_out[2207] = ~layer2_out[3935] | layer2_out[3934];
    assign layer3_out[2208] = layer2_out[4667];
    assign layer3_out[2209] = layer2_out[5094];
    assign layer3_out[2210] = ~layer2_out[3145];
    assign layer3_out[2211] = ~(layer2_out[7653] ^ layer2_out[7654]);
    assign layer3_out[2212] = ~layer2_out[963] | layer2_out[962];
    assign layer3_out[2213] = ~(layer2_out[2757] ^ layer2_out[2758]);
    assign layer3_out[2214] = layer2_out[1429] & layer2_out[1430];
    assign layer3_out[2215] = layer2_out[6058];
    assign layer3_out[2216] = layer2_out[3071];
    assign layer3_out[2217] = layer2_out[4467];
    assign layer3_out[2218] = ~(layer2_out[7551] & layer2_out[7552]);
    assign layer3_out[2219] = ~layer2_out[5651];
    assign layer3_out[2220] = ~layer2_out[6875];
    assign layer3_out[2221] = ~layer2_out[3839];
    assign layer3_out[2222] = ~(layer2_out[5794] & layer2_out[5795]);
    assign layer3_out[2223] = ~layer2_out[7708];
    assign layer3_out[2224] = ~layer2_out[2359] | layer2_out[2358];
    assign layer3_out[2225] = layer2_out[3481];
    assign layer3_out[2226] = ~(layer2_out[4532] & layer2_out[4533]);
    assign layer3_out[2227] = ~layer2_out[6291];
    assign layer3_out[2228] = layer2_out[2383] & ~layer2_out[2384];
    assign layer3_out[2229] = ~(layer2_out[4495] & layer2_out[4496]);
    assign layer3_out[2230] = layer2_out[6708] & ~layer2_out[6707];
    assign layer3_out[2231] = layer2_out[6495] & layer2_out[6496];
    assign layer3_out[2232] = layer2_out[1426] & ~layer2_out[1427];
    assign layer3_out[2233] = layer2_out[2756];
    assign layer3_out[2234] = ~layer2_out[1546];
    assign layer3_out[2235] = layer2_out[7892] ^ layer2_out[7893];
    assign layer3_out[2236] = ~layer2_out[3658];
    assign layer3_out[2237] = layer2_out[5382] & ~layer2_out[5381];
    assign layer3_out[2238] = layer2_out[1229];
    assign layer3_out[2239] = layer2_out[4621];
    assign layer3_out[2240] = ~(layer2_out[5659] & layer2_out[5660]);
    assign layer3_out[2241] = layer2_out[649] & ~layer2_out[648];
    assign layer3_out[2242] = layer2_out[5033];
    assign layer3_out[2243] = ~(layer2_out[938] ^ layer2_out[939]);
    assign layer3_out[2244] = ~(layer2_out[7760] & layer2_out[7761]);
    assign layer3_out[2245] = ~layer2_out[2996] | layer2_out[2995];
    assign layer3_out[2246] = layer2_out[5347];
    assign layer3_out[2247] = ~layer2_out[7585];
    assign layer3_out[2248] = layer2_out[6420] & ~layer2_out[6419];
    assign layer3_out[2249] = layer2_out[1369] | layer2_out[1370];
    assign layer3_out[2250] = ~layer2_out[2925] | layer2_out[2926];
    assign layer3_out[2251] = ~layer2_out[7068];
    assign layer3_out[2252] = layer2_out[4943] | layer2_out[4944];
    assign layer3_out[2253] = ~(layer2_out[3189] | layer2_out[3190]);
    assign layer3_out[2254] = layer2_out[1474] & layer2_out[1475];
    assign layer3_out[2255] = layer2_out[786] & ~layer2_out[785];
    assign layer3_out[2256] = ~layer2_out[4591] | layer2_out[4592];
    assign layer3_out[2257] = ~(layer2_out[6014] ^ layer2_out[6015]);
    assign layer3_out[2258] = layer2_out[6070];
    assign layer3_out[2259] = ~layer2_out[6876] | layer2_out[6877];
    assign layer3_out[2260] = layer2_out[7437];
    assign layer3_out[2261] = ~layer2_out[4931];
    assign layer3_out[2262] = layer2_out[2104] | layer2_out[2105];
    assign layer3_out[2263] = ~layer2_out[2370] | layer2_out[2369];
    assign layer3_out[2264] = ~(layer2_out[3217] ^ layer2_out[3218]);
    assign layer3_out[2265] = layer2_out[1063];
    assign layer3_out[2266] = layer2_out[4506] & ~layer2_out[4505];
    assign layer3_out[2267] = ~layer2_out[1972];
    assign layer3_out[2268] = layer2_out[3054] | layer2_out[3055];
    assign layer3_out[2269] = ~layer2_out[4757];
    assign layer3_out[2270] = layer2_out[1937];
    assign layer3_out[2271] = layer2_out[2649];
    assign layer3_out[2272] = ~layer2_out[2578];
    assign layer3_out[2273] = layer2_out[3140];
    assign layer3_out[2274] = ~layer2_out[1169];
    assign layer3_out[2275] = layer2_out[7747] ^ layer2_out[7748];
    assign layer3_out[2276] = layer2_out[5530] ^ layer2_out[5531];
    assign layer3_out[2277] = ~layer2_out[7623];
    assign layer3_out[2278] = ~layer2_out[6604] | layer2_out[6605];
    assign layer3_out[2279] = layer2_out[7730] | layer2_out[7731];
    assign layer3_out[2280] = layer2_out[540];
    assign layer3_out[2281] = layer2_out[1935];
    assign layer3_out[2282] = ~(layer2_out[5002] ^ layer2_out[5003]);
    assign layer3_out[2283] = ~(layer2_out[7708] | layer2_out[7709]);
    assign layer3_out[2284] = ~layer2_out[3787] | layer2_out[3786];
    assign layer3_out[2285] = layer2_out[2545];
    assign layer3_out[2286] = ~layer2_out[5015] | layer2_out[5014];
    assign layer3_out[2287] = ~layer2_out[3530] | layer2_out[3531];
    assign layer3_out[2288] = layer2_out[7583] & ~layer2_out[7582];
    assign layer3_out[2289] = layer2_out[643] & ~layer2_out[644];
    assign layer3_out[2290] = layer2_out[7888];
    assign layer3_out[2291] = layer2_out[3906] & ~layer2_out[3905];
    assign layer3_out[2292] = layer2_out[4588];
    assign layer3_out[2293] = layer2_out[3923] ^ layer2_out[3924];
    assign layer3_out[2294] = ~layer2_out[1675];
    assign layer3_out[2295] = ~(layer2_out[7560] ^ layer2_out[7561]);
    assign layer3_out[2296] = layer2_out[3278] & layer2_out[3279];
    assign layer3_out[2297] = layer2_out[3654] & ~layer2_out[3655];
    assign layer3_out[2298] = layer2_out[3269] & ~layer2_out[3268];
    assign layer3_out[2299] = layer2_out[4908] | layer2_out[4909];
    assign layer3_out[2300] = layer2_out[5680];
    assign layer3_out[2301] = ~layer2_out[3704];
    assign layer3_out[2302] = ~layer2_out[5374];
    assign layer3_out[2303] = layer2_out[6121] | layer2_out[6122];
    assign layer3_out[2304] = layer2_out[7661];
    assign layer3_out[2305] = ~(layer2_out[2849] | layer2_out[2850]);
    assign layer3_out[2306] = ~layer2_out[740];
    assign layer3_out[2307] = ~(layer2_out[4939] | layer2_out[4940]);
    assign layer3_out[2308] = ~layer2_out[5461] | layer2_out[5460];
    assign layer3_out[2309] = ~(layer2_out[3097] & layer2_out[3098]);
    assign layer3_out[2310] = ~layer2_out[7110] | layer2_out[7111];
    assign layer3_out[2311] = layer2_out[926];
    assign layer3_out[2312] = layer2_out[6382];
    assign layer3_out[2313] = ~(layer2_out[7654] ^ layer2_out[7655]);
    assign layer3_out[2314] = ~layer2_out[6610];
    assign layer3_out[2315] = ~(layer2_out[3234] & layer2_out[3235]);
    assign layer3_out[2316] = layer2_out[4481] & ~layer2_out[4482];
    assign layer3_out[2317] = ~(layer2_out[7522] | layer2_out[7523]);
    assign layer3_out[2318] = ~layer2_out[3210] | layer2_out[3211];
    assign layer3_out[2319] = layer2_out[2249] & ~layer2_out[2248];
    assign layer3_out[2320] = layer2_out[3658] & layer2_out[3659];
    assign layer3_out[2321] = layer2_out[844] | layer2_out[845];
    assign layer3_out[2322] = ~layer2_out[1952];
    assign layer3_out[2323] = layer2_out[7133] & ~layer2_out[7132];
    assign layer3_out[2324] = ~layer2_out[2201];
    assign layer3_out[2325] = ~layer2_out[1477] | layer2_out[1476];
    assign layer3_out[2326] = ~layer2_out[5298] | layer2_out[5299];
    assign layer3_out[2327] = layer2_out[1682];
    assign layer3_out[2328] = ~(layer2_out[7526] ^ layer2_out[7527]);
    assign layer3_out[2329] = layer2_out[2724] | layer2_out[2725];
    assign layer3_out[2330] = layer2_out[323];
    assign layer3_out[2331] = layer2_out[1731];
    assign layer3_out[2332] = layer2_out[1569] & ~layer2_out[1568];
    assign layer3_out[2333] = layer2_out[6258] | layer2_out[6259];
    assign layer3_out[2334] = ~(layer2_out[4475] ^ layer2_out[4476]);
    assign layer3_out[2335] = ~layer2_out[277];
    assign layer3_out[2336] = ~(layer2_out[5515] ^ layer2_out[5516]);
    assign layer3_out[2337] = layer2_out[1379];
    assign layer3_out[2338] = ~(layer2_out[5864] | layer2_out[5865]);
    assign layer3_out[2339] = layer2_out[7208] ^ layer2_out[7209];
    assign layer3_out[2340] = ~layer2_out[2721];
    assign layer3_out[2341] = ~layer2_out[2463];
    assign layer3_out[2342] = layer2_out[5748];
    assign layer3_out[2343] = layer2_out[5923] ^ layer2_out[5924];
    assign layer3_out[2344] = layer2_out[550];
    assign layer3_out[2345] = 1'b0;
    assign layer3_out[2346] = ~(layer2_out[3446] ^ layer2_out[3447]);
    assign layer3_out[2347] = ~(layer2_out[3323] | layer2_out[3324]);
    assign layer3_out[2348] = ~layer2_out[3679];
    assign layer3_out[2349] = ~(layer2_out[6500] & layer2_out[6501]);
    assign layer3_out[2350] = layer2_out[5536];
    assign layer3_out[2351] = ~(layer2_out[958] | layer2_out[959]);
    assign layer3_out[2352] = layer2_out[4562];
    assign layer3_out[2353] = layer2_out[5014];
    assign layer3_out[2354] = layer2_out[2747];
    assign layer3_out[2355] = ~layer2_out[217];
    assign layer3_out[2356] = layer2_out[7776] & layer2_out[7777];
    assign layer3_out[2357] = layer2_out[7143] & ~layer2_out[7144];
    assign layer3_out[2358] = ~(layer2_out[7229] ^ layer2_out[7230]);
    assign layer3_out[2359] = ~layer2_out[4859];
    assign layer3_out[2360] = layer2_out[5273] ^ layer2_out[5274];
    assign layer3_out[2361] = layer2_out[173] & ~layer2_out[172];
    assign layer3_out[2362] = layer2_out[5438];
    assign layer3_out[2363] = layer2_out[992];
    assign layer3_out[2364] = layer2_out[2269];
    assign layer3_out[2365] = ~(layer2_out[4203] & layer2_out[4204]);
    assign layer3_out[2366] = ~layer2_out[5517];
    assign layer3_out[2367] = ~layer2_out[7285] | layer2_out[7284];
    assign layer3_out[2368] = layer2_out[5459] | layer2_out[5460];
    assign layer3_out[2369] = layer2_out[6882] | layer2_out[6883];
    assign layer3_out[2370] = layer2_out[7584] & ~layer2_out[7583];
    assign layer3_out[2371] = layer2_out[2150] ^ layer2_out[2151];
    assign layer3_out[2372] = layer2_out[3449];
    assign layer3_out[2373] = ~layer2_out[1877] | layer2_out[1876];
    assign layer3_out[2374] = ~layer2_out[5884];
    assign layer3_out[2375] = ~layer2_out[3010] | layer2_out[3009];
    assign layer3_out[2376] = layer2_out[7407] & ~layer2_out[7408];
    assign layer3_out[2377] = ~(layer2_out[3175] ^ layer2_out[3176]);
    assign layer3_out[2378] = ~layer2_out[5911];
    assign layer3_out[2379] = layer2_out[2206];
    assign layer3_out[2380] = ~layer2_out[3838] | layer2_out[3839];
    assign layer3_out[2381] = ~layer2_out[5447];
    assign layer3_out[2382] = ~layer2_out[7900] | layer2_out[7899];
    assign layer3_out[2383] = layer2_out[3063];
    assign layer3_out[2384] = ~(layer2_out[1464] ^ layer2_out[1465]);
    assign layer3_out[2385] = ~(layer2_out[1543] | layer2_out[1544]);
    assign layer3_out[2386] = ~layer2_out[265];
    assign layer3_out[2387] = layer2_out[6215];
    assign layer3_out[2388] = layer2_out[2421];
    assign layer3_out[2389] = ~layer2_out[3078];
    assign layer3_out[2390] = ~layer2_out[2897];
    assign layer3_out[2391] = ~layer2_out[7638];
    assign layer3_out[2392] = layer2_out[2247];
    assign layer3_out[2393] = ~layer2_out[4343];
    assign layer3_out[2394] = layer2_out[4518] & ~layer2_out[4519];
    assign layer3_out[2395] = ~layer2_out[4503];
    assign layer3_out[2396] = layer2_out[7112];
    assign layer3_out[2397] = ~layer2_out[621];
    assign layer3_out[2398] = ~(layer2_out[5149] | layer2_out[5150]);
    assign layer3_out[2399] = layer2_out[2135] & ~layer2_out[2136];
    assign layer3_out[2400] = layer2_out[2991] ^ layer2_out[2992];
    assign layer3_out[2401] = layer2_out[4298] ^ layer2_out[4299];
    assign layer3_out[2402] = ~(layer2_out[7131] & layer2_out[7132]);
    assign layer3_out[2403] = ~layer2_out[4984];
    assign layer3_out[2404] = ~layer2_out[3812];
    assign layer3_out[2405] = layer2_out[2892] & ~layer2_out[2893];
    assign layer3_out[2406] = layer2_out[2520];
    assign layer3_out[2407] = ~layer2_out[7322] | layer2_out[7321];
    assign layer3_out[2408] = layer2_out[5803] ^ layer2_out[5804];
    assign layer3_out[2409] = layer2_out[1423] & ~layer2_out[1422];
    assign layer3_out[2410] = ~(layer2_out[4445] & layer2_out[4446]);
    assign layer3_out[2411] = ~layer2_out[4515] | layer2_out[4514];
    assign layer3_out[2412] = ~(layer2_out[1698] ^ layer2_out[1699]);
    assign layer3_out[2413] = ~layer2_out[1156];
    assign layer3_out[2414] = layer2_out[6440] | layer2_out[6441];
    assign layer3_out[2415] = ~(layer2_out[3466] & layer2_out[3467]);
    assign layer3_out[2416] = layer2_out[5923] & ~layer2_out[5922];
    assign layer3_out[2417] = layer2_out[2971];
    assign layer3_out[2418] = layer2_out[7058];
    assign layer3_out[2419] = ~layer2_out[3533];
    assign layer3_out[2420] = ~layer2_out[2100];
    assign layer3_out[2421] = ~layer2_out[3902] | layer2_out[3903];
    assign layer3_out[2422] = ~(layer2_out[3483] & layer2_out[3484]);
    assign layer3_out[2423] = ~layer2_out[5211];
    assign layer3_out[2424] = layer2_out[359] & ~layer2_out[360];
    assign layer3_out[2425] = ~layer2_out[7824];
    assign layer3_out[2426] = layer2_out[1137] & ~layer2_out[1136];
    assign layer3_out[2427] = ~layer2_out[4987];
    assign layer3_out[2428] = ~layer2_out[6767] | layer2_out[6768];
    assign layer3_out[2429] = layer2_out[5711] & ~layer2_out[5712];
    assign layer3_out[2430] = ~(layer2_out[4200] | layer2_out[4201]);
    assign layer3_out[2431] = ~(layer2_out[2148] ^ layer2_out[2149]);
    assign layer3_out[2432] = ~layer2_out[439];
    assign layer3_out[2433] = ~layer2_out[5625];
    assign layer3_out[2434] = ~(layer2_out[2270] | layer2_out[2271]);
    assign layer3_out[2435] = ~layer2_out[5626];
    assign layer3_out[2436] = ~(layer2_out[3885] ^ layer2_out[3886]);
    assign layer3_out[2437] = layer2_out[324];
    assign layer3_out[2438] = ~layer2_out[4688] | layer2_out[4689];
    assign layer3_out[2439] = ~layer2_out[6653];
    assign layer3_out[2440] = ~layer2_out[1233] | layer2_out[1232];
    assign layer3_out[2441] = layer2_out[3549] & ~layer2_out[3548];
    assign layer3_out[2442] = layer2_out[3833];
    assign layer3_out[2443] = ~layer2_out[4818];
    assign layer3_out[2444] = layer2_out[5127] & ~layer2_out[5128];
    assign layer3_out[2445] = layer2_out[494] & ~layer2_out[495];
    assign layer3_out[2446] = ~layer2_out[4648] | layer2_out[4647];
    assign layer3_out[2447] = ~layer2_out[4153];
    assign layer3_out[2448] = ~layer2_out[818];
    assign layer3_out[2449] = ~layer2_out[236] | layer2_out[235];
    assign layer3_out[2450] = layer2_out[1258];
    assign layer3_out[2451] = ~(layer2_out[89] | layer2_out[90]);
    assign layer3_out[2452] = layer2_out[3886] & ~layer2_out[3887];
    assign layer3_out[2453] = layer2_out[3596];
    assign layer3_out[2454] = layer2_out[7969];
    assign layer3_out[2455] = layer2_out[4778];
    assign layer3_out[2456] = layer2_out[6505];
    assign layer3_out[2457] = layer2_out[294] ^ layer2_out[295];
    assign layer3_out[2458] = layer2_out[3111];
    assign layer3_out[2459] = ~layer2_out[1637];
    assign layer3_out[2460] = layer2_out[1886] & ~layer2_out[1885];
    assign layer3_out[2461] = ~layer2_out[7360] | layer2_out[7361];
    assign layer3_out[2462] = layer2_out[7683] & ~layer2_out[7682];
    assign layer3_out[2463] = ~(layer2_out[6239] | layer2_out[6240]);
    assign layer3_out[2464] = ~(layer2_out[2797] & layer2_out[2798]);
    assign layer3_out[2465] = ~(layer2_out[54] | layer2_out[55]);
    assign layer3_out[2466] = layer2_out[5631] & ~layer2_out[5630];
    assign layer3_out[2467] = layer2_out[5825] & ~layer2_out[5826];
    assign layer3_out[2468] = ~layer2_out[4988];
    assign layer3_out[2469] = ~layer2_out[5511];
    assign layer3_out[2470] = ~layer2_out[3473];
    assign layer3_out[2471] = ~layer2_out[2279];
    assign layer3_out[2472] = layer2_out[7633];
    assign layer3_out[2473] = layer2_out[777];
    assign layer3_out[2474] = ~(layer2_out[6705] | layer2_out[6706]);
    assign layer3_out[2475] = layer2_out[6929];
    assign layer3_out[2476] = ~layer2_out[6369] | layer2_out[6368];
    assign layer3_out[2477] = layer2_out[4793] & ~layer2_out[4792];
    assign layer3_out[2478] = layer2_out[704] & ~layer2_out[705];
    assign layer3_out[2479] = ~layer2_out[7795];
    assign layer3_out[2480] = layer2_out[1845];
    assign layer3_out[2481] = layer2_out[6359] | layer2_out[6360];
    assign layer3_out[2482] = ~(layer2_out[6541] | layer2_out[6542]);
    assign layer3_out[2483] = ~(layer2_out[4490] ^ layer2_out[4491]);
    assign layer3_out[2484] = layer2_out[1280];
    assign layer3_out[2485] = layer2_out[5252] ^ layer2_out[5253];
    assign layer3_out[2486] = layer2_out[4126];
    assign layer3_out[2487] = ~layer2_out[7610] | layer2_out[7611];
    assign layer3_out[2488] = ~layer2_out[1983];
    assign layer3_out[2489] = ~(layer2_out[5152] & layer2_out[5153]);
    assign layer3_out[2490] = layer2_out[141] ^ layer2_out[142];
    assign layer3_out[2491] = ~layer2_out[4322];
    assign layer3_out[2492] = ~layer2_out[7006];
    assign layer3_out[2493] = layer2_out[6545];
    assign layer3_out[2494] = layer2_out[4066] ^ layer2_out[4067];
    assign layer3_out[2495] = ~layer2_out[1900];
    assign layer3_out[2496] = layer2_out[5091] | layer2_out[5092];
    assign layer3_out[2497] = ~layer2_out[4151] | layer2_out[4150];
    assign layer3_out[2498] = ~layer2_out[7740];
    assign layer3_out[2499] = layer2_out[7943] ^ layer2_out[7944];
    assign layer3_out[2500] = ~layer2_out[3613];
    assign layer3_out[2501] = ~layer2_out[6513];
    assign layer3_out[2502] = ~layer2_out[2847];
    assign layer3_out[2503] = layer2_out[2281] | layer2_out[2282];
    assign layer3_out[2504] = ~(layer2_out[7179] ^ layer2_out[7180]);
    assign layer3_out[2505] = layer2_out[2790] & ~layer2_out[2791];
    assign layer3_out[2506] = ~(layer2_out[2127] & layer2_out[2128]);
    assign layer3_out[2507] = layer2_out[7009] & layer2_out[7010];
    assign layer3_out[2508] = ~layer2_out[3018] | layer2_out[3017];
    assign layer3_out[2509] = layer2_out[7669] & layer2_out[7670];
    assign layer3_out[2510] = layer2_out[6653];
    assign layer3_out[2511] = ~layer2_out[6175];
    assign layer3_out[2512] = ~(layer2_out[1827] | layer2_out[1828]);
    assign layer3_out[2513] = ~layer2_out[6782] | layer2_out[6783];
    assign layer3_out[2514] = layer2_out[1566];
    assign layer3_out[2515] = ~layer2_out[1192];
    assign layer3_out[2516] = ~layer2_out[692];
    assign layer3_out[2517] = ~layer2_out[1214];
    assign layer3_out[2518] = ~layer2_out[3992];
    assign layer3_out[2519] = layer2_out[7657] ^ layer2_out[7658];
    assign layer3_out[2520] = ~(layer2_out[7183] & layer2_out[7184]);
    assign layer3_out[2521] = layer2_out[6608] | layer2_out[6609];
    assign layer3_out[2522] = layer2_out[2599];
    assign layer3_out[2523] = layer2_out[5351];
    assign layer3_out[2524] = ~layer2_out[6018] | layer2_out[6017];
    assign layer3_out[2525] = ~layer2_out[7877];
    assign layer3_out[2526] = layer2_out[2884] | layer2_out[2885];
    assign layer3_out[2527] = ~(layer2_out[6774] | layer2_out[6775]);
    assign layer3_out[2528] = ~layer2_out[5079] | layer2_out[5080];
    assign layer3_out[2529] = ~layer2_out[7634];
    assign layer3_out[2530] = layer2_out[1778] | layer2_out[1779];
    assign layer3_out[2531] = ~layer2_out[835] | layer2_out[834];
    assign layer3_out[2532] = layer2_out[6387];
    assign layer3_out[2533] = layer2_out[7335] & ~layer2_out[7334];
    assign layer3_out[2534] = ~layer2_out[6000];
    assign layer3_out[2535] = layer2_out[5634];
    assign layer3_out[2536] = layer2_out[1665] | layer2_out[1666];
    assign layer3_out[2537] = 1'b1;
    assign layer3_out[2538] = layer2_out[995];
    assign layer3_out[2539] = ~layer2_out[6863];
    assign layer3_out[2540] = layer2_out[3409];
    assign layer3_out[2541] = ~(layer2_out[4855] | layer2_out[4856]);
    assign layer3_out[2542] = layer2_out[3139] & ~layer2_out[3138];
    assign layer3_out[2543] = layer2_out[7282] & ~layer2_out[7283];
    assign layer3_out[2544] = ~layer2_out[1858];
    assign layer3_out[2545] = layer2_out[6015];
    assign layer3_out[2546] = ~(layer2_out[5349] & layer2_out[5350]);
    assign layer3_out[2547] = layer2_out[5217] | layer2_out[5218];
    assign layer3_out[2548] = layer2_out[5044] & ~layer2_out[5045];
    assign layer3_out[2549] = layer2_out[6243] ^ layer2_out[6244];
    assign layer3_out[2550] = layer2_out[4278];
    assign layer3_out[2551] = layer2_out[2211];
    assign layer3_out[2552] = layer2_out[2205] ^ layer2_out[2206];
    assign layer3_out[2553] = ~layer2_out[251];
    assign layer3_out[2554] = layer2_out[4611] & ~layer2_out[4612];
    assign layer3_out[2555] = ~layer2_out[5352];
    assign layer3_out[2556] = ~layer2_out[3782];
    assign layer3_out[2557] = layer2_out[933];
    assign layer3_out[2558] = layer2_out[649] & layer2_out[650];
    assign layer3_out[2559] = layer2_out[2461] & ~layer2_out[2460];
    assign layer3_out[2560] = ~(layer2_out[3817] | layer2_out[3818]);
    assign layer3_out[2561] = layer2_out[1414] ^ layer2_out[1415];
    assign layer3_out[2562] = layer2_out[4130] & ~layer2_out[4131];
    assign layer3_out[2563] = ~layer2_out[4697];
    assign layer3_out[2564] = ~layer2_out[4182] | layer2_out[4183];
    assign layer3_out[2565] = 1'b1;
    assign layer3_out[2566] = ~layer2_out[957] | layer2_out[956];
    assign layer3_out[2567] = layer2_out[2632] & layer2_out[2633];
    assign layer3_out[2568] = layer2_out[5743];
    assign layer3_out[2569] = layer2_out[596] & layer2_out[597];
    assign layer3_out[2570] = layer2_out[1986];
    assign layer3_out[2571] = layer2_out[1147] & layer2_out[1148];
    assign layer3_out[2572] = ~(layer2_out[3372] ^ layer2_out[3373]);
    assign layer3_out[2573] = 1'b1;
    assign layer3_out[2574] = layer2_out[7092] ^ layer2_out[7093];
    assign layer3_out[2575] = ~(layer2_out[2282] ^ layer2_out[2283]);
    assign layer3_out[2576] = layer2_out[4795] & layer2_out[4796];
    assign layer3_out[2577] = ~(layer2_out[3146] & layer2_out[3147]);
    assign layer3_out[2578] = layer2_out[2160];
    assign layer3_out[2579] = layer2_out[1033];
    assign layer3_out[2580] = ~layer2_out[6196] | layer2_out[6195];
    assign layer3_out[2581] = ~layer2_out[6294] | layer2_out[6293];
    assign layer3_out[2582] = ~layer2_out[1455];
    assign layer3_out[2583] = ~(layer2_out[2625] | layer2_out[2626]);
    assign layer3_out[2584] = layer2_out[1194] & ~layer2_out[1193];
    assign layer3_out[2585] = layer2_out[151] ^ layer2_out[152];
    assign layer3_out[2586] = layer2_out[7168] & ~layer2_out[7169];
    assign layer3_out[2587] = layer2_out[0];
    assign layer3_out[2588] = layer2_out[2473] & layer2_out[2474];
    assign layer3_out[2589] = ~layer2_out[4537];
    assign layer3_out[2590] = layer2_out[555] & ~layer2_out[554];
    assign layer3_out[2591] = layer2_out[6071];
    assign layer3_out[2592] = layer2_out[7588] | layer2_out[7589];
    assign layer3_out[2593] = ~layer2_out[3630] | layer2_out[3631];
    assign layer3_out[2594] = ~(layer2_out[6333] | layer2_out[6334]);
    assign layer3_out[2595] = ~layer2_out[5524] | layer2_out[5523];
    assign layer3_out[2596] = layer2_out[2481];
    assign layer3_out[2597] = layer2_out[2628];
    assign layer3_out[2598] = ~layer2_out[7280];
    assign layer3_out[2599] = layer2_out[7277] ^ layer2_out[7278];
    assign layer3_out[2600] = ~(layer2_out[3442] | layer2_out[3443]);
    assign layer3_out[2601] = 1'b1;
    assign layer3_out[2602] = layer2_out[6186] ^ layer2_out[6187];
    assign layer3_out[2603] = ~(layer2_out[5497] & layer2_out[5498]);
    assign layer3_out[2604] = layer2_out[2675];
    assign layer3_out[2605] = ~(layer2_out[5596] ^ layer2_out[5597]);
    assign layer3_out[2606] = ~layer2_out[2083];
    assign layer3_out[2607] = 1'b1;
    assign layer3_out[2608] = ~layer2_out[1331];
    assign layer3_out[2609] = layer2_out[3789] & ~layer2_out[3788];
    assign layer3_out[2610] = ~(layer2_out[4339] ^ layer2_out[4340]);
    assign layer3_out[2611] = layer2_out[5271];
    assign layer3_out[2612] = layer2_out[6612] & ~layer2_out[6611];
    assign layer3_out[2613] = layer2_out[4209];
    assign layer3_out[2614] = ~(layer2_out[1102] ^ layer2_out[1103]);
    assign layer3_out[2615] = layer2_out[7140] | layer2_out[7141];
    assign layer3_out[2616] = ~layer2_out[443] | layer2_out[442];
    assign layer3_out[2617] = layer2_out[483] | layer2_out[484];
    assign layer3_out[2618] = ~layer2_out[7178];
    assign layer3_out[2619] = ~layer2_out[1453] | layer2_out[1452];
    assign layer3_out[2620] = ~layer2_out[6370];
    assign layer3_out[2621] = ~layer2_out[3940];
    assign layer3_out[2622] = layer2_out[4640];
    assign layer3_out[2623] = ~layer2_out[2743] | layer2_out[2744];
    assign layer3_out[2624] = layer2_out[64];
    assign layer3_out[2625] = layer2_out[5336];
    assign layer3_out[2626] = ~layer2_out[6539] | layer2_out[6540];
    assign layer3_out[2627] = ~(layer2_out[5697] & layer2_out[5698]);
    assign layer3_out[2628] = ~(layer2_out[5492] ^ layer2_out[5493]);
    assign layer3_out[2629] = ~layer2_out[3388] | layer2_out[3389];
    assign layer3_out[2630] = ~layer2_out[565];
    assign layer3_out[2631] = ~layer2_out[1577];
    assign layer3_out[2632] = ~layer2_out[7546] | layer2_out[7545];
    assign layer3_out[2633] = layer2_out[6278];
    assign layer3_out[2634] = ~(layer2_out[5145] | layer2_out[5146]);
    assign layer3_out[2635] = layer2_out[3195] & layer2_out[3196];
    assign layer3_out[2636] = ~layer2_out[4817];
    assign layer3_out[2637] = layer2_out[2285];
    assign layer3_out[2638] = layer2_out[4632] | layer2_out[4633];
    assign layer3_out[2639] = layer2_out[3792] ^ layer2_out[3793];
    assign layer3_out[2640] = layer2_out[3728];
    assign layer3_out[2641] = layer2_out[6207];
    assign layer3_out[2642] = layer2_out[3581] & layer2_out[3582];
    assign layer3_out[2643] = ~layer2_out[2108];
    assign layer3_out[2644] = ~layer2_out[1685];
    assign layer3_out[2645] = layer2_out[4991];
    assign layer3_out[2646] = layer2_out[4020] ^ layer2_out[4021];
    assign layer3_out[2647] = ~layer2_out[6113] | layer2_out[6112];
    assign layer3_out[2648] = layer2_out[821];
    assign layer3_out[2649] = ~(layer2_out[6134] | layer2_out[6135]);
    assign layer3_out[2650] = layer2_out[6674] ^ layer2_out[6675];
    assign layer3_out[2651] = layer2_out[405] & layer2_out[406];
    assign layer3_out[2652] = ~layer2_out[85] | layer2_out[86];
    assign layer3_out[2653] = layer2_out[1515];
    assign layer3_out[2654] = 1'b1;
    assign layer3_out[2655] = layer2_out[3669] & layer2_out[3670];
    assign layer3_out[2656] = layer2_out[5575] & layer2_out[5576];
    assign layer3_out[2657] = layer2_out[4303];
    assign layer3_out[2658] = ~(layer2_out[44] | layer2_out[45]);
    assign layer3_out[2659] = layer2_out[3801] & ~layer2_out[3800];
    assign layer3_out[2660] = layer2_out[4545];
    assign layer3_out[2661] = 1'b0;
    assign layer3_out[2662] = layer2_out[2198] & ~layer2_out[2199];
    assign layer3_out[2663] = ~layer2_out[4117];
    assign layer3_out[2664] = ~layer2_out[6183] | layer2_out[6184];
    assign layer3_out[2665] = ~layer2_out[5223] | layer2_out[5224];
    assign layer3_out[2666] = layer2_out[7247] | layer2_out[7248];
    assign layer3_out[2667] = ~layer2_out[6627] | layer2_out[6626];
    assign layer3_out[2668] = ~(layer2_out[2180] | layer2_out[2181]);
    assign layer3_out[2669] = layer2_out[4241];
    assign layer3_out[2670] = ~(layer2_out[4813] & layer2_out[4814]);
    assign layer3_out[2671] = 1'b1;
    assign layer3_out[2672] = ~(layer2_out[4100] | layer2_out[4101]);
    assign layer3_out[2673] = layer2_out[1960];
    assign layer3_out[2674] = ~layer2_out[1822];
    assign layer3_out[2675] = ~(layer2_out[5875] & layer2_out[5876]);
    assign layer3_out[2676] = layer2_out[1958];
    assign layer3_out[2677] = layer2_out[5120];
    assign layer3_out[2678] = ~layer2_out[7096];
    assign layer3_out[2679] = ~layer2_out[4210];
    assign layer3_out[2680] = layer2_out[7167];
    assign layer3_out[2681] = layer2_out[4394] & layer2_out[4395];
    assign layer3_out[2682] = layer2_out[5733];
    assign layer3_out[2683] = layer2_out[1699] | layer2_out[1700];
    assign layer3_out[2684] = ~layer2_out[5688];
    assign layer3_out[2685] = layer2_out[7166];
    assign layer3_out[2686] = layer2_out[4374];
    assign layer3_out[2687] = layer2_out[1759];
    assign layer3_out[2688] = layer2_out[5429] & ~layer2_out[5428];
    assign layer3_out[2689] = ~(layer2_out[1103] ^ layer2_out[1104]);
    assign layer3_out[2690] = layer2_out[5971] & layer2_out[5972];
    assign layer3_out[2691] = layer2_out[5090] ^ layer2_out[5091];
    assign layer3_out[2692] = ~layer2_out[4757];
    assign layer3_out[2693] = ~(layer2_out[3621] ^ layer2_out[3622]);
    assign layer3_out[2694] = ~layer2_out[5362];
    assign layer3_out[2695] = ~(layer2_out[791] ^ layer2_out[792]);
    assign layer3_out[2696] = ~(layer2_out[41] ^ layer2_out[42]);
    assign layer3_out[2697] = layer2_out[7596] | layer2_out[7597];
    assign layer3_out[2698] = layer2_out[2948];
    assign layer3_out[2699] = 1'b0;
    assign layer3_out[2700] = ~layer2_out[2293];
    assign layer3_out[2701] = ~layer2_out[5475];
    assign layer3_out[2702] = layer2_out[6122] & layer2_out[6123];
    assign layer3_out[2703] = layer2_out[6673] & ~layer2_out[6672];
    assign layer3_out[2704] = 1'b0;
    assign layer3_out[2705] = ~layer2_out[2174];
    assign layer3_out[2706] = layer2_out[6911];
    assign layer3_out[2707] = layer2_out[1612];
    assign layer3_out[2708] = layer2_out[4032];
    assign layer3_out[2709] = layer2_out[3083];
    assign layer3_out[2710] = layer2_out[490];
    assign layer3_out[2711] = ~layer2_out[6174];
    assign layer3_out[2712] = ~layer2_out[7570] | layer2_out[7569];
    assign layer3_out[2713] = layer2_out[4018];
    assign layer3_out[2714] = ~layer2_out[1920];
    assign layer3_out[2715] = ~layer2_out[945];
    assign layer3_out[2716] = ~layer2_out[7085];
    assign layer3_out[2717] = ~layer2_out[4186];
    assign layer3_out[2718] = ~layer2_out[5994];
    assign layer3_out[2719] = layer2_out[5330];
    assign layer3_out[2720] = layer2_out[6315];
    assign layer3_out[2721] = layer2_out[6473];
    assign layer3_out[2722] = layer2_out[2694] | layer2_out[2695];
    assign layer3_out[2723] = ~layer2_out[5222];
    assign layer3_out[2724] = ~layer2_out[4166];
    assign layer3_out[2725] = ~(layer2_out[5498] | layer2_out[5499]);
    assign layer3_out[2726] = layer2_out[820] & ~layer2_out[819];
    assign layer3_out[2727] = layer2_out[6908] ^ layer2_out[6909];
    assign layer3_out[2728] = ~(layer2_out[232] ^ layer2_out[233]);
    assign layer3_out[2729] = layer2_out[7587];
    assign layer3_out[2730] = ~(layer2_out[2894] & layer2_out[2895]);
    assign layer3_out[2731] = ~layer2_out[1461];
    assign layer3_out[2732] = ~layer2_out[745] | layer2_out[746];
    assign layer3_out[2733] = ~layer2_out[3889];
    assign layer3_out[2734] = ~layer2_out[4534];
    assign layer3_out[2735] = ~layer2_out[1102] | layer2_out[1101];
    assign layer3_out[2736] = ~layer2_out[1787];
    assign layer3_out[2737] = layer2_out[4681] & ~layer2_out[4680];
    assign layer3_out[2738] = layer2_out[6010] & ~layer2_out[6011];
    assign layer3_out[2739] = ~(layer2_out[3875] | layer2_out[3876]);
    assign layer3_out[2740] = layer2_out[4419] | layer2_out[4420];
    assign layer3_out[2741] = layer2_out[437] ^ layer2_out[438];
    assign layer3_out[2742] = layer2_out[1118] & ~layer2_out[1119];
    assign layer3_out[2743] = layer2_out[1767] & ~layer2_out[1768];
    assign layer3_out[2744] = ~layer2_out[458];
    assign layer3_out[2745] = layer2_out[2371];
    assign layer3_out[2746] = layer2_out[5203] & ~layer2_out[5202];
    assign layer3_out[2747] = ~layer2_out[808];
    assign layer3_out[2748] = layer2_out[6480] & ~layer2_out[6479];
    assign layer3_out[2749] = ~(layer2_out[7509] & layer2_out[7510]);
    assign layer3_out[2750] = ~(layer2_out[4831] ^ layer2_out[4832]);
    assign layer3_out[2751] = layer2_out[1074] | layer2_out[1075];
    assign layer3_out[2752] = layer2_out[3192];
    assign layer3_out[2753] = layer2_out[5095];
    assign layer3_out[2754] = ~(layer2_out[6110] & layer2_out[6111]);
    assign layer3_out[2755] = layer2_out[6405] & ~layer2_out[6406];
    assign layer3_out[2756] = layer2_out[122] ^ layer2_out[123];
    assign layer3_out[2757] = layer2_out[3292];
    assign layer3_out[2758] = layer2_out[2717] & ~layer2_out[2718];
    assign layer3_out[2759] = ~layer2_out[2467] | layer2_out[2468];
    assign layer3_out[2760] = ~(layer2_out[7141] ^ layer2_out[7142]);
    assign layer3_out[2761] = ~layer2_out[1008];
    assign layer3_out[2762] = layer2_out[1608] & layer2_out[1609];
    assign layer3_out[2763] = layer2_out[1149];
    assign layer3_out[2764] = layer2_out[5289];
    assign layer3_out[2765] = layer2_out[4629] ^ layer2_out[4630];
    assign layer3_out[2766] = ~(layer2_out[3471] ^ layer2_out[3472]);
    assign layer3_out[2767] = layer2_out[2533];
    assign layer3_out[2768] = ~(layer2_out[961] & layer2_out[962]);
    assign layer3_out[2769] = layer2_out[3921] & ~layer2_out[3922];
    assign layer3_out[2770] = layer2_out[1852] & ~layer2_out[1853];
    assign layer3_out[2771] = layer2_out[7758];
    assign layer3_out[2772] = ~layer2_out[1463];
    assign layer3_out[2773] = layer2_out[6203] & ~layer2_out[6204];
    assign layer3_out[2774] = ~layer2_out[6639] | layer2_out[6640];
    assign layer3_out[2775] = ~layer2_out[5759];
    assign layer3_out[2776] = ~layer2_out[7119] | layer2_out[7120];
    assign layer3_out[2777] = layer2_out[2878];
    assign layer3_out[2778] = layer2_out[1835];
    assign layer3_out[2779] = layer2_out[3790] & ~layer2_out[3789];
    assign layer3_out[2780] = ~(layer2_out[5852] | layer2_out[5853]);
    assign layer3_out[2781] = ~(layer2_out[6889] | layer2_out[6890]);
    assign layer3_out[2782] = layer2_out[5218];
    assign layer3_out[2783] = ~(layer2_out[693] | layer2_out[694]);
    assign layer3_out[2784] = 1'b0;
    assign layer3_out[2785] = layer2_out[5703] ^ layer2_out[5704];
    assign layer3_out[2786] = ~layer2_out[1840] | layer2_out[1839];
    assign layer3_out[2787] = layer2_out[6438];
    assign layer3_out[2788] = layer2_out[2712] & ~layer2_out[2711];
    assign layer3_out[2789] = layer2_out[7191];
    assign layer3_out[2790] = layer2_out[7500];
    assign layer3_out[2791] = layer2_out[3353] & ~layer2_out[3354];
    assign layer3_out[2792] = layer2_out[66];
    assign layer3_out[2793] = ~layer2_out[2537];
    assign layer3_out[2794] = layer2_out[3777] ^ layer2_out[3778];
    assign layer3_out[2795] = layer2_out[7336] & ~layer2_out[7335];
    assign layer3_out[2796] = 1'b0;
    assign layer3_out[2797] = ~layer2_out[6705];
    assign layer3_out[2798] = 1'b0;
    assign layer3_out[2799] = ~layer2_out[4332];
    assign layer3_out[2800] = ~layer2_out[3713] | layer2_out[3712];
    assign layer3_out[2801] = ~layer2_out[2703];
    assign layer3_out[2802] = layer2_out[3999] & ~layer2_out[3998];
    assign layer3_out[2803] = ~(layer2_out[7737] ^ layer2_out[7738]);
    assign layer3_out[2804] = layer2_out[7717] | layer2_out[7718];
    assign layer3_out[2805] = ~layer2_out[2409];
    assign layer3_out[2806] = ~(layer2_out[3569] ^ layer2_out[3570]);
    assign layer3_out[2807] = layer2_out[5985] | layer2_out[5986];
    assign layer3_out[2808] = layer2_out[1673] ^ layer2_out[1674];
    assign layer3_out[2809] = 1'b0;
    assign layer3_out[2810] = ~layer2_out[382] | layer2_out[383];
    assign layer3_out[2811] = ~layer2_out[2436];
    assign layer3_out[2812] = layer2_out[4610] | layer2_out[4611];
    assign layer3_out[2813] = layer2_out[6] & ~layer2_out[5];
    assign layer3_out[2814] = layer2_out[3541] & ~layer2_out[3542];
    assign layer3_out[2815] = layer2_out[6530] & ~layer2_out[6531];
    assign layer3_out[2816] = layer2_out[525] | layer2_out[526];
    assign layer3_out[2817] = layer2_out[2774];
    assign layer3_out[2818] = ~layer2_out[5363] | layer2_out[5364];
    assign layer3_out[2819] = ~layer2_out[4972];
    assign layer3_out[2820] = layer2_out[839] & ~layer2_out[838];
    assign layer3_out[2821] = ~layer2_out[1158];
    assign layer3_out[2822] = ~layer2_out[3428];
    assign layer3_out[2823] = ~(layer2_out[2476] ^ layer2_out[2477]);
    assign layer3_out[2824] = layer2_out[5786] & ~layer2_out[5787];
    assign layer3_out[2825] = layer2_out[6806] & ~layer2_out[6805];
    assign layer3_out[2826] = layer2_out[1737];
    assign layer3_out[2827] = layer2_out[7059] & ~layer2_out[7060];
    assign layer3_out[2828] = layer2_out[968];
    assign layer3_out[2829] = ~(layer2_out[147] & layer2_out[148]);
    assign layer3_out[2830] = layer2_out[2888];
    assign layer3_out[2831] = layer2_out[3881] & layer2_out[3882];
    assign layer3_out[2832] = layer2_out[4785] & ~layer2_out[4786];
    assign layer3_out[2833] = ~layer2_out[2082];
    assign layer3_out[2834] = layer2_out[2200];
    assign layer3_out[2835] = ~layer2_out[4457];
    assign layer3_out[2836] = layer2_out[3944];
    assign layer3_out[2837] = layer2_out[4708] ^ layer2_out[4709];
    assign layer3_out[2838] = layer2_out[6034] ^ layer2_out[6035];
    assign layer3_out[2839] = layer2_out[5834];
    assign layer3_out[2840] = layer2_out[5073];
    assign layer3_out[2841] = ~layer2_out[7353] | layer2_out[7354];
    assign layer3_out[2842] = ~(layer2_out[3566] | layer2_out[3567]);
    assign layer3_out[2843] = ~layer2_out[1350];
    assign layer3_out[2844] = ~(layer2_out[6123] | layer2_out[6124]);
    assign layer3_out[2845] = ~(layer2_out[1623] | layer2_out[1624]);
    assign layer3_out[2846] = layer2_out[355] & ~layer2_out[354];
    assign layer3_out[2847] = ~layer2_out[1697];
    assign layer3_out[2848] = layer2_out[4886] & layer2_out[4887];
    assign layer3_out[2849] = layer2_out[1582];
    assign layer3_out[2850] = layer2_out[5929];
    assign layer3_out[2851] = layer2_out[6912] ^ layer2_out[6913];
    assign layer3_out[2852] = ~(layer2_out[2531] ^ layer2_out[2532]);
    assign layer3_out[2853] = ~(layer2_out[780] & layer2_out[781]);
    assign layer3_out[2854] = layer2_out[5785];
    assign layer3_out[2855] = layer2_out[6631];
    assign layer3_out[2856] = layer2_out[6045];
    assign layer3_out[2857] = ~layer2_out[4062];
    assign layer3_out[2858] = layer2_out[1834];
    assign layer3_out[2859] = layer2_out[5193];
    assign layer3_out[2860] = layer2_out[1427];
    assign layer3_out[2861] = layer2_out[3707];
    assign layer3_out[2862] = layer2_out[1987] & ~layer2_out[1988];
    assign layer3_out[2863] = layer2_out[4683];
    assign layer3_out[2864] = layer2_out[4214];
    assign layer3_out[2865] = layer2_out[3066] & layer2_out[3067];
    assign layer3_out[2866] = layer2_out[1344];
    assign layer3_out[2867] = ~layer2_out[97] | layer2_out[96];
    assign layer3_out[2868] = ~layer2_out[1659];
    assign layer3_out[2869] = layer2_out[111];
    assign layer3_out[2870] = layer2_out[6319] | layer2_out[6320];
    assign layer3_out[2871] = layer2_out[2825] & ~layer2_out[2824];
    assign layer3_out[2872] = layer2_out[1269] | layer2_out[1270];
    assign layer3_out[2873] = layer2_out[1335] ^ layer2_out[1336];
    assign layer3_out[2874] = layer2_out[5325];
    assign layer3_out[2875] = layer2_out[1001];
    assign layer3_out[2876] = layer2_out[3644] & layer2_out[3645];
    assign layer3_out[2877] = layer2_out[3960];
    assign layer3_out[2878] = 1'b1;
    assign layer3_out[2879] = layer2_out[3357] & layer2_out[3358];
    assign layer3_out[2880] = ~layer2_out[4170] | layer2_out[4171];
    assign layer3_out[2881] = layer2_out[1683] | layer2_out[1684];
    assign layer3_out[2882] = layer2_out[6533] & layer2_out[6534];
    assign layer3_out[2883] = ~layer2_out[3885];
    assign layer3_out[2884] = layer2_out[242] ^ layer2_out[243];
    assign layer3_out[2885] = ~layer2_out[4630];
    assign layer3_out[2886] = ~layer2_out[6899];
    assign layer3_out[2887] = ~(layer2_out[6133] | layer2_out[6134]);
    assign layer3_out[2888] = layer2_out[1457] & layer2_out[1458];
    assign layer3_out[2889] = layer2_out[7474];
    assign layer3_out[2890] = layer2_out[1409] & ~layer2_out[1408];
    assign layer3_out[2891] = ~layer2_out[5910] | layer2_out[5911];
    assign layer3_out[2892] = layer2_out[4420];
    assign layer3_out[2893] = ~layer2_out[2425];
    assign layer3_out[2894] = layer2_out[4069];
    assign layer3_out[2895] = ~layer2_out[2442];
    assign layer3_out[2896] = ~(layer2_out[1527] ^ layer2_out[1528]);
    assign layer3_out[2897] = ~layer2_out[6918];
    assign layer3_out[2898] = layer2_out[4605] & layer2_out[4606];
    assign layer3_out[2899] = layer2_out[2535] & ~layer2_out[2536];
    assign layer3_out[2900] = layer2_out[591] & ~layer2_out[590];
    assign layer3_out[2901] = ~layer2_out[3825] | layer2_out[3826];
    assign layer3_out[2902] = layer2_out[7559] & ~layer2_out[7560];
    assign layer3_out[2903] = layer2_out[4112];
    assign layer3_out[2904] = layer2_out[5515] & ~layer2_out[5514];
    assign layer3_out[2905] = ~layer2_out[3599];
    assign layer3_out[2906] = layer2_out[5628] & ~layer2_out[5629];
    assign layer3_out[2907] = layer2_out[6126] & layer2_out[6127];
    assign layer3_out[2908] = ~layer2_out[1417];
    assign layer3_out[2909] = ~layer2_out[4957] | layer2_out[4958];
    assign layer3_out[2910] = layer2_out[3361];
    assign layer3_out[2911] = layer2_out[1304] ^ layer2_out[1305];
    assign layer3_out[2912] = layer2_out[4754];
    assign layer3_out[2913] = layer2_out[7472] & ~layer2_out[7471];
    assign layer3_out[2914] = ~layer2_out[949];
    assign layer3_out[2915] = ~layer2_out[2109];
    assign layer3_out[2916] = ~layer2_out[506];
    assign layer3_out[2917] = ~layer2_out[1753] | layer2_out[1752];
    assign layer3_out[2918] = ~layer2_out[4772];
    assign layer3_out[2919] = ~(layer2_out[2238] & layer2_out[2239]);
    assign layer3_out[2920] = layer2_out[1211];
    assign layer3_out[2921] = layer2_out[3032] | layer2_out[3033];
    assign layer3_out[2922] = layer2_out[1380];
    assign layer3_out[2923] = ~(layer2_out[6411] & layer2_out[6412]);
    assign layer3_out[2924] = layer2_out[3498] | layer2_out[3499];
    assign layer3_out[2925] = 1'b1;
    assign layer3_out[2926] = ~(layer2_out[1997] ^ layer2_out[1998]);
    assign layer3_out[2927] = ~(layer2_out[4239] & layer2_out[4240]);
    assign layer3_out[2928] = layer2_out[4284];
    assign layer3_out[2929] = ~layer2_out[1265];
    assign layer3_out[2930] = ~layer2_out[3901];
    assign layer3_out[2931] = layer2_out[6773] ^ layer2_out[6774];
    assign layer3_out[2932] = ~layer2_out[6397] | layer2_out[6396];
    assign layer3_out[2933] = layer2_out[1382];
    assign layer3_out[2934] = ~layer2_out[6099];
    assign layer3_out[2935] = ~layer2_out[5682];
    assign layer3_out[2936] = layer2_out[2641] ^ layer2_out[2642];
    assign layer3_out[2937] = layer2_out[6860] | layer2_out[6861];
    assign layer3_out[2938] = layer2_out[6059];
    assign layer3_out[2939] = layer2_out[2190] & ~layer2_out[2191];
    assign layer3_out[2940] = ~(layer2_out[7099] & layer2_out[7100]);
    assign layer3_out[2941] = layer2_out[42] & ~layer2_out[43];
    assign layer3_out[2942] = ~layer2_out[2941] | layer2_out[2940];
    assign layer3_out[2943] = layer2_out[5588] | layer2_out[5589];
    assign layer3_out[2944] = layer2_out[2265] & layer2_out[2266];
    assign layer3_out[2945] = ~(layer2_out[5722] | layer2_out[5723]);
    assign layer3_out[2946] = layer2_out[6276];
    assign layer3_out[2947] = ~layer2_out[4235] | layer2_out[4234];
    assign layer3_out[2948] = layer2_out[2043] & ~layer2_out[2044];
    assign layer3_out[2949] = ~(layer2_out[1038] | layer2_out[1039]);
    assign layer3_out[2950] = layer2_out[7104] ^ layer2_out[7105];
    assign layer3_out[2951] = layer2_out[5692] & ~layer2_out[5691];
    assign layer3_out[2952] = 1'b1;
    assign layer3_out[2953] = layer2_out[3243] & layer2_out[3244];
    assign layer3_out[2954] = layer2_out[641];
    assign layer3_out[2955] = layer2_out[750];
    assign layer3_out[2956] = ~layer2_out[3034];
    assign layer3_out[2957] = ~(layer2_out[4065] | layer2_out[4066]);
    assign layer3_out[2958] = layer2_out[4666] & ~layer2_out[4667];
    assign layer3_out[2959] = layer2_out[5235] ^ layer2_out[5236];
    assign layer3_out[2960] = layer2_out[1726];
    assign layer3_out[2961] = ~layer2_out[7237] | layer2_out[7236];
    assign layer3_out[2962] = ~layer2_out[2349];
    assign layer3_out[2963] = ~layer2_out[1099] | layer2_out[1098];
    assign layer3_out[2964] = layer2_out[7802] & ~layer2_out[7801];
    assign layer3_out[2965] = layer2_out[6757] | layer2_out[6758];
    assign layer3_out[2966] = 1'b0;
    assign layer3_out[2967] = ~layer2_out[3563];
    assign layer3_out[2968] = layer2_out[1678];
    assign layer3_out[2969] = layer2_out[3734] & ~layer2_out[3733];
    assign layer3_out[2970] = layer2_out[5677] | layer2_out[5678];
    assign layer3_out[2971] = layer2_out[3906] & ~layer2_out[3907];
    assign layer3_out[2972] = layer2_out[6958] | layer2_out[6959];
    assign layer3_out[2973] = ~(layer2_out[4642] | layer2_out[4643]);
    assign layer3_out[2974] = ~layer2_out[552];
    assign layer3_out[2975] = layer2_out[5083];
    assign layer3_out[2976] = ~(layer2_out[4648] & layer2_out[4649]);
    assign layer3_out[2977] = layer2_out[863] | layer2_out[864];
    assign layer3_out[2978] = layer2_out[7660] & ~layer2_out[7661];
    assign layer3_out[2979] = layer2_out[4743];
    assign layer3_out[2980] = 1'b1;
    assign layer3_out[2981] = ~(layer2_out[542] | layer2_out[543]);
    assign layer3_out[2982] = layer2_out[6441] & layer2_out[6442];
    assign layer3_out[2983] = ~(layer2_out[4979] & layer2_out[4980]);
    assign layer3_out[2984] = ~layer2_out[30] | layer2_out[29];
    assign layer3_out[2985] = ~layer2_out[1120] | layer2_out[1121];
    assign layer3_out[2986] = ~(layer2_out[6770] | layer2_out[6771]);
    assign layer3_out[2987] = ~layer2_out[5840] | layer2_out[5839];
    assign layer3_out[2988] = layer2_out[6963];
    assign layer3_out[2989] = ~layer2_out[4924];
    assign layer3_out[2990] = layer2_out[5282];
    assign layer3_out[2991] = layer2_out[7293] & layer2_out[7294];
    assign layer3_out[2992] = ~layer2_out[1342];
    assign layer3_out[2993] = ~layer2_out[386] | layer2_out[385];
    assign layer3_out[2994] = ~layer2_out[5391] | layer2_out[5390];
    assign layer3_out[2995] = layer2_out[1471];
    assign layer3_out[2996] = layer2_out[1797];
    assign layer3_out[2997] = layer2_out[7486] | layer2_out[7487];
    assign layer3_out[2998] = ~(layer2_out[3423] ^ layer2_out[3424]);
    assign layer3_out[2999] = layer2_out[814] | layer2_out[815];
    assign layer3_out[3000] = layer2_out[5374];
    assign layer3_out[3001] = layer2_out[2340] & ~layer2_out[2341];
    assign layer3_out[3002] = 1'b0;
    assign layer3_out[3003] = layer2_out[5600] ^ layer2_out[5601];
    assign layer3_out[3004] = layer2_out[3343] & ~layer2_out[3342];
    assign layer3_out[3005] = layer2_out[3589];
    assign layer3_out[3006] = 1'b0;
    assign layer3_out[3007] = 1'b1;
    assign layer3_out[3008] = ~layer2_out[247] | layer2_out[248];
    assign layer3_out[3009] = ~layer2_out[7428] | layer2_out[7427];
    assign layer3_out[3010] = ~(layer2_out[7922] & layer2_out[7923]);
    assign layer3_out[3011] = ~(layer2_out[3812] | layer2_out[3813]);
    assign layer3_out[3012] = 1'b1;
    assign layer3_out[3013] = layer2_out[4880];
    assign layer3_out[3014] = ~layer2_out[3386];
    assign layer3_out[3015] = layer2_out[7775];
    assign layer3_out[3016] = ~layer2_out[7817];
    assign layer3_out[3017] = layer2_out[6538] | layer2_out[6539];
    assign layer3_out[3018] = layer2_out[1473];
    assign layer3_out[3019] = layer2_out[1141];
    assign layer3_out[3020] = ~layer2_out[1333];
    assign layer3_out[3021] = layer2_out[6899] | layer2_out[6900];
    assign layer3_out[3022] = ~(layer2_out[817] & layer2_out[818]);
    assign layer3_out[3023] = layer2_out[1524];
    assign layer3_out[3024] = ~layer2_out[1011];
    assign layer3_out[3025] = ~layer2_out[5878];
    assign layer3_out[3026] = ~layer2_out[2243];
    assign layer3_out[3027] = 1'b1;
    assign layer3_out[3028] = ~layer2_out[5847];
    assign layer3_out[3029] = ~layer2_out[1869];
    assign layer3_out[3030] = ~layer2_out[3103] | layer2_out[3102];
    assign layer3_out[3031] = ~(layer2_out[801] ^ layer2_out[802]);
    assign layer3_out[3032] = ~layer2_out[6244] | layer2_out[6245];
    assign layer3_out[3033] = ~(layer2_out[705] | layer2_out[706]);
    assign layer3_out[3034] = ~(layer2_out[4354] | layer2_out[4355]);
    assign layer3_out[3035] = 1'b1;
    assign layer3_out[3036] = ~layer2_out[7691] | layer2_out[7692];
    assign layer3_out[3037] = layer2_out[2016];
    assign layer3_out[3038] = layer2_out[5627];
    assign layer3_out[3039] = layer2_out[3029] ^ layer2_out[3030];
    assign layer3_out[3040] = layer2_out[215] ^ layer2_out[216];
    assign layer3_out[3041] = layer2_out[3127] & ~layer2_out[3128];
    assign layer3_out[3042] = layer2_out[6576] | layer2_out[6577];
    assign layer3_out[3043] = ~(layer2_out[7488] ^ layer2_out[7489]);
    assign layer3_out[3044] = layer2_out[3706];
    assign layer3_out[3045] = layer2_out[6589];
    assign layer3_out[3046] = layer2_out[6030];
    assign layer3_out[3047] = layer2_out[2311] & ~layer2_out[2312];
    assign layer3_out[3048] = ~layer2_out[6042];
    assign layer3_out[3049] = ~layer2_out[752];
    assign layer3_out[3050] = layer2_out[6402] & layer2_out[6403];
    assign layer3_out[3051] = ~(layer2_out[2366] ^ layer2_out[2367]);
    assign layer3_out[3052] = layer2_out[392] & ~layer2_out[393];
    assign layer3_out[3053] = layer2_out[2514];
    assign layer3_out[3054] = 1'b1;
    assign layer3_out[3055] = ~layer2_out[6917] | layer2_out[6916];
    assign layer3_out[3056] = ~(layer2_out[472] | layer2_out[473]);
    assign layer3_out[3057] = layer2_out[560] & ~layer2_out[561];
    assign layer3_out[3058] = ~layer2_out[5695];
    assign layer3_out[3059] = layer2_out[3364] & layer2_out[3365];
    assign layer3_out[3060] = ~layer2_out[68];
    assign layer3_out[3061] = layer2_out[6052] & ~layer2_out[6053];
    assign layer3_out[3062] = ~layer2_out[7894];
    assign layer3_out[3063] = ~layer2_out[2356];
    assign layer3_out[3064] = layer2_out[7533] & ~layer2_out[7532];
    assign layer3_out[3065] = layer2_out[2727] ^ layer2_out[2728];
    assign layer3_out[3066] = layer2_out[7828];
    assign layer3_out[3067] = layer2_out[1182] | layer2_out[1183];
    assign layer3_out[3068] = ~(layer2_out[7408] ^ layer2_out[7409]);
    assign layer3_out[3069] = ~layer2_out[5952];
    assign layer3_out[3070] = ~layer2_out[6429];
    assign layer3_out[3071] = layer2_out[3100];
    assign layer3_out[3072] = layer2_out[3582];
    assign layer3_out[3073] = ~layer2_out[4988];
    assign layer3_out[3074] = layer2_out[7805] ^ layer2_out[7806];
    assign layer3_out[3075] = ~layer2_out[1270];
    assign layer3_out[3076] = layer2_out[4139] | layer2_out[4140];
    assign layer3_out[3077] = layer2_out[5827];
    assign layer3_out[3078] = ~layer2_out[5489];
    assign layer3_out[3079] = ~(layer2_out[6170] & layer2_out[6171]);
    assign layer3_out[3080] = layer2_out[6746] & ~layer2_out[6745];
    assign layer3_out[3081] = layer2_out[228];
    assign layer3_out[3082] = layer2_out[329] ^ layer2_out[330];
    assign layer3_out[3083] = 1'b0;
    assign layer3_out[3084] = ~layer2_out[6091] | layer2_out[6092];
    assign layer3_out[3085] = layer2_out[2055] ^ layer2_out[2056];
    assign layer3_out[3086] = ~layer2_out[2886];
    assign layer3_out[3087] = ~layer2_out[4129] | layer2_out[4128];
    assign layer3_out[3088] = layer2_out[3327];
    assign layer3_out[3089] = ~layer2_out[7867];
    assign layer3_out[3090] = layer2_out[2663];
    assign layer3_out[3091] = ~(layer2_out[5398] | layer2_out[5399]);
    assign layer3_out[3092] = ~(layer2_out[7552] & layer2_out[7553]);
    assign layer3_out[3093] = layer2_out[5377];
    assign layer3_out[3094] = layer2_out[1596] & ~layer2_out[1597];
    assign layer3_out[3095] = ~(layer2_out[2992] | layer2_out[2993]);
    assign layer3_out[3096] = ~(layer2_out[7699] & layer2_out[7700]);
    assign layer3_out[3097] = ~layer2_out[5643];
    assign layer3_out[3098] = layer2_out[3702];
    assign layer3_out[3099] = ~layer2_out[5026];
    assign layer3_out[3100] = 1'b0;
    assign layer3_out[3101] = ~(layer2_out[583] ^ layer2_out[584]);
    assign layer3_out[3102] = layer2_out[4769];
    assign layer3_out[3103] = ~layer2_out[2556];
    assign layer3_out[3104] = 1'b1;
    assign layer3_out[3105] = layer2_out[5938] ^ layer2_out[5939];
    assign layer3_out[3106] = ~layer2_out[2365];
    assign layer3_out[3107] = layer2_out[6839] & ~layer2_out[6840];
    assign layer3_out[3108] = ~layer2_out[7536];
    assign layer3_out[3109] = ~layer2_out[2159] | layer2_out[2158];
    assign layer3_out[3110] = ~layer2_out[7287];
    assign layer3_out[3111] = layer2_out[6138] & ~layer2_out[6137];
    assign layer3_out[3112] = ~layer2_out[3514] | layer2_out[3513];
    assign layer3_out[3113] = 1'b1;
    assign layer3_out[3114] = ~layer2_out[2134];
    assign layer3_out[3115] = ~layer2_out[269];
    assign layer3_out[3116] = layer2_out[7228] ^ layer2_out[7229];
    assign layer3_out[3117] = layer2_out[1925];
    assign layer3_out[3118] = ~layer2_out[6316];
    assign layer3_out[3119] = ~layer2_out[3505] | layer2_out[3504];
    assign layer3_out[3120] = ~layer2_out[1357];
    assign layer3_out[3121] = layer2_out[6143] | layer2_out[6144];
    assign layer3_out[3122] = layer2_out[340] ^ layer2_out[341];
    assign layer3_out[3123] = ~layer2_out[5555];
    assign layer3_out[3124] = ~layer2_out[3180] | layer2_out[3181];
    assign layer3_out[3125] = ~layer2_out[7967];
    assign layer3_out[3126] = layer2_out[6923] & layer2_out[6924];
    assign layer3_out[3127] = layer2_out[1432] | layer2_out[1433];
    assign layer3_out[3128] = layer2_out[5070];
    assign layer3_out[3129] = layer2_out[4470] & layer2_out[4471];
    assign layer3_out[3130] = layer2_out[2363] & ~layer2_out[2364];
    assign layer3_out[3131] = ~layer2_out[422];
    assign layer3_out[3132] = layer2_out[2124] & layer2_out[2125];
    assign layer3_out[3133] = ~layer2_out[2731];
    assign layer3_out[3134] = ~(layer2_out[4525] ^ layer2_out[4526]);
    assign layer3_out[3135] = ~(layer2_out[5968] | layer2_out[5969]);
    assign layer3_out[3136] = layer2_out[193] & ~layer2_out[192];
    assign layer3_out[3137] = layer2_out[6007] | layer2_out[6008];
    assign layer3_out[3138] = layer2_out[3068];
    assign layer3_out[3139] = layer2_out[3769] & ~layer2_out[3770];
    assign layer3_out[3140] = ~layer2_out[6655];
    assign layer3_out[3141] = ~layer2_out[6297];
    assign layer3_out[3142] = layer2_out[3741] & ~layer2_out[3740];
    assign layer3_out[3143] = ~layer2_out[6853];
    assign layer3_out[3144] = layer2_out[5991];
    assign layer3_out[3145] = layer2_out[2715] & ~layer2_out[2714];
    assign layer3_out[3146] = layer2_out[1023] ^ layer2_out[1024];
    assign layer3_out[3147] = ~(layer2_out[1309] & layer2_out[1310]);
    assign layer3_out[3148] = ~layer2_out[1962] | layer2_out[1961];
    assign layer3_out[3149] = ~layer2_out[938] | layer2_out[937];
    assign layer3_out[3150] = 1'b1;
    assign layer3_out[3151] = ~layer2_out[7014] | layer2_out[7015];
    assign layer3_out[3152] = ~layer2_out[7652];
    assign layer3_out[3153] = layer2_out[225] | layer2_out[226];
    assign layer3_out[3154] = ~(layer2_out[5198] | layer2_out[5199]);
    assign layer3_out[3155] = layer2_out[7112] & layer2_out[7113];
    assign layer3_out[3156] = ~(layer2_out[4163] | layer2_out[4164]);
    assign layer3_out[3157] = ~(layer2_out[304] ^ layer2_out[305]);
    assign layer3_out[3158] = ~layer2_out[6640] | layer2_out[6641];
    assign layer3_out[3159] = layer2_out[4773] ^ layer2_out[4774];
    assign layer3_out[3160] = ~(layer2_out[4305] & layer2_out[4306]);
    assign layer3_out[3161] = layer2_out[6583];
    assign layer3_out[3162] = layer2_out[81];
    assign layer3_out[3163] = layer2_out[7470] ^ layer2_out[7471];
    assign layer3_out[3164] = layer2_out[795];
    assign layer3_out[3165] = layer2_out[6484];
    assign layer3_out[3166] = layer2_out[7958] ^ layer2_out[7959];
    assign layer3_out[3167] = ~layer2_out[1189] | layer2_out[1190];
    assign layer3_out[3168] = layer2_out[618] & layer2_out[619];
    assign layer3_out[3169] = ~layer2_out[6082];
    assign layer3_out[3170] = ~layer2_out[3982] | layer2_out[3983];
    assign layer3_out[3171] = ~layer2_out[4311];
    assign layer3_out[3172] = ~(layer2_out[4431] & layer2_out[4432]);
    assign layer3_out[3173] = ~layer2_out[749] | layer2_out[748];
    assign layer3_out[3174] = ~(layer2_out[1759] & layer2_out[1760]);
    assign layer3_out[3175] = ~(layer2_out[6791] | layer2_out[6792]);
    assign layer3_out[3176] = ~layer2_out[5378];
    assign layer3_out[3177] = ~layer2_out[6551] | layer2_out[6552];
    assign layer3_out[3178] = ~layer2_out[6078] | layer2_out[6079];
    assign layer3_out[3179] = ~layer2_out[1268] | layer2_out[1269];
    assign layer3_out[3180] = layer2_out[7001] ^ layer2_out[7002];
    assign layer3_out[3181] = ~layer2_out[2254] | layer2_out[2255];
    assign layer3_out[3182] = layer2_out[4730];
    assign layer3_out[3183] = ~(layer2_out[4073] ^ layer2_out[4074]);
    assign layer3_out[3184] = layer2_out[2362] | layer2_out[2363];
    assign layer3_out[3185] = layer2_out[3810];
    assign layer3_out[3186] = layer2_out[1996];
    assign layer3_out[3187] = ~(layer2_out[2446] ^ layer2_out[2447]);
    assign layer3_out[3188] = ~layer2_out[7753];
    assign layer3_out[3189] = layer2_out[3330];
    assign layer3_out[3190] = layer2_out[3428];
    assign layer3_out[3191] = ~layer2_out[6763];
    assign layer3_out[3192] = layer2_out[7641] & ~layer2_out[7640];
    assign layer3_out[3193] = ~layer2_out[5029] | layer2_out[5028];
    assign layer3_out[3194] = ~layer2_out[4740];
    assign layer3_out[3195] = layer2_out[4344] & layer2_out[4345];
    assign layer3_out[3196] = ~layer2_out[2430] | layer2_out[2431];
    assign layer3_out[3197] = ~layer2_out[1495] | layer2_out[1496];
    assign layer3_out[3198] = ~layer2_out[6570];
    assign layer3_out[3199] = layer2_out[3770] & ~layer2_out[3771];
    assign layer3_out[3200] = ~layer2_out[6800] | layer2_out[6801];
    assign layer3_out[3201] = ~layer2_out[2841] | layer2_out[2840];
    assign layer3_out[3202] = layer2_out[5894] ^ layer2_out[5895];
    assign layer3_out[3203] = layer2_out[535] & ~layer2_out[534];
    assign layer3_out[3204] = layer2_out[245] ^ layer2_out[246];
    assign layer3_out[3205] = ~layer2_out[6616] | layer2_out[6617];
    assign layer3_out[3206] = layer2_out[1538] & layer2_out[1539];
    assign layer3_out[3207] = 1'b1;
    assign layer3_out[3208] = ~layer2_out[4142];
    assign layer3_out[3209] = layer2_out[1702] & ~layer2_out[1701];
    assign layer3_out[3210] = ~layer2_out[7515];
    assign layer3_out[3211] = layer2_out[1370] & layer2_out[1371];
    assign layer3_out[3212] = layer2_out[3000] & layer2_out[3001];
    assign layer3_out[3213] = layer2_out[610] ^ layer2_out[611];
    assign layer3_out[3214] = ~layer2_out[1809] | layer2_out[1808];
    assign layer3_out[3215] = layer2_out[5186];
    assign layer3_out[3216] = layer2_out[6245] & ~layer2_out[6246];
    assign layer3_out[3217] = layer2_out[7046] | layer2_out[7047];
    assign layer3_out[3218] = ~(layer2_out[7524] & layer2_out[7525]);
    assign layer3_out[3219] = layer2_out[6691] & ~layer2_out[6690];
    assign layer3_out[3220] = ~layer2_out[7241] | layer2_out[7242];
    assign layer3_out[3221] = layer2_out[5241];
    assign layer3_out[3222] = layer2_out[7786];
    assign layer3_out[3223] = ~(layer2_out[449] & layer2_out[450]);
    assign layer3_out[3224] = layer2_out[5508] & ~layer2_out[5507];
    assign layer3_out[3225] = layer2_out[5256];
    assign layer3_out[3226] = layer2_out[985] | layer2_out[986];
    assign layer3_out[3227] = ~layer2_out[6136];
    assign layer3_out[3228] = ~layer2_out[1202] | layer2_out[1203];
    assign layer3_out[3229] = ~layer2_out[6644];
    assign layer3_out[3230] = 1'b1;
    assign layer3_out[3231] = ~layer2_out[826];
    assign layer3_out[3232] = layer2_out[364] & layer2_out[365];
    assign layer3_out[3233] = layer2_out[4600];
    assign layer3_out[3234] = layer2_out[455];
    assign layer3_out[3235] = ~layer2_out[3702];
    assign layer3_out[3236] = layer2_out[2371];
    assign layer3_out[3237] = ~(layer2_out[4607] | layer2_out[4608]);
    assign layer3_out[3238] = 1'b0;
    assign layer3_out[3239] = ~layer2_out[6018] | layer2_out[6019];
    assign layer3_out[3240] = ~layer2_out[169] | layer2_out[170];
    assign layer3_out[3241] = ~layer2_out[7998];
    assign layer3_out[3242] = layer2_out[3462] ^ layer2_out[3463];
    assign layer3_out[3243] = layer2_out[7936] & layer2_out[7937];
    assign layer3_out[3244] = layer2_out[322] & ~layer2_out[321];
    assign layer3_out[3245] = layer2_out[6166];
    assign layer3_out[3246] = ~layer2_out[5540];
    assign layer3_out[3247] = 1'b1;
    assign layer3_out[3248] = layer2_out[7231];
    assign layer3_out[3249] = layer2_out[1301] & ~layer2_out[1302];
    assign layer3_out[3250] = ~layer2_out[5494];
    assign layer3_out[3251] = layer2_out[1651];
    assign layer3_out[3252] = layer2_out[4926] & ~layer2_out[4927];
    assign layer3_out[3253] = layer2_out[2699] ^ layer2_out[2700];
    assign layer3_out[3254] = ~(layer2_out[4289] & layer2_out[4290]);
    assign layer3_out[3255] = ~layer2_out[1801];
    assign layer3_out[3256] = layer2_out[3170] & ~layer2_out[3171];
    assign layer3_out[3257] = layer2_out[3495];
    assign layer3_out[3258] = layer2_out[2997] & ~layer2_out[2996];
    assign layer3_out[3259] = layer2_out[161];
    assign layer3_out[3260] = layer2_out[5585] & layer2_out[5586];
    assign layer3_out[3261] = layer2_out[4952];
    assign layer3_out[3262] = ~layer2_out[1199] | layer2_out[1198];
    assign layer3_out[3263] = ~layer2_out[345];
    assign layer3_out[3264] = ~(layer2_out[2931] ^ layer2_out[2932]);
    assign layer3_out[3265] = ~layer2_out[3682];
    assign layer3_out[3266] = ~layer2_out[5188] | layer2_out[5189];
    assign layer3_out[3267] = layer2_out[1401] ^ layer2_out[1402];
    assign layer3_out[3268] = layer2_out[6128] ^ layer2_out[6129];
    assign layer3_out[3269] = ~(layer2_out[3065] ^ layer2_out[3066]);
    assign layer3_out[3270] = ~layer2_out[3349];
    assign layer3_out[3271] = ~layer2_out[7612] | layer2_out[7613];
    assign layer3_out[3272] = layer2_out[5699] & ~layer2_out[5698];
    assign layer3_out[3273] = layer2_out[5097] | layer2_out[5098];
    assign layer3_out[3274] = ~(layer2_out[522] & layer2_out[523]);
    assign layer3_out[3275] = layer2_out[2684] & ~layer2_out[2683];
    assign layer3_out[3276] = ~layer2_out[166] | layer2_out[165];
    assign layer3_out[3277] = layer2_out[2441];
    assign layer3_out[3278] = ~layer2_out[2716];
    assign layer3_out[3279] = layer2_out[7289] & ~layer2_out[7288];
    assign layer3_out[3280] = layer2_out[997] & layer2_out[998];
    assign layer3_out[3281] = layer2_out[1018];
    assign layer3_out[3282] = ~layer2_out[3142];
    assign layer3_out[3283] = ~(layer2_out[4071] & layer2_out[4072]);
    assign layer3_out[3284] = layer2_out[2204];
    assign layer3_out[3285] = layer2_out[4736] | layer2_out[4737];
    assign layer3_out[3286] = layer2_out[6560] & layer2_out[6561];
    assign layer3_out[3287] = layer2_out[3321] | layer2_out[3322];
    assign layer3_out[3288] = layer2_out[5130];
    assign layer3_out[3289] = ~layer2_out[2836] | layer2_out[2835];
    assign layer3_out[3290] = ~layer2_out[6321];
    assign layer3_out[3291] = layer2_out[941] & layer2_out[942];
    assign layer3_out[3292] = ~(layer2_out[2507] & layer2_out[2508]);
    assign layer3_out[3293] = layer2_out[6852] & ~layer2_out[6853];
    assign layer3_out[3294] = ~layer2_out[3744];
    assign layer3_out[3295] = ~(layer2_out[1610] | layer2_out[1611]);
    assign layer3_out[3296] = ~(layer2_out[284] | layer2_out[285]);
    assign layer3_out[3297] = ~(layer2_out[7947] ^ layer2_out[7948]);
    assign layer3_out[3298] = ~layer2_out[475] | layer2_out[474];
    assign layer3_out[3299] = layer2_out[6197] | layer2_out[6198];
    assign layer3_out[3300] = ~(layer2_out[5125] ^ layer2_out[5126]);
    assign layer3_out[3301] = layer2_out[5663] | layer2_out[5664];
    assign layer3_out[3302] = ~layer2_out[5059];
    assign layer3_out[3303] = ~layer2_out[4018] | layer2_out[4019];
    assign layer3_out[3304] = ~(layer2_out[5154] ^ layer2_out[5155]);
    assign layer3_out[3305] = layer2_out[4568];
    assign layer3_out[3306] = layer2_out[6380];
    assign layer3_out[3307] = layer2_out[2042];
    assign layer3_out[3308] = ~layer2_out[5994];
    assign layer3_out[3309] = layer2_out[5313] | layer2_out[5314];
    assign layer3_out[3310] = layer2_out[6391] & ~layer2_out[6392];
    assign layer3_out[3311] = ~layer2_out[7251];
    assign layer3_out[3312] = ~layer2_out[1297];
    assign layer3_out[3313] = layer2_out[2729];
    assign layer3_out[3314] = ~layer2_out[6400];
    assign layer3_out[3315] = ~(layer2_out[341] ^ layer2_out[342]);
    assign layer3_out[3316] = ~layer2_out[4719];
    assign layer3_out[3317] = layer2_out[5032];
    assign layer3_out[3318] = ~(layer2_out[7404] & layer2_out[7405]);
    assign layer3_out[3319] = ~layer2_out[2575];
    assign layer3_out[3320] = ~layer2_out[1140] | layer2_out[1139];
    assign layer3_out[3321] = layer2_out[5426] ^ layer2_out[5427];
    assign layer3_out[3322] = ~layer2_out[402];
    assign layer3_out[3323] = layer2_out[4086] & ~layer2_out[4087];
    assign layer3_out[3324] = layer2_out[3816] | layer2_out[3817];
    assign layer3_out[3325] = 1'b0;
    assign layer3_out[3326] = ~(layer2_out[1331] | layer2_out[1332]);
    assign layer3_out[3327] = ~(layer2_out[2831] | layer2_out[2832]);
    assign layer3_out[3328] = ~layer2_out[5699];
    assign layer3_out[3329] = ~layer2_out[3653];
    assign layer3_out[3330] = layer2_out[2126] | layer2_out[2127];
    assign layer3_out[3331] = layer2_out[7659];
    assign layer3_out[3332] = ~layer2_out[5339];
    assign layer3_out[3333] = layer2_out[491] & ~layer2_out[490];
    assign layer3_out[3334] = layer2_out[1596];
    assign layer3_out[3335] = layer2_out[7925] ^ layer2_out[7926];
    assign layer3_out[3336] = layer2_out[509] & ~layer2_out[508];
    assign layer3_out[3337] = ~layer2_out[5821];
    assign layer3_out[3338] = layer2_out[3026];
    assign layer3_out[3339] = ~layer2_out[3304];
    assign layer3_out[3340] = layer2_out[25] | layer2_out[26];
    assign layer3_out[3341] = layer2_out[83];
    assign layer3_out[3342] = layer2_out[4035] & ~layer2_out[4036];
    assign layer3_out[3343] = layer2_out[3381] | layer2_out[3382];
    assign layer3_out[3344] = layer2_out[1129];
    assign layer3_out[3345] = layer2_out[4725];
    assign layer3_out[3346] = layer2_out[6872] & ~layer2_out[6871];
    assign layer3_out[3347] = ~(layer2_out[1392] ^ layer2_out[1393]);
    assign layer3_out[3348] = layer2_out[5162];
    assign layer3_out[3349] = ~layer2_out[7200];
    assign layer3_out[3350] = layer2_out[1755] ^ layer2_out[1756];
    assign layer3_out[3351] = layer2_out[5856];
    assign layer3_out[3352] = ~(layer2_out[3415] & layer2_out[3416]);
    assign layer3_out[3353] = layer2_out[980] | layer2_out[981];
    assign layer3_out[3354] = layer2_out[1916] & layer2_out[1917];
    assign layer3_out[3355] = layer2_out[6501] | layer2_out[6502];
    assign layer3_out[3356] = layer2_out[4000] & layer2_out[4001];
    assign layer3_out[3357] = layer2_out[6416];
    assign layer3_out[3358] = layer2_out[7592];
    assign layer3_out[3359] = ~layer2_out[5773];
    assign layer3_out[3360] = layer2_out[7815] & ~layer2_out[7814];
    assign layer3_out[3361] = ~layer2_out[4910];
    assign layer3_out[3362] = ~layer2_out[4335] | layer2_out[4336];
    assign layer3_out[3363] = layer2_out[5452] & ~layer2_out[5451];
    assign layer3_out[3364] = ~layer2_out[3745] | layer2_out[3746];
    assign layer3_out[3365] = layer2_out[3290];
    assign layer3_out[3366] = layer2_out[1656];
    assign layer3_out[3367] = ~layer2_out[6435];
    assign layer3_out[3368] = layer2_out[6521] ^ layer2_out[6522];
    assign layer3_out[3369] = layer2_out[6120];
    assign layer3_out[3370] = ~layer2_out[323] | layer2_out[322];
    assign layer3_out[3371] = ~layer2_out[5073] | layer2_out[5074];
    assign layer3_out[3372] = ~(layer2_out[880] ^ layer2_out[881]);
    assign layer3_out[3373] = layer2_out[248] ^ layer2_out[249];
    assign layer3_out[3374] = ~layer2_out[2693];
    assign layer3_out[3375] = ~(layer2_out[5063] | layer2_out[5064]);
    assign layer3_out[3376] = layer2_out[1056] ^ layer2_out[1057];
    assign layer3_out[3377] = ~layer2_out[5457] | layer2_out[5456];
    assign layer3_out[3378] = layer2_out[6696] | layer2_out[6697];
    assign layer3_out[3379] = layer2_out[6153];
    assign layer3_out[3380] = ~(layer2_out[7366] | layer2_out[7367]);
    assign layer3_out[3381] = ~layer2_out[4209] | layer2_out[4208];
    assign layer3_out[3382] = layer2_out[1528] & layer2_out[1529];
    assign layer3_out[3383] = ~(layer2_out[6090] & layer2_out[6091]);
    assign layer3_out[3384] = 1'b0;
    assign layer3_out[3385] = layer2_out[1807] & layer2_out[1808];
    assign layer3_out[3386] = ~layer2_out[6949] | layer2_out[6950];
    assign layer3_out[3387] = ~(layer2_out[182] ^ layer2_out[183]);
    assign layer3_out[3388] = ~layer2_out[754];
    assign layer3_out[3389] = ~layer2_out[2335];
    assign layer3_out[3390] = ~layer2_out[4822] | layer2_out[4821];
    assign layer3_out[3391] = ~layer2_out[635];
    assign layer3_out[3392] = ~layer2_out[666];
    assign layer3_out[3393] = ~layer2_out[5816];
    assign layer3_out[3394] = ~(layer2_out[7088] ^ layer2_out[7089]);
    assign layer3_out[3395] = layer2_out[2012];
    assign layer3_out[3396] = layer2_out[5064] & ~layer2_out[5065];
    assign layer3_out[3397] = layer2_out[3820];
    assign layer3_out[3398] = ~layer2_out[7330];
    assign layer3_out[3399] = ~layer2_out[6239];
    assign layer3_out[3400] = layer2_out[7803];
    assign layer3_out[3401] = ~layer2_out[7295];
    assign layer3_out[3402] = layer2_out[2513] | layer2_out[2514];
    assign layer3_out[3403] = ~layer2_out[171];
    assign layer3_out[3404] = ~layer2_out[4755];
    assign layer3_out[3405] = layer2_out[4864] & layer2_out[4865];
    assign layer3_out[3406] = layer2_out[5804];
    assign layer3_out[3407] = ~layer2_out[5632];
    assign layer3_out[3408] = layer2_out[6009];
    assign layer3_out[3409] = layer2_out[7720];
    assign layer3_out[3410] = ~(layer2_out[1116] ^ layer2_out[1117]);
    assign layer3_out[3411] = layer2_out[79] & ~layer2_out[80];
    assign layer3_out[3412] = ~layer2_out[1893];
    assign layer3_out[3413] = ~layer2_out[3508];
    assign layer3_out[3414] = ~(layer2_out[798] ^ layer2_out[799]);
    assign layer3_out[3415] = ~(layer2_out[3666] | layer2_out[3667]);
    assign layer3_out[3416] = ~layer2_out[4081] | layer2_out[4082];
    assign layer3_out[3417] = layer2_out[1755];
    assign layer3_out[3418] = ~layer2_out[840] | layer2_out[839];
    assign layer3_out[3419] = layer2_out[6316] & ~layer2_out[6315];
    assign layer3_out[3420] = ~layer2_out[1719];
    assign layer3_out[3421] = ~layer2_out[7825];
    assign layer3_out[3422] = ~layer2_out[5458] | layer2_out[5459];
    assign layer3_out[3423] = ~layer2_out[6585];
    assign layer3_out[3424] = layer2_out[6922] & ~layer2_out[6921];
    assign layer3_out[3425] = layer2_out[5724];
    assign layer3_out[3426] = ~(layer2_out[3946] | layer2_out[3947]);
    assign layer3_out[3427] = ~(layer2_out[5102] ^ layer2_out[5103]);
    assign layer3_out[3428] = layer2_out[7744] & ~layer2_out[7743];
    assign layer3_out[3429] = ~layer2_out[5143] | layer2_out[5144];
    assign layer3_out[3430] = ~layer2_out[2764] | layer2_out[2765];
    assign layer3_out[3431] = 1'b0;
    assign layer3_out[3432] = ~layer2_out[5562];
    assign layer3_out[3433] = ~layer2_out[4663];
    assign layer3_out[3434] = layer2_out[6992];
    assign layer3_out[3435] = layer2_out[4557] ^ layer2_out[4558];
    assign layer3_out[3436] = layer2_out[7664];
    assign layer3_out[3437] = ~layer2_out[5430];
    assign layer3_out[3438] = ~layer2_out[2217];
    assign layer3_out[3439] = ~(layer2_out[1454] & layer2_out[1455]);
    assign layer3_out[3440] = layer2_out[5802] & layer2_out[5803];
    assign layer3_out[3441] = ~(layer2_out[1707] ^ layer2_out[1708]);
    assign layer3_out[3442] = layer2_out[2427];
    assign layer3_out[3443] = ~layer2_out[4144] | layer2_out[4143];
    assign layer3_out[3444] = ~(layer2_out[1978] | layer2_out[1979]);
    assign layer3_out[3445] = ~layer2_out[120] | layer2_out[119];
    assign layer3_out[3446] = ~(layer2_out[2588] | layer2_out[2589]);
    assign layer3_out[3447] = ~(layer2_out[7195] & layer2_out[7196]);
    assign layer3_out[3448] = ~layer2_out[6867] | layer2_out[6866];
    assign layer3_out[3449] = layer2_out[5250] | layer2_out[5251];
    assign layer3_out[3450] = ~(layer2_out[2583] & layer2_out[2584]);
    assign layer3_out[3451] = layer2_out[629] & ~layer2_out[630];
    assign layer3_out[3452] = layer2_out[6053] ^ layer2_out[6054];
    assign layer3_out[3453] = layer2_out[2120] & layer2_out[2121];
    assign layer3_out[3454] = 1'b0;
    assign layer3_out[3455] = ~layer2_out[7892];
    assign layer3_out[3456] = layer2_out[128] & ~layer2_out[129];
    assign layer3_out[3457] = layer2_out[7500] & layer2_out[7501];
    assign layer3_out[3458] = ~layer2_out[5623] | layer2_out[5622];
    assign layer3_out[3459] = layer2_out[1990];
    assign layer3_out[3460] = layer2_out[2982] | layer2_out[2983];
    assign layer3_out[3461] = ~layer2_out[5219] | layer2_out[5220];
    assign layer3_out[3462] = layer2_out[6989];
    assign layer3_out[3463] = layer2_out[4453] & ~layer2_out[4452];
    assign layer3_out[3464] = ~(layer2_out[5356] & layer2_out[5357]);
    assign layer3_out[3465] = 1'b0;
    assign layer3_out[3466] = layer2_out[4627] & ~layer2_out[4626];
    assign layer3_out[3467] = ~layer2_out[7657];
    assign layer3_out[3468] = layer2_out[600] | layer2_out[601];
    assign layer3_out[3469] = layer2_out[4933] & layer2_out[4934];
    assign layer3_out[3470] = ~layer2_out[142];
    assign layer3_out[3471] = layer2_out[4794] ^ layer2_out[4795];
    assign layer3_out[3472] = ~layer2_out[3913] | layer2_out[3912];
    assign layer3_out[3473] = layer2_out[1037];
    assign layer3_out[3474] = ~layer2_out[504];
    assign layer3_out[3475] = ~layer2_out[1430];
    assign layer3_out[3476] = ~layer2_out[7433] | layer2_out[7434];
    assign layer3_out[3477] = ~(layer2_out[4301] | layer2_out[4302]);
    assign layer3_out[3478] = ~layer2_out[2281];
    assign layer3_out[3479] = layer2_out[2682] ^ layer2_out[2683];
    assign layer3_out[3480] = layer2_out[7228];
    assign layer3_out[3481] = layer2_out[7301] ^ layer2_out[7302];
    assign layer3_out[3482] = 1'b0;
    assign layer3_out[3483] = layer2_out[3843];
    assign layer3_out[3484] = ~layer2_out[4311];
    assign layer3_out[3485] = 1'b1;
    assign layer3_out[3486] = layer2_out[3767] | layer2_out[3768];
    assign layer3_out[3487] = ~layer2_out[7027];
    assign layer3_out[3488] = layer2_out[1599] ^ layer2_out[1600];
    assign layer3_out[3489] = ~layer2_out[2856];
    assign layer3_out[3490] = ~(layer2_out[6934] & layer2_out[6935]);
    assign layer3_out[3491] = layer2_out[5289];
    assign layer3_out[3492] = layer2_out[7161] & ~layer2_out[7162];
    assign layer3_out[3493] = ~layer2_out[4480];
    assign layer3_out[3494] = ~layer2_out[3711];
    assign layer3_out[3495] = layer2_out[2237] | layer2_out[2238];
    assign layer3_out[3496] = 1'b1;
    assign layer3_out[3497] = 1'b0;
    assign layer3_out[3498] = ~layer2_out[2318];
    assign layer3_out[3499] = layer2_out[7871];
    assign layer3_out[3500] = layer2_out[6643] & ~layer2_out[6644];
    assign layer3_out[3501] = layer2_out[5818] & layer2_out[5819];
    assign layer3_out[3502] = ~layer2_out[297];
    assign layer3_out[3503] = ~layer2_out[4063];
    assign layer3_out[3504] = layer2_out[5372];
    assign layer3_out[3505] = layer2_out[5720];
    assign layer3_out[3506] = layer2_out[7226];
    assign layer3_out[3507] = layer2_out[2910] & layer2_out[2911];
    assign layer3_out[3508] = ~layer2_out[6084];
    assign layer3_out[3509] = layer2_out[363];
    assign layer3_out[3510] = layer2_out[7429] & ~layer2_out[7430];
    assign layer3_out[3511] = layer2_out[5399] | layer2_out[5400];
    assign layer3_out[3512] = layer2_out[2163] | layer2_out[2164];
    assign layer3_out[3513] = layer2_out[725] & ~layer2_out[724];
    assign layer3_out[3514] = layer2_out[4415];
    assign layer3_out[3515] = layer2_out[5614] & layer2_out[5615];
    assign layer3_out[3516] = layer2_out[1176];
    assign layer3_out[3517] = layer2_out[6061] ^ layer2_out[6062];
    assign layer3_out[3518] = layer2_out[7193];
    assign layer3_out[3519] = ~layer2_out[1006];
    assign layer3_out[3520] = ~layer2_out[1771];
    assign layer3_out[3521] = layer2_out[2309] & layer2_out[2310];
    assign layer3_out[3522] = ~layer2_out[3433];
    assign layer3_out[3523] = layer2_out[1028] & ~layer2_out[1027];
    assign layer3_out[3524] = ~(layer2_out[7568] ^ layer2_out[7569]);
    assign layer3_out[3525] = layer2_out[2639] ^ layer2_out[2640];
    assign layer3_out[3526] = ~layer2_out[2808];
    assign layer3_out[3527] = layer2_out[4432] | layer2_out[4433];
    assign layer3_out[3528] = layer2_out[92];
    assign layer3_out[3529] = layer2_out[4076];
    assign layer3_out[3530] = ~layer2_out[7332] | layer2_out[7331];
    assign layer3_out[3531] = layer2_out[2374];
    assign layer3_out[3532] = layer2_out[5362];
    assign layer3_out[3533] = ~layer2_out[5222] | layer2_out[5223];
    assign layer3_out[3534] = layer2_out[1551] | layer2_out[1552];
    assign layer3_out[3535] = ~layer2_out[737] | layer2_out[736];
    assign layer3_out[3536] = layer2_out[1429];
    assign layer3_out[3537] = ~layer2_out[1957] | layer2_out[1956];
    assign layer3_out[3538] = layer2_out[3944];
    assign layer3_out[3539] = layer2_out[4005];
    assign layer3_out[3540] = layer2_out[1552] & ~layer2_out[1553];
    assign layer3_out[3541] = layer2_out[2655] | layer2_out[2656];
    assign layer3_out[3542] = layer2_out[4856];
    assign layer3_out[3543] = ~(layer2_out[2780] & layer2_out[2781]);
    assign layer3_out[3544] = ~(layer2_out[1670] | layer2_out[1671]);
    assign layer3_out[3545] = ~layer2_out[2816];
    assign layer3_out[3546] = ~(layer2_out[7157] | layer2_out[7158]);
    assign layer3_out[3547] = layer2_out[1738] | layer2_out[1739];
    assign layer3_out[3548] = layer2_out[4423] & layer2_out[4424];
    assign layer3_out[3549] = ~layer2_out[7739];
    assign layer3_out[3550] = ~layer2_out[7901];
    assign layer3_out[3551] = ~(layer2_out[6502] & layer2_out[6503]);
    assign layer3_out[3552] = ~layer2_out[6161];
    assign layer3_out[3553] = ~layer2_out[5749] | layer2_out[5750];
    assign layer3_out[3554] = ~layer2_out[1480];
    assign layer3_out[3555] = layer2_out[1404] ^ layer2_out[1405];
    assign layer3_out[3556] = layer2_out[898] & layer2_out[899];
    assign layer3_out[3557] = ~layer2_out[6742];
    assign layer3_out[3558] = layer2_out[7279] & ~layer2_out[7278];
    assign layer3_out[3559] = ~layer2_out[4407] | layer2_out[4406];
    assign layer3_out[3560] = ~layer2_out[3617] | layer2_out[3618];
    assign layer3_out[3561] = layer2_out[6448] & layer2_out[6449];
    assign layer3_out[3562] = ~(layer2_out[4836] & layer2_out[4837]);
    assign layer3_out[3563] = layer2_out[6485] ^ layer2_out[6486];
    assign layer3_out[3564] = ~layer2_out[4766] | layer2_out[4765];
    assign layer3_out[3565] = ~layer2_out[1002] | layer2_out[1001];
    assign layer3_out[3566] = ~layer2_out[7504];
    assign layer3_out[3567] = ~(layer2_out[7377] | layer2_out[7378]);
    assign layer3_out[3568] = layer2_out[4776] ^ layer2_out[4777];
    assign layer3_out[3569] = ~(layer2_out[2883] & layer2_out[2884]);
    assign layer3_out[3570] = ~(layer2_out[7646] ^ layer2_out[7647]);
    assign layer3_out[3571] = ~layer2_out[3037] | layer2_out[3036];
    assign layer3_out[3572] = ~layer2_out[1115] | layer2_out[1116];
    assign layer3_out[3573] = ~(layer2_out[6148] & layer2_out[6149]);
    assign layer3_out[3574] = layer2_out[407] | layer2_out[408];
    assign layer3_out[3575] = layer2_out[267] & ~layer2_out[268];
    assign layer3_out[3576] = layer2_out[5866] & ~layer2_out[5865];
    assign layer3_out[3577] = ~layer2_out[644] | layer2_out[645];
    assign layer3_out[3578] = ~layer2_out[3];
    assign layer3_out[3579] = ~(layer2_out[273] ^ layer2_out[274]);
    assign layer3_out[3580] = layer2_out[6922] ^ layer2_out[6923];
    assign layer3_out[3581] = layer2_out[6962];
    assign layer3_out[3582] = layer2_out[755] | layer2_out[756];
    assign layer3_out[3583] = ~(layer2_out[2156] ^ layer2_out[2157]);
    assign layer3_out[3584] = 1'b1;
    assign layer3_out[3585] = ~layer2_out[4491];
    assign layer3_out[3586] = ~layer2_out[3826] | layer2_out[3827];
    assign layer3_out[3587] = layer2_out[5843] ^ layer2_out[5844];
    assign layer3_out[3588] = layer2_out[6128];
    assign layer3_out[3589] = layer2_out[2018] & ~layer2_out[2019];
    assign layer3_out[3590] = ~layer2_out[75];
    assign layer3_out[3591] = layer2_out[5899];
    assign layer3_out[3592] = ~layer2_out[7848] | layer2_out[7847];
    assign layer3_out[3593] = layer2_out[6854] & ~layer2_out[6855];
    assign layer3_out[3594] = ~layer2_out[5312];
    assign layer3_out[3595] = ~layer2_out[555] | layer2_out[556];
    assign layer3_out[3596] = layer2_out[1917] & ~layer2_out[1918];
    assign layer3_out[3597] = layer2_out[7056] & ~layer2_out[7057];
    assign layer3_out[3598] = ~layer2_out[899];
    assign layer3_out[3599] = ~(layer2_out[381] ^ layer2_out[382]);
    assign layer3_out[3600] = layer2_out[256];
    assign layer3_out[3601] = 1'b1;
    assign layer3_out[3602] = layer2_out[6236] | layer2_out[6237];
    assign layer3_out[3603] = ~(layer2_out[1071] ^ layer2_out[1072]);
    assign layer3_out[3604] = layer2_out[6713];
    assign layer3_out[3605] = ~layer2_out[486] | layer2_out[485];
    assign layer3_out[3606] = ~layer2_out[2380] | layer2_out[2379];
    assign layer3_out[3607] = ~layer2_out[3436] | layer2_out[3435];
    assign layer3_out[3608] = ~(layer2_out[403] & layer2_out[404]);
    assign layer3_out[3609] = ~layer2_out[1684];
    assign layer3_out[3610] = ~layer2_out[1096] | layer2_out[1095];
    assign layer3_out[3611] = layer2_out[7050];
    assign layer3_out[3612] = ~layer2_out[7463];
    assign layer3_out[3613] = layer2_out[1076];
    assign layer3_out[3614] = layer2_out[5056] | layer2_out[5057];
    assign layer3_out[3615] = layer2_out[1292] & ~layer2_out[1293];
    assign layer3_out[3616] = layer2_out[1505] & ~layer2_out[1504];
    assign layer3_out[3617] = ~layer2_out[1843];
    assign layer3_out[3618] = ~(layer2_out[3856] ^ layer2_out[3857]);
    assign layer3_out[3619] = layer2_out[3337];
    assign layer3_out[3620] = layer2_out[5873];
    assign layer3_out[3621] = ~layer2_out[5640];
    assign layer3_out[3622] = layer2_out[2139] ^ layer2_out[2140];
    assign layer3_out[3623] = ~layer2_out[6254] | layer2_out[6255];
    assign layer3_out[3624] = layer2_out[2225];
    assign layer3_out[3625] = layer2_out[1814];
    assign layer3_out[3626] = ~layer2_out[1985] | layer2_out[1986];
    assign layer3_out[3627] = layer2_out[2399] & ~layer2_out[2398];
    assign layer3_out[3628] = ~layer2_out[6930] | layer2_out[6931];
    assign layer3_out[3629] = ~(layer2_out[6567] ^ layer2_out[6568]);
    assign layer3_out[3630] = ~layer2_out[4904];
    assign layer3_out[3631] = layer2_out[6693] ^ layer2_out[6694];
    assign layer3_out[3632] = layer2_out[6262] & ~layer2_out[6263];
    assign layer3_out[3633] = layer2_out[7977] ^ layer2_out[7978];
    assign layer3_out[3634] = layer2_out[2431] | layer2_out[2432];
    assign layer3_out[3635] = ~layer2_out[6428] | layer2_out[6427];
    assign layer3_out[3636] = ~(layer2_out[3349] | layer2_out[3350]);
    assign layer3_out[3637] = ~layer2_out[4359];
    assign layer3_out[3638] = layer2_out[3308] & ~layer2_out[3309];
    assign layer3_out[3639] = layer2_out[154];
    assign layer3_out[3640] = ~layer2_out[7225];
    assign layer3_out[3641] = ~(layer2_out[1525] | layer2_out[1526]);
    assign layer3_out[3642] = layer2_out[4198] | layer2_out[4199];
    assign layer3_out[3643] = layer2_out[2894] & ~layer2_out[2893];
    assign layer3_out[3644] = layer2_out[4742] & ~layer2_out[4741];
    assign layer3_out[3645] = layer2_out[7383] & ~layer2_out[7384];
    assign layer3_out[3646] = layer2_out[6225];
    assign layer3_out[3647] = ~(layer2_out[766] ^ layer2_out[767]);
    assign layer3_out[3648] = ~(layer2_out[7430] | layer2_out[7431]);
    assign layer3_out[3649] = 1'b0;
    assign layer3_out[3650] = ~layer2_out[3249];
    assign layer3_out[3651] = layer2_out[5669];
    assign layer3_out[3652] = 1'b0;
    assign layer3_out[3653] = ~layer2_out[2732] | layer2_out[2733];
    assign layer3_out[3654] = layer2_out[3565] | layer2_out[3566];
    assign layer3_out[3655] = layer2_out[7565];
    assign layer3_out[3656] = layer2_out[1751] | layer2_out[1752];
    assign layer3_out[3657] = ~layer2_out[7375] | layer2_out[7376];
    assign layer3_out[3658] = ~layer2_out[5638] | layer2_out[5639];
    assign layer3_out[3659] = layer2_out[7725] | layer2_out[7726];
    assign layer3_out[3660] = layer2_out[4850] ^ layer2_out[4851];
    assign layer3_out[3661] = ~(layer2_out[4460] & layer2_out[4461]);
    assign layer3_out[3662] = layer2_out[164] & layer2_out[165];
    assign layer3_out[3663] = layer2_out[1615] | layer2_out[1616];
    assign layer3_out[3664] = ~(layer2_out[837] ^ layer2_out[838]);
    assign layer3_out[3665] = layer2_out[93] | layer2_out[94];
    assign layer3_out[3666] = ~(layer2_out[7984] & layer2_out[7985]);
    assign layer3_out[3667] = layer2_out[5214];
    assign layer3_out[3668] = layer2_out[7712] & layer2_out[7713];
    assign layer3_out[3669] = layer2_out[761];
    assign layer3_out[3670] = layer2_out[6425] & ~layer2_out[6424];
    assign layer3_out[3671] = ~(layer2_out[4387] ^ layer2_out[4388]);
    assign layer3_out[3672] = ~layer2_out[6156] | layer2_out[6157];
    assign layer3_out[3673] = layer2_out[2770];
    assign layer3_out[3674] = ~(layer2_out[2326] ^ layer2_out[2327]);
    assign layer3_out[3675] = layer2_out[6876] & ~layer2_out[6875];
    assign layer3_out[3676] = layer2_out[2868] & ~layer2_out[2867];
    assign layer3_out[3677] = layer2_out[7402] & layer2_out[7403];
    assign layer3_out[3678] = layer2_out[6010] & ~layer2_out[6009];
    assign layer3_out[3679] = layer2_out[523] ^ layer2_out[524];
    assign layer3_out[3680] = ~layer2_out[5280];
    assign layer3_out[3681] = ~layer2_out[5436];
    assign layer3_out[3682] = ~layer2_out[5929];
    assign layer3_out[3683] = layer2_out[7951] & layer2_out[7952];
    assign layer3_out[3684] = ~layer2_out[7991];
    assign layer3_out[3685] = ~layer2_out[4457];
    assign layer3_out[3686] = ~layer2_out[3368] | layer2_out[3369];
    assign layer3_out[3687] = layer2_out[4671] & layer2_out[4672];
    assign layer3_out[3688] = ~(layer2_out[6728] & layer2_out[6729]);
    assign layer3_out[3689] = ~(layer2_out[2224] | layer2_out[2225]);
    assign layer3_out[3690] = layer2_out[5489] & layer2_out[5490];
    assign layer3_out[3691] = ~layer2_out[3570];
    assign layer3_out[3692] = ~(layer2_out[7207] | layer2_out[7208]);
    assign layer3_out[3693] = ~layer2_out[3434] | layer2_out[3433];
    assign layer3_out[3694] = ~layer2_out[4503];
    assign layer3_out[3695] = layer2_out[6426];
    assign layer3_out[3696] = layer2_out[2250] | layer2_out[2251];
    assign layer3_out[3697] = ~layer2_out[1108];
    assign layer3_out[3698] = ~(layer2_out[1508] | layer2_out[1509]);
    assign layer3_out[3699] = layer2_out[7898];
    assign layer3_out[3700] = ~layer2_out[2028];
    assign layer3_out[3701] = layer2_out[1076] & ~layer2_out[1075];
    assign layer3_out[3702] = layer2_out[3854];
    assign layer3_out[3703] = ~layer2_out[1257] | layer2_out[1258];
    assign layer3_out[3704] = ~layer2_out[668] | layer2_out[667];
    assign layer3_out[3705] = ~layer2_out[7258];
    assign layer3_out[3706] = ~(layer2_out[2822] & layer2_out[2823]);
    assign layer3_out[3707] = layer2_out[1864];
    assign layer3_out[3708] = layer2_out[1688] ^ layer2_out[1689];
    assign layer3_out[3709] = ~layer2_out[5000];
    assign layer3_out[3710] = layer2_out[1426];
    assign layer3_out[3711] = layer2_out[5664] ^ layer2_out[5665];
    assign layer3_out[3712] = ~(layer2_out[2079] | layer2_out[2080]);
    assign layer3_out[3713] = layer2_out[7343] & layer2_out[7344];
    assign layer3_out[3714] = layer2_out[6612] & ~layer2_out[6613];
    assign layer3_out[3715] = layer2_out[3871] & ~layer2_out[3872];
    assign layer3_out[3716] = ~layer2_out[2326] | layer2_out[2325];
    assign layer3_out[3717] = ~layer2_out[7775] | layer2_out[7776];
    assign layer3_out[3718] = layer2_out[7025] & layer2_out[7026];
    assign layer3_out[3719] = ~layer2_out[3252];
    assign layer3_out[3720] = ~(layer2_out[7066] | layer2_out[7067]);
    assign layer3_out[3721] = layer2_out[476] & ~layer2_out[477];
    assign layer3_out[3722] = ~layer2_out[7027];
    assign layer3_out[3723] = layer2_out[2660];
    assign layer3_out[3724] = ~layer2_out[5569] | layer2_out[5568];
    assign layer3_out[3725] = layer2_out[3635] & ~layer2_out[3636];
    assign layer3_out[3726] = layer2_out[1590];
    assign layer3_out[3727] = ~layer2_out[2266];
    assign layer3_out[3728] = layer2_out[5433];
    assign layer3_out[3729] = ~layer2_out[1606] | layer2_out[1605];
    assign layer3_out[3730] = layer2_out[4935];
    assign layer3_out[3731] = layer2_out[1107];
    assign layer3_out[3732] = ~layer2_out[5564];
    assign layer3_out[3733] = ~layer2_out[4229] | layer2_out[4228];
    assign layer3_out[3734] = ~(layer2_out[1622] | layer2_out[1623]);
    assign layer3_out[3735] = layer2_out[1830] | layer2_out[1831];
    assign layer3_out[3736] = ~layer2_out[401];
    assign layer3_out[3737] = layer2_out[2708] ^ layer2_out[2709];
    assign layer3_out[3738] = ~layer2_out[4929];
    assign layer3_out[3739] = ~layer2_out[6590] | layer2_out[6589];
    assign layer3_out[3740] = layer2_out[1491];
    assign layer3_out[3741] = 1'b1;
    assign layer3_out[3742] = layer2_out[5039] ^ layer2_out[5040];
    assign layer3_out[3743] = layer2_out[4487];
    assign layer3_out[3744] = layer2_out[7555] & layer2_out[7556];
    assign layer3_out[3745] = layer2_out[334] & ~layer2_out[333];
    assign layer3_out[3746] = layer2_out[7045];
    assign layer3_out[3747] = layer2_out[4410] & ~layer2_out[4411];
    assign layer3_out[3748] = layer2_out[5182];
    assign layer3_out[3749] = layer2_out[4861];
    assign layer3_out[3750] = ~layer2_out[2050] | layer2_out[2051];
    assign layer3_out[3751] = layer2_out[2132];
    assign layer3_out[3752] = layer2_out[6905] | layer2_out[6906];
    assign layer3_out[3753] = layer2_out[4544] & ~layer2_out[4545];
    assign layer3_out[3754] = ~layer2_out[5067];
    assign layer3_out[3755] = layer2_out[5858];
    assign layer3_out[3756] = layer2_out[5701];
    assign layer3_out[3757] = layer2_out[1017] & layer2_out[1018];
    assign layer3_out[3758] = layer2_out[7672] & layer2_out[7673];
    assign layer3_out[3759] = ~(layer2_out[2045] ^ layer2_out[2046]);
    assign layer3_out[3760] = ~layer2_out[6903] | layer2_out[6902];
    assign layer3_out[3761] = layer2_out[184];
    assign layer3_out[3762] = layer2_out[6729] & ~layer2_out[6730];
    assign layer3_out[3763] = layer2_out[2181] ^ layer2_out[2182];
    assign layer3_out[3764] = ~layer2_out[2209];
    assign layer3_out[3765] = layer2_out[3554] & layer2_out[3555];
    assign layer3_out[3766] = layer2_out[6303];
    assign layer3_out[3767] = layer2_out[2466];
    assign layer3_out[3768] = ~layer2_out[6547];
    assign layer3_out[3769] = layer2_out[1548];
    assign layer3_out[3770] = layer2_out[4595] & layer2_out[4596];
    assign layer3_out[3771] = ~layer2_out[2186];
    assign layer3_out[3772] = ~layer2_out[4265];
    assign layer3_out[3773] = ~layer2_out[2485];
    assign layer3_out[3774] = 1'b0;
    assign layer3_out[3775] = layer2_out[1867];
    assign layer3_out[3776] = ~layer2_out[6776] | layer2_out[6777];
    assign layer3_out[3777] = ~layer2_out[4841] | layer2_out[4840];
    assign layer3_out[3778] = layer2_out[2654] & ~layer2_out[2653];
    assign layer3_out[3779] = ~(layer2_out[1021] ^ layer2_out[1022]);
    assign layer3_out[3780] = layer2_out[4366];
    assign layer3_out[3781] = ~(layer2_out[721] & layer2_out[722]);
    assign layer3_out[3782] = ~layer2_out[2830] | layer2_out[2829];
    assign layer3_out[3783] = layer2_out[2486] ^ layer2_out[2487];
    assign layer3_out[3784] = layer2_out[57];
    assign layer3_out[3785] = ~layer2_out[1306];
    assign layer3_out[3786] = ~layer2_out[3283] | layer2_out[3282];
    assign layer3_out[3787] = ~(layer2_out[3720] ^ layer2_out[3721]);
    assign layer3_out[3788] = ~layer2_out[2562];
    assign layer3_out[3789] = layer2_out[1905] & layer2_out[1906];
    assign layer3_out[3790] = ~layer2_out[3089];
    assign layer3_out[3791] = ~layer2_out[6455];
    assign layer3_out[3792] = layer2_out[5674];
    assign layer3_out[3793] = layer2_out[6204];
    assign layer3_out[3794] = ~layer2_out[1327] | layer2_out[1326];
    assign layer3_out[3795] = layer2_out[1424];
    assign layer3_out[3796] = ~layer2_out[5121] | layer2_out[5122];
    assign layer3_out[3797] = ~layer2_out[1041] | layer2_out[1040];
    assign layer3_out[3798] = layer2_out[4295] & ~layer2_out[4296];
    assign layer3_out[3799] = layer2_out[6712] | layer2_out[6713];
    assign layer3_out[3800] = ~layer2_out[4279] | layer2_out[4280];
    assign layer3_out[3801] = layer2_out[7670];
    assign layer3_out[3802] = ~layer2_out[7358] | layer2_out[7357];
    assign layer3_out[3803] = ~layer2_out[7932];
    assign layer3_out[3804] = ~layer2_out[3537];
    assign layer3_out[3805] = ~layer2_out[709] | layer2_out[708];
    assign layer3_out[3806] = ~layer2_out[1271];
    assign layer3_out[3807] = ~(layer2_out[4739] | layer2_out[4740]);
    assign layer3_out[3808] = ~layer2_out[4263];
    assign layer3_out[3809] = layer2_out[7114];
    assign layer3_out[3810] = layer2_out[4644] ^ layer2_out[4645];
    assign layer3_out[3811] = ~(layer2_out[1587] | layer2_out[1588]);
    assign layer3_out[3812] = layer2_out[1197];
    assign layer3_out[3813] = layer2_out[802] & ~layer2_out[803];
    assign layer3_out[3814] = layer2_out[2572];
    assign layer3_out[3815] = layer2_out[6948] & ~layer2_out[6947];
    assign layer3_out[3816] = layer2_out[6762];
    assign layer3_out[3817] = layer2_out[5886];
    assign layer3_out[3818] = layer2_out[4093] | layer2_out[4094];
    assign layer3_out[3819] = layer2_out[1046] & layer2_out[1047];
    assign layer3_out[3820] = layer2_out[3352] & ~layer2_out[3351];
    assign layer3_out[3821] = ~(layer2_out[2680] ^ layer2_out[2681]);
    assign layer3_out[3822] = layer2_out[6954] | layer2_out[6955];
    assign layer3_out[3823] = layer2_out[1221] ^ layer2_out[1222];
    assign layer3_out[3824] = ~layer2_out[5110] | layer2_out[5109];
    assign layer3_out[3825] = ~layer2_out[2263];
    assign layer3_out[3826] = layer2_out[5621] & layer2_out[5622];
    assign layer3_out[3827] = ~layer2_out[7974];
    assign layer3_out[3828] = ~layer2_out[3690];
    assign layer3_out[3829] = ~layer2_out[3093];
    assign layer3_out[3830] = ~layer2_out[6390];
    assign layer3_out[3831] = layer2_out[3852];
    assign layer3_out[3832] = layer2_out[4306];
    assign layer3_out[3833] = ~layer2_out[3849];
    assign layer3_out[3834] = ~(layer2_out[3729] | layer2_out[3730]);
    assign layer3_out[3835] = ~(layer2_out[1083] ^ layer2_out[1084]);
    assign layer3_out[3836] = layer2_out[5539];
    assign layer3_out[3837] = layer2_out[2454] & ~layer2_out[2455];
    assign layer3_out[3838] = layer2_out[5504];
    assign layer3_out[3839] = ~layer2_out[5701] | layer2_out[5702];
    assign layer3_out[3840] = layer2_out[907];
    assign layer3_out[3841] = 1'b0;
    assign layer3_out[3842] = layer2_out[2347] ^ layer2_out[2348];
    assign layer3_out[3843] = ~layer2_out[3157];
    assign layer3_out[3844] = layer2_out[6021];
    assign layer3_out[3845] = layer2_out[7635] & ~layer2_out[7636];
    assign layer3_out[3846] = ~(layer2_out[5545] | layer2_out[5546]);
    assign layer3_out[3847] = ~layer2_out[7765] | layer2_out[7766];
    assign layer3_out[3848] = layer2_out[5148] & ~layer2_out[5149];
    assign layer3_out[3849] = layer2_out[5662] & ~layer2_out[5663];
    assign layer3_out[3850] = ~(layer2_out[2768] & layer2_out[2769]);
    assign layer3_out[3851] = layer2_out[6942] & ~layer2_out[6943];
    assign layer3_out[3852] = layer2_out[3602] | layer2_out[3603];
    assign layer3_out[3853] = ~(layer2_out[2586] ^ layer2_out[2587]);
    assign layer3_out[3854] = layer2_out[778] ^ layer2_out[779];
    assign layer3_out[3855] = layer2_out[3242] & layer2_out[3243];
    assign layer3_out[3856] = layer2_out[711] | layer2_out[712];
    assign layer3_out[3857] = layer2_out[5589];
    assign layer3_out[3858] = ~layer2_out[1851] | layer2_out[1850];
    assign layer3_out[3859] = layer2_out[2456] & ~layer2_out[2455];
    assign layer3_out[3860] = layer2_out[3561] & ~layer2_out[3560];
    assign layer3_out[3861] = layer2_out[6328] & ~layer2_out[6327];
    assign layer3_out[3862] = ~(layer2_out[1025] ^ layer2_out[1026]);
    assign layer3_out[3863] = ~layer2_out[6301];
    assign layer3_out[3864] = layer2_out[4890] | layer2_out[4891];
    assign layer3_out[3865] = ~layer2_out[5717] | layer2_out[5718];
    assign layer3_out[3866] = layer2_out[5614] & ~layer2_out[5613];
    assign layer3_out[3867] = ~layer2_out[5747] | layer2_out[5746];
    assign layer3_out[3868] = ~layer2_out[2274] | layer2_out[2275];
    assign layer3_out[3869] = ~layer2_out[1955] | layer2_out[1956];
    assign layer3_out[3870] = ~layer2_out[1434];
    assign layer3_out[3871] = layer2_out[1470];
    assign layer3_out[3872] = ~(layer2_out[3291] ^ layer2_out[3292]);
    assign layer3_out[3873] = layer2_out[10];
    assign layer3_out[3874] = layer2_out[3034] ^ layer2_out[3035];
    assign layer3_out[3875] = layer2_out[3989];
    assign layer3_out[3876] = ~(layer2_out[6101] | layer2_out[6102]);
    assign layer3_out[3877] = ~(layer2_out[1598] | layer2_out[1599]);
    assign layer3_out[3878] = layer2_out[942];
    assign layer3_out[3879] = layer2_out[3184] ^ layer2_out[3185];
    assign layer3_out[3880] = ~layer2_out[3482];
    assign layer3_out[3881] = layer2_out[4878] & layer2_out[4879];
    assign layer3_out[3882] = layer2_out[156];
    assign layer3_out[3883] = ~(layer2_out[3192] | layer2_out[3193]);
    assign layer3_out[3884] = ~layer2_out[6780];
    assign layer3_out[3885] = 1'b1;
    assign layer3_out[3886] = ~layer2_out[628] | layer2_out[629];
    assign layer3_out[3887] = ~layer2_out[6475];
    assign layer3_out[3888] = layer2_out[3378];
    assign layer3_out[3889] = ~layer2_out[3855] | layer2_out[3854];
    assign layer3_out[3890] = layer2_out[5934] & layer2_out[5935];
    assign layer3_out[3891] = layer2_out[1914] & layer2_out[1915];
    assign layer3_out[3892] = layer2_out[4367];
    assign layer3_out[3893] = ~layer2_out[447];
    assign layer3_out[3894] = ~layer2_out[1964];
    assign layer3_out[3895] = layer2_out[2620];
    assign layer3_out[3896] = ~(layer2_out[3161] ^ layer2_out[3162]);
    assign layer3_out[3897] = layer2_out[7573] & layer2_out[7574];
    assign layer3_out[3898] = layer2_out[1990];
    assign layer3_out[3899] = ~layer2_out[238];
    assign layer3_out[3900] = ~layer2_out[5269];
    assign layer3_out[3901] = layer2_out[7819] | layer2_out[7820];
    assign layer3_out[3902] = layer2_out[6024] & layer2_out[6025];
    assign layer3_out[3903] = ~(layer2_out[3015] & layer2_out[3016]);
    assign layer3_out[3904] = layer2_out[7000] | layer2_out[7001];
    assign layer3_out[3905] = layer2_out[6977] | layer2_out[6978];
    assign layer3_out[3906] = layer2_out[4800] & layer2_out[4801];
    assign layer3_out[3907] = ~layer2_out[6194];
    assign layer3_out[3908] = layer2_out[5337];
    assign layer3_out[3909] = layer2_out[5767];
    assign layer3_out[3910] = 1'b1;
    assign layer3_out[3911] = ~layer2_out[5017];
    assign layer3_out[3912] = layer2_out[6841] & ~layer2_out[6840];
    assign layer3_out[3913] = ~layer2_out[2709];
    assign layer3_out[3914] = ~(layer2_out[6755] & layer2_out[6756]);
    assign layer3_out[3915] = layer2_out[2412];
    assign layer3_out[3916] = layer2_out[282] & ~layer2_out[283];
    assign layer3_out[3917] = ~(layer2_out[684] | layer2_out[685]);
    assign layer3_out[3918] = ~layer2_out[4475];
    assign layer3_out[3919] = layer2_out[6795] & layer2_out[6796];
    assign layer3_out[3920] = layer2_out[2599];
    assign layer3_out[3921] = layer2_out[2144];
    assign layer3_out[3922] = ~layer2_out[5403];
    assign layer3_out[3923] = layer2_out[2440];
    assign layer3_out[3924] = layer2_out[7361];
    assign layer3_out[3925] = layer2_out[6309] & ~layer2_out[6308];
    assign layer3_out[3926] = ~layer2_out[1570];
    assign layer3_out[3927] = ~(layer2_out[4871] ^ layer2_out[4872]);
    assign layer3_out[3928] = layer2_out[4446] ^ layer2_out[4447];
    assign layer3_out[3929] = layer2_out[3039] & layer2_out[3040];
    assign layer3_out[3930] = ~layer2_out[2222] | layer2_out[2221];
    assign layer3_out[3931] = layer2_out[4696];
    assign layer3_out[3932] = layer2_out[3108] & layer2_out[3109];
    assign layer3_out[3933] = ~layer2_out[7509] | layer2_out[7508];
    assign layer3_out[3934] = layer2_out[2629];
    assign layer3_out[3935] = ~layer2_out[5684];
    assign layer3_out[3936] = layer2_out[5757] & layer2_out[5758];
    assign layer3_out[3937] = ~layer2_out[7325];
    assign layer3_out[3938] = ~(layer2_out[281] ^ layer2_out[282]);
    assign layer3_out[3939] = layer2_out[7939] & ~layer2_out[7938];
    assign layer3_out[3940] = ~layer2_out[4058];
    assign layer3_out[3941] = ~layer2_out[1871] | layer2_out[1870];
    assign layer3_out[3942] = ~(layer2_out[80] | layer2_out[81]);
    assign layer3_out[3943] = ~(layer2_out[1153] ^ layer2_out[1154]);
    assign layer3_out[3944] = ~layer2_out[2092];
    assign layer3_out[3945] = layer2_out[7249];
    assign layer3_out[3946] = ~layer2_out[4372] | layer2_out[4373];
    assign layer3_out[3947] = ~(layer2_out[869] ^ layer2_out[870]);
    assign layer3_out[3948] = layer2_out[2479] & ~layer2_out[2478];
    assign layer3_out[3949] = ~layer2_out[1613];
    assign layer3_out[3950] = layer2_out[4368];
    assign layer3_out[3951] = layer2_out[6275] ^ layer2_out[6276];
    assign layer3_out[3952] = ~layer2_out[1833];
    assign layer3_out[3953] = ~(layer2_out[4111] | layer2_out[4112]);
    assign layer3_out[3954] = ~(layer2_out[7626] ^ layer2_out[7627]);
    assign layer3_out[3955] = ~(layer2_out[1053] | layer2_out[1054]);
    assign layer3_out[3956] = ~layer2_out[5672];
    assign layer3_out[3957] = ~layer2_out[3997];
    assign layer3_out[3958] = ~layer2_out[7401];
    assign layer3_out[3959] = ~(layer2_out[4109] & layer2_out[4110]);
    assign layer3_out[3960] = ~layer2_out[2071] | layer2_out[2072];
    assign layer3_out[3961] = layer2_out[992];
    assign layer3_out[3962] = layer2_out[6361];
    assign layer3_out[3963] = layer2_out[3426];
    assign layer3_out[3964] = layer2_out[7431] & ~layer2_out[7432];
    assign layer3_out[3965] = layer2_out[5972] | layer2_out[5973];
    assign layer3_out[3966] = ~layer2_out[3956];
    assign layer3_out[3967] = ~(layer2_out[686] | layer2_out[687]);
    assign layer3_out[3968] = layer2_out[984];
    assign layer3_out[3969] = ~(layer2_out[4959] ^ layer2_out[4960]);
    assign layer3_out[3970] = layer2_out[4935] & ~layer2_out[4936];
    assign layer3_out[3971] = ~layer2_out[3960] | layer2_out[3959];
    assign layer3_out[3972] = ~layer2_out[7680];
    assign layer3_out[3973] = layer2_out[4868] ^ layer2_out[4869];
    assign layer3_out[3974] = ~layer2_out[4760];
    assign layer3_out[3975] = layer2_out[4586];
    assign layer3_out[3976] = ~(layer2_out[1768] | layer2_out[1769]);
    assign layer3_out[3977] = ~layer2_out[7572];
    assign layer3_out[3978] = ~layer2_out[2954] | layer2_out[2953];
    assign layer3_out[3979] = ~layer2_out[6962];
    assign layer3_out[3980] = 1'b1;
    assign layer3_out[3981] = layer2_out[913] ^ layer2_out[914];
    assign layer3_out[3982] = 1'b1;
    assign layer3_out[3983] = layer2_out[3401];
    assign layer3_out[3984] = ~layer2_out[4526];
    assign layer3_out[3985] = ~layer2_out[5947] | layer2_out[5946];
    assign layer3_out[3986] = 1'b0;
    assign layer3_out[3987] = layer2_out[1175] & ~layer2_out[1174];
    assign layer3_out[3988] = layer2_out[7652] | layer2_out[7653];
    assign layer3_out[3989] = layer2_out[4608] | layer2_out[4609];
    assign layer3_out[3990] = ~layer2_out[2531] | layer2_out[2530];
    assign layer3_out[3991] = layer2_out[7875];
    assign layer3_out[3992] = layer2_out[2453];
    assign layer3_out[3993] = ~layer2_out[4626] | layer2_out[4625];
    assign layer3_out[3994] = layer2_out[4277];
    assign layer3_out[3995] = ~(layer2_out[7941] & layer2_out[7942]);
    assign layer3_out[3996] = ~layer2_out[5897];
    assign layer3_out[3997] = layer2_out[1944];
    assign layer3_out[3998] = ~layer2_out[4428] | layer2_out[4427];
    assign layer3_out[3999] = ~(layer2_out[6925] & layer2_out[6926]);
    assign layer3_out[4000] = ~layer2_out[4301];
    assign layer3_out[4001] = ~(layer2_out[4691] & layer2_out[4692]);
    assign layer3_out[4002] = layer2_out[6343];
    assign layer3_out[4003] = ~layer2_out[7611] | layer2_out[7612];
    assign layer3_out[4004] = ~layer2_out[2918] | layer2_out[2917];
    assign layer3_out[4005] = ~(layer2_out[5524] ^ layer2_out[5525]);
    assign layer3_out[4006] = ~layer2_out[5586] | layer2_out[5587];
    assign layer3_out[4007] = ~layer2_out[4820];
    assign layer3_out[4008] = ~(layer2_out[7844] | layer2_out[7845]);
    assign layer3_out[4009] = ~layer2_out[7945];
    assign layer3_out[4010] = layer2_out[3346];
    assign layer3_out[4011] = ~layer2_out[2170] | layer2_out[2169];
    assign layer3_out[4012] = layer2_out[3266];
    assign layer3_out[4013] = layer2_out[6410];
    assign layer3_out[4014] = ~layer2_out[7895] | layer2_out[7896];
    assign layer3_out[4015] = layer2_out[550];
    assign layer3_out[4016] = ~layer2_out[2701] | layer2_out[2700];
    assign layer3_out[4017] = ~layer2_out[5691] | layer2_out[5690];
    assign layer3_out[4018] = layer2_out[6593];
    assign layer3_out[4019] = ~layer2_out[3756];
    assign layer3_out[4020] = ~layer2_out[197];
    assign layer3_out[4021] = layer2_out[5168];
    assign layer3_out[4022] = ~layer2_out[4676];
    assign layer3_out[4023] = layer2_out[7489] | layer2_out[7490];
    assign layer3_out[4024] = layer2_out[3674] | layer2_out[3675];
    assign layer3_out[4025] = layer2_out[6803];
    assign layer3_out[4026] = ~(layer2_out[346] & layer2_out[347]);
    assign layer3_out[4027] = ~layer2_out[3814];
    assign layer3_out[4028] = ~layer2_out[7429];
    assign layer3_out[4029] = ~layer2_out[1244];
    assign layer3_out[4030] = ~layer2_out[5418];
    assign layer3_out[4031] = layer2_out[6482];
    assign layer3_out[4032] = layer2_out[4513] | layer2_out[4514];
    assign layer3_out[4033] = ~layer2_out[7827] | layer2_out[7826];
    assign layer3_out[4034] = ~layer2_out[5069] | layer2_out[5068];
    assign layer3_out[4035] = layer2_out[7774];
    assign layer3_out[4036] = layer2_out[7723] | layer2_out[7724];
    assign layer3_out[4037] = ~layer2_out[6075];
    assign layer3_out[4038] = ~layer2_out[5191];
    assign layer3_out[4039] = layer2_out[2875] & ~layer2_out[2874];
    assign layer3_out[4040] = ~layer2_out[2902];
    assign layer3_out[4041] = 1'b1;
    assign layer3_out[4042] = layer2_out[4370];
    assign layer3_out[4043] = 1'b0;
    assign layer3_out[4044] = ~(layer2_out[670] ^ layer2_out[671]);
    assign layer3_out[4045] = layer2_out[407];
    assign layer3_out[4046] = ~layer2_out[578];
    assign layer3_out[4047] = ~(layer2_out[6347] ^ layer2_out[6348]);
    assign layer3_out[4048] = layer2_out[4903];
    assign layer3_out[4049] = ~layer2_out[4870];
    assign layer3_out[4050] = layer2_out[6104];
    assign layer3_out[4051] = ~layer2_out[2501];
    assign layer3_out[4052] = layer2_out[118];
    assign layer3_out[4053] = layer2_out[4243];
    assign layer3_out[4054] = layer2_out[981] | layer2_out[982];
    assign layer3_out[4055] = ~(layer2_out[959] ^ layer2_out[960]);
    assign layer3_out[4056] = ~(layer2_out[1603] ^ layer2_out[1604]);
    assign layer3_out[4057] = layer2_out[2740] | layer2_out[2741];
    assign layer3_out[4058] = layer2_out[1185];
    assign layer3_out[4059] = layer2_out[84] & ~layer2_out[83];
    assign layer3_out[4060] = layer2_out[1256] | layer2_out[1257];
    assign layer3_out[4061] = layer2_out[7637];
    assign layer3_out[4062] = ~(layer2_out[5098] & layer2_out[5099]);
    assign layer3_out[4063] = layer2_out[969] & ~layer2_out[968];
    assign layer3_out[4064] = ~(layer2_out[4767] | layer2_out[4768]);
    assign layer3_out[4065] = ~(layer2_out[2479] | layer2_out[2480]);
    assign layer3_out[4066] = layer2_out[870];
    assign layer3_out[4067] = 1'b1;
    assign layer3_out[4068] = ~(layer2_out[1276] & layer2_out[1277]);
    assign layer3_out[4069] = layer2_out[6798];
    assign layer3_out[4070] = layer2_out[6365] & ~layer2_out[6364];
    assign layer3_out[4071] = ~layer2_out[1347];
    assign layer3_out[4072] = ~layer2_out[5272];
    assign layer3_out[4073] = ~layer2_out[5431];
    assign layer3_out[4074] = layer2_out[4936] & ~layer2_out[4937];
    assign layer3_out[4075] = ~layer2_out[464];
    assign layer3_out[4076] = layer2_out[6040] ^ layer2_out[6041];
    assign layer3_out[4077] = layer2_out[5761];
    assign layer3_out[4078] = ~layer2_out[1545] | layer2_out[1546];
    assign layer3_out[4079] = layer2_out[7369] & layer2_out[7370];
    assign layer3_out[4080] = layer2_out[3614] | layer2_out[3615];
    assign layer3_out[4081] = layer2_out[1084] ^ layer2_out[1085];
    assign layer3_out[4082] = ~layer2_out[6655];
    assign layer3_out[4083] = ~layer2_out[2588] | layer2_out[2587];
    assign layer3_out[4084] = layer2_out[5694];
    assign layer3_out[4085] = layer2_out[318] & ~layer2_out[319];
    assign layer3_out[4086] = layer2_out[2973];
    assign layer3_out[4087] = layer2_out[2923];
    assign layer3_out[4088] = layer2_out[7620] & ~layer2_out[7619];
    assign layer3_out[4089] = ~(layer2_out[5318] & layer2_out[5319]);
    assign layer3_out[4090] = ~(layer2_out[1887] ^ layer2_out[1888]);
    assign layer3_out[4091] = ~layer2_out[1735] | layer2_out[1734];
    assign layer3_out[4092] = ~(layer2_out[5526] ^ layer2_out[5527]);
    assign layer3_out[4093] = ~(layer2_out[502] | layer2_out[503]);
    assign layer3_out[4094] = layer2_out[6498];
    assign layer3_out[4095] = layer2_out[3538] & ~layer2_out[3537];
    assign layer3_out[4096] = layer2_out[6972] & layer2_out[6973];
    assign layer3_out[4097] = layer2_out[2342] & ~layer2_out[2343];
    assign layer3_out[4098] = ~layer2_out[3978];
    assign layer3_out[4099] = layer2_out[7518] & layer2_out[7519];
    assign layer3_out[4100] = layer2_out[5869];
    assign layer3_out[4101] = ~(layer2_out[4106] ^ layer2_out[4107]);
    assign layer3_out[4102] = ~(layer2_out[4067] & layer2_out[4068]);
    assign layer3_out[4103] = ~layer2_out[1499];
    assign layer3_out[4104] = ~layer2_out[6933];
    assign layer3_out[4105] = ~layer2_out[2075];
    assign layer3_out[4106] = layer2_out[2761] & ~layer2_out[2762];
    assign layer3_out[4107] = ~(layer2_out[3776] | layer2_out[3777]);
    assign layer3_out[4108] = layer2_out[4404];
    assign layer3_out[4109] = layer2_out[4017];
    assign layer3_out[4110] = layer2_out[1584];
    assign layer3_out[4111] = layer2_out[3403] ^ layer2_out[3404];
    assign layer3_out[4112] = ~(layer2_out[3531] | layer2_out[3532]);
    assign layer3_out[4113] = layer2_out[7269] ^ layer2_out[7270];
    assign layer3_out[4114] = ~layer2_out[1592];
    assign layer3_out[4115] = ~layer2_out[5876];
    assign layer3_out[4116] = ~layer2_out[3858];
    assign layer3_out[4117] = ~layer2_out[460];
    assign layer3_out[4118] = ~layer2_out[1560];
    assign layer3_out[4119] = layer2_out[587] & ~layer2_out[588];
    assign layer3_out[4120] = layer2_out[5671] & layer2_out[5672];
    assign layer3_out[4121] = layer2_out[6068];
    assign layer3_out[4122] = layer2_out[4808] ^ layer2_out[4809];
    assign layer3_out[4123] = ~layer2_out[6535];
    assign layer3_out[4124] = layer2_out[553] & layer2_out[554];
    assign layer3_out[4125] = layer2_out[4003] & ~layer2_out[4004];
    assign layer3_out[4126] = layer2_out[7559] & ~layer2_out[7558];
    assign layer3_out[4127] = ~layer2_out[229];
    assign layer3_out[4128] = layer2_out[4879] & ~layer2_out[4880];
    assign layer3_out[4129] = layer2_out[4135] & ~layer2_out[4136];
    assign layer3_out[4130] = ~layer2_out[2183];
    assign layer3_out[4131] = layer2_out[1760] & ~layer2_out[1761];
    assign layer3_out[4132] = layer2_out[5427];
    assign layer3_out[4133] = ~layer2_out[3755] | layer2_out[3754];
    assign layer3_out[4134] = ~layer2_out[6726];
    assign layer3_out[4135] = ~layer2_out[2761];
    assign layer3_out[4136] = layer2_out[3274];
    assign layer3_out[4137] = layer2_out[1233];
    assign layer3_out[4138] = ~layer2_out[203] | layer2_out[204];
    assign layer3_out[4139] = ~layer2_out[396];
    assign layer3_out[4140] = ~layer2_out[1225];
    assign layer3_out[4141] = layer2_out[3320];
    assign layer3_out[4142] = ~(layer2_out[5094] & layer2_out[5095]);
    assign layer3_out[4143] = ~layer2_out[5470];
    assign layer3_out[4144] = layer2_out[3681] & layer2_out[3682];
    assign layer3_out[4145] = layer2_out[5712] & ~layer2_out[5713];
    assign layer3_out[4146] = layer2_out[7400];
    assign layer3_out[4147] = layer2_out[6837] | layer2_out[6838];
    assign layer3_out[4148] = layer2_out[7171];
    assign layer3_out[4149] = layer2_out[3244];
    assign layer3_out[4150] = layer2_out[4261];
    assign layer3_out[4151] = layer2_out[7800] | layer2_out[7801];
    assign layer3_out[4152] = 1'b0;
    assign layer3_out[4153] = ~(layer2_out[5370] & layer2_out[5371]);
    assign layer3_out[4154] = layer2_out[4232] & ~layer2_out[4233];
    assign layer3_out[4155] = ~(layer2_out[7695] & layer2_out[7696]);
    assign layer3_out[4156] = layer2_out[1649];
    assign layer3_out[4157] = ~(layer2_out[6540] | layer2_out[6541]);
    assign layer3_out[4158] = ~layer2_out[4624];
    assign layer3_out[4159] = layer2_out[2967] & ~layer2_out[2966];
    assign layer3_out[4160] = layer2_out[7349] ^ layer2_out[7350];
    assign layer3_out[4161] = ~(layer2_out[7622] & layer2_out[7623]);
    assign layer3_out[4162] = ~(layer2_out[6781] & layer2_out[6782]);
    assign layer3_out[4163] = ~(layer2_out[1854] | layer2_out[1855]);
    assign layer3_out[4164] = layer2_out[1977] ^ layer2_out[1978];
    assign layer3_out[4165] = ~layer2_out[4206];
    assign layer3_out[4166] = layer2_out[2863];
    assign layer3_out[4167] = ~layer2_out[5509];
    assign layer3_out[4168] = layer2_out[4564];
    assign layer3_out[4169] = ~layer2_out[3370] | layer2_out[3371];
    assign layer3_out[4170] = layer2_out[660] ^ layer2_out[661];
    assign layer3_out[4171] = ~layer2_out[2136];
    assign layer3_out[4172] = ~layer2_out[275] | layer2_out[276];
    assign layer3_out[4173] = layer2_out[6596] & ~layer2_out[6595];
    assign layer3_out[4174] = ~layer2_out[2935];
    assign layer3_out[4175] = layer2_out[2263] & layer2_out[2264];
    assign layer3_out[4176] = ~(layer2_out[7995] | layer2_out[7996]);
    assign layer3_out[4177] = 1'b0;
    assign layer3_out[4178] = layer2_out[5392];
    assign layer3_out[4179] = layer2_out[5629];
    assign layer3_out[4180] = layer2_out[1145] & ~layer2_out[1146];
    assign layer3_out[4181] = layer2_out[7128];
    assign layer3_out[4182] = layer2_out[3245] & layer2_out[3246];
    assign layer3_out[4183] = ~layer2_out[2010] | layer2_out[2009];
    assign layer3_out[4184] = ~layer2_out[535] | layer2_out[536];
    assign layer3_out[4185] = layer2_out[1774] ^ layer2_out[1775];
    assign layer3_out[4186] = ~(layer2_out[1954] | layer2_out[1955]);
    assign layer3_out[4187] = layer2_out[1178] & ~layer2_out[1177];
    assign layer3_out[4188] = layer2_out[2114] & ~layer2_out[2115];
    assign layer3_out[4189] = layer2_out[115] & ~layer2_out[114];
    assign layer3_out[4190] = layer2_out[7124];
    assign layer3_out[4191] = 1'b0;
    assign layer3_out[4192] = layer2_out[1863] & layer2_out[1864];
    assign layer3_out[4193] = layer2_out[5453] & layer2_out[5454];
    assign layer3_out[4194] = ~layer2_out[2188];
    assign layer3_out[4195] = ~layer2_out[2053] | layer2_out[2054];
    assign layer3_out[4196] = ~(layer2_out[2397] | layer2_out[2398]);
    assign layer3_out[4197] = layer2_out[6063] & layer2_out[6064];
    assign layer3_out[4198] = ~layer2_out[3315];
    assign layer3_out[4199] = ~(layer2_out[6648] & layer2_out[6649]);
    assign layer3_out[4200] = layer2_out[5825] & ~layer2_out[5824];
    assign layer3_out[4201] = ~(layer2_out[6335] | layer2_out[6336]);
    assign layer3_out[4202] = ~(layer2_out[3010] & layer2_out[3011]);
    assign layer3_out[4203] = ~layer2_out[7811] | layer2_out[7812];
    assign layer3_out[4204] = ~layer2_out[6748];
    assign layer3_out[4205] = layer2_out[603] & ~layer2_out[602];
    assign layer3_out[4206] = ~layer2_out[1134];
    assign layer3_out[4207] = ~layer2_out[310];
    assign layer3_out[4208] = layer2_out[6762] & layer2_out[6763];
    assign layer3_out[4209] = layer2_out[3765] | layer2_out[3766];
    assign layer3_out[4210] = ~layer2_out[2121] | layer2_out[2122];
    assign layer3_out[4211] = ~(layer2_out[3160] ^ layer2_out[3161]);
    assign layer3_out[4212] = layer2_out[1272] & ~layer2_out[1273];
    assign layer3_out[4213] = ~layer2_out[3096];
    assign layer3_out[4214] = ~layer2_out[4314] | layer2_out[4315];
    assign layer3_out[4215] = layer2_out[6628] & ~layer2_out[6627];
    assign layer3_out[4216] = ~layer2_out[6518] | layer2_out[6517];
    assign layer3_out[4217] = ~layer2_out[5304];
    assign layer3_out[4218] = layer2_out[2399] | layer2_out[2400];
    assign layer3_out[4219] = layer2_out[3925];
    assign layer3_out[4220] = layer2_out[4775];
    assign layer3_out[4221] = ~(layer2_out[2495] | layer2_out[2496]);
    assign layer3_out[4222] = ~layer2_out[4981];
    assign layer3_out[4223] = 1'b0;
    assign layer3_out[4224] = layer2_out[4197] & ~layer2_out[4198];
    assign layer3_out[4225] = ~layer2_out[4422] | layer2_out[4421];
    assign layer3_out[4226] = layer2_out[5141] ^ layer2_out[5142];
    assign layer3_out[4227] = ~layer2_out[6105];
    assign layer3_out[4228] = ~(layer2_out[2739] ^ layer2_out[2740]);
    assign layer3_out[4229] = layer2_out[2685] & ~layer2_out[2684];
    assign layer3_out[4230] = layer2_out[3211];
    assign layer3_out[4231] = layer2_out[5553] ^ layer2_out[5554];
    assign layer3_out[4232] = layer2_out[3866] & ~layer2_out[3867];
    assign layer3_out[4233] = layer2_out[7401];
    assign layer3_out[4234] = layer2_out[1718];
    assign layer3_out[4235] = layer2_out[5980] & ~layer2_out[5979];
    assign layer3_out[4236] = layer2_out[6664];
    assign layer3_out[4237] = ~layer2_out[3328];
    assign layer3_out[4238] = layer2_out[1941] ^ layer2_out[1942];
    assign layer3_out[4239] = ~layer2_out[469];
    assign layer3_out[4240] = layer2_out[7890] | layer2_out[7891];
    assign layer3_out[4241] = layer2_out[2098] & layer2_out[2099];
    assign layer3_out[4242] = layer2_out[1509] | layer2_out[1510];
    assign layer3_out[4243] = layer2_out[2902] & ~layer2_out[2901];
    assign layer3_out[4244] = ~layer2_out[2572] | layer2_out[2571];
    assign layer3_out[4245] = ~(layer2_out[1803] ^ layer2_out[1804]);
    assign layer3_out[4246] = layer2_out[975] | layer2_out[976];
    assign layer3_out[4247] = ~layer2_out[1741];
    assign layer3_out[4248] = layer2_out[789] & ~layer2_out[788];
    assign layer3_out[4249] = ~layer2_out[7506] | layer2_out[7507];
    assign layer3_out[4250] = ~layer2_out[4437];
    assign layer3_out[4251] = layer2_out[5893];
    assign layer3_out[4252] = ~(layer2_out[4911] & layer2_out[4912]);
    assign layer3_out[4253] = ~layer2_out[632];
    assign layer3_out[4254] = ~layer2_out[1220];
    assign layer3_out[4255] = ~layer2_out[2548];
    assign layer3_out[4256] = ~layer2_out[610];
    assign layer3_out[4257] = ~layer2_out[3209] | layer2_out[3208];
    assign layer3_out[4258] = ~layer2_out[5910];
    assign layer3_out[4259] = ~layer2_out[5357];
    assign layer3_out[4260] = ~layer2_out[530] | layer2_out[529];
    assign layer3_out[4261] = layer2_out[6422];
    assign layer3_out[4262] = layer2_out[5797] & ~layer2_out[5798];
    assign layer3_out[4263] = layer2_out[1945] & ~layer2_out[1944];
    assign layer3_out[4264] = ~layer2_out[2800];
    assign layer3_out[4265] = ~(layer2_out[6575] ^ layer2_out[6576]);
    assign layer3_out[4266] = layer2_out[349] | layer2_out[350];
    assign layer3_out[4267] = layer2_out[2098] & ~layer2_out[2097];
    assign layer3_out[4268] = layer2_out[2677];
    assign layer3_out[4269] = layer2_out[3557];
    assign layer3_out[4270] = layer2_out[1199] ^ layer2_out[1200];
    assign layer3_out[4271] = ~layer2_out[5861];
    assign layer3_out[4272] = ~(layer2_out[3158] | layer2_out[3159]);
    assign layer3_out[4273] = ~layer2_out[4247];
    assign layer3_out[4274] = ~(layer2_out[3475] | layer2_out[3476]);
    assign layer3_out[4275] = layer2_out[5140] & layer2_out[5141];
    assign layer3_out[4276] = layer2_out[7577] & ~layer2_out[7576];
    assign layer3_out[4277] = ~layer2_out[3731];
    assign layer3_out[4278] = ~(layer2_out[4851] | layer2_out[4852]);
    assign layer3_out[4279] = layer2_out[7972] & layer2_out[7973];
    assign layer3_out[4280] = layer2_out[2269];
    assign layer3_out[4281] = ~(layer2_out[1965] & layer2_out[1966]);
    assign layer3_out[4282] = ~(layer2_out[7255] & layer2_out[7256]);
    assign layer3_out[4283] = ~layer2_out[5963];
    assign layer3_out[4284] = ~layer2_out[4235];
    assign layer3_out[4285] = layer2_out[1705] ^ layer2_out[1706];
    assign layer3_out[4286] = layer2_out[7299] & layer2_out[7300];
    assign layer3_out[4287] = layer2_out[4962] & layer2_out[4963];
    assign layer3_out[4288] = ~(layer2_out[7816] & layer2_out[7817]);
    assign layer3_out[4289] = layer2_out[6561] & layer2_out[6562];
    assign layer3_out[4290] = layer2_out[3756] & ~layer2_out[3757];
    assign layer3_out[4291] = ~layer2_out[1058];
    assign layer3_out[4292] = ~(layer2_out[7139] ^ layer2_out[7140]);
    assign layer3_out[4293] = ~(layer2_out[3713] & layer2_out[3714]);
    assign layer3_out[4294] = layer2_out[5307] & layer2_out[5308];
    assign layer3_out[4295] = ~(layer2_out[2078] | layer2_out[2079]);
    assign layer3_out[4296] = layer2_out[6486] & ~layer2_out[6487];
    assign layer3_out[4297] = ~layer2_out[4731];
    assign layer3_out[4298] = layer2_out[6178] & layer2_out[6179];
    assign layer3_out[4299] = layer2_out[7103];
    assign layer3_out[4300] = ~layer2_out[1892];
    assign layer3_out[4301] = ~(layer2_out[6033] ^ layer2_out[6034]);
    assign layer3_out[4302] = ~layer2_out[5785];
    assign layer3_out[4303] = ~layer2_out[5689] | layer2_out[5690];
    assign layer3_out[4304] = layer2_out[1299] & ~layer2_out[1300];
    assign layer3_out[4305] = 1'b0;
    assign layer3_out[4306] = layer2_out[713];
    assign layer3_out[4307] = ~layer2_out[3647];
    assign layer3_out[4308] = ~(layer2_out[2046] ^ layer2_out[2047]);
    assign layer3_out[4309] = layer2_out[2925];
    assign layer3_out[4310] = ~layer2_out[4191];
    assign layer3_out[4311] = ~layer2_out[319];
    assign layer3_out[4312] = ~layer2_out[3771];
    assign layer3_out[4313] = layer2_out[952];
    assign layer3_out[4314] = layer2_out[5547] | layer2_out[5548];
    assign layer3_out[4315] = layer2_out[2670] ^ layer2_out[2671];
    assign layer3_out[4316] = layer2_out[5789];
    assign layer3_out[4317] = ~layer2_out[465];
    assign layer3_out[4318] = layer2_out[3718];
    assign layer3_out[4319] = layer2_out[2167];
    assign layer3_out[4320] = layer2_out[4564] | layer2_out[4565];
    assign layer3_out[4321] = ~(layer2_out[4080] & layer2_out[4081]);
    assign layer3_out[4322] = ~layer2_out[6731] | layer2_out[6732];
    assign layer3_out[4323] = 1'b1;
    assign layer3_out[4324] = ~(layer2_out[6850] & layer2_out[6851]);
    assign layer3_out[4325] = ~layer2_out[7555] | layer2_out[7554];
    assign layer3_out[4326] = layer2_out[2216];
    assign layer3_out[4327] = ~layer2_out[4255];
    assign layer3_out[4328] = layer2_out[145] & ~layer2_out[144];
    assign layer3_out[4329] = ~layer2_out[2160];
    assign layer3_out[4330] = ~(layer2_out[3331] ^ layer2_out[3332]);
    assign layer3_out[4331] = layer2_out[4007];
    assign layer3_out[4332] = ~(layer2_out[3272] ^ layer2_out[3273]);
    assign layer3_out[4333] = ~layer2_out[405] | layer2_out[404];
    assign layer3_out[4334] = ~layer2_out[6711];
    assign layer3_out[4335] = layer2_out[2773] ^ layer2_out[2774];
    assign layer3_out[4336] = layer2_out[975];
    assign layer3_out[4337] = layer2_out[2449];
    assign layer3_out[4338] = ~layer2_out[5467];
    assign layer3_out[4339] = ~layer2_out[1639];
    assign layer3_out[4340] = layer2_out[7016];
    assign layer3_out[4341] = layer2_out[1826] ^ layer2_out[1827];
    assign layer3_out[4342] = ~(layer2_out[2826] & layer2_out[2827]);
    assign layer3_out[4343] = layer2_out[6636];
    assign layer3_out[4344] = layer2_out[3322];
    assign layer3_out[4345] = layer2_out[7135];
    assign layer3_out[4346] = layer2_out[7242];
    assign layer3_out[4347] = ~(layer2_out[1448] ^ layer2_out[1449]);
    assign layer3_out[4348] = layer2_out[2905] & ~layer2_out[2904];
    assign layer3_out[4349] = layer2_out[5100] | layer2_out[5101];
    assign layer3_out[4350] = ~layer2_out[52] | layer2_out[51];
    assign layer3_out[4351] = ~(layer2_out[4946] & layer2_out[4947]);
    assign layer3_out[4352] = ~layer2_out[7007];
    assign layer3_out[4353] = layer2_out[3995] ^ layer2_out[3996];
    assign layer3_out[4354] = 1'b0;
    assign layer3_out[4355] = layer2_out[3524] & layer2_out[3525];
    assign layer3_out[4356] = ~layer2_out[7676];
    assign layer3_out[4357] = layer2_out[7476] ^ layer2_out[7477];
    assign layer3_out[4358] = ~(layer2_out[6193] ^ layer2_out[6194]);
    assign layer3_out[4359] = ~layer2_out[3623] | layer2_out[3624];
    assign layer3_out[4360] = ~layer2_out[2314];
    assign layer3_out[4361] = ~(layer2_out[84] | layer2_out[85]);
    assign layer3_out[4362] = ~layer2_out[934];
    assign layer3_out[4363] = layer2_out[6487] ^ layer2_out[6488];
    assign layer3_out[4364] = layer2_out[4078];
    assign layer3_out[4365] = layer2_out[2275] ^ layer2_out[2276];
    assign layer3_out[4366] = layer2_out[888] & layer2_out[889];
    assign layer3_out[4367] = ~layer2_out[3689];
    assign layer3_out[4368] = ~layer2_out[1310];
    assign layer3_out[4369] = ~layer2_out[2772];
    assign layer3_out[4370] = layer2_out[3222] ^ layer2_out[3223];
    assign layer3_out[4371] = layer2_out[6822];
    assign layer3_out[4372] = ~(layer2_out[6945] | layer2_out[6946]);
    assign layer3_out[4373] = layer2_out[2779] ^ layer2_out[2780];
    assign layer3_out[4374] = layer2_out[813] & layer2_out[814];
    assign layer3_out[4375] = ~layer2_out[290] | layer2_out[291];
    assign layer3_out[4376] = ~layer2_out[6036] | layer2_out[6037];
    assign layer3_out[4377] = layer2_out[5933];
    assign layer3_out[4378] = ~(layer2_out[1205] & layer2_out[1206]);
    assign layer3_out[4379] = layer2_out[5049] & ~layer2_out[5050];
    assign layer3_out[4380] = ~layer2_out[7758];
    assign layer3_out[4381] = ~layer2_out[5016];
    assign layer3_out[4382] = layer2_out[6700];
    assign layer3_out[4383] = layer2_out[6537];
    assign layer3_out[4384] = ~layer2_out[6864];
    assign layer3_out[4385] = layer2_out[2061];
    assign layer3_out[4386] = layer2_out[4064] & layer2_out[4065];
    assign layer3_out[4387] = layer2_out[5871];
    assign layer3_out[4388] = layer2_out[5880] & ~layer2_out[5881];
    assign layer3_out[4389] = layer2_out[2488];
    assign layer3_out[4390] = layer2_out[1328] & layer2_out[1329];
    assign layer3_out[4391] = ~(layer2_out[5041] ^ layer2_out[5042]);
    assign layer3_out[4392] = layer2_out[7276] & ~layer2_out[7275];
    assign layer3_out[4393] = ~(layer2_out[2386] | layer2_out[2387]);
    assign layer3_out[4394] = layer2_out[6250];
    assign layer3_out[4395] = layer2_out[2076] & layer2_out[2077];
    assign layer3_out[4396] = layer2_out[1556];
    assign layer3_out[4397] = layer2_out[6496];
    assign layer3_out[4398] = ~layer2_out[4097];
    assign layer3_out[4399] = layer2_out[175] & ~layer2_out[174];
    assign layer3_out[4400] = ~layer2_out[6772];
    assign layer3_out[4401] = ~(layer2_out[3145] | layer2_out[3146]);
    assign layer3_out[4402] = ~layer2_out[2040];
    assign layer3_out[4403] = ~layer2_out[5562];
    assign layer3_out[4404] = layer2_out[7805] & ~layer2_out[7804];
    assign layer3_out[4405] = layer2_out[6913] & ~layer2_out[6914];
    assign layer3_out[4406] = ~(layer2_out[326] & layer2_out[327]);
    assign layer3_out[4407] = ~layer2_out[6527];
    assign layer3_out[4408] = ~(layer2_out[894] & layer2_out[895]);
    assign layer3_out[4409] = ~layer2_out[2202] | layer2_out[2203];
    assign layer3_out[4410] = layer2_out[5997];
    assign layer3_out[4411] = layer2_out[6060] & ~layer2_out[6061];
    assign layer3_out[4412] = ~layer2_out[6416];
    assign layer3_out[4413] = ~layer2_out[4919];
    assign layer3_out[4414] = layer2_out[7200] | layer2_out[7201];
    assign layer3_out[4415] = ~layer2_out[7355] | layer2_out[7356];
    assign layer3_out[4416] = ~(layer2_out[4543] & layer2_out[4544]);
    assign layer3_out[4417] = layer2_out[5571] & layer2_out[5572];
    assign layer3_out[4418] = layer2_out[6751] ^ layer2_out[6752];
    assign layer3_out[4419] = layer2_out[2647];
    assign layer3_out[4420] = ~layer2_out[4866];
    assign layer3_out[4421] = ~(layer2_out[812] ^ layer2_out[813]);
    assign layer3_out[4422] = ~(layer2_out[2432] | layer2_out[2433]);
    assign layer3_out[4423] = ~layer2_out[897];
    assign layer3_out[4424] = ~(layer2_out[3686] & layer2_out[3687]);
    assign layer3_out[4425] = ~layer2_out[2891];
    assign layer3_out[4426] = ~layer2_out[2980] | layer2_out[2981];
    assign layer3_out[4427] = ~(layer2_out[5841] | layer2_out[5842]);
    assign layer3_out[4428] = ~layer2_out[126] | layer2_out[125];
    assign layer3_out[4429] = ~layer2_out[4639];
    assign layer3_out[4430] = ~(layer2_out[876] | layer2_out[877]);
    assign layer3_out[4431] = ~layer2_out[1637];
    assign layer3_out[4432] = ~layer2_out[5817] | layer2_out[5816];
    assign layer3_out[4433] = layer2_out[446];
    assign layer3_out[4434] = layer2_out[435] & ~layer2_out[434];
    assign layer3_out[4435] = layer2_out[1089] & ~layer2_out[1090];
    assign layer3_out[4436] = layer2_out[729] | layer2_out[730];
    assign layer3_out[4437] = ~layer2_out[16];
    assign layer3_out[4438] = ~layer2_out[2645];
    assign layer3_out[4439] = layer2_out[5132];
    assign layer3_out[4440] = layer2_out[1579] & ~layer2_out[1578];
    assign layer3_out[4441] = ~layer2_out[4619] | layer2_out[4620];
    assign layer3_out[4442] = ~(layer2_out[561] & layer2_out[562]);
    assign layer3_out[4443] = ~layer2_out[5883];
    assign layer3_out[4444] = ~layer2_out[6718];
    assign layer3_out[4445] = ~(layer2_out[7271] | layer2_out[7272]);
    assign layer3_out[4446] = ~(layer2_out[3319] | layer2_out[3320]);
    assign layer3_out[4447] = ~(layer2_out[4119] & layer2_out[4120]);
    assign layer3_out[4448] = layer2_out[6610];
    assign layer3_out[4449] = layer2_out[6232];
    assign layer3_out[4450] = layer2_out[7313] ^ layer2_out[7314];
    assign layer3_out[4451] = ~(layer2_out[3584] & layer2_out[3585]);
    assign layer3_out[4452] = layer2_out[7760];
    assign layer3_out[4453] = ~(layer2_out[2612] ^ layer2_out[2613]);
    assign layer3_out[4454] = layer2_out[2737];
    assign layer3_out[4455] = ~layer2_out[4824];
    assign layer3_out[4456] = layer2_out[2630] | layer2_out[2631];
    assign layer3_out[4457] = ~layer2_out[5174] | layer2_out[5173];
    assign layer3_out[4458] = layer2_out[2258] & ~layer2_out[2257];
    assign layer3_out[4459] = layer2_out[2039];
    assign layer3_out[4460] = ~layer2_out[5474] | layer2_out[5473];
    assign layer3_out[4461] = layer2_out[787];
    assign layer3_out[4462] = ~(layer2_out[2651] ^ layer2_out[2652]);
    assign layer3_out[4463] = ~layer2_out[3950] | layer2_out[3949];
    assign layer3_out[4464] = ~layer2_out[502];
    assign layer3_out[4465] = ~layer2_out[3233];
    assign layer3_out[4466] = ~layer2_out[6075];
    assign layer3_out[4467] = ~layer2_out[3665] | layer2_out[3666];
    assign layer3_out[4468] = ~(layer2_out[4211] & layer2_out[4212]);
    assign layer3_out[4469] = ~layer2_out[4471] | layer2_out[4472];
    assign layer3_out[4470] = ~layer2_out[7608];
    assign layer3_out[4471] = layer2_out[1939] & ~layer2_out[1938];
    assign layer3_out[4472] = ~(layer2_out[126] & layer2_out[127]);
    assign layer3_out[4473] = layer2_out[4394] & ~layer2_out[4393];
    assign layer3_out[4474] = layer2_out[576] ^ layer2_out[577];
    assign layer3_out[4475] = layer2_out[1776] & ~layer2_out[1777];
    assign layer3_out[4476] = ~(layer2_out[6022] & layer2_out[6023]);
    assign layer3_out[4477] = layer2_out[7120] | layer2_out[7121];
    assign layer3_out[4478] = layer2_out[1562];
    assign layer3_out[4479] = layer2_out[5754];
    assign layer3_out[4480] = ~layer2_out[312] | layer2_out[313];
    assign layer3_out[4481] = layer2_out[3824] ^ layer2_out[3825];
    assign layer3_out[4482] = ~(layer2_out[1] | layer2_out[2]);
    assign layer3_out[4483] = layer2_out[830];
    assign layer3_out[4484] = ~(layer2_out[3436] & layer2_out[3437]);
    assign layer3_out[4485] = ~layer2_out[7357] | layer2_out[7356];
    assign layer3_out[4486] = ~(layer2_out[5748] ^ layer2_out[5749]);
    assign layer3_out[4487] = layer2_out[3301] & layer2_out[3302];
    assign layer3_out[4488] = layer2_out[5513] | layer2_out[5514];
    assign layer3_out[4489] = ~(layer2_out[3171] | layer2_out[3172]);
    assign layer3_out[4490] = layer2_out[4087];
    assign layer3_out[4491] = ~(layer2_out[906] ^ layer2_out[907]);
    assign layer3_out[4492] = layer2_out[2226] ^ layer2_out[2227];
    assign layer3_out[4493] = ~layer2_out[3800];
    assign layer3_out[4494] = ~(layer2_out[4076] & layer2_out[4077]);
    assign layer3_out[4495] = ~layer2_out[5479];
    assign layer3_out[4496] = ~layer2_out[5518];
    assign layer3_out[4497] = ~layer2_out[615];
    assign layer3_out[4498] = layer2_out[6375];
    assign layer3_out[4499] = ~(layer2_out[1336] & layer2_out[1337]);
    assign layer3_out[4500] = ~layer2_out[6706] | layer2_out[6707];
    assign layer3_out[4501] = ~layer2_out[6715];
    assign layer3_out[4502] = layer2_out[3890];
    assign layer3_out[4503] = ~layer2_out[3226];
    assign layer3_out[4504] = layer2_out[5697] & ~layer2_out[5696];
    assign layer3_out[4505] = ~(layer2_out[5185] | layer2_out[5186]);
    assign layer3_out[4506] = ~(layer2_out[2125] & layer2_out[2126]);
    assign layer3_out[4507] = layer2_out[5231] & ~layer2_out[5230];
    assign layer3_out[4508] = layer2_out[2574];
    assign layer3_out[4509] = ~layer2_out[1559];
    assign layer3_out[4510] = ~(layer2_out[1307] ^ layer2_out[1308]);
    assign layer3_out[4511] = layer2_out[3526] | layer2_out[3527];
    assign layer3_out[4512] = ~layer2_out[7162] | layer2_out[7163];
    assign layer3_out[4513] = ~layer2_out[1316];
    assign layer3_out[4514] = layer2_out[7338];
    assign layer3_out[4515] = layer2_out[7440] & layer2_out[7441];
    assign layer3_out[4516] = ~layer2_out[1082] | layer2_out[1083];
    assign layer3_out[4517] = layer2_out[3060];
    assign layer3_out[4518] = layer2_out[6364];
    assign layer3_out[4519] = ~layer2_out[140];
    assign layer3_out[4520] = layer2_out[2948] & ~layer2_out[2949];
    assign layer3_out[4521] = ~layer2_out[1519];
    assign layer3_out[4522] = layer2_out[2451] ^ layer2_out[2452];
    assign layer3_out[4523] = ~layer2_out[4632] | layer2_out[4631];
    assign layer3_out[4524] = ~layer2_out[1784];
    assign layer3_out[4525] = ~layer2_out[5513] | layer2_out[5512];
    assign layer3_out[4526] = ~layer2_out[1976];
    assign layer3_out[4527] = layer2_out[110];
    assign layer3_out[4528] = ~layer2_out[1929];
    assign layer3_out[4529] = ~layer2_out[3675];
    assign layer3_out[4530] = ~layer2_out[3536];
    assign layer3_out[4531] = ~layer2_out[7908];
    assign layer3_out[4532] = layer2_out[5292] & ~layer2_out[5291];
    assign layer3_out[4533] = layer2_out[3908] & ~layer2_out[3909];
    assign layer3_out[4534] = ~(layer2_out[2560] | layer2_out[2561]);
    assign layer3_out[4535] = layer2_out[2977];
    assign layer3_out[4536] = layer2_out[500] ^ layer2_out[501];
    assign layer3_out[4537] = ~layer2_out[24];
    assign layer3_out[4538] = ~layer2_out[390] | layer2_out[391];
    assign layer3_out[4539] = ~layer2_out[7768] | layer2_out[7767];
    assign layer3_out[4540] = ~(layer2_out[3131] ^ layer2_out[3132]);
    assign layer3_out[4541] = ~layer2_out[5015];
    assign layer3_out[4542] = ~(layer2_out[6970] ^ layer2_out[6971]);
    assign layer3_out[4543] = ~layer2_out[6341] | layer2_out[6340];
    assign layer3_out[4544] = ~layer2_out[2105] | layer2_out[2106];
    assign layer3_out[4545] = ~(layer2_out[5040] | layer2_out[5041]);
    assign layer3_out[4546] = layer2_out[6813] | layer2_out[6814];
    assign layer3_out[4547] = layer2_out[846] | layer2_out[847];
    assign layer3_out[4548] = layer2_out[1252] | layer2_out[1253];
    assign layer3_out[4549] = ~(layer2_out[3193] & layer2_out[3194]);
    assign layer3_out[4550] = ~layer2_out[1619] | layer2_out[1618];
    assign layer3_out[4551] = 1'b0;
    assign layer3_out[4552] = ~layer2_out[5512];
    assign layer3_out[4553] = 1'b0;
    assign layer3_out[4554] = layer2_out[5323] & ~layer2_out[5324];
    assign layer3_out[4555] = layer2_out[3764] & ~layer2_out[3765];
    assign layer3_out[4556] = layer2_out[5482];
    assign layer3_out[4557] = ~layer2_out[4918];
    assign layer3_out[4558] = layer2_out[2253] & layer2_out[2254];
    assign layer3_out[4559] = layer2_out[7967] | layer2_out[7968];
    assign layer3_out[4560] = ~(layer2_out[6483] | layer2_out[6484]);
    assign layer3_out[4561] = layer2_out[331];
    assign layer3_out[4562] = layer2_out[6393] & layer2_out[6394];
    assign layer3_out[4563] = 1'b1;
    assign layer3_out[4564] = ~layer2_out[1387];
    assign layer3_out[4565] = ~layer2_out[3617];
    assign layer3_out[4566] = layer2_out[1441] & ~layer2_out[1442];
    assign layer3_out[4567] = layer2_out[4267] & ~layer2_out[4268];
    assign layer3_out[4568] = ~(layer2_out[2750] & layer2_out[2751]);
    assign layer3_out[4569] = layer2_out[2858] & ~layer2_out[2859];
    assign layer3_out[4570] = ~layer2_out[7853] | layer2_out[7852];
    assign layer3_out[4571] = layer2_out[1196];
    assign layer3_out[4572] = layer2_out[499] ^ layer2_out[500];
    assign layer3_out[4573] = ~layer2_out[790];
    assign layer3_out[4574] = layer2_out[5864];
    assign layer3_out[4575] = layer2_out[3511] & ~layer2_out[3512];
    assign layer3_out[4576] = layer2_out[5163];
    assign layer3_out[4577] = layer2_out[2470] & ~layer2_out[2471];
    assign layer3_out[4578] = ~(layer2_out[7809] ^ layer2_out[7810]);
    assign layer3_out[4579] = layer2_out[5607];
    assign layer3_out[4580] = layer2_out[4440];
    assign layer3_out[4581] = layer2_out[3442];
    assign layer3_out[4582] = ~layer2_out[2152];
    assign layer3_out[4583] = layer2_out[5519];
    assign layer3_out[4584] = ~layer2_out[4354];
    assign layer3_out[4585] = layer2_out[2837] & ~layer2_out[2838];
    assign layer3_out[4586] = ~layer2_out[4551] | layer2_out[4550];
    assign layer3_out[4587] = layer2_out[4384] & ~layer2_out[4385];
    assign layer3_out[4588] = ~layer2_out[427];
    assign layer3_out[4589] = ~layer2_out[7461];
    assign layer3_out[4590] = layer2_out[4621] & layer2_out[4622];
    assign layer3_out[4591] = ~layer2_out[6269];
    assign layer3_out[4592] = ~(layer2_out[6980] ^ layer2_out[6981]);
    assign layer3_out[4593] = layer2_out[5976] & ~layer2_out[5977];
    assign layer3_out[4594] = layer2_out[92] & layer2_out[93];
    assign layer3_out[4595] = layer2_out[4221];
    assign layer3_out[4596] = ~layer2_out[6572] | layer2_out[6573];
    assign layer3_out[4597] = layer2_out[2354] | layer2_out[2355];
    assign layer3_out[4598] = layer2_out[4661] & ~layer2_out[4660];
    assign layer3_out[4599] = ~layer2_out[2154] | layer2_out[2153];
    assign layer3_out[4600] = layer2_out[2004];
    assign layer3_out[4601] = ~layer2_out[4329];
    assign layer3_out[4602] = layer2_out[5394];
    assign layer3_out[4603] = layer2_out[515] & layer2_out[516];
    assign layer3_out[4604] = layer2_out[3816];
    assign layer3_out[4605] = ~layer2_out[2746] | layer2_out[2747];
    assign layer3_out[4606] = layer2_out[2071] & ~layer2_out[2070];
    assign layer3_out[4607] = layer2_out[3089];
    assign layer3_out[4608] = layer2_out[5941] | layer2_out[5942];
    assign layer3_out[4609] = layer2_out[1882];
    assign layer3_out[4610] = layer2_out[5657] ^ layer2_out[5658];
    assign layer3_out[4611] = ~(layer2_out[7201] ^ layer2_out[7202]);
    assign layer3_out[4612] = layer2_out[2895] & ~layer2_out[2896];
    assign layer3_out[4613] = ~layer2_out[4969];
    assign layer3_out[4614] = layer2_out[3961] | layer2_out[3962];
    assign layer3_out[4615] = layer2_out[5746];
    assign layer3_out[4616] = layer2_out[1791] & layer2_out[1792];
    assign layer3_out[4617] = ~layer2_out[4164] | layer2_out[4165];
    assign layer3_out[4618] = ~layer2_out[1135] | layer2_out[1136];
    assign layer3_out[4619] = layer2_out[4815] ^ layer2_out[4816];
    assign layer3_out[4620] = layer2_out[6665] | layer2_out[6666];
    assign layer3_out[4621] = ~layer2_out[7264] | layer2_out[7263];
    assign layer3_out[4622] = ~layer2_out[2876];
    assign layer3_out[4623] = ~layer2_out[630];
    assign layer3_out[4624] = ~layer2_out[7982] | layer2_out[7983];
    assign layer3_out[4625] = layer2_out[3163] | layer2_out[3164];
    assign layer3_out[4626] = layer2_out[7487];
    assign layer3_out[4627] = layer2_out[1294];
    assign layer3_out[4628] = 1'b1;
    assign layer3_out[4629] = layer2_out[4898];
    assign layer3_out[4630] = ~(layer2_out[5499] | layer2_out[5500]);
    assign layer3_out[4631] = layer2_out[2283];
    assign layer3_out[4632] = ~layer2_out[6032];
    assign layer3_out[4633] = layer2_out[1743] & layer2_out[1744];
    assign layer3_out[4634] = layer2_out[4416];
    assign layer3_out[4635] = ~(layer2_out[4360] | layer2_out[4361]);
    assign layer3_out[4636] = ~(layer2_out[2437] & layer2_out[2438]);
    assign layer3_out[4637] = layer2_out[748] & ~layer2_out[747];
    assign layer3_out[4638] = ~layer2_out[4949] | layer2_out[4950];
    assign layer3_out[4639] = layer2_out[6081] & ~layer2_out[6082];
    assign layer3_out[4640] = ~layer2_out[5987];
    assign layer3_out[4641] = layer2_out[7853] & layer2_out[7854];
    assign layer3_out[4642] = ~layer2_out[5506] | layer2_out[5505];
    assign layer3_out[4643] = ~(layer2_out[3514] ^ layer2_out[3515]);
    assign layer3_out[4644] = ~layer2_out[5518];
    assign layer3_out[4645] = ~(layer2_out[3606] ^ layer2_out[3607]);
    assign layer3_out[4646] = layer2_out[1079] & ~layer2_out[1080];
    assign layer3_out[4647] = 1'b1;
    assign layer3_out[4648] = layer2_out[5919];
    assign layer3_out[4649] = ~layer2_out[1411] | layer2_out[1412];
    assign layer3_out[4650] = ~layer2_out[4673];
    assign layer3_out[4651] = layer2_out[7988];
    assign layer3_out[4652] = ~layer2_out[3137];
    assign layer3_out[4653] = ~layer2_out[1373];
    assign layer3_out[4654] = layer2_out[6827];
    assign layer3_out[4655] = ~layer2_out[5111] | layer2_out[5112];
    assign layer3_out[4656] = ~layer2_out[6273] | layer2_out[6274];
    assign layer3_out[4657] = layer2_out[3992];
    assign layer3_out[4658] = layer2_out[1950];
    assign layer3_out[4659] = layer2_out[1014];
    assign layer3_out[4660] = ~(layer2_out[205] ^ layer2_out[206]);
    assign layer3_out[4661] = layer2_out[6832];
    assign layer3_out[4662] = ~(layer2_out[7413] & layer2_out[7414]);
    assign layer3_out[4663] = layer2_out[7008] & layer2_out[7009];
    assign layer3_out[4664] = layer2_out[4749] & ~layer2_out[4750];
    assign layer3_out[4665] = ~(layer2_out[87] | layer2_out[88]);
    assign layer3_out[4666] = ~layer2_out[4718] | layer2_out[4717];
    assign layer3_out[4667] = layer2_out[805] | layer2_out[806];
    assign layer3_out[4668] = layer2_out[6690];
    assign layer3_out[4669] = layer2_out[3627];
    assign layer3_out[4670] = ~layer2_out[4145] | layer2_out[4144];
    assign layer3_out[4671] = layer2_out[266];
    assign layer3_out[4672] = layer2_out[5557];
    assign layer3_out[4673] = layer2_out[6514] | layer2_out[6515];
    assign layer3_out[4674] = layer2_out[4291];
    assign layer3_out[4675] = ~layer2_out[3621];
    assign layer3_out[4676] = layer2_out[4] | layer2_out[5];
    assign layer3_out[4677] = ~(layer2_out[2445] | layer2_out[2446]);
    assign layer3_out[4678] = layer2_out[809] & ~layer2_out[808];
    assign layer3_out[4679] = ~(layer2_out[3595] ^ layer2_out[3596]);
    assign layer3_out[4680] = layer2_out[4554] & ~layer2_out[4553];
    assign layer3_out[4681] = layer2_out[6734] & ~layer2_out[6733];
    assign layer3_out[4682] = layer2_out[1585] & layer2_out[1586];
    assign layer3_out[4683] = ~layer2_out[4662];
    assign layer3_out[4684] = ~(layer2_out[6758] & layer2_out[6759]);
    assign layer3_out[4685] = ~(layer2_out[5550] & layer2_out[5551]);
    assign layer3_out[4686] = ~layer2_out[4751];
    assign layer3_out[4687] = ~(layer2_out[6029] & layer2_out[6030]);
    assign layer3_out[4688] = layer2_out[5814] & ~layer2_out[5813];
    assign layer3_out[4689] = ~layer2_out[2312];
    assign layer3_out[4690] = layer2_out[220] ^ layer2_out[221];
    assign layer3_out[4691] = layer2_out[2814] ^ layer2_out[2815];
    assign layer3_out[4692] = ~layer2_out[5083];
    assign layer3_out[4693] = ~(layer2_out[3352] | layer2_out[3353]);
    assign layer3_out[4694] = ~layer2_out[6562];
    assign layer3_out[4695] = layer2_out[4173];
    assign layer3_out[4696] = layer2_out[7382];
    assign layer3_out[4697] = ~layer2_out[6227];
    assign layer3_out[4698] = ~layer2_out[3137];
    assign layer3_out[4699] = layer2_out[4014] & ~layer2_out[4013];
    assign layer3_out[4700] = ~(layer2_out[772] | layer2_out[773]);
    assign layer3_out[4701] = layer2_out[930] & layer2_out[931];
    assign layer3_out[4702] = ~(layer2_out[2350] & layer2_out[2351]);
    assign layer3_out[4703] = ~layer2_out[3207];
    assign layer3_out[4704] = ~layer2_out[1320] | layer2_out[1319];
    assign layer3_out[4705] = layer2_out[3724] & layer2_out[3725];
    assign layer3_out[4706] = layer2_out[4155] & ~layer2_out[4154];
    assign layer3_out[4707] = ~layer2_out[3125] | layer2_out[3124];
    assign layer3_out[4708] = ~(layer2_out[5364] & layer2_out[5365]);
    assign layer3_out[4709] = layer2_out[6785] & ~layer2_out[6786];
    assign layer3_out[4710] = ~layer2_out[3733] | layer2_out[3732];
    assign layer3_out[4711] = ~layer2_out[5703];
    assign layer3_out[4712] = ~(layer2_out[3523] & layer2_out[3524]);
    assign layer3_out[4713] = layer2_out[868] & ~layer2_out[869];
    assign layer3_out[4714] = layer2_out[4053] ^ layer2_out[4054];
    assign layer3_out[4715] = ~layer2_out[224] | layer2_out[223];
    assign layer3_out[4716] = ~layer2_out[419];
    assign layer3_out[4717] = ~layer2_out[5536];
    assign layer3_out[4718] = layer2_out[6921];
    assign layer3_out[4719] = ~layer2_out[827];
    assign layer3_out[4720] = layer2_out[4955] & layer2_out[4956];
    assign layer3_out[4721] = layer2_out[7520];
    assign layer3_out[4722] = ~layer2_out[2340];
    assign layer3_out[4723] = 1'b0;
    assign layer3_out[4724] = ~(layer2_out[7975] & layer2_out[7976]);
    assign layer3_out[4725] = ~(layer2_out[6344] | layer2_out[6345]);
    assign layer3_out[4726] = layer2_out[4321];
    assign layer3_out[4727] = layer2_out[2887] & ~layer2_out[2888];
    assign layer3_out[4728] = ~(layer2_out[2255] | layer2_out[2256]);
    assign layer3_out[4729] = ~layer2_out[304] | layer2_out[303];
    assign layer3_out[4730] = layer2_out[4262];
    assign layer3_out[4731] = ~layer2_out[2177];
    assign layer3_out[4732] = ~layer2_out[20] | layer2_out[19];
    assign layer3_out[4733] = ~layer2_out[6865];
    assign layer3_out[4734] = layer2_out[2506] & layer2_out[2507];
    assign layer3_out[4735] = ~(layer2_out[7711] & layer2_out[7712]);
    assign layer3_out[4736] = ~layer2_out[2457];
    assign layer3_out[4737] = ~layer2_out[54] | layer2_out[53];
    assign layer3_out[4738] = layer2_out[2050];
    assign layer3_out[4739] = ~(layer2_out[416] ^ layer2_out[417]);
    assign layer3_out[4740] = layer2_out[2621] & ~layer2_out[2620];
    assign layer3_out[4741] = layer2_out[4237] & ~layer2_out[4236];
    assign layer3_out[4742] = ~layer2_out[2779];
    assign layer3_out[4743] = ~(layer2_out[1463] ^ layer2_out[1464]);
    assign layer3_out[4744] = layer2_out[868] & ~layer2_out[867];
    assign layer3_out[4745] = ~layer2_out[5188] | layer2_out[5187];
    assign layer3_out[4746] = ~layer2_out[5653] | layer2_out[5654];
    assign layer3_out[4747] = layer2_out[3867] & ~layer2_out[3868];
    assign layer3_out[4748] = layer2_out[5199] | layer2_out[5200];
    assign layer3_out[4749] = layer2_out[4568];
    assign layer3_out[4750] = ~layer2_out[7090] | layer2_out[7091];
    assign layer3_out[4751] = ~(layer2_out[3489] ^ layer2_out[3490]);
    assign layer3_out[4752] = ~(layer2_out[4519] & layer2_out[4520]);
    assign layer3_out[4753] = layer2_out[7152] | layer2_out[7153];
    assign layer3_out[4754] = layer2_out[6897] & layer2_out[6898];
    assign layer3_out[4755] = ~(layer2_out[6732] | layer2_out[6733]);
    assign layer3_out[4756] = layer2_out[2245] | layer2_out[2246];
    assign layer3_out[4757] = ~layer2_out[3491] | layer2_out[3492];
    assign layer3_out[4758] = ~layer2_out[233];
    assign layer3_out[4759] = layer2_out[4132] & ~layer2_out[4131];
    assign layer3_out[4760] = layer2_out[7156] ^ layer2_out[7157];
    assign layer3_out[4761] = layer2_out[7267];
    assign layer3_out[4762] = ~layer2_out[2713];
    assign layer3_out[4763] = layer2_out[5581] & layer2_out[5582];
    assign layer3_out[4764] = ~layer2_out[6872] | layer2_out[6873];
    assign layer3_out[4765] = ~(layer2_out[2775] | layer2_out[2776]);
    assign layer3_out[4766] = ~layer2_out[5570];
    assign layer3_out[4767] = ~layer2_out[2839];
    assign layer3_out[4768] = layer2_out[1238];
    assign layer3_out[4769] = layer2_out[4774];
    assign layer3_out[4770] = layer2_out[4547];
    assign layer3_out[4771] = layer2_out[1875];
    assign layer3_out[4772] = ~layer2_out[5077];
    assign layer3_out[4773] = ~layer2_out[1948] | layer2_out[1949];
    assign layer3_out[4774] = layer2_out[2022] & ~layer2_out[2021];
    assign layer3_out[4775] = ~layer2_out[2594];
    assign layer3_out[4776] = ~layer2_out[3203] | layer2_out[3202];
    assign layer3_out[4777] = ~layer2_out[7526] | layer2_out[7525];
    assign layer3_out[4778] = layer2_out[2014];
    assign layer3_out[4779] = 1'b0;
    assign layer3_out[4780] = ~layer2_out[3166];
    assign layer3_out[4781] = layer2_out[4541];
    assign layer3_out[4782] = ~layer2_out[4982];
    assign layer3_out[4783] = ~layer2_out[4811];
    assign layer3_out[4784] = ~(layer2_out[6798] & layer2_out[6799]);
    assign layer3_out[4785] = ~layer2_out[7786];
    assign layer3_out[4786] = ~layer2_out[182] | layer2_out[181];
    assign layer3_out[4787] = ~layer2_out[389];
    assign layer3_out[4788] = ~layer2_out[3950] | layer2_out[3951];
    assign layer3_out[4789] = ~(layer2_out[177] & layer2_out[178]);
    assign layer3_out[4790] = layer2_out[1178];
    assign layer3_out[4791] = layer2_out[1602] & ~layer2_out[1603];
    assign layer3_out[4792] = layer2_out[78] & layer2_out[79];
    assign layer3_out[4793] = layer2_out[6011];
    assign layer3_out[4794] = ~layer2_out[3002];
    assign layer3_out[4795] = layer2_out[520];
    assign layer3_out[4796] = layer2_out[2885] & ~layer2_out[2886];
    assign layer3_out[4797] = ~layer2_out[7498] | layer2_out[7497];
    assign layer3_out[4798] = layer2_out[5034];
    assign layer3_out[4799] = layer2_out[2602] & ~layer2_out[2601];
    assign layer3_out[4800] = ~(layer2_out[5565] ^ layer2_out[5566]);
    assign layer3_out[4801] = ~(layer2_out[6600] | layer2_out[6601]);
    assign layer3_out[4802] = layer2_out[6135] | layer2_out[6136];
    assign layer3_out[4803] = ~layer2_out[2194];
    assign layer3_out[4804] = layer2_out[691] & ~layer2_out[690];
    assign layer3_out[4805] = ~layer2_out[2142];
    assign layer3_out[4806] = layer2_out[7158];
    assign layer3_out[4807] = layer2_out[3965] ^ layer2_out[3966];
    assign layer3_out[4808] = layer2_out[642] ^ layer2_out[643];
    assign layer3_out[4809] = ~layer2_out[742];
    assign layer3_out[4810] = layer2_out[879] ^ layer2_out[880];
    assign layer3_out[4811] = ~layer2_out[737];
    assign layer3_out[4812] = ~(layer2_out[4606] ^ layer2_out[4607]);
    assign layer3_out[4813] = ~(layer2_out[2622] & layer2_out[2623]);
    assign layer3_out[4814] = ~(layer2_out[387] ^ layer2_out[388]);
    assign layer3_out[4815] = layer2_out[299];
    assign layer3_out[4816] = ~(layer2_out[3254] ^ layer2_out[3255]);
    assign layer3_out[4817] = layer2_out[1617] | layer2_out[1618];
    assign layer3_out[4818] = ~(layer2_out[4008] & layer2_out[4009]);
    assign layer3_out[4819] = layer2_out[4333] & ~layer2_out[4334];
    assign layer3_out[4820] = ~layer2_out[7304];
    assign layer3_out[4821] = 1'b0;
    assign layer3_out[4822] = layer2_out[2061];
    assign layer3_out[4823] = layer2_out[1991];
    assign layer3_out[4824] = layer2_out[4188] & ~layer2_out[4189];
    assign layer3_out[4825] = layer2_out[1890];
    assign layer3_out[4826] = ~(layer2_out[7557] | layer2_out[7558]);
    assign layer3_out[4827] = layer2_out[4374];
    assign layer3_out[4828] = 1'b0;
    assign layer3_out[4829] = ~layer2_out[6820];
    assign layer3_out[4830] = layer2_out[7948] ^ layer2_out[7949];
    assign layer3_out[4831] = layer2_out[6857] | layer2_out[6858];
    assign layer3_out[4832] = ~layer2_out[2271];
    assign layer3_out[4833] = layer2_out[4752] ^ layer2_out[4753];
    assign layer3_out[4834] = 1'b1;
    assign layer3_out[4835] = layer2_out[2107];
    assign layer3_out[4836] = layer2_out[2786];
    assign layer3_out[4837] = layer2_out[680] | layer2_out[681];
    assign layer3_out[4838] = ~layer2_out[5009];
    assign layer3_out[4839] = ~layer2_out[3993];
    assign layer3_out[4840] = layer2_out[722];
    assign layer3_out[4841] = ~(layer2_out[5637] | layer2_out[5638]);
    assign layer3_out[4842] = ~(layer2_out[7137] ^ layer2_out[7138]);
    assign layer3_out[4843] = layer2_out[709];
    assign layer3_out[4844] = layer2_out[6827];
    assign layer3_out[4845] = ~layer2_out[1902];
    assign layer3_out[4846] = layer2_out[3984];
    assign layer3_out[4847] = layer2_out[4154];
    assign layer3_out[4848] = ~layer2_out[4901] | layer2_out[4900];
    assign layer3_out[4849] = layer2_out[7491] | layer2_out[7492];
    assign layer3_out[4850] = layer2_out[625] ^ layer2_out[626];
    assign layer3_out[4851] = layer2_out[7762] & layer2_out[7763];
    assign layer3_out[4852] = ~(layer2_out[5665] | layer2_out[5666]);
    assign layer3_out[4853] = layer2_out[3619] & ~layer2_out[3618];
    assign layer3_out[4854] = layer2_out[4699] & ~layer2_out[4700];
    assign layer3_out[4855] = layer2_out[3121] & ~layer2_out[3120];
    assign layer3_out[4856] = layer2_out[3306] ^ layer2_out[3307];
    assign layer3_out[4857] = ~layer2_out[7682];
    assign layer3_out[4858] = layer2_out[1810] ^ layer2_out[1811];
    assign layer3_out[4859] = layer2_out[948] & ~layer2_out[949];
    assign layer3_out[4860] = ~layer2_out[4575];
    assign layer3_out[4861] = layer2_out[7023] & ~layer2_out[7022];
    assign layer3_out[4862] = layer2_out[5828] & ~layer2_out[5829];
    assign layer3_out[4863] = layer2_out[6224] & ~layer2_out[6225];
    assign layer3_out[4864] = layer2_out[804] & ~layer2_out[805];
    assign layer3_out[4865] = layer2_out[2086] & ~layer2_out[2087];
    assign layer3_out[4866] = layer2_out[6796] | layer2_out[6797];
    assign layer3_out[4867] = layer2_out[1277];
    assign layer3_out[4868] = ~layer2_out[1574];
    assign layer3_out[4869] = ~(layer2_out[7072] ^ layer2_out[7073]);
    assign layer3_out[4870] = ~layer2_out[5906];
    assign layer3_out[4871] = ~layer2_out[5849] | layer2_out[5848];
    assign layer3_out[4872] = ~layer2_out[3955];
    assign layer3_out[4873] = layer2_out[1391] & ~layer2_out[1392];
    assign layer3_out[4874] = layer2_out[7735];
    assign layer3_out[4875] = layer2_out[5438] & ~layer2_out[5439];
    assign layer3_out[4876] = layer2_out[1044];
    assign layer3_out[4877] = layer2_out[3153];
    assign layer3_out[4878] = layer2_out[4604] & ~layer2_out[4603];
    assign layer3_out[4879] = layer2_out[5800] & ~layer2_out[5799];
    assign layer3_out[4880] = layer2_out[537] & ~layer2_out[536];
    assign layer3_out[4881] = ~layer2_out[607] | layer2_out[606];
    assign layer3_out[4882] = layer2_out[6760] & layer2_out[6761];
    assign layer3_out[4883] = ~(layer2_out[1099] & layer2_out[1100]);
    assign layer3_out[4884] = layer2_out[2138];
    assign layer3_out[4885] = ~layer2_out[1985];
    assign layer3_out[4886] = 1'b1;
    assign layer3_out[4887] = ~layer2_out[701];
    assign layer3_out[4888] = ~(layer2_out[3639] | layer2_out[3640]);
    assign layer3_out[4889] = layer2_out[1530] & ~layer2_out[1529];
    assign layer3_out[4890] = ~(layer2_out[4875] | layer2_out[4876]);
    assign layer3_out[4891] = layer2_out[5713] ^ layer2_out[5714];
    assign layer3_out[4892] = layer2_out[4293] & ~layer2_out[4294];
    assign layer3_out[4893] = layer2_out[7092];
    assign layer3_out[4894] = layer2_out[5709];
    assign layer3_out[4895] = layer2_out[6460];
    assign layer3_out[4896] = ~(layer2_out[6109] ^ layer2_out[6110]);
    assign layer3_out[4897] = ~layer2_out[5376];
    assign layer3_out[4898] = ~(layer2_out[7434] & layer2_out[7435]);
    assign layer3_out[4899] = layer2_out[4846];
    assign layer3_out[4900] = ~layer2_out[5809] | layer2_out[5808];
    assign layer3_out[4901] = ~(layer2_out[3608] ^ layer2_out[3609]);
    assign layer3_out[4902] = layer2_out[680] & ~layer2_out[679];
    assign layer3_out[4903] = layer2_out[3377] & ~layer2_out[3376];
    assign layer3_out[4904] = layer2_out[5276] | layer2_out[5277];
    assign layer3_out[4905] = layer2_out[4551] & layer2_out[4552];
    assign layer3_out[4906] = ~layer2_out[5190];
    assign layer3_out[4907] = ~layer2_out[6013];
    assign layer3_out[4908] = ~layer2_out[1325] | layer2_out[1326];
    assign layer3_out[4909] = ~layer2_out[7246];
    assign layer3_out[4910] = ~layer2_out[782];
    assign layer3_out[4911] = ~layer2_out[2499] | layer2_out[2498];
    assign layer3_out[4912] = layer2_out[1218];
    assign layer3_out[4913] = layer2_out[3281];
    assign layer3_out[4914] = ~layer2_out[5443];
    assign layer3_out[4915] = layer2_out[2798] | layer2_out[2799];
    assign layer3_out[4916] = ~layer2_out[3930] | layer2_out[3929];
    assign layer3_out[4917] = ~(layer2_out[7032] ^ layer2_out[7033]);
    assign layer3_out[4918] = layer2_out[3295];
    assign layer3_out[4919] = layer2_out[5481] & ~layer2_out[5480];
    assign layer3_out[4920] = layer2_out[7813] & ~layer2_out[7812];
    assign layer3_out[4921] = 1'b0;
    assign layer3_out[4922] = layer2_out[1421] & ~layer2_out[1420];
    assign layer3_out[4923] = ~(layer2_out[7854] | layer2_out[7855]);
    assign layer3_out[4924] = layer2_out[6139] ^ layer2_out[6140];
    assign layer3_out[4925] = ~layer2_out[2083];
    assign layer3_out[4926] = ~layer2_out[2691];
    assign layer3_out[4927] = 1'b0;
    assign layer3_out[4928] = layer2_out[4916];
    assign layer3_out[4929] = 1'b0;
    assign layer3_out[4930] = layer2_out[5001] ^ layer2_out[5002];
    assign layer3_out[4931] = layer2_out[6330];
    assign layer3_out[4932] = ~(layer2_out[3821] & layer2_out[3822]);
    assign layer3_out[4933] = layer2_out[1728] & layer2_out[1729];
    assign layer3_out[4934] = ~layer2_out[7119];
    assign layer3_out[4935] = layer2_out[5533] & ~layer2_out[5532];
    assign layer3_out[4936] = ~layer2_out[7455] | layer2_out[7454];
    assign layer3_out[4937] = ~layer2_out[6621];
    assign layer3_out[4938] = layer2_out[3020] ^ layer2_out[3021];
    assign layer3_out[4939] = layer2_out[2483] | layer2_out[2484];
    assign layer3_out[4940] = layer2_out[4520] ^ layer2_out[4521];
    assign layer3_out[4941] = layer2_out[5424];
    assign layer3_out[4942] = ~layer2_out[1071] | layer2_out[1070];
    assign layer3_out[4943] = ~layer2_out[2452];
    assign layer3_out[4944] = ~layer2_out[4772] | layer2_out[4773];
    assign layer3_out[4945] = layer2_out[7993];
    assign layer3_out[4946] = layer2_out[3221];
    assign layer3_out[4947] = layer2_out[5846];
    assign layer3_out[4948] = 1'b0;
    assign layer3_out[4949] = ~layer2_out[5260];
    assign layer3_out[4950] = layer2_out[608] & ~layer2_out[609];
    assign layer3_out[4951] = ~(layer2_out[7494] | layer2_out[7495]);
    assign layer3_out[4952] = ~(layer2_out[507] ^ layer2_out[508]);
    assign layer3_out[4953] = layer2_out[5618];
    assign layer3_out[4954] = layer2_out[4517];
    assign layer3_out[4955] = ~(layer2_out[1100] | layer2_out[1101]);
    assign layer3_out[4956] = layer2_out[3172] & layer2_out[3173];
    assign layer3_out[4957] = ~(layer2_out[7396] & layer2_out[7397]);
    assign layer3_out[4958] = layer2_out[4442];
    assign layer3_out[4959] = layer2_out[444];
    assign layer3_out[4960] = layer2_out[6662];
    assign layer3_out[4961] = 1'b0;
    assign layer3_out[4962] = ~(layer2_out[2522] & layer2_out[2523]);
    assign layer3_out[4963] = layer2_out[7249];
    assign layer3_out[4964] = layer2_out[6591] & layer2_out[6592];
    assign layer3_out[4965] = ~layer2_out[1839];
    assign layer3_out[4966] = layer2_out[3796] & layer2_out[3797];
    assign layer3_out[4967] = ~layer2_out[3851] | layer2_out[3850];
    assign layer3_out[4968] = layer2_out[612];
    assign layer3_out[4969] = ~(layer2_out[6422] ^ layer2_out[6423]);
    assign layer3_out[4970] = ~(layer2_out[6025] ^ layer2_out[6026]);
    assign layer3_out[4971] = ~layer2_out[7970];
    assign layer3_out[4972] = ~layer2_out[1918];
    assign layer3_out[4973] = layer2_out[5047];
    assign layer3_out[4974] = ~(layer2_out[2958] ^ layer2_out[2959]);
    assign layer3_out[4975] = ~(layer2_out[2974] & layer2_out[2975]);
    assign layer3_out[4976] = ~layer2_out[2034] | layer2_out[2033];
    assign layer3_out[4977] = ~(layer2_out[1969] | layer2_out[1970]);
    assign layer3_out[4978] = ~layer2_out[6043] | layer2_out[6042];
    assign layer3_out[4979] = layer2_out[1542] & ~layer2_out[1541];
    assign layer3_out[4980] = layer2_out[5198];
    assign layer3_out[4981] = layer2_out[7041];
    assign layer3_out[4982] = ~layer2_out[3496];
    assign layer3_out[4983] = layer2_out[3302] | layer2_out[3303];
    assign layer3_out[4984] = layer2_out[3466] & ~layer2_out[3465];
    assign layer3_out[4985] = ~layer2_out[5967];
    assign layer3_out[4986] = ~layer2_out[775];
    assign layer3_out[4987] = ~layer2_out[199];
    assign layer3_out[4988] = layer2_out[6352] & ~layer2_out[6353];
    assign layer3_out[4989] = ~layer2_out[1728] | layer2_out[1727];
    assign layer3_out[4990] = layer2_out[7271] & ~layer2_out[7270];
    assign layer3_out[4991] = ~layer2_out[7019] | layer2_out[7020];
    assign layer3_out[4992] = layer2_out[7029];
    assign layer3_out[4993] = layer2_out[1255] | layer2_out[1256];
    assign layer3_out[4994] = layer2_out[5243];
    assign layer3_out[4995] = ~(layer2_out[5105] | layer2_out[5106]);
    assign layer3_out[4996] = ~layer2_out[707];
    assign layer3_out[4997] = layer2_out[6468] | layer2_out[6469];
    assign layer3_out[4998] = ~layer2_out[7796] | layer2_out[7797];
    assign layer3_out[4999] = ~(layer2_out[7051] | layer2_out[7052]);
    assign layer3_out[5000] = ~(layer2_out[3109] | layer2_out[3110]);
    assign layer3_out[5001] = layer2_out[7598] ^ layer2_out[7599];
    assign layer3_out[5002] = ~layer2_out[772];
    assign layer3_out[5003] = ~layer2_out[5147] | layer2_out[5146];
    assign layer3_out[5004] = ~layer2_out[918];
    assign layer3_out[5005] = layer2_out[5322];
    assign layer3_out[5006] = ~layer2_out[7662] | layer2_out[7663];
    assign layer3_out[5007] = layer2_out[2678] | layer2_out[2679];
    assign layer3_out[5008] = layer2_out[5823] & ~layer2_out[5822];
    assign layer3_out[5009] = ~layer2_out[3975] | layer2_out[3974];
    assign layer3_out[5010] = layer2_out[4687];
    assign layer3_out[5011] = layer2_out[3385] & ~layer2_out[3386];
    assign layer3_out[5012] = ~layer2_out[7815];
    assign layer3_out[5013] = layer2_out[6464] ^ layer2_out[6465];
    assign layer3_out[5014] = ~layer2_out[3809];
    assign layer3_out[5015] = layer2_out[4777];
    assign layer3_out[5016] = layer2_out[861];
    assign layer3_out[5017] = layer2_out[3942] & layer2_out[3943];
    assign layer3_out[5018] = layer2_out[1226] & layer2_out[1227];
    assign layer3_out[5019] = layer2_out[1652];
    assign layer3_out[5020] = layer2_out[6619];
    assign layer3_out[5021] = ~layer2_out[1626];
    assign layer3_out[5022] = layer2_out[5196] & layer2_out[5197];
    assign layer3_out[5023] = ~layer2_out[4347];
    assign layer3_out[5024] = ~layer2_out[5903];
    assign layer3_out[5025] = layer2_out[3932] & ~layer2_out[3931];
    assign layer3_out[5026] = 1'b1;
    assign layer3_out[5027] = ~layer2_out[2462];
    assign layer3_out[5028] = ~(layer2_out[1773] ^ layer2_out[1774]);
    assign layer3_out[5029] = layer2_out[3123] & ~layer2_out[3124];
    assign layer3_out[5030] = layer2_out[1709] & ~layer2_out[1708];
    assign layer3_out[5031] = layer2_out[4161] & layer2_out[4162];
    assign layer3_out[5032] = layer2_out[6848] ^ layer2_out[6849];
    assign layer3_out[5033] = ~layer2_out[7287];
    assign layer3_out[5034] = layer2_out[5167] & ~layer2_out[5166];
    assign layer3_out[5035] = ~layer2_out[5112] | layer2_out[5113];
    assign layer3_out[5036] = layer2_out[1750] & ~layer2_out[1749];
    assign layer3_out[5037] = layer2_out[1880] ^ layer2_out[1881];
    assign layer3_out[5038] = ~layer2_out[3191];
    assign layer3_out[5039] = 1'b1;
    assign layer3_out[5040] = layer2_out[3221];
    assign layer3_out[5041] = layer2_out[512] | layer2_out[513];
    assign layer3_out[5042] = layer2_out[4930] & ~layer2_out[4929];
    assign layer3_out[5043] = ~layer2_out[1286];
    assign layer3_out[5044] = ~(layer2_out[6671] ^ layer2_out[6672]);
    assign layer3_out[5045] = layer2_out[6701];
    assign layer3_out[5046] = ~(layer2_out[3458] & layer2_out[3459]);
    assign layer3_out[5047] = layer2_out[2976];
    assign layer3_out[5048] = layer2_out[2830] | layer2_out[2831];
    assign layer3_out[5049] = ~layer2_out[7873] | layer2_out[7874];
    assign layer3_out[5050] = layer2_out[2960];
    assign layer3_out[5051] = layer2_out[7932] | layer2_out[7933];
    assign layer3_out[5052] = ~(layer2_out[7302] ^ layer2_out[7303]);
    assign layer3_out[5053] = ~layer2_out[1532];
    assign layer3_out[5054] = ~layer2_out[6901];
    assign layer3_out[5055] = ~layer2_out[2834] | layer2_out[2833];
    assign layer3_out[5056] = layer2_out[1771] | layer2_out[1772];
    assign layer3_out[5057] = ~layer2_out[1119];
    assign layer3_out[5058] = layer2_out[293];
    assign layer3_out[5059] = layer2_out[515];
    assign layer3_out[5060] = layer2_out[6065] ^ layer2_out[6066];
    assign layer3_out[5061] = layer2_out[872] & layer2_out[873];
    assign layer3_out[5062] = 1'b1;
    assign layer3_out[5063] = layer2_out[7352] ^ layer2_out[7353];
    assign layer3_out[5064] = layer2_out[6738];
    assign layer3_out[5065] = ~(layer2_out[4270] & layer2_out[4271]);
    assign layer3_out[5066] = ~layer2_out[7342] | layer2_out[7341];
    assign layer3_out[5067] = ~(layer2_out[2541] ^ layer2_out[2542]);
    assign layer3_out[5068] = layer2_out[3746] | layer2_out[3747];
    assign layer3_out[5069] = layer2_out[2232];
    assign layer3_out[5070] = ~layer2_out[4026];
    assign layer3_out[5071] = ~layer2_out[988];
    assign layer3_out[5072] = ~layer2_out[3028];
    assign layer3_out[5073] = layer2_out[2421];
    assign layer3_out[5074] = ~(layer2_out[2177] & layer2_out[2178]);
    assign layer3_out[5075] = ~(layer2_out[1519] & layer2_out[1520]);
    assign layer3_out[5076] = ~layer2_out[1436] | layer2_out[1437];
    assign layer3_out[5077] = ~layer2_out[4888];
    assign layer3_out[5078] = ~layer2_out[871] | layer2_out[872];
    assign layer3_out[5079] = ~layer2_out[4140];
    assign layer3_out[5080] = layer2_out[6433];
    assign layer3_out[5081] = 1'b1;
    assign layer3_out[5082] = layer2_out[2565] & layer2_out[2566];
    assign layer3_out[5083] = ~layer2_out[7565];
    assign layer3_out[5084] = layer2_out[5800] & ~layer2_out[5801];
    assign layer3_out[5085] = layer2_out[6517];
    assign layer3_out[5086] = ~layer2_out[3918];
    assign layer3_out[5087] = ~layer2_out[7414];
    assign layer3_out[5088] = layer2_out[4501] & ~layer2_out[4500];
    assign layer3_out[5089] = ~layer2_out[367] | layer2_out[368];
    assign layer3_out[5090] = layer2_out[5353];
    assign layer3_out[5091] = layer2_out[3970];
    assign layer3_out[5092] = layer2_out[3112];
    assign layer3_out[5093] = layer2_out[1524];
    assign layer3_out[5094] = ~(layer2_out[301] & layer2_out[302]);
    assign layer3_out[5095] = layer2_out[5469] & ~layer2_out[5468];
    assign layer3_out[5096] = layer2_out[7300] & ~layer2_out[7301];
    assign layer3_out[5097] = layer2_out[528] ^ layer2_out[529];
    assign layer3_out[5098] = layer2_out[1490];
    assign layer3_out[5099] = layer2_out[682] & ~layer2_out[681];
    assign layer3_out[5100] = layer2_out[733] & layer2_out[734];
    assign layer3_out[5101] = ~layer2_out[2001];
    assign layer3_out[5102] = ~layer2_out[2794] | layer2_out[2793];
    assign layer3_out[5103] = ~layer2_out[5891] | layer2_out[5890];
    assign layer3_out[5104] = ~layer2_out[1062] | layer2_out[1063];
    assign layer3_out[5105] = ~(layer2_out[541] ^ layer2_out[542]);
    assign layer3_out[5106] = layer2_out[1251];
    assign layer3_out[5107] = ~(layer2_out[7044] ^ layer2_out[7045]);
    assign layer3_out[5108] = ~(layer2_out[828] ^ layer2_out[829]);
    assign layer3_out[5109] = ~layer2_out[5817];
    assign layer3_out[5110] = layer2_out[7933] & ~layer2_out[7934];
    assign layer3_out[5111] = layer2_out[7394];
    assign layer3_out[5112] = layer2_out[3807] & ~layer2_out[3806];
    assign layer3_out[5113] = ~(layer2_out[5831] ^ layer2_out[5832]);
    assign layer3_out[5114] = layer2_out[4055];
    assign layer3_out[5115] = layer2_out[3148];
    assign layer3_out[5116] = ~layer2_out[4760];
    assign layer3_out[5117] = layer2_out[4397] & ~layer2_out[4398];
    assign layer3_out[5118] = layer2_out[2961];
    assign layer3_out[5119] = layer2_out[4179];
    assign layer3_out[5120] = ~(layer2_out[2808] & layer2_out[2809]);
    assign layer3_out[5121] = layer2_out[3778] | layer2_out[3779];
    assign layer3_out[5122] = ~layer2_out[1607] | layer2_out[1606];
    assign layer3_out[5123] = layer2_out[3035] | layer2_out[3036];
    assign layer3_out[5124] = layer2_out[4395] & ~layer2_out[4396];
    assign layer3_out[5125] = layer2_out[1981];
    assign layer3_out[5126] = ~(layer2_out[6324] ^ layer2_out[6325]);
    assign layer3_out[5127] = layer2_out[121] & layer2_out[122];
    assign layer3_out[5128] = ~layer2_out[3276] | layer2_out[3275];
    assign layer3_out[5129] = ~(layer2_out[6870] ^ layer2_out[6871]);
    assign layer3_out[5130] = ~(layer2_out[1515] | layer2_out[1516]);
    assign layer3_out[5131] = layer2_out[6650];
    assign layer3_out[5132] = ~layer2_out[2706];
    assign layer3_out[5133] = ~layer2_out[3205] | layer2_out[3204];
    assign layer3_out[5134] = ~layer2_out[3504];
    assign layer3_out[5135] = layer2_out[1788];
    assign layer3_out[5136] = layer2_out[7534] & ~layer2_out[7533];
    assign layer3_out[5137] = ~layer2_out[1822] | layer2_out[1823];
    assign layer3_out[5138] = layer2_out[7095];
    assign layer3_out[5139] = ~layer2_out[1581] | layer2_out[1582];
    assign layer3_out[5140] = ~layer2_out[5708];
    assign layer3_out[5141] = layer2_out[1144];
    assign layer3_out[5142] = layer2_out[6771] & layer2_out[6772];
    assign layer3_out[5143] = ~layer2_out[3593] | layer2_out[3592];
    assign layer3_out[5144] = ~(layer2_out[2676] | layer2_out[2677]);
    assign layer3_out[5145] = layer2_out[412] | layer2_out[413];
    assign layer3_out[5146] = layer2_out[6401];
    assign layer3_out[5147] = layer2_out[1605];
    assign layer3_out[5148] = ~layer2_out[3378];
    assign layer3_out[5149] = ~(layer2_out[178] & layer2_out[179]);
    assign layer3_out[5150] = layer2_out[1260] & layer2_out[1261];
    assign layer3_out[5151] = ~(layer2_out[5836] ^ layer2_out[5837]);
    assign layer3_out[5152] = layer2_out[6964] | layer2_out[6965];
    assign layer3_out[5153] = ~layer2_out[5191];
    assign layer3_out[5154] = layer2_out[3589] & ~layer2_out[3588];
    assign layer3_out[5155] = layer2_out[5772] ^ layer2_out[5773];
    assign layer3_out[5156] = ~(layer2_out[6256] ^ layer2_out[6257]);
    assign layer3_out[5157] = layer2_out[2168];
    assign layer3_out[5158] = ~(layer2_out[661] | layer2_out[662]);
    assign layer3_out[5159] = layer2_out[780];
    assign layer3_out[5160] = ~(layer2_out[7706] | layer2_out[7707]);
    assign layer3_out[5161] = layer2_out[136];
    assign layer3_out[5162] = layer2_out[6267] & ~layer2_out[6268];
    assign layer3_out[5163] = layer2_out[585];
    assign layer3_out[5164] = ~(layer2_out[1032] ^ layer2_out[1033]);
    assign layer3_out[5165] = layer2_out[7638];
    assign layer3_out[5166] = ~layer2_out[6287] | layer2_out[6286];
    assign layer3_out[5167] = ~(layer2_out[5788] ^ layer2_out[5789]);
    assign layer3_out[5168] = 1'b0;
    assign layer3_out[5169] = layer2_out[3257];
    assign layer3_out[5170] = layer2_out[7752] ^ layer2_out[7753];
    assign layer3_out[5171] = ~layer2_out[2327];
    assign layer3_out[5172] = layer2_out[7073] | layer2_out[7074];
    assign layer3_out[5173] = layer2_out[383] ^ layer2_out[384];
    assign layer3_out[5174] = ~layer2_out[3648];
    assign layer3_out[5175] = ~layer2_out[761] | layer2_out[762];
    assign layer3_out[5176] = ~(layer2_out[5004] | layer2_out[5005]);
    assign layer3_out[5177] = ~layer2_out[3050];
    assign layer3_out[5178] = layer2_out[6100];
    assign layer3_out[5179] = layer2_out[1397];
    assign layer3_out[5180] = 1'b0;
    assign layer3_out[5181] = ~(layer2_out[150] ^ layer2_out[151]);
    assign layer3_out[5182] = ~(layer2_out[1829] ^ layer2_out[1830]);
    assign layer3_out[5183] = layer2_out[7978] | layer2_out[7979];
    assign layer3_out[5184] = ~layer2_out[6229];
    assign layer3_out[5185] = ~(layer2_out[3044] ^ layer2_out[3045]);
    assign layer3_out[5186] = ~layer2_out[6046] | layer2_out[6047];
    assign layer3_out[5187] = ~(layer2_out[7881] | layer2_out[7882]);
    assign layer3_out[5188] = ~layer2_out[1921] | layer2_out[1922];
    assign layer3_out[5189] = ~(layer2_out[6429] & layer2_out[6430]);
    assign layer3_out[5190] = ~layer2_out[4380] | layer2_out[4381];
    assign layer3_out[5191] = ~layer2_out[4253];
    assign layer3_out[5192] = ~(layer2_out[468] ^ layer2_out[469]);
    assign layer3_out[5193] = 1'b1;
    assign layer3_out[5194] = ~layer2_out[3056] | layer2_out[3055];
    assign layer3_out[5195] = ~layer2_out[6173];
    assign layer3_out[5196] = 1'b0;
    assign layer3_out[5197] = layer2_out[1164];
    assign layer3_out[5198] = ~layer2_out[1502];
    assign layer3_out[5199] = layer2_out[5696] & ~layer2_out[5695];
    assign layer3_out[5200] = ~layer2_out[1602] | layer2_out[1601];
    assign layer3_out[5201] = layer2_out[7916];
    assign layer3_out[5202] = layer2_out[7297];
    assign layer3_out[5203] = layer2_out[5308] & layer2_out[5309];
    assign layer3_out[5204] = layer2_out[4596] & layer2_out[4597];
    assign layer3_out[5205] = layer2_out[1388];
    assign layer3_out[5206] = layer2_out[1454];
    assign layer3_out[5207] = layer2_out[2669];
    assign layer3_out[5208] = layer2_out[6740];
    assign layer3_out[5209] = layer2_out[2818] & layer2_out[2819];
    assign layer3_out[5210] = layer2_out[954] ^ layer2_out[955];
    assign layer3_out[5211] = ~layer2_out[6994];
    assign layer3_out[5212] = layer2_out[7423];
    assign layer3_out[5213] = ~layer2_out[1416];
    assign layer3_out[5214] = ~layer2_out[2090] | layer2_out[2089];
    assign layer3_out[5215] = layer2_out[7349] & ~layer2_out[7348];
    assign layer3_out[5216] = ~(layer2_out[6967] & layer2_out[6968]);
    assign layer3_out[5217] = ~layer2_out[5103];
    assign layer3_out[5218] = layer2_out[5858];
    assign layer3_out[5219] = layer2_out[3304] ^ layer2_out[3305];
    assign layer3_out[5220] = layer2_out[4417];
    assign layer3_out[5221] = ~layer2_out[7742];
    assign layer3_out[5222] = layer2_out[335];
    assign layer3_out[5223] = layer2_out[4163] & ~layer2_out[4162];
    assign layer3_out[5224] = layer2_out[1713];
    assign layer3_out[5225] = ~(layer2_out[1682] ^ layer2_out[1683]);
    assign layer3_out[5226] = ~layer2_out[3846] | layer2_out[3845];
    assign layer3_out[5227] = ~layer2_out[4085];
    assign layer3_out[5228] = ~(layer2_out[31] & layer2_out[32]);
    assign layer3_out[5229] = layer2_out[7387] & layer2_out[7388];
    assign layer3_out[5230] = layer2_out[4484] & layer2_out[4485];
    assign layer3_out[5231] = ~layer2_out[5752];
    assign layer3_out[5232] = ~layer2_out[3418];
    assign layer3_out[5233] = 1'b1;
    assign layer3_out[5234] = layer2_out[1437];
    assign layer3_out[5235] = ~(layer2_out[6444] & layer2_out[6445]);
    assign layer3_out[5236] = layer2_out[4505] & ~layer2_out[4504];
    assign layer3_out[5237] = layer2_out[260] ^ layer2_out[261];
    assign layer3_out[5238] = layer2_out[348] | layer2_out[349];
    assign layer3_out[5239] = ~layer2_out[280];
    assign layer3_out[5240] = 1'b1;
    assign layer3_out[5241] = layer2_out[7240] & layer2_out[7241];
    assign layer3_out[5242] = layer2_out[1441];
    assign layer3_out[5243] = layer2_out[2106] & ~layer2_out[2107];
    assign layer3_out[5244] = layer2_out[6048];
    assign layer3_out[5245] = layer2_out[1851] ^ layer2_out[1852];
    assign layer3_out[5246] = ~layer2_out[4129] | layer2_out[4130];
    assign layer3_out[5247] = ~layer2_out[4849];
    assign layer3_out[5248] = layer2_out[5828];
    assign layer3_out[5249] = layer2_out[1709] & layer2_out[1710];
    assign layer3_out[5250] = ~layer2_out[5759];
    assign layer3_out[5251] = ~layer2_out[2032] | layer2_out[2031];
    assign layer3_out[5252] = layer2_out[6070] & ~layer2_out[6071];
    assign layer3_out[5253] = ~layer2_out[4590];
    assign layer3_out[5254] = ~(layer2_out[1764] ^ layer2_out[1765]);
    assign layer3_out[5255] = layer2_out[7076] & ~layer2_out[7075];
    assign layer3_out[5256] = 1'b1;
    assign layer3_out[5257] = layer2_out[4705];
    assign layer3_out[5258] = ~layer2_out[2529];
    assign layer3_out[5259] = layer2_out[4562];
    assign layer3_out[5260] = ~(layer2_out[6005] | layer2_out[6006]);
    assign layer3_out[5261] = ~(layer2_out[3847] | layer2_out[3848]);
    assign layer3_out[5262] = ~layer2_out[2235] | layer2_out[2234];
    assign layer3_out[5263] = layer2_out[1908] & ~layer2_out[1909];
    assign layer3_out[5264] = ~layer2_out[3198] | layer2_out[3199];
    assign layer3_out[5265] = layer2_out[4533] & ~layer2_out[4534];
    assign layer3_out[5266] = layer2_out[3230] & ~layer2_out[3231];
    assign layer3_out[5267] = layer2_out[1015] & layer2_out[1016];
    assign layer3_out[5268] = layer2_out[765] & ~layer2_out[766];
    assign layer3_out[5269] = ~layer2_out[3663];
    assign layer3_out[5270] = layer2_out[2583];
    assign layer3_out[5271] = ~layer2_out[6235];
    assign layer3_out[5272] = ~layer2_out[1998] | layer2_out[1999];
    assign layer3_out[5273] = layer2_out[262] & layer2_out[263];
    assign layer3_out[5274] = 1'b1;
    assign layer3_out[5275] = layer2_out[7164] & layer2_out[7165];
    assign layer3_out[5276] = layer2_out[746] & ~layer2_out[747];
    assign layer3_out[5277] = ~layer2_out[1334];
    assign layer3_out[5278] = layer2_out[4913];
    assign layer3_out[5279] = layer2_out[2907] ^ layer2_out[2908];
    assign layer3_out[5280] = 1'b1;
    assign layer3_out[5281] = layer2_out[1646] & layer2_out[1647];
    assign layer3_out[5282] = ~(layer2_out[852] & layer2_out[853]);
    assign layer3_out[5283] = ~layer2_out[3247];
    assign layer3_out[5284] = layer2_out[6915] ^ layer2_out[6916];
    assign layer3_out[5285] = ~layer2_out[763] | layer2_out[764];
    assign layer3_out[5286] = layer2_out[1248];
    assign layer3_out[5287] = ~layer2_out[7746];
    assign layer3_out[5288] = ~layer2_out[2196] | layer2_out[2195];
    assign layer3_out[5289] = layer2_out[6289];
    assign layer3_out[5290] = layer2_out[3754];
    assign layer3_out[5291] = layer2_out[7148] ^ layer2_out[7149];
    assign layer3_out[5292] = layer2_out[2938] ^ layer2_out[2939];
    assign layer3_out[5293] = ~layer2_out[237] | layer2_out[238];
    assign layer3_out[5294] = ~layer2_out[5570];
    assign layer3_out[5295] = ~(layer2_out[1840] & layer2_out[1841]);
    assign layer3_out[5296] = ~layer2_out[3372];
    assign layer3_out[5297] = layer2_out[1750];
    assign layer3_out[5298] = layer2_out[3567] & ~layer2_out[3568];
    assign layer3_out[5299] = layer2_out[5902] & layer2_out[5903];
    assign layer3_out[5300] = layer2_out[2485];
    assign layer3_out[5301] = layer2_out[1365];
    assign layer3_out[5302] = ~layer2_out[4204];
    assign layer3_out[5303] = layer2_out[1586];
    assign layer3_out[5304] = layer2_out[852] & ~layer2_out[851];
    assign layer3_out[5305] = layer2_out[3862] & layer2_out[3863];
    assign layer3_out[5306] = ~(layer2_out[7946] & layer2_out[7947]);
    assign layer3_out[5307] = ~layer2_out[7700];
    assign layer3_out[5308] = ~(layer2_out[4288] & layer2_out[4289]);
    assign layer3_out[5309] = ~(layer2_out[3603] | layer2_out[3604]);
    assign layer3_out[5310] = ~layer2_out[157];
    assign layer3_out[5311] = layer2_out[2233];
    assign layer3_out[5312] = layer2_out[278] & layer2_out[279];
    assign layer3_out[5313] = layer2_out[1054] & ~layer2_out[1055];
    assign layer3_out[5314] = layer2_out[7380] & ~layer2_out[7381];
    assign layer3_out[5315] = ~layer2_out[468];
    assign layer3_out[5316] = ~layer2_out[1563];
    assign layer3_out[5317] = ~layer2_out[1398] | layer2_out[1397];
    assign layer3_out[5318] = layer2_out[2570];
    assign layer3_out[5319] = ~layer2_out[13];
    assign layer3_out[5320] = ~layer2_out[5124];
    assign layer3_out[5321] = ~layer2_out[2735];
    assign layer3_out[5322] = ~layer2_out[4019] | layer2_out[4020];
    assign layer3_out[5323] = layer2_out[4482] & layer2_out[4483];
    assign layer3_out[5324] = ~layer2_out[887];
    assign layer3_out[5325] = 1'b0;
    assign layer3_out[5326] = layer2_out[1315];
    assign layer3_out[5327] = ~(layer2_out[1164] ^ layer2_out[1165]);
    assign layer3_out[5328] = layer2_out[1109] | layer2_out[1110];
    assign layer3_out[5329] = ~(layer2_out[6212] | layer2_out[6213]);
    assign layer3_out[5330] = layer2_out[945];
    assign layer3_out[5331] = layer2_out[2004];
    assign layer3_out[5332] = ~layer2_out[3678] | layer2_out[3677];
    assign layer3_out[5333] = layer2_out[1499] ^ layer2_out[1500];
    assign layer3_out[5334] = ~(layer2_out[479] | layer2_out[480]);
    assign layer3_out[5335] = layer2_out[2057];
    assign layer3_out[5336] = 1'b1;
    assign layer3_out[5337] = ~(layer2_out[4786] | layer2_out[4787]);
    assign layer3_out[5338] = ~(layer2_out[966] & layer2_out[967]);
    assign layer3_out[5339] = layer2_out[7031] & layer2_out[7032];
    assign layer3_out[5340] = layer2_out[5065];
    assign layer3_out[5341] = layer2_out[3283] ^ layer2_out[3284];
    assign layer3_out[5342] = ~layer2_out[3559];
    assign layer3_out[5343] = ~layer2_out[5754] | layer2_out[5753];
    assign layer3_out[5344] = layer2_out[155] & layer2_out[156];
    assign layer3_out[5345] = ~(layer2_out[7836] ^ layer2_out[7837]);
    assign layer3_out[5346] = layer2_out[1713] & ~layer2_out[1712];
    assign layer3_out[5347] = layer2_out[6365] | layer2_out[6366];
    assign layer3_out[5348] = ~(layer2_out[6563] | layer2_out[6564]);
    assign layer3_out[5349] = 1'b1;
    assign layer3_out[5350] = layer2_out[6119];
    assign layer3_out[5351] = ~layer2_out[2865];
    assign layer3_out[5352] = ~layer2_out[4684];
    assign layer3_out[5353] = ~layer2_out[4810];
    assign layer3_out[5354] = ~layer2_out[3780];
    assign layer3_out[5355] = layer2_out[2308];
    assign layer3_out[5356] = layer2_out[5544];
    assign layer3_out[5357] = ~layer2_out[3475] | layer2_out[3474];
    assign layer3_out[5358] = layer2_out[5113];
    assign layer3_out[5359] = ~layer2_out[1836] | layer2_out[1835];
    assign layer3_out[5360] = layer2_out[380];
    assign layer3_out[5361] = ~(layer2_out[3083] | layer2_out[3084]);
    assign layer3_out[5362] = layer2_out[6461] & layer2_out[6462];
    assign layer3_out[5363] = layer2_out[6062] | layer2_out[6063];
    assign layer3_out[5364] = layer2_out[59] & ~layer2_out[60];
    assign layer3_out[5365] = ~layer2_out[2140];
    assign layer3_out[5366] = layer2_out[5259];
    assign layer3_out[5367] = layer2_out[4124];
    assign layer3_out[5368] = layer2_out[7683];
    assign layer3_out[5369] = layer2_out[4517] & layer2_out[4518];
    assign layer3_out[5370] = ~(layer2_out[7835] & layer2_out[7836]);
    assign layer3_out[5371] = ~layer2_out[3176];
    assign layer3_out[5372] = layer2_out[7719];
    assign layer3_out[5373] = ~layer2_out[5315] | layer2_out[5316];
    assign layer3_out[5374] = layer2_out[7155];
    assign layer3_out[5375] = layer2_out[5578] & ~layer2_out[5577];
    assign layer3_out[5376] = layer2_out[6118];
    assign layer3_out[5377] = layer2_out[6725];
    assign layer3_out[5378] = layer2_out[6146];
    assign layer3_out[5379] = layer2_out[2176];
    assign layer3_out[5380] = ~layer2_out[2008];
    assign layer3_out[5381] = ~(layer2_out[6506] & layer2_out[6507]);
    assign layer3_out[5382] = ~(layer2_out[239] | layer2_out[240]);
    assign layer3_out[5383] = ~layer2_out[7580] | layer2_out[7581];
    assign layer3_out[5384] = layer2_out[7957] | layer2_out[7958];
    assign layer3_out[5385] = ~(layer2_out[7064] | layer2_out[7065]);
    assign layer3_out[5386] = layer2_out[5579];
    assign layer3_out[5387] = ~layer2_out[2378] | layer2_out[2379];
    assign layer3_out[5388] = layer2_out[2373];
    assign layer3_out[5389] = layer2_out[7667];
    assign layer3_out[5390] = ~(layer2_out[2674] & layer2_out[2675]);
    assign layer3_out[5391] = ~(layer2_out[2138] ^ layer2_out[2139]);
    assign layer3_out[5392] = ~layer2_out[6002] | layer2_out[6003];
    assign layer3_out[5393] = ~(layer2_out[7994] | layer2_out[7995]);
    assign layer3_out[5394] = layer2_out[5055] & ~layer2_out[5056];
    assign layer3_out[5395] = ~layer2_out[6159] | layer2_out[6160];
    assign layer3_out[5396] = ~layer2_out[7613] | layer2_out[7614];
    assign layer3_out[5397] = ~layer2_out[6521] | layer2_out[6520];
    assign layer3_out[5398] = ~layer2_out[5485];
    assign layer3_out[5399] = layer2_out[4069] & ~layer2_out[4070];
    assign layer3_out[5400] = ~layer2_out[1356];
    assign layer3_out[5401] = ~(layer2_out[3440] & layer2_out[3441]);
    assign layer3_out[5402] = ~layer2_out[4832] | layer2_out[4833];
    assign layer3_out[5403] = layer2_out[6499];
    assign layer3_out[5404] = layer2_out[3801] ^ layer2_out[3802];
    assign layer3_out[5405] = layer2_out[4015] ^ layer2_out[4016];
    assign layer3_out[5406] = ~layer2_out[6900];
    assign layer3_out[5407] = layer2_out[5162];
    assign layer3_out[5408] = ~layer2_out[2655] | layer2_out[2654];
    assign layer3_out[5409] = ~layer2_out[2026];
    assign layer3_out[5410] = ~layer2_out[7126];
    assign layer3_out[5411] = ~layer2_out[4402];
    assign layer3_out[5412] = layer2_out[6944] | layer2_out[6945];
    assign layer3_out[5413] = ~layer2_out[6294] | layer2_out[6295];
    assign layer3_out[5414] = layer2_out[328];
    assign layer3_out[5415] = layer2_out[1240] & ~layer2_out[1241];
    assign layer3_out[5416] = ~layer2_out[2804];
    assign layer3_out[5417] = ~layer2_out[5633] | layer2_out[5632];
    assign layer3_out[5418] = ~layer2_out[1438] | layer2_out[1439];
    assign layer3_out[5419] = ~layer2_out[7575] | layer2_out[7574];
    assign layer3_out[5420] = ~(layer2_out[1049] & layer2_out[1050]);
    assign layer3_out[5421] = ~(layer2_out[3823] ^ layer2_out[3824]);
    assign layer3_out[5422] = ~(layer2_out[6255] | layer2_out[6256]);
    assign layer3_out[5423] = layer2_out[5604] | layer2_out[5605];
    assign layer3_out[5424] = layer2_out[2404];
    assign layer3_out[5425] = ~(layer2_out[7359] | layer2_out[7360]);
    assign layer3_out[5426] = ~(layer2_out[1398] ^ layer2_out[1399]);
    assign layer3_out[5427] = layer2_out[5538];
    assign layer3_out[5428] = layer2_out[5788];
    assign layer3_out[5429] = layer2_out[4912];
    assign layer3_out[5430] = layer2_out[3881] & ~layer2_out[3880];
    assign layer3_out[5431] = layer2_out[488];
    assign layer3_out[5432] = ~layer2_out[2267] | layer2_out[2268];
    assign layer3_out[5433] = ~layer2_out[7466];
    assign layer3_out[5434] = layer2_out[6491] | layer2_out[6492];
    assign layer3_out[5435] = ~layer2_out[5563] | layer2_out[5564];
    assign layer3_out[5436] = ~layer2_out[6966];
    assign layer3_out[5437] = layer2_out[5078] ^ layer2_out[5079];
    assign layer3_out[5438] = layer2_out[5085];
    assign layer3_out[5439] = ~(layer2_out[3389] ^ layer2_out[3390]);
    assign layer3_out[5440] = ~layer2_out[4135] | layer2_out[4134];
    assign layer3_out[5441] = layer2_out[5808];
    assign layer3_out[5442] = layer2_out[5779] & layer2_out[5780];
    assign layer3_out[5443] = ~layer2_out[38];
    assign layer3_out[5444] = ~layer2_out[7939];
    assign layer3_out[5445] = ~(layer2_out[6553] & layer2_out[6554]);
    assign layer3_out[5446] = layer2_out[4132];
    assign layer3_out[5447] = ~layer2_out[6776] | layer2_out[6775];
    assign layer3_out[5448] = ~layer2_out[73] | layer2_out[74];
    assign layer3_out[5449] = ~(layer2_out[6208] ^ layer2_out[6209]);
    assign layer3_out[5450] = layer2_out[7382] & layer2_out[7383];
    assign layer3_out[5451] = layer2_out[4435];
    assign layer3_out[5452] = layer2_out[882];
    assign layer3_out[5453] = ~(layer2_out[2815] & layer2_out[2816]);
    assign layer3_out[5454] = layer2_out[452] & ~layer2_out[451];
    assign layer3_out[5455] = layer2_out[3019] ^ layer2_out[3020];
    assign layer3_out[5456] = ~layer2_out[3607];
    assign layer3_out[5457] = ~(layer2_out[7911] | layer2_out[7912]);
    assign layer3_out[5458] = layer2_out[6085] & layer2_out[6086];
    assign layer3_out[5459] = ~layer2_out[3584];
    assign layer3_out[5460] = ~layer2_out[4091] | layer2_out[4090];
    assign layer3_out[5461] = ~(layer2_out[7952] ^ layer2_out[7953]);
    assign layer3_out[5462] = ~(layer2_out[2310] & layer2_out[2311]);
    assign layer3_out[5463] = layer2_out[7603] | layer2_out[7604];
    assign layer3_out[5464] = layer2_out[5583];
    assign layer3_out[5465] = ~layer2_out[7743];
    assign layer3_out[5466] = layer2_out[1185];
    assign layer3_out[5467] = ~layer2_out[3155];
    assign layer3_out[5468] = ~layer2_out[3672] | layer2_out[3671];
    assign layer3_out[5469] = ~layer2_out[7900] | layer2_out[7901];
    assign layer3_out[5470] = layer2_out[6785] & ~layer2_out[6784];
    assign layer3_out[5471] = ~(layer2_out[6535] ^ layer2_out[6536]);
    assign layer3_out[5472] = ~(layer2_out[4651] | layer2_out[4652]);
    assign layer3_out[5473] = layer2_out[6578] | layer2_out[6579];
    assign layer3_out[5474] = ~(layer2_out[7823] | layer2_out[7824]);
    assign layer3_out[5475] = ~layer2_out[180];
    assign layer3_out[5476] = layer2_out[3834] & ~layer2_out[3835];
    assign layer3_out[5477] = ~layer2_out[7694] | layer2_out[7693];
    assign layer3_out[5478] = layer2_out[4529] ^ layer2_out[4530];
    assign layer3_out[5479] = ~(layer2_out[4733] | layer2_out[4734]);
    assign layer3_out[5480] = ~(layer2_out[7391] | layer2_out[7392]);
    assign layer3_out[5481] = ~(layer2_out[4597] & layer2_out[4598]);
    assign layer3_out[5482] = layer2_out[4265] | layer2_out[4266];
    assign layer3_out[5483] = layer2_out[1903];
    assign layer3_out[5484] = ~(layer2_out[1096] | layer2_out[1097]);
    assign layer3_out[5485] = ~layer2_out[2750];
    assign layer3_out[5486] = ~layer2_out[6965];
    assign layer3_out[5487] = layer2_out[7865] ^ layer2_out[7866];
    assign layer3_out[5488] = layer2_out[3766] & layer2_out[3767];
    assign layer3_out[5489] = layer2_out[5752];
    assign layer3_out[5490] = ~layer2_out[4263] | layer2_out[4262];
    assign layer3_out[5491] = ~layer2_out[462];
    assign layer3_out[5492] = ~layer2_out[832];
    assign layer3_out[5493] = ~(layer2_out[2396] | layer2_out[2397]);
    assign layer3_out[5494] = layer2_out[6940] & layer2_out[6941];
    assign layer3_out[5495] = layer2_out[7675] & layer2_out[7676];
    assign layer3_out[5496] = ~layer2_out[3510] | layer2_out[3511];
    assign layer3_out[5497] = ~layer2_out[946];
    assign layer3_out[5498] = ~layer2_out[5284];
    assign layer3_out[5499] = layer2_out[987] | layer2_out[988];
    assign layer3_out[5500] = ~layer2_out[3917];
    assign layer3_out[5501] = ~layer2_out[4045] | layer2_out[4046];
    assign layer3_out[5502] = layer2_out[7069] ^ layer2_out[7070];
    assign layer3_out[5503] = ~layer2_out[1156];
    assign layer3_out[5504] = layer2_out[5152];
    assign layer3_out[5505] = layer2_out[3103];
    assign layer3_out[5506] = ~(layer2_out[339] ^ layer2_out[340]);
    assign layer3_out[5507] = layer2_out[6821] & ~layer2_out[6820];
    assign layer3_out[5508] = ~layer2_out[3738] | layer2_out[3737];
    assign layer3_out[5509] = ~(layer2_out[3086] & layer2_out[3087]);
    assign layer3_out[5510] = ~layer2_out[4295];
    assign layer3_out[5511] = layer2_out[2980];
    assign layer3_out[5512] = layer2_out[7309] ^ layer2_out[7310];
    assign layer3_out[5513] = ~(layer2_out[986] & layer2_out[987]);
    assign layer3_out[5514] = layer2_out[6228];
    assign layer3_out[5515] = layer2_out[147];
    assign layer3_out[5516] = layer2_out[6317] & layer2_out[6318];
    assign layer3_out[5517] = ~layer2_out[7385];
    assign layer3_out[5518] = 1'b1;
    assign layer3_out[5519] = layer2_out[4054] | layer2_out[4055];
    assign layer3_out[5520] = ~layer2_out[1548];
    assign layer3_out[5521] = layer2_out[8];
    assign layer3_out[5522] = ~layer2_out[2048];
    assign layer3_out[5523] = ~layer2_out[4038] | layer2_out[4039];
    assign layer3_out[5524] = layer2_out[3558] ^ layer2_out[3559];
    assign layer3_out[5525] = layer2_out[6272];
    assign layer3_out[5526] = layer2_out[3716] & ~layer2_out[3717];
    assign layer3_out[5527] = ~(layer2_out[477] ^ layer2_out[478]);
    assign layer3_out[5528] = ~layer2_out[7851] | layer2_out[7852];
    assign layer3_out[5529] = ~layer2_out[770];
    assign layer3_out[5530] = ~layer2_out[7922];
    assign layer3_out[5531] = ~layer2_out[557] | layer2_out[556];
    assign layer3_out[5532] = ~layer2_out[3947];
    assign layer3_out[5533] = layer2_out[2536] ^ layer2_out[2537];
    assign layer3_out[5534] = 1'b0;
    assign layer3_out[5535] = ~(layer2_out[3964] ^ layer2_out[3965]);
    assign layer3_out[5536] = layer2_out[5237] & ~layer2_out[5238];
    assign layer3_out[5537] = ~layer2_out[1238];
    assign layer3_out[5538] = layer2_out[2777] | layer2_out[2778];
    assign layer3_out[5539] = layer2_out[7791] | layer2_out[7792];
    assign layer3_out[5540] = layer2_out[5305];
    assign layer3_out[5541] = ~layer2_out[859];
    assign layer3_out[5542] = ~layer2_out[7578];
    assign layer3_out[5543] = ~layer2_out[3388];
    assign layer3_out[5544] = layer2_out[7323] ^ layer2_out[7324];
    assign layer3_out[5545] = ~layer2_out[4149] | layer2_out[4150];
    assign layer3_out[5546] = ~(layer2_out[4758] ^ layer2_out[4759]);
    assign layer3_out[5547] = ~layer2_out[4997] | layer2_out[4996];
    assign layer3_out[5548] = ~layer2_out[4738] | layer2_out[4739];
    assign layer3_out[5549] = ~layer2_out[1246] | layer2_out[1247];
    assign layer3_out[5550] = layer2_out[5761];
    assign layer3_out[5551] = ~(layer2_out[7783] & layer2_out[7784]);
    assign layer3_out[5552] = layer2_out[5675] ^ layer2_out[5676];
    assign layer3_out[5553] = ~(layer2_out[758] | layer2_out[759]);
    assign layer3_out[5554] = ~(layer2_out[2704] | layer2_out[2705]);
    assign layer3_out[5555] = ~layer2_out[3087];
    assign layer3_out[5556] = layer2_out[2088];
    assign layer3_out[5557] = ~(layer2_out[5010] | layer2_out[5011]);
    assign layer3_out[5558] = layer2_out[2521] & ~layer2_out[2522];
    assign layer3_out[5559] = layer2_out[5866];
    assign layer3_out[5560] = layer2_out[7729] & ~layer2_out[7730];
    assign layer3_out[5561] = layer2_out[5339];
    assign layer3_out[5562] = layer2_out[2567] & ~layer2_out[2568];
    assign layer3_out[5563] = ~(layer2_out[7684] & layer2_out[7685]);
    assign layer3_out[5564] = ~layer2_out[425];
    assign layer3_out[5565] = layer2_out[4167] | layer2_out[4168];
    assign layer3_out[5566] = ~layer2_out[1483] | layer2_out[1484];
    assign layer3_out[5567] = layer2_out[4977] & ~layer2_out[4976];
    assign layer3_out[5568] = layer2_out[2945] | layer2_out[2946];
    assign layer3_out[5569] = layer2_out[3578];
    assign layer3_out[5570] = layer2_out[3869] & ~layer2_out[3870];
    assign layer3_out[5571] = layer2_out[7223];
    assign layer3_out[5572] = ~layer2_out[7139] | layer2_out[7138];
    assign layer3_out[5573] = ~layer2_out[7644];
    assign layer3_out[5574] = layer2_out[7326] & ~layer2_out[7325];
    assign layer3_out[5575] = layer2_out[3651] & ~layer2_out[3652];
    assign layer3_out[5576] = ~layer2_out[5226] | layer2_out[5225];
    assign layer3_out[5577] = ~(layer2_out[5005] ^ layer2_out[5006]);
    assign layer3_out[5578] = layer2_out[6048] & ~layer2_out[6049];
    assign layer3_out[5579] = ~layer2_out[4361];
    assign layer3_out[5580] = layer2_out[5841];
    assign layer3_out[5581] = 1'b0;
    assign layer3_out[5582] = layer2_out[2252];
    assign layer3_out[5583] = layer2_out[5424];
    assign layer3_out[5584] = ~layer2_out[4807];
    assign layer3_out[5585] = layer2_out[6377] & ~layer2_out[6376];
    assign layer3_out[5586] = ~(layer2_out[1792] & layer2_out[1793]);
    assign layer3_out[5587] = ~layer2_out[4464];
    assign layer3_out[5588] = ~layer2_out[3880];
    assign layer3_out[5589] = ~layer2_out[823];
    assign layer3_out[5590] = ~layer2_out[61];
    assign layer3_out[5591] = ~layer2_out[1854] | layer2_out[1853];
    assign layer3_out[5592] = ~(layer2_out[1348] | layer2_out[1349]);
    assign layer3_out[5593] = ~layer2_out[7328];
    assign layer3_out[5594] = layer2_out[1246];
    assign layer3_out[5595] = layer2_out[573] & ~layer2_out[574];
    assign layer3_out[5596] = layer2_out[7150];
    assign layer3_out[5597] = ~layer2_out[4921];
    assign layer3_out[5598] = ~(layer2_out[858] & layer2_out[859]);
    assign layer3_out[5599] = ~layer2_out[7755];
    assign layer3_out[5600] = 1'b1;
    assign layer3_out[5601] = ~layer2_out[158] | layer2_out[159];
    assign layer3_out[5602] = ~(layer2_out[3156] & layer2_out[3157]);
    assign layer3_out[5603] = layer2_out[4042];
    assign layer3_out[5604] = ~(layer2_out[3393] ^ layer2_out[3394]);
    assign layer3_out[5605] = layer2_out[4002] | layer2_out[4003];
    assign layer3_out[5606] = layer2_out[2551] & ~layer2_out[2552];
    assign layer3_out[5607] = ~layer2_out[4837];
    assign layer3_out[5608] = ~layer2_out[4321] | layer2_out[4322];
    assign layer3_out[5609] = layer2_out[4883] & layer2_out[4884];
    assign layer3_out[5610] = layer2_out[4341] ^ layer2_out[4342];
    assign layer3_out[5611] = layer2_out[6917] ^ layer2_out[6918];
    assign layer3_out[5612] = ~layer2_out[7114] | layer2_out[7115];
    assign layer3_out[5613] = layer2_out[6951] & ~layer2_out[6952];
    assign layer3_out[5614] = ~layer2_out[5965];
    assign layer3_out[5615] = layer2_out[7291] & ~layer2_out[7290];
    assign layer3_out[5616] = layer2_out[2197] | layer2_out[2198];
    assign layer3_out[5617] = layer2_out[3600] & layer2_out[3601];
    assign layer3_out[5618] = 1'b0;
    assign layer3_out[5619] = ~(layer2_out[6842] | layer2_out[6843]);
    assign layer3_out[5620] = ~layer2_out[378];
    assign layer3_out[5621] = ~layer2_out[2950];
    assign layer3_out[5622] = layer2_out[1051];
    assign layer3_out[5623] = layer2_out[925];
    assign layer3_out[5624] = layer2_out[1048] | layer2_out[1049];
    assign layer3_out[5625] = ~layer2_out[2488];
    assign layer3_out[5626] = layer2_out[6979];
    assign layer3_out[5627] = ~layer2_out[5649];
    assign layer3_out[5628] = layer2_out[7698] | layer2_out[7699];
    assign layer3_out[5629] = ~layer2_out[422];
    assign layer3_out[5630] = ~(layer2_out[2718] & layer2_out[2719]);
    assign layer3_out[5631] = layer2_out[837];
    assign layer3_out[5632] = ~layer2_out[2260];
    assign layer3_out[5633] = layer2_out[3406] & ~layer2_out[3407];
    assign layer3_out[5634] = layer2_out[697];
    assign layer3_out[5635] = ~layer2_out[6079];
    assign layer3_out[5636] = ~layer2_out[2956];
    assign layer3_out[5637] = layer2_out[1374] ^ layer2_out[1375];
    assign layer3_out[5638] = layer2_out[3381] & ~layer2_out[3380];
    assign layer3_out[5639] = ~layer2_out[2927];
    assign layer3_out[5640] = layer2_out[6648];
    assign layer3_out[5641] = layer2_out[3685];
    assign layer3_out[5642] = layer2_out[7879] & ~layer2_out[7880];
    assign layer3_out[5643] = ~layer2_out[432];
    assign layer3_out[5644] = layer2_out[102] | layer2_out[103];
    assign layer3_out[5645] = ~layer2_out[4559];
    assign layer3_out[5646] = ~(layer2_out[2471] & layer2_out[2472]);
    assign layer3_out[5647] = layer2_out[1723] & ~layer2_out[1724];
    assign layer3_out[5648] = layer2_out[5692] & ~layer2_out[5693];
    assign layer3_out[5649] = layer2_out[3544] & ~layer2_out[3545];
    assign layer3_out[5650] = layer2_out[6448];
    assign layer3_out[5651] = ~layer2_out[2628];
    assign layer3_out[5652] = ~layer2_out[5072] | layer2_out[5071];
    assign layer3_out[5653] = ~layer2_out[6623];
    assign layer3_out[5654] = ~layer2_out[219];
    assign layer3_out[5655] = ~layer2_out[314];
    assign layer3_out[5656] = layer2_out[4292];
    assign layer3_out[5657] = ~(layer2_out[6896] | layer2_out[6897]);
    assign layer3_out[5658] = layer2_out[4994];
    assign layer3_out[5659] = ~(layer2_out[6914] & layer2_out[6915]);
    assign layer3_out[5660] = ~layer2_out[6281] | layer2_out[6280];
    assign layer3_out[5661] = layer2_out[5739] ^ layer2_out[5740];
    assign layer3_out[5662] = layer2_out[4874] & ~layer2_out[4873];
    assign layer3_out[5663] = ~layer2_out[116] | layer2_out[117];
    assign layer3_out[5664] = layer2_out[4715];
    assign layer3_out[5665] = ~layer2_out[444];
    assign layer3_out[5666] = layer2_out[7057];
    assign layer3_out[5667] = ~(layer2_out[3552] & layer2_out[3553]);
    assign layer3_out[5668] = ~layer2_out[5916];
    assign layer3_out[5669] = layer2_out[6464] & ~layer2_out[6463];
    assign layer3_out[5670] = layer2_out[4539] & layer2_out[4540];
    assign layer3_out[5671] = 1'b0;
    assign layer3_out[5672] = ~layer2_out[7602] | layer2_out[7601];
    assign layer3_out[5673] = ~layer2_out[5574];
    assign layer3_out[5674] = layer2_out[2540];
    assign layer3_out[5675] = ~(layer2_out[7316] | layer2_out[7317]);
    assign layer3_out[5676] = layer2_out[961];
    assign layer3_out[5677] = ~(layer2_out[1565] & layer2_out[1566]);
    assign layer3_out[5678] = layer2_out[4095] | layer2_out[4096];
    assign layer3_out[5679] = 1'b1;
    assign layer3_out[5680] = layer2_out[5021] & ~layer2_out[5022];
    assign layer3_out[5681] = ~(layer2_out[7153] & layer2_out[7154]);
    assign layer3_out[5682] = layer2_out[69] & ~layer2_out[70];
    assign layer3_out[5683] = ~(layer2_out[2428] | layer2_out[2429]);
    assign layer3_out[5684] = layer2_out[4413] | layer2_out[4414];
    assign layer3_out[5685] = ~layer2_out[7685];
    assign layer3_out[5686] = ~(layer2_out[688] & layer2_out[689]);
    assign layer3_out[5687] = layer2_out[6001] & layer2_out[6002];
    assign layer3_out[5688] = ~layer2_out[218];
    assign layer3_out[5689] = 1'b0;
    assign layer3_out[5690] = layer2_out[7575];
    assign layer3_out[5691] = ~layer2_out[7284] | layer2_out[7283];
    assign layer3_out[5692] = ~layer2_out[1194];
    assign layer3_out[5693] = ~layer2_out[4560];
    assign layer3_out[5694] = layer2_out[5153] & ~layer2_out[5154];
    assign layer3_out[5695] = layer2_out[7405] | layer2_out[7406];
    assign layer3_out[5696] = ~layer2_out[2497] | layer2_out[2496];
    assign layer3_out[5697] = layer2_out[7837];
    assign layer3_out[5698] = layer2_out[7924] & ~layer2_out[7925];
    assign layer3_out[5699] = ~layer2_out[1912];
    assign layer3_out[5700] = layer2_out[6339] & layer2_out[6340];
    assign layer3_out[5701] = layer2_out[3299] & ~layer2_out[3300];
    assign layer3_out[5702] = ~(layer2_out[6044] & layer2_out[6045]);
    assign layer3_out[5703] = layer2_out[5533] ^ layer2_out[5534];
    assign layer3_out[5704] = layer2_out[1754];
    assign layer3_out[5705] = layer2_out[6832] & ~layer2_out[6833];
    assign layer3_out[5706] = layer2_out[6026];
    assign layer3_out[5707] = 1'b0;
    assign layer3_out[5708] = layer2_out[6210] & ~layer2_out[6211];
    assign layer3_out[5709] = layer2_out[4259];
    assign layer3_out[5710] = layer2_out[1872];
    assign layer3_out[5711] = ~(layer2_out[7459] & layer2_out[7460]);
    assign layer3_out[5712] = ~(layer2_out[6108] ^ layer2_out[6109]);
    assign layer3_out[5713] = ~layer2_out[4341] | layer2_out[4340];
    assign layer3_out[5714] = layer2_out[6465] & layer2_out[6466];
    assign layer3_out[5715] = layer2_out[1967] ^ layer2_out[1968];
    assign layer3_out[5716] = ~(layer2_out[1253] ^ layer2_out[1254]);
    assign layer3_out[5717] = layer2_out[5943] & ~layer2_out[5944];
    assign layer3_out[5718] = layer2_out[2983] | layer2_out[2984];
    assign layer3_out[5719] = ~(layer2_out[5009] ^ layer2_out[5010]);
    assign layer3_out[5720] = ~(layer2_out[3938] & layer2_out[3939]);
    assign layer3_out[5721] = layer2_out[2392];
    assign layer3_out[5722] = layer2_out[2104] & ~layer2_out[2103];
    assign layer3_out[5723] = ~layer2_out[1197];
    assign layer3_out[5724] = ~(layer2_out[1672] & layer2_out[1673]);
    assign layer3_out[5725] = layer2_out[4968] | layer2_out[4969];
    assign layer3_out[5726] = ~(layer2_out[4802] & layer2_out[4803]);
    assign layer3_out[5727] = layer2_out[4535] | layer2_out[4536];
    assign layer3_out[5728] = layer2_out[2235] ^ layer2_out[2236];
    assign layer3_out[5729] = ~layer2_out[526];
    assign layer3_out[5730] = ~layer2_out[5850];
    assign layer3_out[5731] = layer2_out[4571] | layer2_out[4572];
    assign layer3_out[5732] = ~layer2_out[7573] | layer2_out[7572];
    assign layer3_out[5733] = layer2_out[5326] & layer2_out[5327];
    assign layer3_out[5734] = layer2_out[4428] & layer2_out[4429];
    assign layer3_out[5735] = ~(layer2_out[6213] | layer2_out[6214]);
    assign layer3_out[5736] = layer2_out[5504] & ~layer2_out[5503];
    assign layer3_out[5737] = ~layer2_out[4763];
    assign layer3_out[5738] = ~layer2_out[4160] | layer2_out[4159];
    assign layer3_out[5739] = ~(layer2_out[5966] & layer2_out[5967]);
    assign layer3_out[5740] = layer2_out[3652] | layer2_out[3653];
    assign layer3_out[5741] = ~(layer2_out[1994] | layer2_out[1995]);
    assign layer3_out[5742] = layer2_out[1658] ^ layer2_out[1659];
    assign layer3_out[5743] = ~layer2_out[4961] | layer2_out[4960];
    assign layer3_out[5744] = layer2_out[1869] & ~layer2_out[1868];
    assign layer3_out[5745] = ~layer2_out[4892];
    assign layer3_out[5746] = ~(layer2_out[2933] & layer2_out[2934]);
    assign layer3_out[5747] = ~layer2_out[5854] | layer2_out[5853];
    assign layer3_out[5748] = ~(layer2_out[6823] | layer2_out[6824]);
    assign layer3_out[5749] = ~(layer2_out[1130] | layer2_out[1131]);
    assign layer3_out[5750] = ~(layer2_out[3699] | layer2_out[3700]);
    assign layer3_out[5751] = layer2_out[6345];
    assign layer3_out[5752] = layer2_out[3] & layer2_out[4];
    assign layer3_out[5753] = ~layer2_out[4704];
    assign layer3_out[5754] = layer2_out[137] & ~layer2_out[136];
    assign layer3_out[5755] = ~(layer2_out[520] ^ layer2_out[521]);
    assign layer3_out[5756] = ~layer2_out[3723] | layer2_out[3724];
    assign layer3_out[5757] = layer2_out[6822];
    assign layer3_out[5758] = ~(layer2_out[6400] | layer2_out[6401]);
    assign layer3_out[5759] = 1'b0;
    assign layer3_out[5760] = layer2_out[4736] & ~layer2_out[4735];
    assign layer3_out[5761] = ~layer2_out[3931];
    assign layer3_out[5762] = layer2_out[129];
    assign layer3_out[5763] = ~layer2_out[5490] | layer2_out[5491];
    assign layer3_out[5764] = layer2_out[3061] ^ layer2_out[3062];
    assign layer3_out[5765] = layer2_out[31];
    assign layer3_out[5766] = ~layer2_out[5169];
    assign layer3_out[5767] = layer2_out[531] & ~layer2_out[532];
    assign layer3_out[5768] = layer2_out[6335];
    assign layer3_out[5769] = layer2_out[4669];
    assign layer3_out[5770] = layer2_out[7464] & ~layer2_out[7463];
    assign layer3_out[5771] = layer2_out[5484];
    assign layer3_out[5772] = layer2_out[5256] ^ layer2_out[5257];
    assign layer3_out[5773] = layer2_out[1097] & ~layer2_out[1098];
    assign layer3_out[5774] = ~layer2_out[616] | layer2_out[617];
    assign layer3_out[5775] = ~(layer2_out[7926] ^ layer2_out[7927]);
    assign layer3_out[5776] = layer2_out[5387];
    assign layer3_out[5777] = ~layer2_out[3024];
    assign layer3_out[5778] = ~layer2_out[1396];
    assign layer3_out[5779] = layer2_out[143] & layer2_out[144];
    assign layer3_out[5780] = ~(layer2_out[90] ^ layer2_out[91]);
    assign layer3_out[5781] = 1'b0;
    assign layer3_out[5782] = layer2_out[3599];
    assign layer3_out[5783] = layer2_out[2157];
    assign layer3_out[5784] = ~layer2_out[5974];
    assign layer3_out[5785] = layer2_out[2927] | layer2_out[2928];
    assign layer3_out[5786] = ~layer2_out[7704];
    assign layer3_out[5787] = ~(layer2_out[7351] | layer2_out[7352]);
    assign layer3_out[5788] = layer2_out[5115] & ~layer2_out[5114];
    assign layer3_out[5789] = ~layer2_out[3956];
    assign layer3_out[5790] = ~layer2_out[1410] | layer2_out[1411];
    assign layer3_out[5791] = 1'b1;
    assign layer3_out[5792] = ~layer2_out[6432];
    assign layer3_out[5793] = ~layer2_out[2946] | layer2_out[2947];
    assign layer3_out[5794] = layer2_out[5608] | layer2_out[5609];
    assign layer3_out[5795] = layer2_out[2503] & layer2_out[2504];
    assign layer3_out[5796] = ~layer2_out[7791];
    assign layer3_out[5797] = layer2_out[2214];
    assign layer3_out[5798] = ~layer2_out[5676] | layer2_out[5677];
    assign layer3_out[5799] = layer2_out[6834];
    assign layer3_out[5800] = layer2_out[7609];
    assign layer3_out[5801] = layer2_out[3525];
    assign layer3_out[5802] = layer2_out[5331] & ~layer2_out[5332];
    assign layer3_out[5803] = layer2_out[7303] | layer2_out[7304];
    assign layer3_out[5804] = layer2_out[2223];
    assign layer3_out[5805] = layer2_out[2656];
    assign layer3_out[5806] = ~(layer2_out[6467] ^ layer2_out[6468]);
    assign layer3_out[5807] = ~layer2_out[6055] | layer2_out[6054];
    assign layer3_out[5808] = layer2_out[367] & ~layer2_out[366];
    assign layer3_out[5809] = ~layer2_out[7211];
    assign layer3_out[5810] = 1'b0;
    assign layer3_out[5811] = ~layer2_out[5179];
    assign layer3_out[5812] = layer2_out[4396] | layer2_out[4397];
    assign layer3_out[5813] = ~layer2_out[843] | layer2_out[842];
    assign layer3_out[5814] = layer2_out[3279];
    assign layer3_out[5815] = layer2_out[1031];
    assign layer3_out[5816] = ~layer2_out[7427];
    assign layer3_out[5817] = layer2_out[6692];
    assign layer3_out[5818] = layer2_out[1449];
    assign layer3_out[5819] = ~layer2_out[7145];
    assign layer3_out[5820] = ~layer2_out[2090] | layer2_out[2091];
    assign layer3_out[5821] = layer2_out[952] & ~layer2_out[953];
    assign layer3_out[5822] = layer2_out[1717] ^ layer2_out[1718];
    assign layer3_out[5823] = ~layer2_out[3461];
    assign layer3_out[5824] = ~layer2_out[5403] | layer2_out[5402];
    assign layer3_out[5825] = layer2_out[5711] & ~layer2_out[5710];
    assign layer3_out[5826] = layer2_out[5740] | layer2_out[5741];
    assign layer3_out[5827] = ~(layer2_out[7184] ^ layer2_out[7185]);
    assign layer3_out[5828] = layer2_out[183];
    assign layer3_out[5829] = layer2_out[4388] & ~layer2_out[4389];
    assign layer3_out[5830] = layer2_out[3811];
    assign layer3_out[5831] = layer2_out[5384];
    assign layer3_out[5832] = layer2_out[5819] | layer2_out[5820];
    assign layer3_out[5833] = ~(layer2_out[6986] ^ layer2_out[6987]);
    assign layer3_out[5834] = layer2_out[7954] ^ layer2_out[7955];
    assign layer3_out[5835] = ~layer2_out[4523];
    assign layer3_out[5836] = ~layer2_out[5262] | layer2_out[5261];
    assign layer3_out[5837] = layer2_out[2116] & layer2_out[2117];
    assign layer3_out[5838] = ~layer2_out[2784];
    assign layer3_out[5839] = layer2_out[7437];
    assign layer3_out[5840] = layer2_out[3149];
    assign layer3_out[5841] = layer2_out[2942] & ~layer2_out[2943];
    assign layer3_out[5842] = layer2_out[7651] & ~layer2_out[7650];
    assign layer3_out[5843] = ~layer2_out[936];
    assign layer3_out[5844] = layer2_out[7129] & ~layer2_out[7128];
    assign layer3_out[5845] = ~(layer2_out[5601] ^ layer2_out[5602]);
    assign layer3_out[5846] = ~layer2_out[6349] | layer2_out[6350];
    assign layer3_out[5847] = layer2_out[7578] & ~layer2_out[7579];
    assign layer3_out[5848] = layer2_out[5765] & layer2_out[5766];
    assign layer3_out[5849] = ~layer2_out[2986] | layer2_out[2987];
    assign layer3_out[5850] = ~layer2_out[7123];
    assign layer3_out[5851] = ~(layer2_out[5551] ^ layer2_out[5552]);
    assign layer3_out[5852] = ~layer2_out[7393];
    assign layer3_out[5853] = ~layer2_out[5674] | layer2_out[5675];
    assign layer3_out[5854] = ~(layer2_out[4970] | layer2_out[4971]);
    assign layer3_out[5855] = 1'b0;
    assign layer3_out[5856] = ~layer2_out[289];
    assign layer3_out[5857] = layer2_out[130];
    assign layer3_out[5858] = ~layer2_out[7802];
    assign layer3_out[5859] = ~(layer2_out[1999] | layer2_out[2000]);
    assign layer3_out[5860] = ~(layer2_out[5343] | layer2_out[5344]);
    assign layer3_out[5861] = layer2_out[7674] & layer2_out[7675];
    assign layer3_out[5862] = ~layer2_out[3718] | layer2_out[3717];
    assign layer3_out[5863] = ~layer2_out[3174];
    assign layer3_out[5864] = layer2_out[6252] & ~layer2_out[6251];
    assign layer3_out[5865] = layer2_out[2987];
    assign layer3_out[5866] = layer2_out[6525];
    assign layer3_out[5867] = ~layer2_out[210];
    assign layer3_out[5868] = ~(layer2_out[5953] & layer2_out[5954]);
    assign layer3_out[5869] = layer2_out[5209] & ~layer2_out[5210];
    assign layer3_out[5870] = ~layer2_out[3640];
    assign layer3_out[5871] = layer2_out[665] & ~layer2_out[664];
    assign layer3_out[5872] = layer2_out[7993];
    assign layer3_out[5873] = ~layer2_out[6749] | layer2_out[6750];
    assign layer3_out[5874] = layer2_out[2167] & layer2_out[2168];
    assign layer3_out[5875] = 1'b0;
    assign layer3_out[5876] = ~(layer2_out[2297] & layer2_out[2298]);
    assign layer3_out[5877] = ~layer2_out[7078];
    assign layer3_out[5878] = layer2_out[4823] & ~layer2_out[4822];
    assign layer3_out[5879] = ~layer2_out[7522];
    assign layer3_out[5880] = ~layer2_out[2461];
    assign layer3_out[5881] = layer2_out[1418];
    assign layer3_out[5882] = layer2_out[5896] & ~layer2_out[5897];
    assign layer3_out[5883] = layer2_out[7265] & ~layer2_out[7264];
    assign layer3_out[5884] = layer2_out[4268] | layer2_out[4269];
    assign layer3_out[5885] = layer2_out[6531] & layer2_out[6532];
    assign layer3_out[5886] = layer2_out[5782] ^ layer2_out[5783];
    assign layer3_out[5887] = ~layer2_out[6184];
    assign layer3_out[5888] = layer2_out[2806] & ~layer2_out[2805];
    assign layer3_out[5889] = ~layer2_out[254];
    assign layer3_out[5890] = ~layer2_out[5838];
    assign layer3_out[5891] = layer2_out[4681];
    assign layer3_out[5892] = ~layer2_out[1163];
    assign layer3_out[5893] = layer2_out[632] & ~layer2_out[631];
    assign layer3_out[5894] = ~(layer2_out[4023] | layer2_out[4024]);
    assign layer3_out[5895] = ~layer2_out[3022];
    assign layer3_out[5896] = layer2_out[7906];
    assign layer3_out[5897] = ~layer2_out[132];
    assign layer3_out[5898] = layer2_out[1177];
    assign layer3_out[5899] = layer2_out[1817] & layer2_out[1818];
    assign layer3_out[5900] = layer2_out[6954] & ~layer2_out[6953];
    assign layer3_out[5901] = layer2_out[3807] & layer2_out[3808];
    assign layer3_out[5902] = layer2_out[5541] ^ layer2_out[5542];
    assign layer3_out[5903] = layer2_out[1872];
    assign layer3_out[5904] = ~(layer2_out[7671] & layer2_out[7672]);
    assign layer3_out[5905] = ~layer2_out[7022];
    assign layer3_out[5906] = layer2_out[6211] & layer2_out[6212];
    assign layer3_out[5907] = ~layer2_out[7549] | layer2_out[7550];
    assign layer3_out[5908] = layer2_out[451];
    assign layer3_out[5909] = ~layer2_out[6249];
    assign layer3_out[5910] = layer2_out[3178];
    assign layer3_out[5911] = ~(layer2_out[3694] ^ layer2_out[3695]);
    assign layer3_out[5912] = layer2_out[3392];
    assign layer3_out[5913] = 1'b1;
    assign layer3_out[5914] = ~layer2_out[1361];
    assign layer3_out[5915] = ~layer2_out[7333];
    assign layer3_out[5916] = ~layer2_out[1029];
    assign layer3_out[5917] = layer2_out[7568];
    assign layer3_out[5918] = layer2_out[6835];
    assign layer3_out[5919] = layer2_out[3416];
    assign layer3_out[5920] = layer2_out[6723];
    assign layer3_out[5921] = layer2_out[2118];
    assign layer3_out[5922] = ~layer2_out[7089];
    assign layer3_out[5923] = layer2_out[4945] | layer2_out[4946];
    assign layer3_out[5924] = layer2_out[809];
    assign layer3_out[5925] = ~layer2_out[4788] | layer2_out[4787];
    assign layer3_out[5926] = ~layer2_out[6816];
    assign layer3_out[5927] = ~(layer2_out[4242] | layer2_out[4243]);
    assign layer3_out[5928] = ~layer2_out[3314];
    assign layer3_out[5929] = ~layer2_out[4233];
    assign layer3_out[5930] = layer2_out[7453] & ~layer2_out[7454];
    assign layer3_out[5931] = layer2_out[3090] & layer2_out[3091];
    assign layer3_out[5932] = ~layer2_out[1573];
    assign layer3_out[5933] = ~layer2_out[6544];
    assign layer3_out[5934] = ~(layer2_out[1806] ^ layer2_out[1807]);
    assign layer3_out[5935] = layer2_out[1152];
    assign layer3_out[5936] = ~layer2_out[440];
    assign layer3_out[5937] = ~layer2_out[6942];
    assign layer3_out[5938] = ~layer2_out[3064] | layer2_out[3063];
    assign layer3_out[5939] = layer2_out[3643];
    assign layer3_out[5940] = ~layer2_out[1503] | layer2_out[1504];
    assign layer3_out[5941] = ~layer2_out[5440] | layer2_out[5441];
    assign layer3_out[5942] = ~layer2_out[4743];
    assign layer3_out[5943] = 1'b1;
    assign layer3_out[5944] = layer2_out[4872] & ~layer2_out[4873];
    assign layer3_out[5945] = layer2_out[426] ^ layer2_out[427];
    assign layer3_out[5946] = ~layer2_out[5107];
    assign layer3_out[5947] = ~layer2_out[7108];
    assign layer3_out[5948] = ~(layer2_out[5157] ^ layer2_out[5158]);
    assign layer3_out[5949] = layer2_out[7843] & layer2_out[7844];
    assign layer3_out[5950] = ~(layer2_out[1766] & layer2_out[1767]);
    assign layer3_out[5951] = ~(layer2_out[6685] | layer2_out[6686]);
    assign layer3_out[5952] = layer2_out[2279];
    assign layer3_out[5953] = ~(layer2_out[6619] & layer2_out[6620]);
    assign layer3_out[5954] = ~layer2_out[1668];
    assign layer3_out[5955] = ~layer2_out[190] | layer2_out[189];
    assign layer3_out[5956] = ~layer2_out[1343];
    assign layer3_out[5957] = ~layer2_out[257];
    assign layer3_out[5958] = ~(layer2_out[6884] & layer2_out[6885]);
    assign layer3_out[5959] = layer2_out[5508] | layer2_out[5509];
    assign layer3_out[5960] = layer2_out[5411] | layer2_out[5412];
    assign layer3_out[5961] = ~layer2_out[7204];
    assign layer3_out[5962] = ~layer2_out[3928];
    assign layer3_out[5963] = layer2_out[3975];
    assign layer3_out[5964] = ~layer2_out[7013];
    assign layer3_out[5965] = layer2_out[6332] & ~layer2_out[6331];
    assign layer3_out[5966] = ~layer2_out[4656] | layer2_out[4655];
    assign layer3_out[5967] = ~(layer2_out[7013] ^ layer2_out[7014]);
    assign layer3_out[5968] = layer2_out[5134] & layer2_out[5135];
    assign layer3_out[5969] = ~layer2_out[1825];
    assign layer3_out[5970] = ~(layer2_out[6873] & layer2_out[6874]);
    assign layer3_out[5971] = layer2_out[3909];
    assign layer3_out[5972] = ~layer2_out[14];
    assign layer3_out[5973] = layer2_out[3023];
    assign layer3_out[5974] = layer2_out[1042] & ~layer2_out[1043];
    assign layer3_out[5975] = layer2_out[5432];
    assign layer3_out[5976] = layer2_out[6168] & layer2_out[6169];
    assign layer3_out[5977] = ~(layer2_out[7766] ^ layer2_out[7767]);
    assign layer3_out[5978] = ~layer2_out[5127];
    assign layer3_out[5979] = ~layer2_out[5645];
    assign layer3_out[5980] = ~layer2_out[806];
    assign layer3_out[5981] = ~(layer2_out[4692] | layer2_out[4693]);
    assign layer3_out[5982] = layer2_out[3424];
    assign layer3_out[5983] = layer2_out[3293] ^ layer2_out[3294];
    assign layer3_out[5984] = ~layer2_out[4470];
    assign layer3_out[5985] = layer2_out[3430] & ~layer2_out[3429];
    assign layer3_out[5986] = ~layer2_out[6031] | layer2_out[6032];
    assign layer3_out[5987] = ~layer2_out[3437];
    assign layer3_out[5988] = layer2_out[3267] & ~layer2_out[3268];
    assign layer3_out[5989] = layer2_out[5240];
    assign layer3_out[5990] = 1'b1;
    assign layer3_out[5991] = layer2_out[3046];
    assign layer3_out[5992] = ~(layer2_out[4839] & layer2_out[4840]);
    assign layer3_out[5993] = layer2_out[3604] & ~layer2_out[3605];
    assign layer3_out[5994] = ~layer2_out[4964] | layer2_out[4963];
    assign layer3_out[5995] = layer2_out[7548] & ~layer2_out[7549];
    assign layer3_out[5996] = layer2_out[1254] & layer2_out[1255];
    assign layer3_out[5997] = ~(layer2_out[3680] & layer2_out[3681]);
    assign layer3_out[5998] = layer2_out[5448];
    assign layer3_out[5999] = ~(layer2_out[1899] | layer2_out[1900]);
    assign layer3_out[6000] = ~layer2_out[7986];
    assign layer3_out[6001] = layer2_out[5457];
    assign layer3_out[6002] = layer2_out[3669];
    assign layer3_out[6003] = layer2_out[5310] | layer2_out[5311];
    assign layer3_out[6004] = ~layer2_out[2790];
    assign layer3_out[6005] = layer2_out[7914] & layer2_out[7915];
    assign layer3_out[6006] = ~layer2_out[7733];
    assign layer3_out[6007] = ~(layer2_out[2095] & layer2_out[2096]);
    assign layer3_out[6008] = layer2_out[1585];
    assign layer3_out[6009] = ~(layer2_out[6066] | layer2_out[6067]);
    assign layer3_out[6010] = layer2_out[5975];
    assign layer3_out[6011] = ~layer2_out[1181];
    assign layer3_out[6012] = ~layer2_out[858];
    assign layer3_out[6013] = layer2_out[457] & ~layer2_out[456];
    assign layer3_out[6014] = ~layer2_out[4384];
    assign layer3_out[6015] = layer2_out[4099] & layer2_out[4100];
    assign layer3_out[6016] = ~layer2_out[6877];
    assign layer3_out[6017] = ~(layer2_out[5542] & layer2_out[5543]);
    assign layer3_out[6018] = layer2_out[4498] & ~layer2_out[4497];
    assign layer3_out[6019] = ~(layer2_out[3576] ^ layer2_out[3577]);
    assign layer3_out[6020] = ~layer2_out[5129] | layer2_out[5128];
    assign layer3_out[6021] = ~layer2_out[4286];
    assign layer3_out[6022] = ~(layer2_out[4798] | layer2_out[4799]);
    assign layer3_out[6023] = ~layer2_out[5661];
    assign layer3_out[6024] = ~(layer2_out[7456] ^ layer2_out[7457]);
    assign layer3_out[6025] = layer2_out[4401];
    assign layer3_out[6026] = ~layer2_out[3638];
    assign layer3_out[6027] = ~layer2_out[7531] | layer2_out[7530];
    assign layer3_out[6028] = layer2_out[4952];
    assign layer3_out[6029] = layer2_out[5027];
    assign layer3_out[6030] = ~layer2_out[2154];
    assign layer3_out[6031] = ~layer2_out[2306] | layer2_out[2307];
    assign layer3_out[6032] = ~layer2_out[5116];
    assign layer3_out[6033] = ~layer2_out[2560];
    assign layer3_out[6034] = ~(layer2_out[1689] & layer2_out[1690]);
    assign layer3_out[6035] = ~layer2_out[3344];
    assign layer3_out[6036] = layer2_out[315] & layer2_out[316];
    assign layer3_out[6037] = layer2_out[3235] & ~layer2_out[3236];
    assign layer3_out[6038] = layer2_out[3773];
    assign layer3_out[6039] = ~layer2_out[4804];
    assign layer3_out[6040] = ~(layer2_out[2618] ^ layer2_out[2619]);
    assign layer3_out[6041] = ~(layer2_out[3053] | layer2_out[3054]);
    assign layer3_out[6042] = layer2_out[5266] ^ layer2_out[5267];
    assign layer3_out[6043] = layer2_out[7403] & ~layer2_out[7404];
    assign layer3_out[6044] = layer2_out[7903];
    assign layer3_out[6045] = layer2_out[3201];
    assign layer3_out[6046] = ~layer2_out[640] | layer2_out[639];
    assign layer3_out[6047] = ~layer2_out[5360] | layer2_out[5361];
    assign layer3_out[6048] = ~(layer2_out[1703] ^ layer2_out[1704]);
    assign layer3_out[6049] = ~layer2_out[395];
    assign layer3_out[6050] = ~(layer2_out[5368] | layer2_out[5369]);
    assign layer3_out[6051] = layer2_out[3129] ^ layer2_out[3130];
    assign layer3_out[6052] = ~(layer2_out[2520] & layer2_out[2521]);
    assign layer3_out[6053] = layer2_out[4914];
    assign layer3_out[6054] = layer2_out[3272];
    assign layer3_out[6055] = ~layer2_out[4254] | layer2_out[4255];
    assign layer3_out[6056] = layer2_out[1236] ^ layer2_out[1237];
    assign layer3_out[6057] = ~(layer2_out[2634] | layer2_out[2635]);
    assign layer3_out[6058] = layer2_out[5220];
    assign layer3_out[6059] = ~(layer2_out[2970] & layer2_out[2971]);
    assign layer3_out[6060] = layer2_out[1290] & layer2_out[1291];
    assign layer3_out[6061] = ~layer2_out[941];
    assign layer3_out[6062] = ~(layer2_out[1400] | layer2_out[1401]);
    assign layer3_out[6063] = layer2_out[6323] | layer2_out[6324];
    assign layer3_out[6064] = layer2_out[197];
    assign layer3_out[6065] = ~(layer2_out[3836] & layer2_out[3837]);
    assign layer3_out[6066] = ~(layer2_out[7673] & layer2_out[7674]);
    assign layer3_out[6067] = layer2_out[409] & ~layer2_out[410];
    assign layer3_out[6068] = ~(layer2_out[3624] | layer2_out[3625]);
    assign layer3_out[6069] = layer2_out[5738] & ~layer2_out[5737];
    assign layer3_out[6070] = ~(layer2_out[2024] & layer2_out[2025]);
    assign layer3_out[6071] = ~layer2_out[3463];
    assign layer3_out[6072] = layer2_out[2023] ^ layer2_out[2024];
    assign layer3_out[6073] = layer2_out[2494] & ~layer2_out[2495];
    assign layer3_out[6074] = ~layer2_out[1535];
    assign layer3_out[6075] = ~layer2_out[4567] | layer2_out[4566];
    assign layer3_out[6076] = layer2_out[4654] | layer2_out[4655];
    assign layer3_out[6077] = ~layer2_out[691] | layer2_out[692];
    assign layer3_out[6078] = ~(layer2_out[6035] ^ layer2_out[6036]);
    assign layer3_out[6079] = layer2_out[848];
    assign layer3_out[6080] = layer2_out[2301];
    assign layer3_out[6081] = layer2_out[1577] & ~layer2_out[1576];
    assign layer3_out[6082] = ~layer2_out[4106] | layer2_out[4105];
    assign layer3_out[6083] = layer2_out[5671];
    assign layer3_out[6084] = layer2_out[2036];
    assign layer3_out[6085] = layer2_out[923] & layer2_out[924];
    assign layer3_out[6086] = layer2_out[1570];
    assign layer3_out[6087] = ~layer2_out[7442] | layer2_out[7441];
    assign layer3_out[6088] = layer2_out[5012] | layer2_out[5013];
    assign layer3_out[6089] = layer2_out[4828] ^ layer2_out[4829];
    assign layer3_out[6090] = ~layer2_out[4444] | layer2_out[4443];
    assign layer3_out[6091] = ~(layer2_out[2911] & layer2_out[2912]);
    assign layer3_out[6092] = layer2_out[3736] ^ layer2_out[3737];
    assign layer3_out[6093] = layer2_out[6750] & ~layer2_out[6751];
    assign layer3_out[6094] = ~(layer2_out[6260] | layer2_out[6261]);
    assign layer3_out[6095] = layer2_out[4891] ^ layer2_out[4892];
    assign layer3_out[6096] = ~layer2_out[4548];
    assign layer3_out[6097] = layer2_out[7181] & ~layer2_out[7180];
    assign layer3_out[6098] = 1'b0;
    assign layer3_out[6099] = ~(layer2_out[1382] | layer2_out[1383]);
    assign layer3_out[6100] = ~(layer2_out[7458] | layer2_out[7459]);
    assign layer3_out[6101] = ~layer2_out[2592] | layer2_out[2593];
    assign layer3_out[6102] = layer2_out[710] & ~layer2_out[711];
    assign layer3_out[6103] = ~layer2_out[2194];
    assign layer3_out[6104] = ~(layer2_out[5405] | layer2_out[5406]);
    assign layer3_out[6105] = layer2_out[598] & layer2_out[599];
    assign layer3_out[6106] = ~(layer2_out[7289] | layer2_out[7290]);
    assign layer3_out[6107] = layer2_out[7691] & ~layer2_out[7690];
    assign layer3_out[6108] = ~layer2_out[4748];
    assign layer3_out[6109] = ~layer2_out[446];
    assign layer3_out[6110] = layer2_out[3635];
    assign layer3_out[6111] = layer2_out[4814] & ~layer2_out[4815];
    assign layer3_out[6112] = layer2_out[2609] ^ layer2_out[2610];
    assign layer3_out[6113] = layer2_out[7692];
    assign layer3_out[6114] = ~(layer2_out[1423] ^ layer2_out[1424]);
    assign layer3_out[6115] = layer2_out[6940] & ~layer2_out[6939];
    assign layer3_out[6116] = ~layer2_out[3162] | layer2_out[3163];
    assign layer3_out[6117] = ~(layer2_out[7529] | layer2_out[7530]);
    assign layer3_out[6118] = ~layer2_out[6447] | layer2_out[6446];
    assign layer3_out[6119] = ~layer2_out[2472];
    assign layer3_out[6120] = layer2_out[6381];
    assign layer3_out[6121] = ~layer2_out[7983];
    assign layer3_out[6122] = ~layer2_out[246];
    assign layer3_out[6123] = layer2_out[7390];
    assign layer3_out[6124] = ~layer2_out[5916];
    assign layer3_out[6125] = layer2_out[6960];
    assign layer3_out[6126] = layer2_out[973] & ~layer2_out[972];
    assign layer3_out[6127] = layer2_out[4764] & layer2_out[4765];
    assign layer3_out[6128] = ~layer2_out[4194] | layer2_out[4193];
    assign layer3_out[6129] = layer2_out[6295];
    assign layer3_out[6130] = layer2_out[1068] & ~layer2_out[1069];
    assign layer3_out[6131] = ~layer2_out[5383] | layer2_out[5382];
    assign layer3_out[6132] = ~layer2_out[489] | layer2_out[488];
    assign layer3_out[6133] = ~layer2_out[6555] | layer2_out[6554];
    assign layer3_out[6134] = ~layer2_out[6642];
    assign layer3_out[6135] = ~(layer2_out[2607] ^ layer2_out[2608]);
    assign layer3_out[6136] = ~layer2_out[2178] | layer2_out[2179];
    assign layer3_out[6137] = ~(layer2_out[4367] & layer2_out[4368]);
    assign layer3_out[6138] = layer2_out[4884];
    assign layer3_out[6139] = ~layer2_out[2616];
    assign layer3_out[6140] = ~(layer2_out[6237] | layer2_out[6238]);
    assign layer3_out[6141] = layer2_out[4138];
    assign layer3_out[6142] = ~layer2_out[4575] | layer2_out[4576];
    assign layer3_out[6143] = layer2_out[719] ^ layer2_out[720];
    assign layer3_out[6144] = layer2_out[3758] & ~layer2_out[3757];
    assign layer3_out[6145] = layer2_out[5043] & ~layer2_out[5042];
    assign layer3_out[6146] = 1'b0;
    assign layer3_out[6147] = layer2_out[3790] ^ layer2_out[3791];
    assign layer3_out[6148] = ~layer2_out[5998];
    assign layer3_out[6149] = layer2_out[6088];
    assign layer3_out[6150] = layer2_out[3200] & ~layer2_out[3199];
    assign layer3_out[6151] = ~layer2_out[670];
    assign layer3_out[6152] = layer2_out[3864] & ~layer2_out[3865];
    assign layer3_out[6153] = ~layer2_out[5386];
    assign layer3_out[6154] = layer2_out[243] ^ layer2_out[244];
    assign layer3_out[6155] = ~layer2_out[1181];
    assign layer3_out[6156] = ~layer2_out[3972] | layer2_out[3971];
    assign layer3_out[6157] = layer2_out[7782];
    assign layer3_out[6158] = layer2_out[2069] | layer2_out[2070];
    assign layer3_out[6159] = layer2_out[311] ^ layer2_out[312];
    assign layer3_out[6160] = ~(layer2_out[1244] & layer2_out[1245]);
    assign layer3_out[6161] = ~(layer2_out[94] & layer2_out[95]);
    assign layer3_out[6162] = 1'b0;
    assign layer3_out[6163] = layer2_out[3517];
    assign layer3_out[6164] = layer2_out[2845];
    assign layer3_out[6165] = layer2_out[824] ^ layer2_out[825];
    assign layer3_out[6166] = ~layer2_out[4613];
    assign layer3_out[6167] = layer2_out[1958];
    assign layer3_out[6168] = layer2_out[1679] | layer2_out[1680];
    assign layer3_out[6169] = layer2_out[5415] & ~layer2_out[5416];
    assign layer3_out[6170] = ~layer2_out[2871] | layer2_out[2872];
    assign layer3_out[6171] = ~(layer2_out[3891] ^ layer2_out[3892]);
    assign layer3_out[6172] = ~layer2_out[5236] | layer2_out[5237];
    assign layer3_out[6173] = layer2_out[5075] ^ layer2_out[5076];
    assign layer3_out[6174] = layer2_out[7481];
    assign layer3_out[6175] = layer2_out[5948];
    assign layer3_out[6176] = ~layer2_out[3862];
    assign layer3_out[6177] = ~(layer2_out[3430] & layer2_out[3431]);
    assign layer3_out[6178] = ~layer2_out[2404];
    assign layer3_out[6179] = ~layer2_out[3264];
    assign layer3_out[6180] = ~layer2_out[3208];
    assign layer3_out[6181] = layer2_out[2413] & ~layer2_out[2412];
    assign layer3_out[6182] = layer2_out[7490] & layer2_out[7491];
    assign layer3_out[6183] = ~layer2_out[5567];
    assign layer3_out[6184] = layer2_out[895] & layer2_out[896];
    assign layer3_out[6185] = ~layer2_out[2390];
    assign layer3_out[6186] = layer2_out[990] & ~layer2_out[991];
    assign layer3_out[6187] = layer2_out[1633];
    assign layer3_out[6188] = 1'b1;
    assign layer3_out[6189] = ~layer2_out[5210];
    assign layer3_out[6190] = ~(layer2_out[3898] | layer2_out[3899]);
    assign layer3_out[6191] = layer2_out[2963] & ~layer2_out[2962];
    assign layer3_out[6192] = layer2_out[4250];
    assign layer3_out[6193] = ~layer2_out[6458];
    assign layer3_out[6194] = layer2_out[7750];
    assign layer3_out[6195] = layer2_out[4522];
    assign layer3_out[6196] = layer2_out[4023];
    assign layer3_out[6197] = ~layer2_out[3086] | layer2_out[3085];
    assign layer3_out[6198] = layer2_out[4258] ^ layer2_out[4259];
    assign layer3_out[6199] = ~layer2_out[3501] | layer2_out[3500];
    assign layer3_out[6200] = layer2_out[97];
    assign layer3_out[6201] = ~layer2_out[2696];
    assign layer3_out[6202] = layer2_out[6592];
    assign layer3_out[6203] = layer2_out[5992];
    assign layer3_out[6204] = 1'b0;
    assign layer3_out[6205] = layer2_out[5616] & ~layer2_out[5617];
    assign layer3_out[6206] = layer2_out[3872] & ~layer2_out[3873];
    assign layer3_out[6207] = ~layer2_out[7296];
    assign layer3_out[6208] = ~(layer2_out[6278] ^ layer2_out[6279]);
    assign layer3_out[6209] = layer2_out[1859] & layer2_out[1860];
    assign layer3_out[6210] = ~layer2_out[264] | layer2_out[265];
    assign layer3_out[6211] = layer2_out[3499] & layer2_out[3500];
    assign layer3_out[6212] = layer2_out[6217] & layer2_out[6218];
    assign layer3_out[6213] = ~(layer2_out[2534] & layer2_out[2535]);
    assign layer3_out[6214] = layer2_out[2297];
    assign layer3_out[6215] = layer2_out[6178] & ~layer2_out[6177];
    assign layer3_out[6216] = ~layer2_out[3327] | layer2_out[3326];
    assign layer3_out[6217] = ~layer2_out[2563];
    assign layer3_out[6218] = ~layer2_out[3239];
    assign layer3_out[6219] = layer2_out[4780];
    assign layer3_out[6220] = layer2_out[4578] | layer2_out[4579];
    assign layer3_out[6221] = layer2_out[2357] & layer2_out[2358];
    assign layer3_out[6222] = layer2_out[5593];
    assign layer3_out[6223] = layer2_out[7996] | layer2_out[7997];
    assign layer3_out[6224] = layer2_out[4990];
    assign layer3_out[6225] = layer2_out[2351];
    assign layer3_out[6226] = layer2_out[133];
    assign layer3_out[6227] = layer2_out[1993];
    assign layer3_out[6228] = layer2_out[2091] | layer2_out[2092];
    assign layer3_out[6229] = ~layer2_out[6449] | layer2_out[6450];
    assign layer3_out[6230] = ~layer2_out[1846];
    assign layer3_out[6231] = ~layer2_out[5739] | layer2_out[5738];
    assign layer3_out[6232] = ~layer2_out[6355] | layer2_out[6356];
    assign layer3_out[6233] = ~layer2_out[5215];
    assign layer3_out[6234] = ~layer2_out[7596];
    assign layer3_out[6235] = layer2_out[212];
    assign layer3_out[6236] = layer2_out[6150] & layer2_out[6151];
    assign layer3_out[6237] = ~layer2_out[5560] | layer2_out[5559];
    assign layer3_out[6238] = ~(layer2_out[1733] & layer2_out[1734]);
    assign layer3_out[6239] = ~layer2_out[1020];
    assign layer3_out[6240] = layer2_out[3094] & ~layer2_out[3093];
    assign layer3_out[6241] = layer2_out[2661] & ~layer2_out[2660];
    assign layer3_out[6242] = ~layer2_out[1339];
    assign layer3_out[6243] = ~layer2_out[5139];
    assign layer3_out[6244] = ~(layer2_out[6004] ^ layer2_out[6005]);
    assign layer3_out[6245] = 1'b0;
    assign layer3_out[6246] = layer2_out[3117];
    assign layer3_out[6247] = layer2_out[5043];
    assign layer3_out[6248] = layer2_out[3112] & ~layer2_out[3113];
    assign layer3_out[6249] = layer2_out[391] | layer2_out[392];
    assign layer3_out[6250] = ~layer2_out[6494];
    assign layer3_out[6251] = ~layer2_out[1193];
    assign layer3_out[6252] = layer2_out[7748];
    assign layer3_out[6253] = ~layer2_out[5683] | layer2_out[5682];
    assign layer3_out[6254] = ~layer2_out[4524] | layer2_out[4525];
    assign layer3_out[6255] = ~layer2_out[7309] | layer2_out[7308];
    assign layer3_out[6256] = layer2_out[6625] | layer2_out[6626];
    assign layer3_out[6257] = layer2_out[7929] & ~layer2_out[7928];
    assign layer3_out[6258] = ~(layer2_out[3325] | layer2_out[3326]);
    assign layer3_out[6259] = ~(layer2_out[2288] | layer2_out[2289]);
    assign layer3_out[6260] = ~(layer2_out[7339] | layer2_out[7340]);
    assign layer3_out[6261] = ~(layer2_out[1746] ^ layer2_out[1747]);
    assign layer3_out[6262] = layer2_out[4215] | layer2_out[4216];
    assign layer3_out[6263] = layer2_out[4812] & ~layer2_out[4813];
    assign layer3_out[6264] = layer2_out[3396];
    assign layer3_out[6265] = layer2_out[2349];
    assign layer3_out[6266] = ~(layer2_out[2657] ^ layer2_out[2658]);
    assign layer3_out[6267] = layer2_out[6698] & ~layer2_out[6697];
    assign layer3_out[6268] = ~layer2_out[7923];
    assign layer3_out[6269] = ~layer2_out[7347] | layer2_out[7348];
    assign layer3_out[6270] = layer2_out[3556];
    assign layer3_out[6271] = layer2_out[5482] | layer2_out[5483];
    assign layer3_out[6272] = ~layer2_out[1538];
    assign layer3_out[6273] = layer2_out[3895] & layer2_out[3896];
    assign layer3_out[6274] = ~(layer2_out[1621] & layer2_out[1622]);
    assign layer3_out[6275] = ~layer2_out[3376] | layer2_out[3375];
    assign layer3_out[6276] = ~(layer2_out[4941] & layer2_out[4942]);
    assign layer3_out[6277] = ~layer2_out[6702] | layer2_out[6703];
    assign layer3_out[6278] = layer2_out[552];
    assign layer3_out[6279] = layer2_out[2843] & layer2_out[2844];
    assign layer3_out[6280] = ~layer2_out[1486];
    assign layer3_out[6281] = layer2_out[3346];
    assign layer3_out[6282] = ~layer2_out[204] | layer2_out[205];
    assign layer3_out[6283] = layer2_out[6509];
    assign layer3_out[6284] = ~layer2_out[6348];
    assign layer3_out[6285] = ~layer2_out[4790];
    assign layer3_out[6286] = ~layer2_out[4867];
    assign layer3_out[6287] = ~layer2_out[3815] | layer2_out[3814];
    assign layer3_out[6288] = layer2_out[3394] & layer2_out[3395];
    assign layer3_out[6289] = ~layer2_out[138];
    assign layer3_out[6290] = layer2_out[1046] & ~layer2_out[1045];
    assign layer3_out[6291] = layer2_out[6755];
    assign layer3_out[6292] = ~(layer2_out[7397] & layer2_out[7398]);
    assign layer3_out[6293] = layer2_out[3704] & ~layer2_out[3703];
    assign layer3_out[6294] = layer2_out[4965] & layer2_out[4966];
    assign layer3_out[6295] = layer2_out[4275];
    assign layer3_out[6296] = layer2_out[4056];
    assign layer3_out[6297] = layer2_out[3359];
    assign layer3_out[6298] = 1'b1;
    assign layer3_out[6299] = layer2_out[2698] & layer2_out[2699];
    assign layer3_out[6300] = layer2_out[5184] ^ layer2_out[5185];
    assign layer3_out[6301] = layer2_out[7053];
    assign layer3_out[6302] = layer2_out[7354] | layer2_out[7355];
    assign layer3_out[6303] = ~layer2_out[7023] | layer2_out[7024];
    assign layer3_out[6304] = 1'b0;
    assign layer3_out[6305] = ~layer2_out[4097];
    assign layer3_out[6306] = ~layer2_out[5879];
    assign layer3_out[6307] = layer2_out[683] ^ layer2_out[684];
    assign layer3_out[6308] = layer2_out[6524] & ~layer2_out[6523];
    assign layer3_out[6309] = ~(layer2_out[1363] | layer2_out[1364]);
    assign layer3_out[6310] = ~layer2_out[2634] | layer2_out[2633];
    assign layer3_out[6311] = layer2_out[3904] | layer2_out[3905];
    assign layer3_out[6312] = layer2_out[7910];
    assign layer3_out[6313] = ~layer2_out[6357];
    assign layer3_out[6314] = ~layer2_out[5535];
    assign layer3_out[6315] = layer2_out[2360] ^ layer2_out[2361];
    assign layer3_out[6316] = ~(layer2_out[6077] | layer2_out[6078]);
    assign layer3_out[6317] = ~layer2_out[7715] | layer2_out[7716];
    assign layer3_out[6318] = layer2_out[5830] | layer2_out[5831];
    assign layer3_out[6319] = layer2_out[2388];
    assign layer3_out[6320] = layer2_out[2503] & ~layer2_out[2502];
    assign layer3_out[6321] = ~layer2_out[6492] | layer2_out[6493];
    assign layer3_out[6322] = ~layer2_out[3966];
    assign layer3_out[6323] = ~layer2_out[2570];
    assign layer3_out[6324] = layer2_out[1339];
    assign layer3_out[6325] = ~(layer2_out[6804] & layer2_out[6805]);
    assign layer3_out[6326] = layer2_out[4238];
    assign layer3_out[6327] = ~layer2_out[2065];
    assign layer3_out[6328] = layer2_out[6989];
    assign layer3_out[6329] = layer2_out[6016] & ~layer2_out[6017];
    assign layer3_out[6330] = layer2_out[6263] | layer2_out[6264];
    assign layer3_out[6331] = ~(layer2_out[2481] | layer2_out[2482]);
    assign layer3_out[6332] = ~layer2_out[5648];
    assign layer3_out[6333] = ~layer2_out[3493];
    assign layer3_out[6334] = ~layer2_out[190] | layer2_out[191];
    assign layer3_out[6335] = ~layer2_out[5666];
    assign layer3_out[6336] = layer2_out[7829] | layer2_out[7830];
    assign layer3_out[6337] = ~layer2_out[831] | layer2_out[832];
    assign layer3_out[6338] = ~layer2_out[2038];
    assign layer3_out[6339] = ~layer2_out[4158];
    assign layer3_out[6340] = layer2_out[6641] ^ layer2_out[6642];
    assign layer3_out[6341] = layer2_out[4782] ^ layer2_out[4783];
    assign layer3_out[6342] = ~layer2_out[4894] | layer2_out[4893];
    assign layer3_out[6343] = ~(layer2_out[7620] & layer2_out[7621]);
    assign layer3_out[6344] = ~layer2_out[6332];
    assign layer3_out[6345] = ~(layer2_out[4744] | layer2_out[4745]);
    assign layer3_out[6346] = layer2_out[885] & layer2_out[886];
    assign layer3_out[6347] = layer2_out[6892];
    assign layer3_out[6348] = layer2_out[3467] & layer2_out[3468];
    assign layer3_out[6349] = ~layer2_out[2112];
    assign layer3_out[6350] = 1'b0;
    assign layer3_out[6351] = ~layer2_out[3122];
    assign layer3_out[6352] = layer2_out[252];
    assign layer3_out[6353] = layer2_out[7868] | layer2_out[7869];
    assign layer3_out[6354] = ~layer2_out[1820];
    assign layer3_out[6355] = layer2_out[594];
    assign layer3_out[6356] = layer2_out[2469] ^ layer2_out[2470];
    assign layer3_out[6357] = layer2_out[6115] & layer2_out[6116];
    assign layer3_out[6358] = ~layer2_out[4060];
    assign layer3_out[6359] = ~layer2_out[1506] | layer2_out[1505];
    assign layer3_out[6360] = layer2_out[4932] ^ layer2_out[4933];
    assign layer3_out[6361] = layer2_out[1823] & ~layer2_out[1824];
    assign layer3_out[6362] = layer2_out[6470] | layer2_out[6471];
    assign layer3_out[6363] = layer2_out[7053] | layer2_out[7054];
    assign layer3_out[6364] = ~(layer2_out[5295] | layer2_out[5296]);
    assign layer3_out[6365] = ~layer2_out[6168];
    assign layer3_out[6366] = layer2_out[2391];
    assign layer3_out[6367] = ~(layer2_out[6688] & layer2_out[6689]);
    assign layer3_out[6368] = layer2_out[4720] | layer2_out[4721];
    assign layer3_out[6369] = ~(layer2_out[2918] ^ layer2_out[2919]);
    assign layer3_out[6370] = layer2_out[1060];
    assign layer3_out[6371] = layer2_out[4126] & layer2_out[4127];
    assign layer3_out[6372] = 1'b1;
    assign layer3_out[6373] = ~layer2_out[919];
    assign layer3_out[6374] = ~layer2_out[6173];
    assign layer3_out[6375] = layer2_out[4727];
    assign layer3_out[6376] = layer2_out[7062] | layer2_out[7063];
    assign layer3_out[6377] = ~layer2_out[6661];
    assign layer3_out[6378] = layer2_out[6366] | layer2_out[6367];
    assign layer3_out[6379] = layer2_out[274] & layer2_out[275];
    assign layer3_out[6380] = layer2_out[5140] & ~layer2_out[5139];
    assign layer3_out[6381] = layer2_out[1972] ^ layer2_out[1973];
    assign layer3_out[6382] = 1'b0;
    assign layer3_out[6383] = layer2_out[1920] & ~layer2_out[1919];
    assign layer3_out[6384] = layer2_out[5579] & ~layer2_out[5578];
    assign layer3_out[6385] = layer2_out[4582] | layer2_out[4583];
    assign layer3_out[6386] = ~layer2_out[2334] | layer2_out[2333];
    assign layer3_out[6387] = ~(layer2_out[1962] | layer2_out[1963]);
    assign layer3_out[6388] = ~layer2_out[6138];
    assign layer3_out[6389] = ~(layer2_out[6985] & layer2_out[6986]);
    assign layer3_out[6390] = layer2_out[5254];
    assign layer3_out[6391] = ~layer2_out[454];
    assign layer3_out[6392] = layer2_out[56];
    assign layer3_out[6393] = ~layer2_out[3894];
    assign layer3_out[6394] = layer2_out[118] | layer2_out[119];
    assign layer3_out[6395] = ~layer2_out[5133] | layer2_out[5134];
    assign layer3_out[6396] = layer2_out[4036] | layer2_out[4037];
    assign layer3_out[6397] = layer2_out[953] & layer2_out[954];
    assign layer3_out[6398] = layer2_out[7071];
    assign layer3_out[6399] = ~layer2_out[7980];
    assign layer3_out[6400] = ~(layer2_out[2751] & layer2_out[2752]);
    assign layer3_out[6401] = layer2_out[259] ^ layer2_out[260];
    assign layer3_out[6402] = layer2_out[59];
    assign layer3_out[6403] = ~(layer2_out[1477] & layer2_out[1478]);
    assign layer3_out[6404] = ~layer2_out[912];
    assign layer3_out[6405] = layer2_out[2602] & layer2_out[2603];
    assign layer3_out[6406] = layer2_out[1170] ^ layer2_out[1171];
    assign layer3_out[6407] = ~(layer2_out[7986] & layer2_out[7987]);
    assign layer3_out[6408] = layer2_out[177];
    assign layer3_out[6409] = ~layer2_out[2649];
    assign layer3_out[6410] = ~layer2_out[854];
    assign layer3_out[6411] = layer2_out[3587] ^ layer2_out[3588];
    assign layer3_out[6412] = layer2_out[7417];
    assign layer3_out[6413] = layer2_out[6117] & ~layer2_out[6118];
    assign layer3_out[6414] = ~(layer2_out[1549] ^ layer2_out[1550]);
    assign layer3_out[6415] = ~layer2_out[6599];
    assign layer3_out[6416] = layer2_out[262];
    assign layer3_out[6417] = ~(layer2_out[6740] | layer2_out[6741]);
    assign layer3_out[6418] = layer2_out[6664];
    assign layer3_out[6419] = layer2_out[7329] & ~layer2_out[7328];
    assign layer3_out[6420] = ~(layer2_out[6708] ^ layer2_out[6709]);
    assign layer3_out[6421] = ~layer2_out[1662];
    assign layer3_out[6422] = ~(layer2_out[4047] & layer2_out[4048]);
    assign layer3_out[6423] = ~layer2_out[200];
    assign layer3_out[6424] = layer2_out[2491];
    assign layer3_out[6425] = layer2_out[4927] & layer2_out[4928];
    assign layer3_out[6426] = ~(layer2_out[5358] & layer2_out[5359]);
    assign layer3_out[6427] = layer2_out[1860] & ~layer2_out[1861];
    assign layer3_out[6428] = layer2_out[5917] ^ layer2_out[5918];
    assign layer3_out[6429] = layer2_out[3783] & ~layer2_out[3782];
    assign layer3_out[6430] = layer2_out[6508] | layer2_out[6509];
    assign layer3_out[6431] = ~(layer2_out[2693] | layer2_out[2694]);
    assign layer3_out[6432] = ~(layer2_out[3216] | layer2_out[3217]);
    assign layer3_out[6433] = ~layer2_out[1848] | layer2_out[1847];
    assign layer3_out[6434] = layer2_out[6584] & layer2_out[6585];
    assign layer3_out[6435] = layer2_out[3914] & layer2_out[3915];
    assign layer3_out[6436] = layer2_out[4133];
    assign layer3_out[6437] = ~(layer2_out[4098] & layer2_out[4099]);
    assign layer3_out[6438] = layer2_out[2019] & ~layer2_out[2020];
    assign layer3_out[6439] = layer2_out[7019] & ~layer2_out[7018];
    assign layer3_out[6440] = layer2_out[2132] & ~layer2_out[2131];
    assign layer3_out[6441] = layer2_out[3610];
    assign layer3_out[6442] = layer2_out[4501] & layer2_out[4502];
    assign layer3_out[6443] = layer2_out[3898];
    assign layer3_out[6444] = layer2_out[4109];
    assign layer3_out[6445] = layer2_out[3845];
    assign layer3_out[6446] = ~layer2_out[7413] | layer2_out[7412];
    assign layer3_out[6447] = 1'b0;
    assign layer3_out[6448] = layer2_out[4709];
    assign layer3_out[6449] = layer2_out[7332] | layer2_out[7333];
    assign layer3_out[6450] = 1'b1;
    assign layer3_out[6451] = layer2_out[3775] | layer2_out[3776];
    assign layer3_out[6452] = layer2_out[716] & ~layer2_out[715];
    assign layer3_out[6453] = ~layer2_out[5495];
    assign layer3_out[6454] = layer2_out[1655];
    assign layer3_out[6455] = layer2_out[3345] & ~layer2_out[3344];
    assign layer3_out[6456] = layer2_out[1288];
    assign layer3_out[6457] = layer2_out[3179] | layer2_out[3180];
    assign layer3_out[6458] = layer2_out[1970] & layer2_out[1971];
    assign layer3_out[6459] = ~layer2_out[7424];
    assign layer3_out[6460] = ~layer2_out[1815];
    assign layer3_out[6461] = ~(layer2_out[5319] ^ layer2_out[5320]);
    assign layer3_out[6462] = ~layer2_out[6188];
    assign layer3_out[6463] = ~layer2_out[6388];
    assign layer3_out[6464] = layer2_out[2414];
    assign layer3_out[6465] = ~layer2_out[1695];
    assign layer3_out[6466] = ~layer2_out[1134];
    assign layer3_out[6467] = ~(layer2_out[7606] & layer2_out[7607]);
    assign layer3_out[6468] = ~(layer2_out[6667] | layer2_out[6668]);
    assign layer3_out[6469] = ~layer2_out[34] | layer2_out[33];
    assign layer3_out[6470] = 1'b0;
    assign layer3_out[6471] = ~(layer2_out[6129] & layer2_out[6130]);
    assign layer3_out[6472] = 1'b0;
    assign layer3_out[6473] = layer2_out[5439] & layer2_out[5440];
    assign layer3_out[6474] = layer2_out[2020] | layer2_out[2021];
    assign layer3_out[6475] = ~layer2_out[718];
    assign layer3_out[6476] = ~(layer2_out[4887] & layer2_out[4888]);
    assign layer3_out[6477] = ~(layer2_out[7087] & layer2_out[7088]);
    assign layer3_out[6478] = ~layer2_out[647];
    assign layer3_out[6479] = ~layer2_out[7545];
    assign layer3_out[6480] = ~layer2_out[3973];
    assign layer3_out[6481] = layer2_out[7501] & layer2_out[7502];
    assign layer3_out[6482] = ~layer2_out[475];
    assign layer3_out[6483] = layer2_out[4403] | layer2_out[4404];
    assign layer3_out[6484] = layer2_out[7170];
    assign layer3_out[6485] = ~layer2_out[2944];
    assign layer3_out[6486] = ~layer2_out[7262] | layer2_out[7263];
    assign layer3_out[6487] = layer2_out[1263];
    assign layer3_out[6488] = 1'b0;
    assign layer3_out[6489] = ~layer2_out[3864];
    assign layer3_out[6490] = layer2_out[4644] & ~layer2_out[4643];
    assign layer3_out[6491] = layer2_out[6608];
    assign layer3_out[6492] = layer2_out[4072] & layer2_out[4073];
    assign layer3_out[6493] = layer2_out[7364] & layer2_out[7365];
    assign layer3_out[6494] = ~layer2_out[1435];
    assign layer3_out[6495] = layer2_out[2866] | layer2_out[2867];
    assign layer3_out[6496] = layer2_out[1901] ^ layer2_out[1902];
    assign layer3_out[6497] = ~layer2_out[4464] | layer2_out[4463];
    assign layer3_out[6498] = layer2_out[3735] & ~layer2_out[3734];
    assign layer3_out[6499] = ~layer2_out[7183] | layer2_out[7182];
    assign layer3_out[6500] = ~layer2_out[3665] | layer2_out[3664];
    assign layer3_out[6501] = layer2_out[2396];
    assign layer3_out[6502] = layer2_out[6394] ^ layer2_out[6395];
    assign layer3_out[6503] = ~layer2_out[756];
    assign layer3_out[6504] = ~layer2_out[2284] | layer2_out[2285];
    assign layer3_out[6505] = layer2_out[4583] & ~layer2_out[4584];
    assign layer3_out[6506] = ~layer2_out[1907];
    assign layer3_out[6507] = layer2_out[5955] & layer2_out[5956];
    assign layer3_out[6508] = ~layer2_out[998] | layer2_out[999];
    assign layer3_out[6509] = layer2_out[1544];
    assign layer3_out[6510] = ~layer2_out[7262];
    assign layer3_out[6511] = layer2_out[7540] | layer2_out[7541];
    assign layer3_out[6512] = layer2_out[674] | layer2_out[675];
    assign layer3_out[6513] = ~layer2_out[2767];
    assign layer3_out[6514] = layer2_out[7078] & layer2_out[7079];
    assign layer3_out[6515] = layer2_out[347];
    assign layer3_out[6516] = ~layer2_out[936] | layer2_out[937];
    assign layer3_out[6517] = ~layer2_out[7100] | layer2_out[7101];
    assign layer3_out[6518] = ~layer2_out[3860];
    assign layer3_out[6519] = layer2_out[2901] & ~layer2_out[2900];
    assign layer3_out[6520] = layer2_out[2796];
    assign layer3_out[6521] = ~layer2_out[2085];
    assign layer3_out[6522] = ~layer2_out[4783] | layer2_out[4784];
    assign layer3_out[6523] = layer2_out[6284] & ~layer2_out[6285];
    assign layer3_out[6524] = layer2_out[753] ^ layer2_out[754];
    assign layer3_out[6525] = layer2_out[4653] ^ layer2_out[4654];
    assign layer3_out[6526] = layer2_out[769] & ~layer2_out[770];
    assign layer3_out[6527] = layer2_out[864] & layer2_out[865];
    assign layer3_out[6528] = ~layer2_out[100];
    assign layer3_out[6529] = layer2_out[6756] & layer2_out[6757];
    assign layer3_out[6530] = layer2_out[3637];
    assign layer3_out[6531] = ~layer2_out[7646];
    assign layer3_out[6532] = layer2_out[1019];
    assign layer3_out[6533] = layer2_out[3498];
    assign layer3_out[6534] = ~(layer2_out[5549] | layer2_out[5550]);
    assign layer3_out[6535] = layer2_out[1420];
    assign layer3_out[6536] = ~layer2_out[4391];
    assign layer3_out[6537] = ~layer2_out[1745] | layer2_out[1746];
    assign layer3_out[6538] = ~(layer2_out[6634] & layer2_out[6635]);
    assign layer3_out[6539] = layer2_out[2424] & ~layer2_out[2423];
    assign layer3_out[6540] = layer2_out[338] & layer2_out[339];
    assign layer3_out[6541] = ~layer2_out[2447] | layer2_out[2448];
    assign layer3_out[6542] = ~(layer2_out[7688] | layer2_out[7689]);
    assign layer3_out[6543] = ~layer2_out[1359] | layer2_out[1358];
    assign layer3_out[6544] = ~layer2_out[667] | layer2_out[666];
    assign layer3_out[6545] = ~(layer2_out[2210] ^ layer2_out[2211]);
    assign layer3_out[6546] = ~(layer2_out[3382] ^ layer2_out[3383]);
    assign layer3_out[6547] = layer2_out[7514] ^ layer2_out[7515];
    assign layer3_out[6548] = layer2_out[7498] & layer2_out[7499];
    assign layer3_out[6549] = 1'b1;
    assign layer3_out[6550] = ~layer2_out[1138];
    assign layer3_out[6551] = layer2_out[6151] | layer2_out[6152];
    assign layer3_out[6552] = ~layer2_out[418] | layer2_out[419];
    assign layer3_out[6553] = ~(layer2_out[7689] ^ layer2_out[7690]);
    assign layer3_out[6554] = ~layer2_out[4014];
    assign layer3_out[6555] = ~(layer2_out[1930] ^ layer2_out[1931]);
    assign layer3_out[6556] = ~layer2_out[4540] | layer2_out[4541];
    assign layer3_out[6557] = ~layer2_out[5991];
    assign layer3_out[6558] = layer2_out[970] & ~layer2_out[971];
    assign layer3_out[6559] = ~(layer2_out[1320] & layer2_out[1321]);
    assign layer3_out[6560] = ~layer2_out[7751] | layer2_out[7750];
    assign layer3_out[6561] = ~layer2_out[6056];
    assign layer3_out[6562] = ~layer2_out[2394];
    assign layer3_out[6563] = layer2_out[3692] & ~layer2_out[3693];
    assign layer3_out[6564] = ~layer2_out[394];
    assign layer3_out[6565] = layer2_out[5341] ^ layer2_out[5342];
    assign layer3_out[6566] = ~(layer2_out[5345] | layer2_out[5346]);
    assign layer3_out[6567] = layer2_out[1802] & layer2_out[1803];
    assign layer3_out[6568] = ~(layer2_out[6851] | layer2_out[6852]);
    assign layer3_out[6569] = layer2_out[1988] | layer2_out[1989];
    assign layer3_out[6570] = ~layer2_out[2565];
    assign layer3_out[6571] = ~layer2_out[424] | layer2_out[425];
    assign layer3_out[6572] = layer2_out[103];
    assign layer3_out[6573] = layer2_out[105];
    assign layer3_out[6574] = layer2_out[7035] | layer2_out[7036];
    assign layer3_out[6575] = ~layer2_out[164];
    assign layer3_out[6576] = ~layer2_out[318];
    assign layer3_out[6577] = layer2_out[4177];
    assign layer3_out[6578] = ~(layer2_out[850] ^ layer2_out[851]);
    assign layer3_out[6579] = layer2_out[5160] | layer2_out[5161];
    assign layer3_out[6580] = 1'b0;
    assign layer3_out[6581] = layer2_out[5768];
    assign layer3_out[6582] = ~layer2_out[4119] | layer2_out[4118];
    assign layer3_out[6583] = ~(layer2_out[4617] ^ layer2_out[4618]);
    assign layer3_out[6584] = ~layer2_out[4996] | layer2_out[4995];
    assign layer3_out[6585] = layer2_out[3714];
    assign layer3_out[6586] = ~(layer2_out[7793] | layer2_out[7794]);
    assign layer3_out[6587] = layer2_out[3336] & ~layer2_out[3335];
    assign layer3_out[6588] = ~layer2_out[3195];
    assign layer3_out[6589] = ~layer2_out[2084] | layer2_out[2085];
    assign layer3_out[6590] = ~layer2_out[1856] | layer2_out[1857];
    assign layer3_out[6591] = ~layer2_out[1895] | layer2_out[1896];
    assign layer3_out[6592] = layer2_out[6695];
    assign layer3_out[6593] = layer2_out[6153] & layer2_out[6154];
    assign layer3_out[6594] = layer2_out[2792] ^ layer2_out[2793];
    assign layer3_out[6595] = ~layer2_out[3334];
    assign layer3_out[6596] = ~(layer2_out[3125] & layer2_out[3126]);
    assign layer3_out[6597] = layer2_out[2529] & layer2_out[2530];
    assign layer3_out[6598] = ~layer2_out[2595];
    assign layer3_out[6599] = ~layer2_out[4469];
    assign layer3_out[6600] = layer2_out[6130] & ~layer2_out[6131];
    assign layer3_out[6601] = ~layer2_out[7792];
    assign layer3_out[6602] = ~layer2_out[7714];
    assign layer3_out[6603] = ~layer2_out[5560] | layer2_out[5561];
    assign layer3_out[6604] = layer2_out[5260] | layer2_out[5261];
    assign layer3_out[6605] = layer2_out[4272];
    assign layer3_out[6606] = ~(layer2_out[5635] & layer2_out[5636]);
    assign layer3_out[6607] = layer2_out[3727] & ~layer2_out[3726];
    assign layer3_out[6608] = layer2_out[1190] & layer2_out[1191];
    assign layer3_out[6609] = ~layer2_out[5892] | layer2_out[5891];
    assign layer3_out[6610] = layer2_out[7004];
    assign layer3_out[6611] = layer2_out[4376];
    assign layer3_out[6612] = ~layer2_out[2782];
    assign layer3_out[6613] = layer2_out[351] | layer2_out[352];
    assign layer3_out[6614] = ~(layer2_out[6737] ^ layer2_out[6738]);
    assign layer3_out[6615] = ~layer2_out[996] | layer2_out[997];
    assign layer3_out[6616] = ~(layer2_out[731] & layer2_out[732]);
    assign layer3_out[6617] = layer2_out[3181] & layer2_out[3182];
    assign layer3_out[6618] = ~layer2_out[7163];
    assign layer3_out[6619] = layer2_out[6363] & ~layer2_out[6362];
    assign layer3_out[6620] = ~layer2_out[4419];
    assign layer3_out[6621] = ~(layer2_out[2873] ^ layer2_out[2874]);
    assign layer3_out[6622] = ~layer2_out[4949];
    assign layer3_out[6623] = layer2_out[6146] & layer2_out[6147];
    assign layer3_out[6624] = ~(layer2_out[7129] & layer2_out[7130]);
    assign layer3_out[6625] = ~layer2_out[1067];
    assign layer3_out[6626] = ~layer2_out[5249];
    assign layer3_out[6627] = layer2_out[7510] | layer2_out[7511];
    assign layer3_out[6628] = ~layer2_out[7005];
    assign layer3_out[6629] = ~(layer2_out[3641] & layer2_out[3642]);
    assign layer3_out[6630] = layer2_out[6414];
    assign layer3_out[6631] = ~layer2_out[752];
    assign layer3_out[6632] = ~layer2_out[5999];
    assign layer3_out[6633] = layer2_out[2880] & ~layer2_out[2881];
    assign layer3_out[6634] = layer2_out[7315] & ~layer2_out[7316];
    assign layer3_out[6635] = ~layer2_out[4323];
    assign layer3_out[6636] = ~(layer2_out[1203] | layer2_out[1204]);
    assign layer3_out[6637] = ~layer2_out[3295] | layer2_out[3296];
    assign layer3_out[6638] = layer2_out[7480];
    assign layer3_out[6639] = layer2_out[4669] & layer2_out[4670];
    assign layer3_out[6640] = layer2_out[4922] & ~layer2_out[4921];
    assign layer3_out[6641] = layer2_out[4442] & ~layer2_out[4443];
    assign layer3_out[6642] = ~layer2_out[1242];
    assign layer3_out[6643] = layer2_out[2333];
    assign layer3_out[6644] = ~layer2_out[1537] | layer2_out[1536];
    assign layer3_out[6645] = layer2_out[3487] | layer2_out[3488];
    assign layer3_out[6646] = layer2_out[2490] | layer2_out[2491];
    assign layer3_out[6647] = layer2_out[5613];
    assign layer3_out[6648] = ~layer2_out[3684];
    assign layer3_out[6649] = ~(layer2_out[4386] & layer2_out[4387]);
    assign layer3_out[6650] = layer2_out[5837] | layer2_out[5838];
    assign layer3_out[6651] = layer2_out[3840];
    assign layer3_out[6652] = layer2_out[6807] & ~layer2_out[6808];
    assign layer3_out[6653] = ~layer2_out[2557] | layer2_out[2556];
    assign layer3_out[6654] = layer2_out[7108];
    assign layer3_out[6655] = layer2_out[792];
    assign layer3_out[6656] = ~layer2_out[2444] | layer2_out[2443];
    assign layer3_out[6657] = layer2_out[3232];
    assign layer3_out[6658] = ~(layer2_out[5450] & layer2_out[5451]);
    assign layer3_out[6659] = layer2_out[4029];
    assign layer3_out[6660] = ~layer2_out[4574] | layer2_out[4573];
    assign layer3_out[6661] = ~layer2_out[6906];
    assign layer3_out[6662] = ~layer2_out[7071] | layer2_out[7072];
    assign layer3_out[6663] = layer2_out[2187];
    assign layer3_out[6664] = layer2_out[6098] & ~layer2_out[6099];
    assign layer3_out[6665] = layer2_out[2002] & ~layer2_out[2001];
    assign layer3_out[6666] = layer2_out[5036];
    assign layer3_out[6667] = ~layer2_out[7483] | layer2_out[7484];
    assign layer3_out[6668] = layer2_out[6890];
    assign layer3_out[6669] = ~layer2_out[3785];
    assign layer3_out[6670] = ~layer2_out[1926];
    assign layer3_out[6671] = layer2_out[687] | layer2_out[688];
    assign layer3_out[6672] = layer2_out[3420] | layer2_out[3421];
    assign layer3_out[6673] = layer2_out[5365];
    assign layer3_out[6674] = ~(layer2_out[2624] | layer2_out[2625]);
    assign layer3_out[6675] = ~(layer2_out[2380] | layer2_out[2381]);
    assign layer3_out[6676] = layer2_out[2635] & layer2_out[2636];
    assign layer3_out[6677] = layer2_out[663] & ~layer2_out[664];
    assign layer3_out[6678] = ~layer2_out[3796] | layer2_out[3795];
    assign layer3_out[6679] = ~layer2_out[6564];
    assign layer3_out[6680] = ~layer2_out[5088];
    assign layer3_out[6681] = layer2_out[4083] & layer2_out[4084];
    assign layer3_out[6682] = ~layer2_out[3298];
    assign layer3_out[6683] = ~layer2_out[6594] | layer2_out[6595];
    assign layer3_out[6684] = layer2_out[892] & layer2_out[893];
    assign layer3_out[6685] = ~layer2_out[3269] | layer2_out[3270];
    assign layer3_out[6686] = 1'b0;
    assign layer3_out[6687] = ~layer2_out[2554];
    assign layer3_out[6688] = layer2_out[5116] | layer2_out[5117];
    assign layer3_out[6689] = ~layer2_out[4393];
    assign layer3_out[6690] = ~(layer2_out[5176] & layer2_out[5177]);
    assign layer3_out[6691] = layer2_out[525];
    assign layer3_out[6692] = ~layer2_out[5956];
    assign layer3_out[6693] = ~layer2_out[7240] | layer2_out[7239];
    assign layer3_out[6694] = ~layer2_out[7502];
    assign layer3_out[6695] = ~layer2_out[7904] | layer2_out[7905];
    assign layer3_out[6696] = ~layer2_out[411] | layer2_out[410];
    assign layer3_out[6697] = layer2_out[1735];
    assign layer3_out[6698] = ~(layer2_out[4094] | layer2_out[4095]);
    assign layer3_out[6699] = layer2_out[1212] ^ layer2_out[1213];
    assign layer3_out[6700] = ~layer2_out[7468] | layer2_out[7467];
    assign layer3_out[6701] = layer2_out[5854];
    assign layer3_out[6702] = ~layer2_out[5275];
    assign layer3_out[6703] = layer2_out[5599];
    assign layer3_out[6704] = ~(layer2_out[2186] ^ layer2_out[2187]);
    assign layer3_out[6705] = layer2_out[7186];
    assign layer3_out[6706] = ~(layer2_out[924] ^ layer2_out[925]);
    assign layer3_out[6707] = layer2_out[5688];
    assign layer3_out[6708] = layer2_out[4707] & layer2_out[4708];
    assign layer3_out[6709] = layer2_out[3620];
    assign layer3_out[6710] = layer2_out[5669];
    assign layer3_out[6711] = layer2_out[3274];
    assign layer3_out[6712] = ~layer2_out[3517];
    assign layer3_out[6713] = layer2_out[306] ^ layer2_out[307];
    assign layer3_out[6714] = ~layer2_out[1531] | layer2_out[1530];
    assign layer3_out[6715] = layer2_out[3041] | layer2_out[3042];
    assign layer3_out[6716] = ~(layer2_out[6881] & layer2_out[6882]);
    assign layer3_out[6717] = ~layer2_out[7395] | layer2_out[7396];
    assign layer3_out[6718] = layer2_out[209] ^ layer2_out[210];
    assign layer3_out[6719] = ~layer2_out[1723] | layer2_out[1722];
    assign layer3_out[6720] = ~layer2_out[6304];
    assign layer3_out[6721] = ~layer2_out[7566];
    assign layer3_out[6722] = ~layer2_out[6695];
    assign layer3_out[6723] = ~layer2_out[7512];
    assign layer3_out[6724] = layer2_out[1466];
    assign layer3_out[6725] = ~layer2_out[1040];
    assign layer3_out[6726] = ~layer2_out[7942];
    assign layer3_out[6727] = layer2_out[1513] | layer2_out[1514];
    assign layer3_out[6728] = layer2_out[5081] ^ layer2_out[5082];
    assign layer3_out[6729] = layer2_out[4070] & layer2_out[4071];
    assign layer3_out[6730] = ~layer2_out[453] | layer2_out[452];
    assign layer3_out[6731] = ~layer2_out[4247];
    assign layer3_out[6732] = 1'b0;
    assign layer3_out[6733] = layer2_out[123];
    assign layer3_out[6734] = ~layer2_out[6716];
    assign layer3_out[6735] = ~(layer2_out[7976] & layer2_out[7977]);
    assign layer3_out[6736] = layer2_out[5593] ^ layer2_out[5594];
    assign layer3_out[6737] = layer2_out[5522];
    assign layer3_out[6738] = layer2_out[2929] ^ layer2_out[2930];
    assign layer3_out[6739] = layer2_out[3399] & layer2_out[3400];
    assign layer3_out[6740] = layer2_out[1562] ^ layer2_out[1563];
    assign layer3_out[6741] = layer2_out[2394] & layer2_out[2395];
    assign layer3_out[6742] = layer2_out[7543] & layer2_out[7544];
    assign layer3_out[6743] = layer2_out[5546] ^ layer2_out[5547];
    assign layer3_out[6744] = layer2_out[7215] & layer2_out[7216];
    assign layer3_out[6745] = layer2_out[1794] & ~layer2_out[1793];
    assign layer3_out[6746] = ~layer2_out[4422];
    assign layer3_out[6747] = layer2_out[4901] & layer2_out[4902];
    assign layer3_out[6748] = ~(layer2_out[1028] ^ layer2_out[1029]);
    assign layer3_out[6749] = 1'b1;
    assign layer3_out[6750] = ~layer2_out[3287];
    assign layer3_out[6751] = ~(layer2_out[175] | layer2_out[176]);
    assign layer3_out[6752] = ~layer2_out[6682];
    assign layer3_out[6753] = layer2_out[1722];
    assign layer3_out[6754] = ~layer2_out[6478];
    assign layer3_out[6755] = layer2_out[2645];
    assign layer3_out[6756] = ~layer2_out[4252];
    assign layer3_out[6757] = layer2_out[4479] & ~layer2_out[4480];
    assign layer3_out[6758] = ~layer2_out[4605];
    assign layer3_out[6759] = layer2_out[1422];
    assign layer3_out[6760] = ~layer2_out[4625];
    assign layer3_out[6761] = layer2_out[3856];
    assign layer3_out[6762] = ~layer2_out[7178];
    assign layer3_out[6763] = layer2_out[2054] & ~layer2_out[2055];
    assign layer3_out[6764] = 1'b1;
    assign layer3_out[6765] = ~layer2_out[1973];
    assign layer3_out[6766] = layer2_out[6572];
    assign layer3_out[6767] = ~(layer2_out[2249] ^ layer2_out[2250]);
    assign layer3_out[6768] = 1'b1;
    assign layer3_out[6769] = layer2_out[3003] | layer2_out[3004];
    assign layer3_out[6770] = ~(layer2_out[6810] & layer2_out[6811]);
    assign layer3_out[6771] = layer2_out[7857] & ~layer2_out[7858];
    assign layer3_out[6772] = ~layer2_out[5413];
    assign layer3_out[6773] = ~layer2_out[2749];
    assign layer3_out[6774] = ~(layer2_out[6903] & layer2_out[6904]);
    assign layer3_out[6775] = layer2_out[1712] & ~layer2_out[1711];
    assign layer3_out[6776] = layer2_out[5958] & ~layer2_out[5959];
    assign layer3_out[6777] = ~layer2_out[6666] | layer2_out[6667];
    assign layer3_out[6778] = layer2_out[27] ^ layer2_out[28];
    assign layer3_out[6779] = ~layer2_out[6396];
    assign layer3_out[6780] = ~layer2_out[6596] | layer2_out[6597];
    assign layer3_out[6781] = layer2_out[7415] & layer2_out[7416];
    assign layer3_out[6782] = ~layer2_out[703];
    assign layer3_out[6783] = layer2_out[6719] ^ layer2_out[6720];
    assign layer3_out[6784] = 1'b1;
    assign layer3_out[6785] = ~layer2_out[7055];
    assign layer3_out[6786] = layer2_out[4351] & ~layer2_out[4350];
    assign layer3_out[6787] = layer2_out[3986];
    assign layer3_out[6788] = layer2_out[916] | layer2_out[917];
    assign layer3_out[6789] = ~layer2_out[4569];
    assign layer3_out[6790] = layer2_out[1923] & ~layer2_out[1922];
    assign layer3_out[6791] = layer2_out[4060] | layer2_out[4061];
    assign layer3_out[6792] = layer2_out[873] | layer2_out[874];
    assign layer3_out[6793] = layer2_out[1539] & ~layer2_out[1540];
    assign layer3_out[6794] = layer2_out[1000];
    assign layer3_out[6795] = layer2_out[4116];
    assign layer3_out[6796] = ~(layer2_out[3843] ^ layer2_out[3844]);
    assign layer3_out[6797] = layer2_out[6368];
    assign layer3_out[6798] = ~layer2_out[7931];
    assign layer3_out[6799] = layer2_out[3611];
    assign layer3_out[6800] = layer2_out[1934] & ~layer2_out[1933];
    assign layer3_out[6801] = layer2_out[2669];
    assign layer3_out[6802] = layer2_out[7198];
    assign layer3_out[6803] = ~layer2_out[909] | layer2_out[908];
    assign layer3_out[6804] = ~(layer2_out[4763] | layer2_out[4764]);
    assign layer3_out[6805] = ~layer2_out[7106];
    assign layer3_out[6806] = ~layer2_out[4051];
    assign layer3_out[6807] = ~layer2_out[6933];
    assign layer3_out[6808] = layer2_out[6162];
    assign layer3_out[6809] = ~layer2_out[6743] | layer2_out[6744];
    assign layer3_out[6810] = layer2_out[1391];
    assign layer3_out[6811] = ~layer2_out[2183];
    assign layer3_out[6812] = layer2_out[1393] | layer2_out[1394];
    assign layer3_out[6813] = ~layer2_out[7679] | layer2_out[7680];
    assign layer3_out[6814] = layer2_out[1386] & ~layer2_out[1385];
    assign layer3_out[6815] = 1'b0;
    assign layer3_out[6816] = ~(layer2_out[2686] | layer2_out[2687]);
    assign layer3_out[6817] = layer2_out[6457];
    assign layer3_out[6818] = layer2_out[1444] & ~layer2_out[1445];
    assign layer3_out[6819] = ~layer2_out[62] | layer2_out[63];
    assign layer3_out[6820] = ~(layer2_out[2286] | layer2_out[2287]);
    assign layer3_out[6821] = layer2_out[7839];
    assign layer3_out[6822] = ~layer2_out[4327];
    assign layer3_out[6823] = ~(layer2_out[4947] ^ layer2_out[4948]);
    assign layer3_out[6824] = ~(layer2_out[7917] | layer2_out[7918]);
    assign layer3_out[6825] = ~layer2_out[6975] | layer2_out[6976];
    assign layer3_out[6826] = ~layer2_out[5271];
    assign layer3_out[6827] = ~(layer2_out[7858] ^ layer2_out[7859]);
    assign layer3_out[6828] = ~layer2_out[3585];
    assign layer3_out[6829] = ~(layer2_out[7024] ^ layer2_out[7025]);
    assign layer3_out[6830] = 1'b1;
    assign layer3_out[6831] = layer2_out[3316];
    assign layer3_out[6832] = ~(layer2_out[2707] ^ layer2_out[2708]);
    assign layer3_out[6833] = layer2_out[7523] ^ layer2_out[7524];
    assign layer3_out[6834] = ~layer2_out[5776] | layer2_out[5775];
    assign layer3_out[6835] = ~layer2_out[5548] | layer2_out[5549];
    assign layer3_out[6836] = ~layer2_out[671];
    assign layer3_out[6837] = layer2_out[2356];
    assign layer3_out[6838] = ~layer2_out[376];
    assign layer3_out[6839] = layer2_out[1782] & ~layer2_out[1781];
    assign layer3_out[6840] = layer2_out[6794] & ~layer2_out[6793];
    assign layer3_out[6841] = ~layer2_out[6314];
    assign layer3_out[6842] = layer2_out[3633] & ~layer2_out[3634];
    assign layer3_out[6843] = layer2_out[5465];
    assign layer3_out[6844] = layer2_out[6264];
    assign layer3_out[6845] = ~layer2_out[4712];
    assign layer3_out[6846] = ~layer2_out[4409] | layer2_out[4410];
    assign layer3_out[6847] = ~(layer2_out[7855] ^ layer2_out[7856]);
    assign layer3_out[6848] = ~layer2_out[4711] | layer2_out[4712];
    assign layer3_out[6849] = layer2_out[7015] | layer2_out[7016];
    assign layer3_out[6850] = layer2_out[7963] & ~layer2_out[7962];
    assign layer3_out[6851] = layer2_out[2650];
    assign layer3_out[6852] = ~(layer2_out[6192] | layer2_out[6193]);
    assign layer3_out[6853] = ~layer2_out[5731];
    assign layer3_out[6854] = ~(layer2_out[1947] & layer2_out[1948]);
    assign layer3_out[6855] = layer2_out[3047] & ~layer2_out[3048];
    assign layer3_out[6856] = ~(layer2_out[4284] ^ layer2_out[4285]);
    assign layer3_out[6857] = layer2_out[5522] & ~layer2_out[5521];
    assign layer3_out[6858] = ~layer2_out[107];
    assign layer3_out[6859] = ~layer2_out[2943];
    assign layer3_out[6860] = layer2_out[3256] & ~layer2_out[3257];
    assign layer3_out[6861] = ~layer2_out[2615] | layer2_out[2614];
    assign layer3_out[6862] = ~layer2_out[1296] | layer2_out[1295];
    assign layer3_out[6863] = layer2_out[4512];
    assign layer3_out[6864] = ~(layer2_out[1634] & layer2_out[1635]);
    assign layer3_out[6865] = layer2_out[1057];
    assign layer3_out[6866] = ~layer2_out[5836] | layer2_out[5835];
    assign layer3_out[6867] = layer2_out[7424];
    assign layer3_out[6868] = layer2_out[5619];
    assign layer3_out[6869] = layer2_out[6566];
    assign layer3_out[6870] = layer2_out[5914];
    assign layer3_out[6871] = layer2_out[7718];
    assign layer3_out[6872] = ~layer2_out[7936];
    assign layer3_out[6873] = layer2_out[3761];
    assign layer3_out[6874] = layer2_out[480] ^ layer2_out[481];
    assign layer3_out[6875] = ~(layer2_out[7267] ^ layer2_out[7268]);
    assign layer3_out[6876] = layer2_out[2213] | layer2_out[2214];
    assign layer3_out[6877] = ~(layer2_out[6305] ^ layer2_out[6306]);
    assign layer3_out[6878] = layer2_out[4137];
    assign layer3_out[6879] = layer2_out[5157];
    assign layer3_out[6880] = ~(layer2_out[5714] ^ layer2_out[5715]);
    assign layer3_out[6881] = layer2_out[4453] ^ layer2_out[4454];
    assign layer3_out[6882] = layer2_out[5621] & ~layer2_out[5620];
    assign layer3_out[6883] = ~(layer2_out[6390] & layer2_out[6391]);
    assign layer3_out[6884] = ~(layer2_out[7834] ^ layer2_out[7835]);
    assign layer3_out[6885] = ~layer2_out[7842] | layer2_out[7841];
    assign layer3_out[6886] = ~(layer2_out[7797] & layer2_out[7798]);
    assign layer3_out[6887] = ~layer2_out[5774] | layer2_out[5775];
    assign layer3_out[6888] = ~layer2_out[5721] | layer2_out[5722];
    assign layer3_out[6889] = layer2_out[2063] & ~layer2_out[2062];
    assign layer3_out[6890] = ~(layer2_out[2859] & layer2_out[2860]);
    assign layer3_out[6891] = ~layer2_out[1642];
    assign layer3_out[6892] = layer2_out[1315];
    assign layer3_out[6893] = ~layer2_out[4811];
    assign layer3_out[6894] = layer2_out[1923] | layer2_out[1924];
    assign layer3_out[6895] = layer2_out[2796] & ~layer2_out[2797];
    assign layer3_out[6896] = layer2_out[3420];
    assign layer3_out[6897] = layer2_out[2742] | layer2_out[2743];
    assign layer3_out[6898] = layer2_out[6581] & ~layer2_out[6580];
    assign layer3_out[6899] = ~(layer2_out[6904] & layer2_out[6905]);
    assign layer3_out[6900] = layer2_out[4028];
    assign layer3_out[6901] = ~layer2_out[4205] | layer2_out[4206];
    assign layer3_out[6902] = ~layer2_out[2220];
    assign layer3_out[6903] = layer2_out[7160] | layer2_out[7161];
    assign layer3_out[6904] = ~layer2_out[5445];
    assign layer3_out[6905] = ~(layer2_out[558] & layer2_out[559]);
    assign layer3_out[6906] = layer2_out[4408] & ~layer2_out[4407];
    assign layer3_out[6907] = ~layer2_out[6490] | layer2_out[6491];
    assign layer3_out[6908] = 1'b0;
    assign layer3_out[6909] = ~layer2_out[5943] | layer2_out[5942];
    assign layer3_out[6910] = layer2_out[5230] & ~layer2_out[5229];
    assign layer3_out[6911] = layer2_out[3049];
    assign layer3_out[6912] = layer2_out[5267] & ~layer2_out[5268];
    assign layer3_out[6913] = ~layer2_out[5862] | layer2_out[5861];
    assign layer3_out[6914] = ~(layer2_out[2658] & layer2_out[2659]);
    assign layer3_out[6915] = layer2_out[2506];
    assign layer3_out[6916] = ~layer2_out[1107];
    assign layer3_out[6917] = ~layer2_out[7614] | layer2_out[7615];
    assign layer3_out[6918] = ~layer2_out[5806];
    assign layer3_out[6919] = ~layer2_out[7506];
    assign layer3_out[6920] = layer2_out[3849];
    assign layer3_out[6921] = layer2_out[1127] & layer2_out[1128];
    assign layer3_out[6922] = layer2_out[2130];
    assign layer3_out[6923] = layer2_out[7604] ^ layer2_out[7605];
    assign layer3_out[6924] = layer2_out[732] | layer2_out[733];
    assign layer3_out[6925] = layer2_out[915];
    assign layer3_out[6926] = ~layer2_out[5231];
    assign layer3_out[6927] = layer2_out[7294] & ~layer2_out[7295];
    assign layer3_out[6928] = layer2_out[7618] & ~layer2_out[7617];
    assign layer3_out[6929] = ~layer2_out[5233] | layer2_out[5232];
    assign layer3_out[6930] = ~layer2_out[1542] | layer2_out[1543];
    assign layer3_out[6931] = 1'b0;
    assign layer3_out[6932] = ~(layer2_out[7953] | layer2_out[7954]);
    assign layer3_out[6933] = ~(layer2_out[7860] | layer2_out[7861]);
    assign layer3_out[6934] = layer2_out[6752] & layer2_out[6753];
    assign layer3_out[6935] = ~layer2_out[2153];
    assign layer3_out[6936] = ~layer2_out[1893] | layer2_out[1894];
    assign layer3_out[6937] = ~layer2_out[7582] | layer2_out[7581];
    assign layer3_out[6938] = ~layer2_out[6325];
    assign layer3_out[6939] = ~(layer2_out[7274] & layer2_out[7275]);
    assign layer3_out[6940] = ~layer2_out[4241];
    assign layer3_out[6941] = layer2_out[3476];
    assign layer3_out[6942] = layer2_out[2525];
    assign layer3_out[6943] = layer2_out[5805];
    assign layer3_out[6944] = ~layer2_out[5045];
    assign layer3_out[6945] = ~(layer2_out[614] & layer2_out[615]);
    assign layer3_out[6946] = layer2_out[1730];
    assign layer3_out[6947] = ~layer2_out[3656] | layer2_out[3657];
    assign layer3_out[6948] = layer2_out[4958] & layer2_out[4959];
    assign layer3_out[6949] = ~layer2_out[5216];
    assign layer3_out[6950] = ~layer2_out[4973] | layer2_out[4972];
    assign layer3_out[6951] = layer2_out[7444] & ~layer2_out[7443];
    assign layer3_out[6952] = ~layer2_out[1014];
    assign layer3_out[6953] = ~(layer2_out[2203] ^ layer2_out[2204]);
    assign layer3_out[6954] = layer2_out[5384];
    assign layer3_out[6955] = ~(layer2_out[7511] ^ layer2_out[7512]);
    assign layer3_out[6956] = ~layer2_out[6768];
    assign layer3_out[6957] = ~layer2_out[5342] | layer2_out[5343];
    assign layer3_out[6958] = layer2_out[4981] ^ layer2_out[4982];
    assign layer3_out[6959] = ~(layer2_out[3214] ^ layer2_out[3215]);
    assign layer3_out[6960] = layer2_out[5555];
    assign layer3_out[6961] = layer2_out[7445] & ~layer2_out[7446];
    assign layer3_out[6962] = ~(layer2_out[1285] | layer2_out[1286]);
    assign layer3_out[6963] = layer2_out[1330] & ~layer2_out[1329];
    assign layer3_out[6964] = ~(layer2_out[7981] ^ layer2_out[7982]);
    assign layer3_out[6965] = 1'b0;
    assign layer3_out[6966] = ~layer2_out[7861];
    assign layer3_out[6967] = layer2_out[6104] & ~layer2_out[6105];
    assign layer3_out[6968] = ~(layer2_out[3953] | layer2_out[3954]);
    assign layer3_out[6969] = layer2_out[2029];
    assign layer3_out[6970] = layer2_out[7845];
    assign layer3_out[6971] = layer2_out[5887];
    assign layer3_out[6972] = layer2_out[4985] & layer2_out[4986];
    assign layer3_out[6973] = layer2_out[7828] | layer2_out[7829];
    assign layer3_out[6974] = ~layer2_out[3820];
    assign layer3_out[6975] = ~(layer2_out[1278] & layer2_out[1279]);
    assign layer3_out[6976] = ~layer2_out[6736];
    assign layer3_out[6977] = layer2_out[430] & layer2_out[431];
    assign layer3_out[6978] = ~layer2_out[6645];
    assign layer3_out[6979] = ~layer2_out[6236];
    assign layer3_out[6980] = ~layer2_out[4550];
    assign layer3_out[6981] = ~layer2_out[2073] | layer2_out[2072];
    assign layer3_out[6982] = layer2_out[2381] ^ layer2_out[2382];
    assign layer3_out[6983] = layer2_out[1148] ^ layer2_out[1149];
    assign layer3_out[6984] = ~layer2_out[7362];
    assign layer3_out[6985] = layer2_out[5954];
    assign layer3_out[6986] = layer2_out[1964];
    assign layer3_out[6987] = layer2_out[7666];
    assign layer3_out[6988] = ~layer2_out[1235];
    assign layer3_out[6989] = layer2_out[4677] & ~layer2_out[4678];
    assign layer3_out[6990] = ~layer2_out[653] | layer2_out[654];
    assign layer3_out[6991] = ~layer2_out[1132] | layer2_out[1131];
    assign layer3_out[6992] = ~(layer2_out[6073] | layer2_out[6074]);
    assign layer3_out[6993] = ~(layer2_out[6552] & layer2_out[6553]);
    assign layer3_out[6994] = ~layer2_out[7678];
    assign layer3_out[6995] = layer2_out[2052] & ~layer2_out[2053];
    assign layer3_out[6996] = layer2_out[1571];
    assign layer3_out[6997] = ~layer2_out[7822] | layer2_out[7823];
    assign layer3_out[6998] = ~layer2_out[904];
    assign layer3_out[6999] = ~layer2_out[6972] | layer2_out[6971];
    assign layer3_out[7000] = ~(layer2_out[2475] | layer2_out[2476]);
    assign layer3_out[7001] = ~(layer2_out[3398] & layer2_out[3399]);
    assign layer3_out[7002] = layer2_out[7388] ^ layer2_out[7389];
    assign layer3_out[7003] = ~(layer2_out[7217] | layer2_out[7218]);
    assign layer3_out[7004] = layer2_out[5763];
    assign layer3_out[7005] = ~layer2_out[2034];
    assign layer3_out[7006] = layer2_out[4448];
    assign layer3_out[7007] = ~layer2_out[6435] | layer2_out[6436];
    assign layer3_out[7008] = ~layer2_out[3519];
    assign layer3_out[7009] = ~(layer2_out[4379] ^ layer2_out[4380]);
    assign layer3_out[7010] = layer2_out[2907];
    assign layer3_out[7011] = ~(layer2_out[582] | layer2_out[583]);
    assign layer3_out[7012] = layer2_out[3510] & ~layer2_out[3509];
    assign layer3_out[7013] = layer2_out[3984] | layer2_out[3985];
    assign layer3_out[7014] = layer2_out[1522];
    assign layer3_out[7015] = layer2_out[1816] ^ layer2_out[1817];
    assign layer3_out[7016] = layer2_out[120] | layer2_out[121];
    assign layer3_out[7017] = ~layer2_out[6424] | layer2_out[6423];
    assign layer3_out[7018] = ~layer2_out[6781];
    assign layer3_out[7019] = layer2_out[4617] & ~layer2_out[4616];
    assign layer3_out[7020] = ~layer2_out[5964];
    assign layer3_out[7021] = ~(layer2_out[6818] ^ layer2_out[6819]);
    assign layer3_out[7022] = ~(layer2_out[6322] & layer2_out[6323]);
    assign layer3_out[7023] = layer2_out[1210];
    assign layer3_out[7024] = layer2_out[1632];
    assign layer3_out[7025] = ~(layer2_out[4833] | layer2_out[4834]);
    assign layer3_out[7026] = layer2_out[796] & layer2_out[797];
    assign layer3_out[7027] = layer2_out[6968];
    assign layer3_out[7028] = ~layer2_out[2245];
    assign layer3_out[7029] = ~layer2_out[6310];
    assign layer3_out[7030] = ~(layer2_out[3118] & layer2_out[3119]);
    assign layer3_out[7031] = layer2_out[1239] ^ layer2_out[1240];
    assign layer3_out[7032] = ~(layer2_out[6602] ^ layer2_out[6603]);
    assign layer3_out[7033] = layer2_out[2016] ^ layer2_out[2017];
    assign layer3_out[7034] = ~(layer2_out[5037] | layer2_out[5038]);
    assign layer3_out[7035] = ~layer2_out[1368];
    assign layer3_out[7036] = ~layer2_out[4671];
    assign layer3_out[7037] = ~layer2_out[3917];
    assign layer3_out[7038] = layer2_out[7527];
    assign layer3_out[7039] = layer2_out[4885] & layer2_out[4886];
    assign layer3_out[7040] = layer2_out[3970] ^ layer2_out[3971];
    assign layer3_out[7041] = layer2_out[163] & ~layer2_out[162];
    assign layer3_out[7042] = layer2_out[5780];
    assign layer3_out[7043] = ~layer2_out[7213];
    assign layer3_out[7044] = 1'b0;
    assign layer3_out[7045] = layer2_out[1042];
    assign layer3_out[7046] = 1'b1;
    assign layer3_out[7047] = layer2_out[3945] & ~layer2_out[3946];
    assign layer3_out[7048] = ~layer2_out[188] | layer2_out[189];
    assign layer3_out[7049] = ~(layer2_out[3659] & layer2_out[3660]);
    assign layer3_out[7050] = 1'b0;
    assign layer3_out[7051] = ~layer2_out[6247];
    assign layer3_out[7052] = ~layer2_out[252];
    assign layer3_out[7053] = ~layer2_out[7359];
    assign layer3_out[7054] = ~(layer2_out[6765] & layer2_out[6766]);
    assign layer3_out[7055] = ~(layer2_out[4439] | layer2_out[4440]);
    assign layer3_out[7056] = layer2_out[3005];
    assign layer3_out[7057] = ~layer2_out[6525] | layer2_out[6526];
    assign layer3_out[7058] = layer2_out[5953] & ~layer2_out[5952];
    assign layer3_out[7059] = ~(layer2_out[2745] & layer2_out[2746]);
    assign layer3_out[7060] = layer2_out[7018];
    assign layer3_out[7061] = ~layer2_out[5321] | layer2_out[5320];
    assign layer3_out[7062] = layer2_out[678];
    assign layer3_out[7063] = layer2_out[6251];
    assign layer3_out[7064] = ~layer2_out[4466] | layer2_out[4465];
    assign layer3_out[7065] = layer2_out[2787] & ~layer2_out[2786];
    assign layer3_out[7066] = ~layer2_out[2052];
    assign layer3_out[7067] = ~layer2_out[6936] | layer2_out[6937];
    assign layer3_out[7068] = ~(layer2_out[179] | layer2_out[180]);
    assign layer3_out[7069] = ~layer2_out[5612];
    assign layer3_out[7070] = ~layer2_out[6300] | layer2_out[6299];
    assign layer3_out[7071] = ~layer2_out[2680] | layer2_out[2679];
    assign layer3_out[7072] = 1'b0;
    assign layer3_out[7073] = layer2_out[6679] & layer2_out[6680];
    assign layer3_out[7074] = ~(layer2_out[6342] | layer2_out[6343]);
    assign layer3_out[7075] = ~(layer2_out[2988] | layer2_out[2989]);
    assign layer3_out[7076] = ~(layer2_out[4554] | layer2_out[4555]);
    assign layer3_out[7077] = layer2_out[5718];
    assign layer3_out[7078] = ~layer2_out[6296] | layer2_out[6297];
    assign layer3_out[7079] = ~layer2_out[6618] | layer2_out[6617];
    assign layer3_out[7080] = layer2_out[1938];
    assign layer3_out[7081] = ~layer2_out[2608];
    assign layer3_out[7082] = ~layer2_out[2497];
    assign layer3_out[7083] = layer2_out[4565];
    assign layer3_out[7084] = layer2_out[5900] ^ layer2_out[5901];
    assign layer3_out[7085] = layer2_out[26];
    assign layer3_out[7086] = layer2_out[5051] | layer2_out[5052];
    assign layer3_out[7087] = ~layer2_out[7420] | layer2_out[7419];
    assign layer3_out[7088] = ~layer2_out[620];
    assign layer3_out[7089] = ~layer2_out[287];
    assign layer3_out[7090] = layer2_out[4187] & ~layer2_out[4188];
    assign layer3_out[7091] = layer2_out[3932];
    assign layer3_out[7092] = layer2_out[47];
    assign layer3_out[7093] = ~(layer2_out[2921] & layer2_out[2922]);
    assign layer3_out[7094] = ~layer2_out[2928];
    assign layer3_out[7095] = ~layer2_out[7640];
    assign layer3_out[7096] = ~layer2_out[6953] | layer2_out[6952];
    assign layer3_out[7097] = ~(layer2_out[4674] ^ layer2_out[4675]);
    assign layer3_out[7098] = ~layer2_out[3832];
    assign layer3_out[7099] = ~layer2_out[6600] | layer2_out[6599];
    assign layer3_out[7100] = ~layer2_out[6038] | layer2_out[6039];
    assign layer3_out[7101] = layer2_out[4199] & layer2_out[4200];
    assign layer3_out[7102] = layer2_out[2261];
    assign layer3_out[7103] = layer2_out[6412] | layer2_out[6413];
    assign layer3_out[7104] = ~layer2_out[5176];
    assign layer3_out[7105] = layer2_out[1283];
    assign layer3_out[7106] = ~layer2_out[4725] | layer2_out[4724];
    assign layer3_out[7107] = layer2_out[2990];
    assign layer3_out[7108] = layer2_out[7197] & layer2_out[7198];
    assign layer3_out[7109] = layer2_out[4636] | layer2_out[4637];
    assign layer3_out[7110] = layer2_out[7193] | layer2_out[7194];
    assign layer3_out[7111] = ~layer2_out[310] | layer2_out[311];
    assign layer3_out[7112] = 1'b0;
    assign layer3_out[7113] = layer2_out[5734] & ~layer2_out[5733];
    assign layer3_out[7114] = ~layer2_out[2130];
    assign layer3_out[7115] = ~layer2_out[4425] | layer2_out[4424];
    assign layer3_out[7116] = ~layer2_out[6039];
    assign layer3_out[7117] = layer2_out[5239] & ~layer2_out[5238];
    assign layer3_out[7118] = ~(layer2_out[148] | layer2_out[149]);
    assign layer3_out[7119] = ~layer2_out[3051] | layer2_out[3052];
    assign layer3_out[7120] = ~layer2_out[566];
    assign layer3_out[7121] = ~(layer2_out[2631] & layer2_out[2632]);
    assign layer3_out[7122] = layer2_out[5724] & ~layer2_out[5725];
    assign layer3_out[7123] = layer2_out[3590] ^ layer2_out[3591];
    assign layer3_out[7124] = layer2_out[3310];
    assign layer3_out[7125] = layer2_out[720] & ~layer2_out[721];
    assign layer3_out[7126] = ~layer2_out[4038] | layer2_out[4037];
    assign layer3_out[7127] = layer2_out[5287] | layer2_out[5288];
    assign layer3_out[7128] = layer2_out[6522];
    assign layer3_out[7129] = layer2_out[2032] | layer2_out[2033];
    assign layer3_out[7130] = layer2_out[727] ^ layer2_out[728];
    assign layer3_out[7131] = 1'b1;
    assign layer3_out[7132] = layer2_out[1787] & ~layer2_out[1786];
    assign layer3_out[7133] = ~layer2_out[3060];
    assign layer3_out[7134] = ~layer2_out[320] | layer2_out[321];
    assign layer3_out[7135] = layer2_out[2068] | layer2_out[2069];
    assign layer3_out[7136] = layer2_out[3934];
    assign layer3_out[7137] = ~layer2_out[639] | layer2_out[638];
    assign layer3_out[7138] = layer2_out[3565];
    assign layer3_out[7139] = layer2_out[4312] | layer2_out[4313];
    assign layer3_out[7140] = layer2_out[4899] ^ layer2_out[4900];
    assign layer3_out[7141] = ~(layer2_out[4299] | layer2_out[4300]);
    assign layer3_out[7142] = ~layer2_out[4508];
    assign layer3_out[7143] = layer2_out[3445] & layer2_out[3446];
    assign layer3_out[7144] = layer2_out[338] & ~layer2_out[337];
    assign layer3_out[7145] = layer2_out[1169] ^ layer2_out[1170];
    assign layer3_out[7146] = layer2_out[168];
    assign layer3_out[7147] = layer2_out[6721] & ~layer2_out[6720];
    assign layer3_out[7148] = ~layer2_out[6248];
    assign layer3_out[7149] = ~(layer2_out[1844] & layer2_out[1845]);
    assign layer3_out[7150] = ~(layer2_out[1113] ^ layer2_out[1114]);
    assign layer3_out[7151] = layer2_out[5820] ^ layer2_out[5821];
    assign layer3_out[7152] = layer2_out[4342] ^ layer2_out[4343];
    assign layer3_out[7153] = layer2_out[313];
    assign layer3_out[7154] = layer2_out[5287] & ~layer2_out[5286];
    assign layer3_out[7155] = layer2_out[6928];
    assign layer3_out[7156] = layer2_out[3897];
    assign layer3_out[7157] = ~(layer2_out[236] ^ layer2_out[237]);
    assign layer3_out[7158] = ~layer2_out[6107] | layer2_out[6108];
    assign layer3_out[7159] = layer2_out[3448] ^ layer2_out[3449];
    assign layer3_out[7160] = layer2_out[6951];
    assign layer3_out[7161] = layer2_out[6240] ^ layer2_out[6241];
    assign layer3_out[7162] = ~layer2_out[6831] | layer2_out[6830];
    assign layer3_out[7163] = layer2_out[3958] | layer2_out[3959];
    assign layer3_out[7164] = layer2_out[743];
    assign layer3_out[7165] = layer2_out[3417] & layer2_out[3418];
    assign layer3_out[7166] = layer2_out[5333] & ~layer2_out[5334];
    assign layer3_out[7167] = ~(layer2_out[1780] & layer2_out[1781]);
    assign layer3_out[7168] = ~layer2_out[4991];
    assign layer3_out[7169] = ~layer2_out[7106] | layer2_out[7105];
    assign layer3_out[7170] = ~(layer2_out[296] ^ layer2_out[297]);
    assign layer3_out[7171] = layer2_out[1512] & layer2_out[1513];
    assign layer3_out[7172] = ~(layer2_out[3605] & layer2_out[3606]);
    assign layer3_out[7173] = ~layer2_out[3204];
    assign layer3_out[7174] = ~layer2_out[545] | layer2_out[546];
    assign layer3_out[7175] = ~layer2_out[6446];
    assign layer3_out[7176] = layer2_out[2544] & ~layer2_out[2543];
    assign layer3_out[7177] = layer2_out[3297] & ~layer2_out[3296];
    assign layer3_out[7178] = layer2_out[13];
    assign layer3_out[7179] = layer2_out[7570];
    assign layer3_out[7180] = ~(layer2_out[3794] | layer2_out[3795]);
    assign layer3_out[7181] = layer2_out[1626];
    assign layer3_out[7182] = ~layer2_out[6529];
    assign layer3_out[7183] = ~(layer2_out[4315] & layer2_out[4316]);
    assign layer3_out[7184] = ~layer2_out[3465];
    assign layer3_out[7185] = layer2_out[1877] ^ layer2_out[1878];
    assign layer3_out[7186] = layer2_out[984];
    assign layer3_out[7187] = layer2_out[2685] & ~layer2_out[2686];
    assign layer3_out[7188] = layer2_out[161] & ~layer2_out[160];
    assign layer3_out[7189] = layer2_out[6606] & ~layer2_out[6607];
    assign layer3_out[7190] = layer2_out[283];
    assign layer3_out[7191] = layer2_out[504] & ~layer2_out[503];
    assign layer3_out[7192] = ~layer2_out[3883];
    assign layer3_out[7193] = ~layer2_out[572] | layer2_out[571];
    assign layer3_out[7194] = ~layer2_out[1216] | layer2_out[1217];
    assign layer3_out[7195] = ~layer2_out[1934];
    assign layer3_out[7196] = layer2_out[1645] & layer2_out[1646];
    assign layer3_out[7197] = layer2_out[7081];
    assign layer3_out[7198] = ~layer2_out[5019];
    assign layer3_out[7199] = ~(layer2_out[5022] | layer2_out[5023]);
    assign layer3_out[7200] = ~(layer2_out[624] ^ layer2_out[625]);
    assign layer3_out[7201] = layer2_out[2018] & ~layer2_out[2017];
    assign layer3_out[7202] = ~layer2_out[6158];
    assign layer3_out[7203] = layer2_out[5726];
    assign layer3_out[7204] = ~layer2_out[6206] | layer2_out[6205];
    assign layer3_out[7205] = ~layer2_out[6164];
    assign layer3_out[7206] = layer2_out[568];
    assign layer3_out[7207] = layer2_out[1690];
    assign layer3_out[7208] = layer2_out[49] | layer2_out[50];
    assign layer3_out[7209] = ~(layer2_out[891] ^ layer2_out[892]);
    assign layer3_out[7210] = layer2_out[2042] & ~layer2_out[2041];
    assign layer3_out[7211] = layer2_out[5727] & ~layer2_out[5728];
    assign layer3_out[7212] = layer2_out[5484] ^ layer2_out[5485];
    assign layer3_out[7213] = layer2_out[4101];
    assign layer3_out[7214] = ~layer2_out[714];
    assign layer3_out[7215] = layer2_out[4877] ^ layer2_out[4878];
    assign layer3_out[7216] = ~(layer2_out[7202] & layer2_out[7203]);
    assign layer3_out[7217] = layer2_out[7663] & ~layer2_out[7664];
    assign layer3_out[7218] = ~(layer2_out[777] & layer2_out[778]);
    assign layer3_out[7219] = 1'b1;
    assign layer3_out[7220] = layer2_out[1748];
    assign layer3_out[7221] = layer2_out[3247];
    assign layer3_out[7222] = ~(layer2_out[4492] & layer2_out[4493]);
    assign layer3_out[7223] = ~layer2_out[2852];
    assign layer3_out[7224] = ~(layer2_out[1412] | layer2_out[1413]);
    assign layer3_out[7225] = ~layer2_out[4957];
    assign layer3_out[7226] = layer2_out[4678] & layer2_out[4679];
    assign layer3_out[7227] = ~(layer2_out[4039] & layer2_out[4040]);
    assign layer3_out[7228] = ~layer2_out[6984];
    assign layer3_out[7229] = layer2_out[2161] ^ layer2_out[2162];
    assign layer3_out[7230] = ~(layer2_out[4918] | layer2_out[4919]);
    assign layer3_out[7231] = layer2_out[5927];
    assign layer3_out[7232] = layer2_out[3259] | layer2_out[3260];
    assign layer3_out[7233] = layer2_out[7960] ^ layer2_out[7961];
    assign layer3_out[7234] = ~(layer2_out[1366] | layer2_out[1367]);
    assign layer3_out[7235] = ~layer2_out[6983] | layer2_out[6982];
    assign layer3_out[7236] = layer2_out[5791];
    assign layer3_out[7237] = layer2_out[5058];
    assign layer3_out[7238] = layer2_out[4904] ^ layer2_out[4905];
    assign layer3_out[7239] = ~layer2_out[3094] | layer2_out[3095];
    assign layer3_out[7240] = layer2_out[1106];
    assign layer3_out[7241] = layer2_out[725] & ~layer2_out[726];
    assign layer3_out[7242] = layer2_out[3186] & layer2_out[3187];
    assign layer3_out[7243] = ~layer2_out[2878];
    assign layer3_out[7244] = layer2_out[7043] & layer2_out[7044];
    assign layer3_out[7245] = layer2_out[6064];
    assign layer3_out[7246] = ~layer2_out[4328];
    assign layer3_out[7247] = ~(layer2_out[7808] | layer2_out[7809]);
    assign layer3_out[7248] = 1'b0;
    assign layer3_out[7249] = layer2_out[2294];
    assign layer3_out[7250] = ~(layer2_out[193] ^ layer2_out[194]);
    assign layer3_out[7251] = layer2_out[957] & layer2_out[958];
    assign layer3_out[7252] = layer2_out[4938];
    assign layer3_out[7253] = layer2_out[4483];
    assign layer3_out[7254] = ~(layer2_out[3625] & layer2_out[3626]);
    assign layer3_out[7255] = 1'b1;
    assign layer3_out[7256] = ~layer2_out[7011];
    assign layer3_out[7257] = layer2_out[201];
    assign layer3_out[7258] = ~(layer2_out[6548] | layer2_out[6549]);
    assign layer3_out[7259] = ~layer2_out[5685];
    assign layer3_out[7260] = layer2_out[4523];
    assign layer3_out[7261] = layer2_out[5862] ^ layer2_out[5863];
    assign layer3_out[7262] = ~(layer2_out[6373] ^ layer2_out[6374]);
    assign layer3_out[7263] = layer2_out[6407] & ~layer2_out[6406];
    assign layer3_out[7264] = ~(layer2_out[4057] | layer2_out[4058]);
    assign layer3_out[7265] = layer2_out[1597];
    assign layer3_out[7266] = ~(layer2_out[1765] ^ layer2_out[1766]);
    assign layer3_out[7267] = layer2_out[7495];
    assign layer3_out[7268] = layer2_out[4166] | layer2_out[4167];
    assign layer3_out[7269] = 1'b1;
    assign layer3_out[7270] = layer2_out[5587];
    assign layer3_out[7271] = ~layer2_out[7136] | layer2_out[7137];
    assign layer3_out[7272] = ~layer2_out[7912];
    assign layer3_out[7273] = layer2_out[108];
    assign layer3_out[7274] = layer2_out[5164];
    assign layer3_out[7275] = layer2_out[877];
    assign layer3_out[7276] = ~(layer2_out[1556] & layer2_out[1557]);
    assign layer3_out[7277] = layer2_out[728] ^ layer2_out[729];
    assign layer3_out[7278] = ~(layer2_out[5661] & layer2_out[5662]);
    assign layer3_out[7279] = ~layer2_out[6357];
    assign layer3_out[7280] = layer2_out[5138];
    assign layer3_out[7281] = ~layer2_out[2230];
    assign layer3_out[7282] = ~layer2_out[4408] | layer2_out[4409];
    assign layer3_out[7283] = ~(layer2_out[3187] ^ layer2_out[3188]);
    assign layer3_out[7284] = ~layer2_out[6801];
    assign layer3_out[7285] = layer2_out[4370];
    assign layer3_out[7286] = layer2_out[3485] | layer2_out[3486];
    assign layer3_out[7287] = layer2_out[1843] & ~layer2_out[1844];
    assign layer3_out[7288] = layer2_out[4828] & ~layer2_out[4827];
    assign layer3_out[7289] = layer2_out[5918] ^ layer2_out[5919];
    assign layer3_out[7290] = ~layer2_out[2524];
    assign layer3_out[7291] = layer2_out[3922];
    assign layer3_out[7292] = ~(layer2_out[6188] ^ layer2_out[6189]);
    assign layer3_out[7293] = ~(layer2_out[3527] ^ layer2_out[3528]);
    assign layer3_out[7294] = layer2_out[1064] ^ layer2_out[1065];
    assign layer3_out[7295] = layer2_out[6603];
    assign layer3_out[7296] = layer2_out[2916] & ~layer2_out[2917];
    assign layer3_out[7297] = ~layer2_out[1152];
    assign layer3_out[7298] = ~layer2_out[6669];
    assign layer3_out[7299] = ~layer2_out[7579];
    assign layer3_out[7300] = layer2_out[7714] | layer2_out[7715];
    assign layer3_out[7301] = 1'b0;
    assign layer3_out[7302] = ~layer2_out[6392];
    assign layer3_out[7303] = layer2_out[7175] | layer2_out[7176];
    assign layer3_out[7304] = layer2_out[4352];
    assign layer3_out[7305] = layer2_out[386];
    assign layer3_out[7306] = ~(layer2_out[1297] | layer2_out[1298]);
    assign layer3_out[7307] = layer2_out[7466] ^ layer2_out[7467];
    assign layer3_out[7308] = ~(layer2_out[1655] & layer2_out[1656]);
    assign layer3_out[7309] = ~layer2_out[41];
    assign layer3_out[7310] = layer2_out[3976];
    assign layer3_out[7311] = ~layer2_out[4531];
    assign layer3_out[7312] = layer2_out[5735] ^ layer2_out[5736];
    assign layer3_out[7313] = layer2_out[2304];
    assign layer3_out[7314] = layer2_out[7541] & layer2_out[7542];
    assign layer3_out[7315] = ~(layer2_out[6620] ^ layer2_out[6621]);
    assign layer3_out[7316] = ~(layer2_out[6709] & layer2_out[6710]);
    assign layer3_out[7317] = ~layer2_out[878];
    assign layer3_out[7318] = layer2_out[7906];
    assign layer3_out[7319] = layer2_out[7299] & ~layer2_out[7298];
    assign layer3_out[7320] = ~layer2_out[4043];
    assign layer3_out[7321] = ~layer2_out[316];
    assign layer3_out[7322] = layer2_out[7211] & ~layer2_out[7210];
    assign layer3_out[7323] = ~layer2_out[6087] | layer2_out[6086];
    assign layer3_out[7324] = ~layer2_out[3921] | layer2_out[3920];
    assign layer3_out[7325] = ~layer2_out[6482];
    assign layer3_out[7326] = ~layer2_out[5469];
    assign layer3_out[7327] = ~layer2_out[727] | layer2_out[726];
    assign layer3_out[7328] = layer2_out[4724];
    assign layer3_out[7329] = layer2_out[3284] & ~layer2_out[3285];
    assign layer3_out[7330] = ~(layer2_out[2604] | layer2_out[2605]);
    assign layer3_out[7331] = ~layer2_out[911];
    assign layer3_out[7332] = 1'b1;
    assign layer3_out[7333] = ~layer2_out[1862];
    assign layer3_out[7334] = layer2_out[3308] & ~layer2_out[3307];
    assign layer3_out[7335] = ~(layer2_out[4494] ^ layer2_out[4495]);
    assign layer3_out[7336] = ~layer2_out[4615] | layer2_out[4616];
    assign layer3_out[7337] = ~layer2_out[6457];
    assign layer3_out[7338] = ~(layer2_out[7687] & layer2_out[7688]);
    assign layer3_out[7339] = ~layer2_out[1332];
    assign layer3_out[7340] = layer2_out[914] & ~layer2_out[915];
    assign layer3_out[7341] = layer2_out[2738] & layer2_out[2739];
    assign layer3_out[7342] = layer2_out[4695];
    assign layer3_out[7343] = layer2_out[211];
    assign layer3_out[7344] = ~layer2_out[1087];
    assign layer3_out[7345] = layer2_out[2400] ^ layer2_out[2401];
    assign layer3_out[7346] = layer2_out[2468] & layer2_out[2469];
    assign layer3_out[7347] = ~layer2_out[2116];
    assign layer3_out[7348] = ~layer2_out[6171] | layer2_out[6172];
    assign layer3_out[7349] = ~layer2_out[1004];
    assign layer3_out[7350] = ~layer2_out[6999];
    assign layer3_out[7351] = layer2_out[621] & ~layer2_out[620];
    assign layer3_out[7352] = ~layer2_out[3594];
    assign layer3_out[7353] = layer2_out[3774] ^ layer2_out[3775];
    assign layer3_out[7354] = ~(layer2_out[7880] & layer2_out[7881]);
    assign layer3_out[7355] = layer2_out[7484] ^ layer2_out[7485];
    assign layer3_out[7356] = ~(layer2_out[4862] ^ layer2_out[4863]);
    assign layer3_out[7357] = layer2_out[866];
    assign layer3_out[7358] = layer2_out[3996] & layer2_out[3997];
    assign layer3_out[7359] = ~layer2_out[1069];
    assign layer3_out[7360] = layer2_out[4968];
    assign layer3_out[7361] = layer2_out[2184];
    assign layer3_out[7362] = layer2_out[7763] ^ layer2_out[7764];
    assign layer3_out[7363] = ~(layer2_out[6843] ^ layer2_out[6844]);
    assign layer3_out[7364] = layer2_out[4510];
    assign layer3_out[7365] = layer2_out[4610];
    assign layer3_out[7366] = ~layer2_out[2873] | layer2_out[2872];
    assign layer3_out[7367] = layer2_out[6573] | layer2_out[6574];
    assign layer3_out[7368] = ~layer2_out[7037] | layer2_out[7036];
    assign layer3_out[7369] = ~(layer2_out[7260] | layer2_out[7261]);
    assign layer3_out[7370] = ~layer2_out[1780];
    assign layer3_out[7371] = 1'b1;
    assign layer3_out[7372] = layer2_out[4816] ^ layer2_out[4817];
    assign layer3_out[7373] = ~layer2_out[1187] | layer2_out[1188];
    assign layer3_out[7374] = layer2_out[5625] & ~layer2_out[5624];
    assign layer3_out[7375] = ~layer2_out[3502];
    assign layer3_out[7376] = layer2_out[4858];
    assign layer3_out[7377] = 1'b0;
    assign layer3_out[7378] = ~(layer2_out[411] ^ layer2_out[412]);
    assign layer3_out[7379] = ~layer2_out[6791];
    assign layer3_out[7380] = layer2_out[6746] & ~layer2_out[6747];
    assign layer3_out[7381] = ~layer2_out[213] | layer2_out[214];
    assign layer3_out[7382] = ~layer2_out[6088];
    assign layer3_out[7383] = layer2_out[65] & ~layer2_out[64];
    assign layer3_out[7384] = layer2_out[6476] ^ layer2_out[6477];
    assign layer3_out[7385] = layer2_out[417];
    assign layer3_out[7386] = ~(layer2_out[4147] ^ layer2_out[4148]);
    assign layer3_out[7387] = ~layer2_out[7956];
    assign layer3_out[7388] = layer2_out[5333] & ~layer2_out[5332];
    assign layer3_out[7389] = ~(layer2_out[6659] ^ layer2_out[6660]);
    assign layer3_out[7390] = layer2_out[2600] | layer2_out[2601];
    assign layer3_out[7391] = layer2_out[2771] ^ layer2_out[2772];
    assign layer3_out[7392] = ~layer2_out[2553];
    assign layer3_out[7393] = ~layer2_out[518];
    assign layer3_out[7394] = layer2_out[116];
    assign layer3_out[7395] = layer2_out[3132];
    assign layer3_out[7396] = layer2_out[6848] & ~layer2_out[6847];
    assign layer3_out[7397] = ~layer2_out[1975];
    assign layer3_out[7398] = ~(layer2_out[3001] | layer2_out[3002]);
    assign layer3_out[7399] = layer2_out[7990];
    assign layer3_out[7400] = ~(layer2_out[2664] & layer2_out[2665]);
    assign layer3_out[7401] = ~layer2_out[4572];
    assign layer3_out[7402] = layer2_out[2915] & layer2_out[2916];
    assign layer3_out[7403] = ~layer2_out[7959] | layer2_out[7960];
    assign layer3_out[7404] = layer2_out[3803];
    assign layer3_out[7405] = layer2_out[2227] & ~layer2_out[2228];
    assign layer3_out[7406] = layer2_out[4665];
    assign layer3_out[7407] = layer2_out[1139];
    assign layer3_out[7408] = ~layer2_out[7260] | layer2_out[7259];
    assign layer3_out[7409] = ~layer2_out[3306];
    assign layer3_out[7410] = ~(layer2_out[2272] | layer2_out[2273]);
    assign layer3_out[7411] = layer2_out[5193];
    assign layer3_out[7412] = ~layer2_out[2758];
    assign layer3_out[7413] = ~layer2_out[486];
    assign layer3_out[7414] = layer2_out[7318];
    assign layer3_out[7415] = layer2_out[6587];
    assign layer3_out[7416] = layer2_out[6838] & layer2_out[6839];
    assign layer3_out[7417] = ~(layer2_out[6329] | layer2_out[6330]);
    assign layer3_out[7418] = ~(layer2_out[3099] & layer2_out[3100]);
    assign layer3_out[7419] = ~layer2_out[5145];
    assign layer3_out[7420] = layer2_out[4251] | layer2_out[4252];
    assign layer3_out[7421] = ~(layer2_out[4826] ^ layer2_out[4827]);
    assign layer3_out[7422] = ~layer2_out[3151];
    assign layer3_out[7423] = layer2_out[1160];
    assign layer3_out[7424] = layer2_out[7468] & ~layer2_out[7469];
    assign layer3_out[7425] = layer2_out[6537] & ~layer2_out[6536];
    assign layer3_out[7426] = ~layer2_out[5444];
    assign layer3_out[7427] = layer2_out[2876];
    assign layer3_out[7428] = ~(layer2_out[7232] ^ layer2_out[7233]);
    assign layer3_out[7429] = layer2_out[6290] & layer2_out[6291];
    assign layer3_out[7430] = layer2_out[5006];
    assign layer3_out[7431] = layer2_out[1354] | layer2_out[1355];
    assign layer3_out[7432] = ~layer2_out[6634] | layer2_out[6633];
    assign layer3_out[7433] = layer2_out[1093] & layer2_out[1094];
    assign layer3_out[7434] = ~(layer2_out[7871] | layer2_out[7872]);
    assign layer3_out[7435] = layer2_out[4124] & layer2_out[4125];
    assign layer3_out[7436] = ~layer2_out[1324];
    assign layer3_out[7437] = layer2_out[2636] & layer2_out[2637];
    assign layer3_out[7438] = ~layer2_out[7190];
    assign layer3_out[7439] = ~layer2_out[5880] | layer2_out[5879];
    assign layer3_out[7440] = layer2_out[3532] | layer2_out[3533];
    assign layer3_out[7441] = layer2_out[4033];
    assign layer3_out[7442] = ~layer2_out[6451];
    assign layer3_out[7443] = layer2_out[6354] ^ layer2_out[6355];
    assign layer3_out[7444] = layer2_out[611] ^ layer2_out[612];
    assign layer3_out[7445] = layer2_out[3185] | layer2_out[3186];
    assign layer3_out[7446] = layer2_out[2549];
    assign layer3_out[7447] = layer2_out[169];
    assign layer3_out[7448] = layer2_out[7736] & ~layer2_out[7737];
    assign layer3_out[7449] = layer2_out[4646];
    assign layer3_out[7450] = ~layer2_out[5684];
    assign layer3_out[7451] = ~layer2_out[559];
    assign layer3_out[7452] = ~layer2_out[6142];
    assign layer3_out[7453] = layer2_out[2102] | layer2_out[2103];
    assign layer3_out[7454] = layer2_out[5477] & ~layer2_out[5478];
    assign layer3_out[7455] = layer2_out[6629] ^ layer2_out[6630];
    assign layer3_out[7456] = ~layer2_out[2835];
    assign layer3_out[7457] = ~(layer2_out[5234] & layer2_out[5235]);
    assign layer3_out[7458] = ~(layer2_out[744] & layer2_out[745]);
    assign layer3_out[7459] = ~layer2_out[1105];
    assign layer3_out[7460] = layer2_out[795] | layer2_out[796];
    assign layer3_out[7461] = layer2_out[3529];
    assign layer3_out[7462] = ~layer2_out[6093] | layer2_out[6094];
    assign layer3_out[7463] = layer2_out[5591];
    assign layer3_out[7464] = ~(layer2_out[7447] & layer2_out[7448]);
    assign layer3_out[7465] = layer2_out[5419] & layer2_out[5420];
    assign layer3_out[7466] = layer2_out[369];
    assign layer3_out[7467] = layer2_out[4309] & ~layer2_out[4308];
    assign layer3_out[7468] = ~layer2_out[7250] | layer2_out[7251];
    assign layer3_out[7469] = layer2_out[6242];
    assign layer3_out[7470] = ~(layer2_out[2719] & layer2_out[2720]);
    assign layer3_out[7471] = ~(layer2_out[1520] & layer2_out[1521]);
    assign layer3_out[7472] = layer2_out[7123] | layer2_out[7124];
    assign layer3_out[7473] = layer2_out[3311];
    assign layer3_out[7474] = layer2_out[1993] & layer2_out[1994];
    assign layer3_out[7475] = layer2_out[1616] & ~layer2_out[1617];
    assign layer3_out[7476] = layer2_out[932];
    assign layer3_out[7477] = ~layer2_out[2787];
    assign layer3_out[7478] = ~layer2_out[7447] | layer2_out[7446];
    assign layer3_out[7479] = layer2_out[7665] | layer2_out[7666];
    assign layer3_out[7480] = layer2_out[2763] ^ layer2_out[2764];
    assign layer3_out[7481] = layer2_out[5463] & ~layer2_out[5462];
    assign layer3_out[7482] = layer2_out[7723] & ~layer2_out[7722];
    assign layer3_out[7483] = layer2_out[6378];
    assign layer3_out[7484] = layer2_out[4297] ^ layer2_out[4298];
    assign layer3_out[7485] = layer2_out[6050] ^ layer2_out[6051];
    assign layer3_out[7486] = ~layer2_out[7196];
    assign layer3_out[7487] = layer2_out[4992] | layer2_out[4993];
    assign layer3_out[7488] = layer2_out[7591];
    assign layer3_out[7489] = ~layer2_out[2123];
    assign layer3_out[7490] = ~layer2_out[1124];
    assign layer3_out[7491] = layer2_out[3397] & layer2_out[3398];
    assign layer3_out[7492] = layer2_out[768];
    assign layer3_out[7493] = ~layer2_out[6076];
    assign layer3_out[7494] = layer2_out[255] | layer2_out[256];
    assign layer3_out[7495] = layer2_out[3460];
    assign layer3_out[7496] = 1'b1;
    assign layer3_out[7497] = ~layer2_out[2008];
    assign layer3_out[7498] = ~layer2_out[6438];
    assign layer3_out[7499] = ~layer2_out[883] | layer2_out[884];
    assign layer3_out[7500] = ~(layer2_out[3818] & layer2_out[3819]);
    assign layer3_out[7501] = layer2_out[5158];
    assign layer3_out[7502] = layer2_out[2753];
    assign layer3_out[7503] = layer2_out[4183] ^ layer2_out[4184];
    assign layer3_out[7504] = ~layer2_out[7548] | layer2_out[7547];
    assign layer3_out[7505] = 1'b0;
    assign layer3_out[7506] = layer2_out[2329] & layer2_out[2330];
    assign layer3_out[7507] = layer2_out[5110] & ~layer2_out[5111];
    assign layer3_out[7508] = ~layer2_out[531];
    assign layer3_out[7509] = ~(layer2_out[6374] & layer2_out[6375]);
    assign layer3_out[7510] = ~layer2_out[5278] | layer2_out[5277];
    assign layer3_out[7511] = ~layer2_out[5757];
    assign layer3_out[7512] = ~(layer2_out[4555] ^ layer2_out[4556]);
    assign layer3_out[7513] = layer2_out[2064];
    assign layer3_out[7514] = layer2_out[5155] & layer2_out[5156];
    assign layer3_out[7515] = layer2_out[6241];
    assign layer3_out[7516] = layer2_out[1905];
    assign layer3_out[7517] = ~(layer2_out[52] ^ layer2_out[53]);
    assign layer3_out[7518] = ~layer2_out[2730] | layer2_out[2729];
    assign layer3_out[7519] = ~layer2_out[558] | layer2_out[557];
    assign layer3_out[7520] = layer2_out[6574] & ~layer2_out[6575];
    assign layer3_out[7521] = layer2_out[2010];
    assign layer3_out[7522] = ~layer2_out[5194] | layer2_out[5195];
    assign layer3_out[7523] = layer2_out[1672];
    assign layer3_out[7524] = layer2_out[4665] & ~layer2_out[4666];
    assign layer3_out[7525] = ~layer2_out[7883];
    assign layer3_out[7526] = ~layer2_out[5377];
    assign layer3_out[7527] = layer2_out[7843] & ~layer2_out[7842];
    assign layer3_out[7528] = layer2_out[3748] | layer2_out[3749];
    assign layer3_out[7529] = layer2_out[580];
    assign layer3_out[7530] = ~(layer2_out[272] & layer2_out[273]);
    assign layer3_out[7531] = layer2_out[3488] ^ layer2_out[3489];
    assign layer3_out[7532] = ~layer2_out[1384] | layer2_out[1385];
    assign layer3_out[7533] = layer2_out[7608];
    assign layer3_out[7534] = layer2_out[438] & ~layer2_out[439];
    assign layer3_out[7535] = ~layer2_out[4089];
    assign layer3_out[7536] = ~layer2_out[7594];
    assign layer3_out[7537] = ~(layer2_out[1789] ^ layer2_out[1790]);
    assign layer3_out[7538] = layer2_out[7011] & ~layer2_out[7010];
    assign layer3_out[7539] = ~(layer2_out[5135] | layer2_out[5136]);
    assign layer3_out[7540] = ~layer2_out[4733];
    assign layer3_out[7541] = layer2_out[3710] & layer2_out[3711];
    assign layer3_out[7542] = layer2_out[6179] & ~layer2_out[6180];
    assign layer3_out[7543] = ~(layer2_out[6097] ^ layer2_out[6098]);
    assign layer3_out[7544] = layer2_out[4412];
    assign layer3_out[7545] = ~layer2_out[3213];
    assign layer3_out[7546] = ~(layer2_out[1534] ^ layer2_out[1535]);
    assign layer3_out[7547] = layer2_out[7716];
    assign layer3_out[7548] = ~layer2_out[3758];
    assign layer3_out[7549] = layer2_out[1686];
    assign layer3_out[7550] = layer2_out[7628];
    assign layer3_out[7551] = layer2_out[2372] & ~layer2_out[2373];
    assign layer3_out[7552] = ~layer2_out[5328] | layer2_out[5327];
    assign layer3_out[7553] = layer2_out[7188];
    assign layer3_out[7554] = layer2_out[2389];
    assign layer3_out[7555] = layer2_out[2143] | layer2_out[2144];
    assign layer3_out[7556] = layer2_out[127];
    assign layer3_out[7557] = ~(layer2_out[3545] & layer2_out[3546]);
    assign layer3_out[7558] = layer2_out[2970];
    assign layer3_out[7559] = layer2_out[4449];
    assign layer3_out[7560] = layer2_out[573];
    assign layer3_out[7561] = layer2_out[4363];
    assign layer3_out[7562] = layer2_out[2968] | layer2_out[2969];
    assign layer3_out[7563] = layer2_out[498] ^ layer2_out[499];
    assign layer3_out[7564] = ~(layer2_out[7306] ^ layer2_out[7307]);
    assign layer3_out[7565] = ~layer2_out[5454];
    assign layer3_out[7566] = layer2_out[3829];
    assign layer3_out[7567] = ~(layer2_out[2364] | layer2_out[2365]);
    assign layer3_out[7568] = layer2_out[1264] | layer2_out[1265];
    assign layer3_out[7569] = ~layer2_out[6350];
    assign layer3_out[7570] = layer2_out[5925] | layer2_out[5926];
    assign layer3_out[7571] = ~(layer2_out[7234] & layer2_out[7235]);
    assign layer3_out[7572] = ~layer2_out[3212] | layer2_out[3213];
    assign layer3_out[7573] = ~layer2_out[379];
    assign layer3_out[7574] = layer2_out[1223] & ~layer2_out[1224];
    assign layer3_out[7575] = layer2_out[768];
    assign layer3_out[7576] = layer2_out[3493];
    assign layer3_out[7577] = ~layer2_out[1732];
    assign layer3_out[7578] = layer2_out[5294];
    assign layer3_out[7579] = layer2_out[4953] & ~layer2_out[4954];
    assign layer3_out[7580] = ~(layer2_out[6432] ^ layer2_out[6433]);
    assign layer3_out[7581] = layer2_out[4855];
    assign layer3_out[7582] = layer2_out[244];
    assign layer3_out[7583] = layer2_out[3742] & ~layer2_out[3741];
    assign layer3_out[7584] = layer2_out[6613];
    assign layer3_out[7585] = ~layer2_out[4858];
    assign layer3_out[7586] = layer2_out[3469] & ~layer2_out[3468];
    assign layer3_out[7587] = layer2_out[10];
    assign layer3_out[7588] = layer2_out[5784] & ~layer2_out[5783];
    assign layer3_out[7589] = ~(layer2_out[6623] & layer2_out[6624]);
    assign layer3_out[7590] = layer2_out[7084] & layer2_out[7085];
    assign layer3_out[7591] = ~layer2_out[3043];
    assign layer3_out[7592] = 1'b0;
    assign layer3_out[7593] = layer2_out[2343];
    assign layer3_out[7594] = ~layer2_out[3895];
    assign layer3_out[7595] = layer2_out[1399];
    assign layer3_out[7596] = layer2_out[5038] & layer2_out[5039];
    assign layer3_out[7597] = ~layer2_out[7588];
    assign layer3_out[7598] = layer2_out[7762];
    assign layer3_out[7599] = ~layer2_out[6728];
    assign layer3_out[7600] = ~(layer2_out[7438] ^ layer2_out[7439]);
    assign layer3_out[7601] = ~(layer2_out[2753] & layer2_out[2754]);
    assign layer3_out[7602] = layer2_out[7629] | layer2_out[7630];
    assign layer3_out[7603] = layer2_out[7956];
    assign layer3_out[7604] = ~layer2_out[3241] | layer2_out[3240];
    assign layer3_out[7605] = layer2_out[1361] & ~layer2_out[1362];
    assign layer3_out[7606] = 1'b0;
    assign layer3_out[7607] = layer2_out[6632] ^ layer2_out[6633];
    assign layer3_out[7608] = layer2_out[2418];
    assign layer3_out[7609] = layer2_out[4975] ^ layer2_out[4976];
    assign layer3_out[7610] = ~layer2_out[6580];
    assign layer3_out[7611] = ~layer2_out[4848] | layer2_out[4849];
    assign layer3_out[7612] = ~layer2_out[3359] | layer2_out[3360];
    assign layer3_out[7613] = ~layer2_out[5178];
    assign layer3_out[7614] = ~layer2_out[3506];
    assign layer3_out[7615] = ~layer2_out[2210] | layer2_out[2209];
    assign layer3_out[7616] = ~(layer2_out[3743] | layer2_out[3744]);
    assign layer3_out[7617] = layer2_out[4994];
    assign layer3_out[7618] = ~layer2_out[7864];
    assign layer3_out[7619] = layer2_out[86] & ~layer2_out[87];
    assign layer3_out[7620] = ~(layer2_out[4399] ^ layer2_out[4400]);
    assign layer3_out[7621] = layer2_out[3936] ^ layer2_out[3937];
    assign layer3_out[7622] = ~(layer2_out[4701] ^ layer2_out[4702]);
    assign layer3_out[7623] = layer2_out[5610];
    assign layer3_out[7624] = ~(layer2_out[5420] & layer2_out[5421]);
    assign layer3_out[7625] = ~(layer2_out[4841] ^ layer2_out[4842]);
    assign layer3_out[7626] = ~layer2_out[6982] | layer2_out[6981];
    assign layer3_out[7627] = layer2_out[4800];
    assign layer3_out[7628] = ~layer2_out[3642] | layer2_out[3643];
    assign layer3_out[7629] = layer2_out[5647];
    assign layer3_out[7630] = layer2_out[4213] & ~layer2_out[4214];
    assign layer3_out[7631] = layer2_out[279] ^ layer2_out[280];
    assign layer3_out[7632] = ~(layer2_out[7379] ^ layer2_out[7380]);
    assign layer3_out[7633] = layer2_out[4376];
    assign layer3_out[7634] = ~layer2_out[3367];
    assign layer3_out[7635] = layer2_out[2592] & ~layer2_out[2591];
    assign layer3_out[7636] = ~layer2_out[3496];
    assign layer3_out[7637] = layer2_out[5520] & layer2_out[5521];
    assign layer3_out[7638] = ~(layer2_out[1161] & layer2_out[1162]);
    assign layer3_out[7639] = ~layer2_out[2298];
    assign layer3_out[7640] = layer2_out[4943];
    assign layer3_out[7641] = ~layer2_out[1144];
    assign layer3_out[7642] = ~layer2_out[3650] | layer2_out[3651];
    assign layer3_out[7643] = layer2_out[372];
    assign layer3_out[7644] = ~(layer2_out[7033] | layer2_out[7034]);
    assign layer3_out[7645] = layer2_out[4281];
    assign layer3_out[7646] = ~layer2_out[3009];
    assign layer3_out[7647] = ~(layer2_out[7507] ^ layer2_out[7508]);
    assign layer3_out[7648] = ~layer2_out[669];
    assign layer3_out[7649] = ~(layer2_out[7047] & layer2_out[7048]);
    assign layer3_out[7650] = layer2_out[4224] ^ layer2_out[4225];
    assign layer3_out[7651] = ~layer2_out[2978];
    assign layer3_out[7652] = ~(layer2_out[5422] ^ layer2_out[5423]);
    assign layer3_out[7653] = ~layer2_out[5981] | layer2_out[5980];
    assign layer3_out[7654] = layer2_out[6488];
    assign layer3_out[7655] = ~(layer2_out[3300] ^ layer2_out[3301]);
    assign layer3_out[7656] = 1'b0;
    assign layer3_out[7657] = layer2_out[6319];
    assign layer3_out[7658] = ~layer2_out[436];
    assign layer3_out[7659] = layer2_out[7452] & layer2_out[7453];
    assign layer3_out[7660] = layer2_out[966];
    assign layer3_out[7661] = ~(layer2_out[2518] | layer2_out[2519]);
    assign layer3_out[7662] = layer2_out[4570] & ~layer2_out[4571];
    assign layer3_out[7663] = ~(layer2_out[7451] | layer2_out[7452]);
    assign layer3_out[7664] = ~(layer2_out[5573] ^ layer2_out[5574]);
    assign layer3_out[7665] = ~layer2_out[6587];
    assign layer3_out[7666] = ~(layer2_out[1078] & layer2_out[1079]);
    assign layer3_out[7667] = ~layer2_out[1023];
    assign layer3_out[7668] = ~(layer2_out[6786] & layer2_out[6787]);
    assign layer3_out[7669] = layer2_out[2060];
    assign layer3_out[7670] = ~(layer2_out[2179] | layer2_out[2180]);
    assign layer3_out[7671] = layer2_out[7312] & layer2_out[7313];
    assign layer3_out[7672] = layer2_out[1204];
    assign layer3_out[7673] = ~(layer2_out[712] | layer2_out[713]);
    assign layer3_out[7674] = layer2_out[638];
    assign layer3_out[7675] = layer2_out[2361];
    assign layer3_out[7676] = ~layer2_out[3910];
    assign layer3_out[7677] = layer2_out[679] & ~layer2_out[678];
    assign layer3_out[7678] = ~layer2_out[7975];
    assign layer3_out[7679] = ~(layer2_out[455] & layer2_out[456]);
    assign layer3_out[7680] = layer2_out[2990] ^ layer2_out[2991];
    assign layer3_out[7681] = layer2_out[6004];
    assign layer3_out[7682] = ~(layer2_out[6730] & layer2_out[6731]);
    assign layer3_out[7683] = layer2_out[7644];
    assign layer3_out[7684] = 1'b1;
    assign layer3_out[7685] = ~layer2_out[6176] | layer2_out[6177];
    assign layer3_out[7686] = ~(layer2_out[7731] ^ layer2_out[7732]);
    assign layer3_out[7687] = ~(layer2_out[5314] | layer2_out[5315]);
    assign layer3_out[7688] = layer2_out[4120] & ~layer2_out[4121];
    assign layer3_out[7689] = layer2_out[1895];
    assign layer3_out[7690] = ~(layer2_out[3553] | layer2_out[3554]);
    assign layer3_out[7691] = ~layer2_out[5024] | layer2_out[5023];
    assign layer3_out[7692] = ~layer2_out[5716];
    assign layer3_out[7693] = layer2_out[3613];
    assign layer3_out[7694] = ~(layer2_out[7049] & layer2_out[7050]);
    assign layer3_out[7695] = ~layer2_out[12];
    assign layer3_out[7696] = layer2_out[4437] & ~layer2_out[4436];
    assign layer3_out[7697] = layer2_out[1551];
    assign layer3_out[7698] = 1'b0;
    assign layer3_out[7699] = ~layer2_out[166] | layer2_out[167];
    assign layer3_out[7700] = layer2_out[1060];
    assign layer3_out[7701] = layer2_out[159] | layer2_out[160];
    assign layer3_out[7702] = layer2_out[5099] & layer2_out[5100];
    assign layer3_out[7703] = layer2_out[371];
    assign layer3_out[7704] = layer2_out[5080];
    assign layer3_out[7705] = ~layer2_out[4226];
    assign layer3_out[7706] = layer2_out[5719];
    assign layer3_out[7707] = ~(layer2_out[3362] | layer2_out[3363]);
    assign layer3_out[7708] = ~layer2_out[232];
    assign layer3_out[7709] = 1'b0;
    assign layer3_out[7710] = layer2_out[4452];
    assign layer3_out[7711] = ~layer2_out[2253];
    assign layer3_out[7712] = ~layer2_out[3833] | layer2_out[3832];
    assign layer3_out[7713] = ~(layer2_out[4175] | layer2_out[4176]);
    assign layer3_out[7714] = layer2_out[4796];
    assign layer3_out[7715] = layer2_out[4364];
    assign layer3_out[7716] = ~layer2_out[1307] | layer2_out[1306];
    assign layer3_out[7717] = ~(layer2_out[2951] & layer2_out[2952]);
    assign layer3_out[7718] = ~layer2_out[4196];
    assign layer3_out[7719] = layer2_out[2824];
    assign layer3_out[7720] = ~layer2_out[4663] | layer2_out[4662];
    assign layer3_out[7721] = 1'b0;
    assign layer3_out[7722] = layer2_out[6598] & ~layer2_out[6597];
    assign layer3_out[7723] = layer2_out[7633];
    assign layer3_out[7724] = 1'b1;
    assign layer3_out[7725] = ~(layer2_out[4217] | layer2_out[4218]);
    assign layer3_out[7726] = layer2_out[152];
    assign layer3_out[7727] = ~layer2_out[4718];
    assign layer3_out[7728] = ~layer2_out[4314];
    assign layer3_out[7729] = ~layer2_out[1267];
    assign layer3_out[7730] = layer2_out[6867] & layer2_out[6868];
    assign layer3_out[7731] = ~layer2_out[4703];
    assign layer3_out[7732] = layer2_out[5302];
    assign layer3_out[7733] = layer2_out[2691];
    assign layer3_out[7734] = layer2_out[5776] ^ layer2_out[5777];
    assign layer3_out[7735] = 1'b0;
    assign layer3_out[7736] = 1'b1;
    assign layer3_out[7737] = ~(layer2_out[1035] | layer2_out[1036]);
    assign layer3_out[7738] = layer2_out[5247];
    assign layer3_out[7739] = ~layer2_out[1283];
    assign layer3_out[7740] = layer2_out[6856] ^ layer2_out[6857];
    assign layer3_out[7741] = layer2_out[1879] ^ layer2_out[1880];
    assign layer3_out[7742] = layer2_out[1311];
    assign layer3_out[7743] = ~layer2_out[2231] | layer2_out[2232];
    assign layer3_out[7744] = layer2_out[7789] & layer2_out[7790];
    assign layer3_out[7745] = ~layer2_out[5624];
    assign layer3_out[7746] = ~layer2_out[7214];
    assign layer3_out[7747] = layer2_out[4940] & layer2_out[4941];
    assign layer3_out[7748] = ~(layer2_out[5433] ^ layer2_out[5434]);
    assign layer3_out[7749] = ~layer2_out[2329];
    assign layer3_out[7750] = ~layer2_out[4490];
    assign layer3_out[7751] = ~layer2_out[3215];
    assign layer3_out[7752] = layer2_out[1693];
    assign layer3_out[7753] = ~(layer2_out[5251] & layer2_out[5252]);
    assign layer3_out[7754] = ~layer2_out[6272];
    assign layer3_out[7755] = ~layer2_out[1383];
    assign layer3_out[7756] = layer2_out[1968] | layer2_out[1969];
    assign layer3_out[7757] = ~layer2_out[306] | layer2_out[305];
    assign layer3_out[7758] = ~(layer2_out[241] | layer2_out[242]);
    assign layer3_out[7759] = layer2_out[6515];
    assign layer3_out[7760] = ~layer2_out[7697];
    assign layer3_out[7761] = ~layer2_out[3632] | layer2_out[3631];
    assign layer3_out[7762] = layer2_out[1883] & ~layer2_out[1882];
    assign layer3_out[7763] = layer2_out[4186] | layer2_out[4187];
    assign layer3_out[7764] = ~layer2_out[2781];
    assign layer3_out[7765] = ~(layer2_out[5984] | layer2_out[5985]);
    assign layer3_out[7766] = layer2_out[3290];
    assign layer3_out[7767] = ~(layer2_out[7876] & layer2_out[7877]);
    assign layer3_out[7768] = ~(layer2_out[4034] | layer2_out[4035]);
    assign layer3_out[7769] = layer2_out[3723];
    assign layer3_out[7770] = layer2_out[35];
    assign layer3_out[7771] = layer2_out[241];
    assign layer3_out[7772] = ~(layer2_out[5607] & layer2_out[5608]);
    assign layer3_out[7773] = layer2_out[2273] & layer2_out[2274];
    assign layer3_out[7774] = ~layer2_out[1831] | layer2_out[1832];
    assign layer3_out[7775] = ~layer2_out[3285] | layer2_out[3286];
    assign layer3_out[7776] = layer2_out[1352];
    assign layer3_out[7777] = layer2_out[7876];
    assign layer3_out[7778] = ~layer2_out[7591];
    assign layer3_out[7779] = ~layer2_out[6301];
    assign layer3_out[7780] = layer2_out[4710] | layer2_out[4711];
    assign layer3_out[7781] = layer2_out[6430];
    assign layer3_out[7782] = ~(layer2_out[1371] | layer2_out[1372]);
    assign layer3_out[7783] = ~layer2_out[5730];
    assign layer3_out[7784] = layer2_out[7117];
    assign layer3_out[7785] = layer2_out[594] ^ layer2_out[595];
    assign layer3_out[7786] = layer2_out[101] & ~layer2_out[102];
    assign layer3_out[7787] = layer2_out[1207];
    assign layer3_out[7788] = layer2_out[2029] & layer2_out[2030];
    assign layer3_out[7789] = layer2_out[1209] & ~layer2_out[1208];
    assign layer3_out[7790] = layer2_out[3422];
    assign layer3_out[7791] = ~layer2_out[6583];
    assign layer3_out[7792] = ~layer2_out[730];
    assign layer3_out[7793] = ~layer2_out[5725];
    assign layer3_out[7794] = ~layer2_out[40] | layer2_out[39];
    assign layer3_out[7795] = layer2_out[2540];
    assign layer3_out[7796] = ~(layer2_out[7310] ^ layer2_out[7311]);
    assign layer3_out[7797] = ~layer2_out[2146];
    assign layer3_out[7798] = layer2_out[7602] ^ layer2_out[7603];
    assign layer3_out[7799] = layer2_out[3209];
    assign layer3_out[7800] = ~layer2_out[6399];
    assign layer3_out[7801] = ~(layer2_out[2408] & layer2_out[2409]);
    assign layer3_out[7802] = ~layer2_out[2196] | layer2_out[2197];
    assign layer3_out[7803] = layer2_out[4473];
    assign layer3_out[7804] = ~(layer2_out[300] & layer2_out[301]);
    assign layer3_out[7805] = layer2_out[7166] & layer2_out[7167];
    assign layer3_out[7806] = ~layer2_out[6369];
    assign layer3_out[7807] = ~layer2_out[6661] | layer2_out[6660];
    assign layer3_out[7808] = layer2_out[943] ^ layer2_out[944];
    assign layer3_out[7809] = layer2_out[6326] & layer2_out[6327];
    assign layer3_out[7810] = ~(layer2_out[2517] ^ layer2_out[2518]);
    assign layer3_out[7811] = ~layer2_out[2870] | layer2_out[2871];
    assign layer3_out[7812] = ~layer2_out[3064];
    assign layer3_out[7813] = layer2_out[1664] ^ layer2_out[1665];
    assign layer3_out[7814] = layer2_out[270] | layer2_out[271];
    assign layer3_out[7815] = ~(layer2_out[7368] & layer2_out[7369]);
    assign layer3_out[7816] = layer2_out[5020] & ~layer2_out[5019];
    assign layer3_out[7817] = ~layer2_out[2316] | layer2_out[2317];
    assign layer3_out[7818] = ~layer2_out[1775] | layer2_out[1776];
    assign layer3_out[7819] = ~layer2_out[7989] | layer2_out[7988];
    assign layer3_out[7820] = ~(layer2_out[5130] ^ layer2_out[5131]);
    assign layer3_out[7821] = ~(layer2_out[6987] ^ layer2_out[6988]);
    assign layer3_out[7822] = ~layer2_out[4185];
    assign layer3_out[7823] = ~layer2_out[461];
    assign layer3_out[7824] = ~layer2_out[1889] | layer2_out[1890];
    assign layer3_out[7825] = ~(layer2_out[6155] | layer2_out[6156]);
    assign layer3_out[7826] = ~(layer2_out[1898] | layer2_out[1899]);
    assign layer3_out[7827] = layer2_out[2804] ^ layer2_out[2805];
    assign layer3_out[7828] = layer2_out[4190];
    assign layer3_out[7829] = ~layer2_out[2562] | layer2_out[2561];
    assign layer3_out[7830] = ~layer2_out[646] | layer2_out[645];
    assign layer3_out[7831] = ~layer2_out[1858];
    assign layer3_out[7832] = layer2_out[214] & ~layer2_out[215];
    assign layer3_out[7833] = ~(layer2_out[5686] & layer2_out[5687]);
    assign layer3_out[7834] = layer2_out[7813] & ~layer2_out[7814];
    assign layer3_out[7835] = ~layer2_out[7060];
    assign layer3_out[7836] = layer2_out[4152];
    assign layer3_out[7837] = ~(layer2_out[6379] & layer2_out[6380]);
    assign layer3_out[7838] = layer2_out[3735];
    assign layer3_out[7839] = ~(layer2_out[2623] & layer2_out[2624]);
    assign layer3_out[7840] = layer2_out[6371] ^ layer2_out[6372];
    assign layer3_out[7841] = ~layer2_out[3646];
    assign layer3_out[7842] = layer2_out[1446];
    assign layer3_out[7843] = ~layer2_out[589];
    assign layer3_out[7844] = ~layer2_out[6616];
    assign layer3_out[7845] = ~layer2_out[6408];
    assign layer3_out[7846] = ~(layer2_out[1742] ^ layer2_out[1743]);
    assign layer3_out[7847] = ~layer2_out[7169];
    assign layer3_out[7848] = ~layer2_out[7345];
    assign layer3_out[7849] = layer2_out[1580] & layer2_out[1581];
    assign layer3_out[7850] = ~layer2_out[6470] | layer2_out[6469];
    assign layer3_out[7851] = 1'b1;
    assign layer3_out[7852] = ~layer2_out[1533];
    assign layer3_out[7853] = layer2_out[1640];
    assign layer3_out[7854] = layer2_out[6090];
    assign layer3_out[7855] = ~(layer2_out[3113] ^ layer2_out[3114]);
    assign layer3_out[7856] = ~(layer2_out[5340] ^ layer2_out[5341]);
    assign layer3_out[7857] = layer2_out[7273] & ~layer2_out[7272];
    assign layer3_out[7858] = ~layer2_out[6426];
    assign layer3_out[7859] = layer2_out[3783] & layer2_out[3784];
    assign layer3_out[7860] = layer2_out[3968] & layer2_out[3969];
    assign layer3_out[7861] = ~(layer2_out[4978] & layer2_out[4979]);
    assign layer3_out[7862] = layer2_out[5577];
    assign layer3_out[7863] = ~layer2_out[3129];
    assign layer3_out[7864] = ~layer2_out[2647];
    assign layer3_out[7865] = ~layer2_out[3153];
    assign layer3_out[7866] = layer2_out[875];
    assign layer3_out[7867] = ~layer2_out[2292];
    assign layer3_out[7868] = layer2_out[7457] | layer2_out[7458];
    assign layer3_out[7869] = ~layer2_out[947] | layer2_out[948];
    assign layer3_out[7870] = ~layer2_out[6895];
    assign layer3_out[7871] = layer2_out[1800] ^ layer2_out[1801];
    assign layer3_out[7872] = ~(layer2_out[1848] | layer2_out[1849]);
    assign layer3_out[7873] = layer2_out[2667] & ~layer2_out[2666];
    assign layer3_out[7874] = ~(layer2_out[6083] | layer2_out[6084]);
    assign layer3_out[7875] = ~(layer2_out[5034] | layer2_out[5035]);
    assign layer3_out[7876] = layer2_out[4507];
    assign layer3_out[7877] = ~(layer2_out[1435] ^ layer2_out[1436]);
    assign layer3_out[7878] = ~layer2_out[1849];
    assign layer3_out[7879] = layer2_out[6460] | layer2_out[6461];
    assign layer3_out[7880] = ~(layer2_out[4329] ^ layer2_out[4330]);
    assign layer3_out[7881] = layer2_out[1227] & ~layer2_out[1228];
    assign layer3_out[7882] = ~layer2_out[6789];
    assign layer3_out[7883] = layer2_out[4043] | layer2_out[4044];
    assign layer3_out[7884] = ~(layer2_out[4496] & layer2_out[4497]);
    assign layer3_out[7885] = ~(layer2_out[95] & layer2_out[96]);
    assign layer3_out[7886] = ~layer2_out[5950];
    assign layer3_out[7887] = 1'b1;
    assign layer3_out[7888] = ~(layer2_out[2716] | layer2_out[2717]);
    assign layer3_out[7889] = layer2_out[5012] & ~layer2_out[5011];
    assign layer3_out[7890] = layer2_out[956];
    assign layer3_out[7891] = ~(layer2_out[7149] & layer2_out[7150]);
    assign layer3_out[7892] = layer2_out[34];
    assign layer3_out[7893] = ~(layer2_out[5957] & layer2_out[5958]);
    assign layer3_out[7894] = ~layer2_out[4398];
    assign layer3_out[7895] = 1'b1;
    assign layer3_out[7896] = layer2_out[4618];
    assign layer3_out[7897] = layer2_out[4922] ^ layer2_out[4923];
    assign layer3_out[7898] = ~layer2_out[6676];
    assign layer3_out[7899] = ~(layer2_out[3951] & layer2_out[3952]);
    assign layer3_out[7900] = ~(layer2_out[7738] | layer2_out[7739]);
    assign layer3_out[7901] = layer2_out[4182];
    assign layer3_out[7902] = layer2_out[3853];
    assign layer3_out[7903] = layer2_out[5874];
    assign layer3_out[7904] = ~layer2_out[6861];
    assign layer3_out[7905] = layer2_out[784];
    assign layer3_out[7906] = ~layer2_out[3540];
    assign layer3_out[7907] = layer2_out[4382];
    assign layer3_out[7908] = layer2_out[5472] & layer2_out[5473];
    assign layer3_out[7909] = ~layer2_out[1266] | layer2_out[1267];
    assign layer3_out[7910] = layer2_out[5888] & layer2_out[5889];
    assign layer3_out[7911] = layer2_out[595] & ~layer2_out[596];
    assign layer3_out[7912] = layer2_out[1218] & ~layer2_out[1217];
    assign layer3_out[7913] = ~layer2_out[5381] | layer2_out[5380];
    assign layer3_out[7914] = layer2_out[3361] | layer2_out[3362];
    assign layer3_out[7915] = ~layer2_out[3026];
    assign layer3_out[7916] = layer2_out[4659];
    assign layer3_out[7917] = layer2_out[5086];
    assign layer3_out[7918] = ~layer2_out[7173] | layer2_out[7172];
    assign layer3_out[7919] = ~layer2_out[1295] | layer2_out[1294];
    assign layer3_out[7920] = layer2_out[5867] & ~layer2_out[5868];
    assign layer3_out[7921] = ~layer2_out[3797];
    assign layer3_out[7922] = ~layer2_out[7962];
    assign layer3_out[7923] = layer2_out[5297] & ~layer2_out[5298];
    assign layer3_out[7924] = layer2_out[4983] & ~layer2_out[4984];
    assign layer3_out[7925] = layer2_out[2512];
    assign layer3_out[7926] = layer2_out[1056];
    assign layer3_out[7927] = layer2_out[373];
    assign layer3_out[7928] = layer2_out[7642] & ~layer2_out[7641];
    assign layer3_out[7929] = 1'b1;
    assign layer3_out[7930] = ~layer2_out[3188];
    assign layer3_out[7931] = layer2_out[3941];
    assign layer3_out[7932] = layer2_out[4357] & ~layer2_out[4356];
    assign layer3_out[7933] = ~layer2_out[4092] | layer2_out[4093];
    assign layer3_out[7934] = layer2_out[2801] & ~layer2_out[2802];
    assign layer3_out[7935] = layer2_out[965] & ~layer2_out[964];
    assign layer3_out[7936] = layer2_out[7919] ^ layer2_out[7920];
    assign layer3_out[7937] = ~layer2_out[6550];
    assign layer3_out[7938] = layer2_out[2526] & layer2_out[2527];
    assign layer3_out[7939] = layer2_out[6288];
    assign layer3_out[7940] = ~layer2_out[5978];
    assign layer3_out[7941] = layer2_out[6908];
    assign layer3_out[7942] = layer2_out[3263];
    assign layer3_out[7943] = layer2_out[4923];
    assign layer3_out[7944] = layer2_out[5983] | layer2_out[5984];
    assign layer3_out[7945] = ~layer2_out[4539] | layer2_out[4538];
    assign layer3_out[7946] = ~layer2_out[4897] | layer2_out[4896];
    assign layer3_out[7947] = ~layer2_out[498];
    assign layer3_out[7948] = layer2_out[7647] | layer2_out[7648];
    assign layer3_out[7949] = layer2_out[2406] | layer2_out[2407];
    assign layer3_out[7950] = layer2_out[3594] | layer2_out[3595];
    assign layer3_out[7951] = layer2_out[2003];
    assign layer3_out[7952] = ~layer2_out[5245] | layer2_out[5244];
    assign layer3_out[7953] = ~(layer2_out[5359] ^ layer2_out[5360]);
    assign layer3_out[7954] = layer2_out[2850] | layer2_out[2851];
    assign layer3_out[7955] = ~(layer2_out[112] & layer2_out[113]);
    assign layer3_out[7956] = ~layer2_out[2353];
    assign layer3_out[7957] = layer2_out[4876] | layer2_out[4877];
    assign layer3_out[7958] = ~layer2_out[3031] | layer2_out[3030];
    assign layer3_out[7959] = 1'b0;
    assign layer3_out[7960] = ~layer2_out[816] | layer2_out[817];
    assign layer3_out[7961] = layer2_out[3410] | layer2_out[3411];
    assign layer3_out[7962] = layer2_out[1327] ^ layer2_out[1328];
    assign layer3_out[7963] = layer2_out[6759] ^ layer2_out[6760];
    assign layer3_out[7964] = ~layer2_out[2201];
    assign layer3_out[7965] = ~(layer2_out[7054] | layer2_out[7055]);
    assign layer3_out[7966] = 1'b0;
    assign layer3_out[7967] = layer2_out[5366] & ~layer2_out[5367];
    assign layer3_out[7968] = layer2_out[6845] & ~layer2_out[6844];
    assign layer3_out[7969] = ~layer2_out[191];
    assign layer3_out[7970] = layer2_out[6223] & layer2_out[6224];
    assign layer3_out[7971] = layer2_out[4615];
    assign layer3_out[7972] = layer2_out[634];
    assign layer3_out[7973] = ~(layer2_out[5636] | layer2_out[5637]);
    assign layer3_out[7974] = layer2_out[2613] & ~layer2_out[2614];
    assign layer3_out[7975] = ~(layer2_out[6261] ^ layer2_out[6262]);
    assign layer3_out[7976] = ~(layer2_out[7780] | layer2_out[7781]);
    assign layer3_out[7977] = layer2_out[6223];
    assign layer3_out[7978] = layer2_out[5705];
    assign layer3_out[7979] = ~layer2_out[4835] | layer2_out[4834];
    assign layer3_out[7980] = ~layer2_out[4738];
    assign layer3_out[7981] = layer2_out[6504];
    assign layer3_out[7982] = 1'b0;
    assign layer3_out[7983] = ~layer2_out[6389];
    assign layer3_out[7984] = layer2_out[1450];
    assign layer3_out[7985] = ~layer2_out[512];
    assign layer3_out[7986] = ~(layer2_out[1061] | layer2_out[1062]);
    assign layer3_out[7987] = ~layer2_out[7206];
    assign layer3_out[7988] = layer2_out[7146] & ~layer2_out[7145];
    assign layer3_out[7989] = ~layer2_out[547] | layer2_out[548];
    assign layer3_out[7990] = layer2_out[866] & ~layer2_out[867];
    assign layer3_out[7991] = layer2_out[187];
    assign layer3_out[7992] = ~layer2_out[5843] | layer2_out[5842];
    assign layer3_out[7993] = layer2_out[7269];
    assign layer3_out[7994] = ~layer2_out[5441];
    assign layer3_out[7995] = layer2_out[4477] | layer2_out[4478];
    assign layer3_out[7996] = ~layer2_out[2931];
    assign layer3_out[7997] = layer2_out[7863] & ~layer2_out[7862];
    assign layer3_out[7998] = ~layer2_out[7769] | layer2_out[7768];
    assign layer3_out[7999] = layer2_out[1511] & ~layer2_out[1510];
    assign layer4_out[0] = layer3_out[5269] ^ layer3_out[5270];
    assign layer4_out[1] = layer3_out[4675];
    assign layer4_out[2] = layer3_out[1933];
    assign layer4_out[3] = ~(layer3_out[3701] ^ layer3_out[3702]);
    assign layer4_out[4] = ~(layer3_out[5641] | layer3_out[5642]);
    assign layer4_out[5] = layer3_out[7831] & ~layer3_out[7830];
    assign layer4_out[6] = ~(layer3_out[1973] ^ layer3_out[1974]);
    assign layer4_out[7] = layer3_out[5045];
    assign layer4_out[8] = layer3_out[913] & ~layer3_out[914];
    assign layer4_out[9] = ~layer3_out[5145] | layer3_out[5146];
    assign layer4_out[10] = ~(layer3_out[930] ^ layer3_out[931]);
    assign layer4_out[11] = ~layer3_out[3112];
    assign layer4_out[12] = ~(layer3_out[6984] | layer3_out[6985]);
    assign layer4_out[13] = ~layer3_out[150];
    assign layer4_out[14] = ~(layer3_out[3518] ^ layer3_out[3519]);
    assign layer4_out[15] = layer3_out[7776] & ~layer3_out[7775];
    assign layer4_out[16] = layer3_out[7819] & ~layer3_out[7820];
    assign layer4_out[17] = layer3_out[4302];
    assign layer4_out[18] = layer3_out[6772] & ~layer3_out[6771];
    assign layer4_out[19] = layer3_out[4347];
    assign layer4_out[20] = ~(layer3_out[6635] | layer3_out[6636]);
    assign layer4_out[21] = ~(layer3_out[6317] & layer3_out[6318]);
    assign layer4_out[22] = ~(layer3_out[3820] ^ layer3_out[3821]);
    assign layer4_out[23] = layer3_out[2331] | layer3_out[2332];
    assign layer4_out[24] = ~layer3_out[5055] | layer3_out[5054];
    assign layer4_out[25] = ~layer3_out[280];
    assign layer4_out[26] = layer3_out[2922] & ~layer3_out[2923];
    assign layer4_out[27] = ~layer3_out[6467] | layer3_out[6468];
    assign layer4_out[28] = ~layer3_out[533] | layer3_out[532];
    assign layer4_out[29] = ~(layer3_out[1494] | layer3_out[1495]);
    assign layer4_out[30] = ~layer3_out[2039] | layer3_out[2040];
    assign layer4_out[31] = ~layer3_out[679];
    assign layer4_out[32] = layer3_out[7984] | layer3_out[7985];
    assign layer4_out[33] = ~layer3_out[4076];
    assign layer4_out[34] = layer3_out[2298];
    assign layer4_out[35] = layer3_out[2214] ^ layer3_out[2215];
    assign layer4_out[36] = layer3_out[3226] & ~layer3_out[3225];
    assign layer4_out[37] = layer3_out[7988] | layer3_out[7989];
    assign layer4_out[38] = layer3_out[5417] & ~layer3_out[5418];
    assign layer4_out[39] = ~(layer3_out[2621] | layer3_out[2622]);
    assign layer4_out[40] = layer3_out[1662];
    assign layer4_out[41] = ~(layer3_out[3013] & layer3_out[3014]);
    assign layer4_out[42] = layer3_out[5981] | layer3_out[5982];
    assign layer4_out[43] = ~(layer3_out[1513] ^ layer3_out[1514]);
    assign layer4_out[44] = layer3_out[3361] ^ layer3_out[3362];
    assign layer4_out[45] = layer3_out[1016] & layer3_out[1017];
    assign layer4_out[46] = ~(layer3_out[3160] & layer3_out[3161]);
    assign layer4_out[47] = layer3_out[1517] | layer3_out[1518];
    assign layer4_out[48] = ~layer3_out[2220] | layer3_out[2221];
    assign layer4_out[49] = ~(layer3_out[2557] & layer3_out[2558]);
    assign layer4_out[50] = layer3_out[836] ^ layer3_out[837];
    assign layer4_out[51] = layer3_out[1327] ^ layer3_out[1328];
    assign layer4_out[52] = ~(layer3_out[6335] & layer3_out[6336]);
    assign layer4_out[53] = layer3_out[3091];
    assign layer4_out[54] = ~layer3_out[4466];
    assign layer4_out[55] = ~(layer3_out[3095] ^ layer3_out[3096]);
    assign layer4_out[56] = ~layer3_out[977] | layer3_out[978];
    assign layer4_out[57] = ~layer3_out[3015];
    assign layer4_out[58] = ~(layer3_out[2841] & layer3_out[2842]);
    assign layer4_out[59] = layer3_out[903] & layer3_out[904];
    assign layer4_out[60] = ~layer3_out[3730];
    assign layer4_out[61] = ~(layer3_out[4307] ^ layer3_out[4308]);
    assign layer4_out[62] = ~(layer3_out[3249] | layer3_out[3250]);
    assign layer4_out[63] = ~layer3_out[5611] | layer3_out[5612];
    assign layer4_out[64] = ~layer3_out[1507];
    assign layer4_out[65] = ~(layer3_out[998] ^ layer3_out[999]);
    assign layer4_out[66] = layer3_out[6890];
    assign layer4_out[67] = layer3_out[6963];
    assign layer4_out[68] = ~(layer3_out[6769] & layer3_out[6770]);
    assign layer4_out[69] = layer3_out[3758] | layer3_out[3759];
    assign layer4_out[70] = layer3_out[4132] & layer3_out[4133];
    assign layer4_out[71] = ~(layer3_out[6170] & layer3_out[6171]);
    assign layer4_out[72] = layer3_out[6004] | layer3_out[6005];
    assign layer4_out[73] = ~layer3_out[6501];
    assign layer4_out[74] = ~layer3_out[4486];
    assign layer4_out[75] = ~layer3_out[5726] | layer3_out[5725];
    assign layer4_out[76] = layer3_out[6218] & ~layer3_out[6217];
    assign layer4_out[77] = layer3_out[6360];
    assign layer4_out[78] = ~(layer3_out[2579] ^ layer3_out[2580]);
    assign layer4_out[79] = ~layer3_out[4228];
    assign layer4_out[80] = ~layer3_out[5381];
    assign layer4_out[81] = layer3_out[2608];
    assign layer4_out[82] = layer3_out[565] ^ layer3_out[566];
    assign layer4_out[83] = layer3_out[6054] & layer3_out[6055];
    assign layer4_out[84] = ~(layer3_out[5767] & layer3_out[5768]);
    assign layer4_out[85] = layer3_out[5427];
    assign layer4_out[86] = layer3_out[4196] & ~layer3_out[4197];
    assign layer4_out[87] = ~layer3_out[3974];
    assign layer4_out[88] = ~(layer3_out[6370] | layer3_out[6371]);
    assign layer4_out[89] = layer3_out[1450] & ~layer3_out[1449];
    assign layer4_out[90] = ~layer3_out[1053] | layer3_out[1054];
    assign layer4_out[91] = layer3_out[6492] & ~layer3_out[6493];
    assign layer4_out[92] = ~layer3_out[6376];
    assign layer4_out[93] = layer3_out[7436];
    assign layer4_out[94] = layer3_out[2244];
    assign layer4_out[95] = layer3_out[1540];
    assign layer4_out[96] = ~(layer3_out[7979] ^ layer3_out[7980]);
    assign layer4_out[97] = layer3_out[6498] ^ layer3_out[6499];
    assign layer4_out[98] = layer3_out[842] | layer3_out[843];
    assign layer4_out[99] = layer3_out[455];
    assign layer4_out[100] = layer3_out[5835];
    assign layer4_out[101] = ~layer3_out[6430] | layer3_out[6431];
    assign layer4_out[102] = ~(layer3_out[2633] | layer3_out[2634]);
    assign layer4_out[103] = layer3_out[3406];
    assign layer4_out[104] = ~(layer3_out[3370] ^ layer3_out[3371]);
    assign layer4_out[105] = layer3_out[5171] & ~layer3_out[5172];
    assign layer4_out[106] = layer3_out[5047] ^ layer3_out[5048];
    assign layer4_out[107] = ~(layer3_out[4670] ^ layer3_out[4671]);
    assign layer4_out[108] = layer3_out[1709] & ~layer3_out[1708];
    assign layer4_out[109] = layer3_out[6616] & ~layer3_out[6617];
    assign layer4_out[110] = layer3_out[2259] & ~layer3_out[2260];
    assign layer4_out[111] = layer3_out[7341];
    assign layer4_out[112] = layer3_out[5951] ^ layer3_out[5952];
    assign layer4_out[113] = ~layer3_out[7215];
    assign layer4_out[114] = layer3_out[2096];
    assign layer4_out[115] = layer3_out[6453];
    assign layer4_out[116] = layer3_out[3440] | layer3_out[3441];
    assign layer4_out[117] = ~layer3_out[6933];
    assign layer4_out[118] = layer3_out[1074] ^ layer3_out[1075];
    assign layer4_out[119] = layer3_out[507];
    assign layer4_out[120] = ~layer3_out[6318] | layer3_out[6319];
    assign layer4_out[121] = ~layer3_out[1438];
    assign layer4_out[122] = ~(layer3_out[6519] | layer3_out[6520]);
    assign layer4_out[123] = ~layer3_out[3821];
    assign layer4_out[124] = 1'b1;
    assign layer4_out[125] = ~layer3_out[2017];
    assign layer4_out[126] = layer3_out[3752] & ~layer3_out[3753];
    assign layer4_out[127] = layer3_out[2146] & ~layer3_out[2145];
    assign layer4_out[128] = ~layer3_out[2627];
    assign layer4_out[129] = ~layer3_out[4737];
    assign layer4_out[130] = ~(layer3_out[2506] & layer3_out[2507]);
    assign layer4_out[131] = ~layer3_out[2832];
    assign layer4_out[132] = ~layer3_out[3954] | layer3_out[3955];
    assign layer4_out[133] = layer3_out[2529];
    assign layer4_out[134] = ~(layer3_out[3949] & layer3_out[3950]);
    assign layer4_out[135] = ~layer3_out[1157];
    assign layer4_out[136] = ~(layer3_out[3392] & layer3_out[3393]);
    assign layer4_out[137] = ~(layer3_out[4652] | layer3_out[4653]);
    assign layer4_out[138] = ~(layer3_out[7090] ^ layer3_out[7091]);
    assign layer4_out[139] = layer3_out[1225];
    assign layer4_out[140] = layer3_out[4010];
    assign layer4_out[141] = ~layer3_out[7783];
    assign layer4_out[142] = layer3_out[4564];
    assign layer4_out[143] = ~layer3_out[7005];
    assign layer4_out[144] = ~(layer3_out[7125] | layer3_out[7126]);
    assign layer4_out[145] = ~(layer3_out[4051] ^ layer3_out[4052]);
    assign layer4_out[146] = layer3_out[4979] & layer3_out[4980];
    assign layer4_out[147] = ~layer3_out[5231];
    assign layer4_out[148] = ~(layer3_out[3962] ^ layer3_out[3963]);
    assign layer4_out[149] = ~layer3_out[5835] | layer3_out[5834];
    assign layer4_out[150] = ~(layer3_out[6753] & layer3_out[6754]);
    assign layer4_out[151] = layer3_out[2696];
    assign layer4_out[152] = layer3_out[4028] & layer3_out[4029];
    assign layer4_out[153] = layer3_out[493];
    assign layer4_out[154] = ~layer3_out[646];
    assign layer4_out[155] = layer3_out[2821] ^ layer3_out[2822];
    assign layer4_out[156] = ~layer3_out[6907];
    assign layer4_out[157] = ~layer3_out[6474];
    assign layer4_out[158] = layer3_out[4504] & ~layer3_out[4505];
    assign layer4_out[159] = layer3_out[1784] ^ layer3_out[1785];
    assign layer4_out[160] = ~layer3_out[2352] | layer3_out[2351];
    assign layer4_out[161] = layer3_out[124] | layer3_out[125];
    assign layer4_out[162] = layer3_out[4408];
    assign layer4_out[163] = ~(layer3_out[3297] ^ layer3_out[3298]);
    assign layer4_out[164] = ~layer3_out[4148];
    assign layer4_out[165] = ~(layer3_out[3637] | layer3_out[3638]);
    assign layer4_out[166] = ~layer3_out[4674];
    assign layer4_out[167] = ~layer3_out[3281];
    assign layer4_out[168] = ~(layer3_out[1262] & layer3_out[1263]);
    assign layer4_out[169] = ~layer3_out[1710];
    assign layer4_out[170] = 1'b0;
    assign layer4_out[171] = ~(layer3_out[822] ^ layer3_out[823]);
    assign layer4_out[172] = layer3_out[3284] & ~layer3_out[3283];
    assign layer4_out[173] = ~(layer3_out[77] ^ layer3_out[78]);
    assign layer4_out[174] = layer3_out[7418] & ~layer3_out[7419];
    assign layer4_out[175] = layer3_out[326] & layer3_out[327];
    assign layer4_out[176] = ~layer3_out[3173];
    assign layer4_out[177] = ~layer3_out[1856];
    assign layer4_out[178] = layer3_out[6395] & layer3_out[6396];
    assign layer4_out[179] = ~(layer3_out[1186] & layer3_out[1187]);
    assign layer4_out[180] = layer3_out[4303] ^ layer3_out[4304];
    assign layer4_out[181] = ~(layer3_out[3964] & layer3_out[3965]);
    assign layer4_out[182] = ~layer3_out[5556];
    assign layer4_out[183] = ~layer3_out[7266] | layer3_out[7267];
    assign layer4_out[184] = layer3_out[6611] ^ layer3_out[6612];
    assign layer4_out[185] = ~(layer3_out[4288] ^ layer3_out[4289]);
    assign layer4_out[186] = layer3_out[7057] & ~layer3_out[7056];
    assign layer4_out[187] = ~(layer3_out[7651] & layer3_out[7652]);
    assign layer4_out[188] = ~(layer3_out[2732] | layer3_out[2733]);
    assign layer4_out[189] = layer3_out[5265];
    assign layer4_out[190] = ~(layer3_out[5313] & layer3_out[5314]);
    assign layer4_out[191] = layer3_out[3587] | layer3_out[3588];
    assign layer4_out[192] = layer3_out[7138];
    assign layer4_out[193] = ~layer3_out[6627] | layer3_out[6626];
    assign layer4_out[194] = layer3_out[3505];
    assign layer4_out[195] = ~layer3_out[3365] | layer3_out[3366];
    assign layer4_out[196] = layer3_out[2044];
    assign layer4_out[197] = ~(layer3_out[694] & layer3_out[695]);
    assign layer4_out[198] = ~layer3_out[2900] | layer3_out[2901];
    assign layer4_out[199] = layer3_out[3080] ^ layer3_out[3081];
    assign layer4_out[200] = layer3_out[2917];
    assign layer4_out[201] = ~layer3_out[6185];
    assign layer4_out[202] = layer3_out[2810];
    assign layer4_out[203] = layer3_out[2801];
    assign layer4_out[204] = layer3_out[25];
    assign layer4_out[205] = ~layer3_out[403];
    assign layer4_out[206] = layer3_out[6752] & layer3_out[6753];
    assign layer4_out[207] = ~layer3_out[1202];
    assign layer4_out[208] = ~(layer3_out[1419] ^ layer3_out[1420]);
    assign layer4_out[209] = ~(layer3_out[3766] ^ layer3_out[3767]);
    assign layer4_out[210] = ~layer3_out[934] | layer3_out[935];
    assign layer4_out[211] = layer3_out[202] & layer3_out[203];
    assign layer4_out[212] = ~layer3_out[7291];
    assign layer4_out[213] = layer3_out[444] | layer3_out[445];
    assign layer4_out[214] = ~layer3_out[7657];
    assign layer4_out[215] = layer3_out[3989] & layer3_out[3990];
    assign layer4_out[216] = layer3_out[5573];
    assign layer4_out[217] = layer3_out[2613];
    assign layer4_out[218] = layer3_out[984] & layer3_out[985];
    assign layer4_out[219] = layer3_out[6076];
    assign layer4_out[220] = ~layer3_out[5124];
    assign layer4_out[221] = layer3_out[4974] & ~layer3_out[4975];
    assign layer4_out[222] = ~(layer3_out[5161] & layer3_out[5162]);
    assign layer4_out[223] = ~layer3_out[2959] | layer3_out[2960];
    assign layer4_out[224] = layer3_out[1690];
    assign layer4_out[225] = ~(layer3_out[1236] ^ layer3_out[1237]);
    assign layer4_out[226] = layer3_out[2122];
    assign layer4_out[227] = layer3_out[7186] & ~layer3_out[7187];
    assign layer4_out[228] = ~(layer3_out[1515] ^ layer3_out[1516]);
    assign layer4_out[229] = layer3_out[2956];
    assign layer4_out[230] = ~(layer3_out[2057] ^ layer3_out[2058]);
    assign layer4_out[231] = ~(layer3_out[4420] | layer3_out[4421]);
    assign layer4_out[232] = ~layer3_out[7184];
    assign layer4_out[233] = layer3_out[7979];
    assign layer4_out[234] = layer3_out[3756] & ~layer3_out[3757];
    assign layer4_out[235] = layer3_out[6832] ^ layer3_out[6833];
    assign layer4_out[236] = layer3_out[7593] & ~layer3_out[7592];
    assign layer4_out[237] = layer3_out[4844] ^ layer3_out[4845];
    assign layer4_out[238] = ~(layer3_out[6639] ^ layer3_out[6640]);
    assign layer4_out[239] = ~layer3_out[151];
    assign layer4_out[240] = ~(layer3_out[4804] ^ layer3_out[4805]);
    assign layer4_out[241] = layer3_out[5485];
    assign layer4_out[242] = ~layer3_out[7974];
    assign layer4_out[243] = ~layer3_out[1393] | layer3_out[1394];
    assign layer4_out[244] = layer3_out[5074];
    assign layer4_out[245] = ~layer3_out[6588];
    assign layer4_out[246] = ~layer3_out[2947];
    assign layer4_out[247] = layer3_out[3548] & layer3_out[3549];
    assign layer4_out[248] = layer3_out[3313] ^ layer3_out[3314];
    assign layer4_out[249] = layer3_out[4164] | layer3_out[4165];
    assign layer4_out[250] = layer3_out[101] | layer3_out[102];
    assign layer4_out[251] = ~layer3_out[5335];
    assign layer4_out[252] = ~layer3_out[434] | layer3_out[435];
    assign layer4_out[253] = layer3_out[1051] & ~layer3_out[1050];
    assign layer4_out[254] = layer3_out[2619] & layer3_out[2620];
    assign layer4_out[255] = layer3_out[5127];
    assign layer4_out[256] = layer3_out[4609] & ~layer3_out[4610];
    assign layer4_out[257] = ~layer3_out[4909] | layer3_out[4910];
    assign layer4_out[258] = layer3_out[2781] ^ layer3_out[2782];
    assign layer4_out[259] = layer3_out[4633];
    assign layer4_out[260] = ~layer3_out[3564] | layer3_out[3563];
    assign layer4_out[261] = layer3_out[3775];
    assign layer4_out[262] = ~layer3_out[2015] | layer3_out[2016];
    assign layer4_out[263] = layer3_out[1522];
    assign layer4_out[264] = layer3_out[4547] & layer3_out[4548];
    assign layer4_out[265] = layer3_out[3540] ^ layer3_out[3541];
    assign layer4_out[266] = layer3_out[6874];
    assign layer4_out[267] = ~(layer3_out[6884] & layer3_out[6885]);
    assign layer4_out[268] = layer3_out[324];
    assign layer4_out[269] = ~layer3_out[6158] | layer3_out[6157];
    assign layer4_out[270] = ~layer3_out[5241];
    assign layer4_out[271] = ~layer3_out[1554];
    assign layer4_out[272] = layer3_out[1871];
    assign layer4_out[273] = ~layer3_out[6736];
    assign layer4_out[274] = ~layer3_out[2405];
    assign layer4_out[275] = layer3_out[4375] & ~layer3_out[4374];
    assign layer4_out[276] = ~(layer3_out[2306] & layer3_out[2307]);
    assign layer4_out[277] = layer3_out[5128] & layer3_out[5129];
    assign layer4_out[278] = layer3_out[1633] & layer3_out[1634];
    assign layer4_out[279] = layer3_out[426] & ~layer3_out[427];
    assign layer4_out[280] = layer3_out[5151];
    assign layer4_out[281] = ~layer3_out[3155];
    assign layer4_out[282] = ~layer3_out[6078] | layer3_out[6077];
    assign layer4_out[283] = layer3_out[4789] | layer3_out[4790];
    assign layer4_out[284] = ~(layer3_out[7907] | layer3_out[7908]);
    assign layer4_out[285] = layer3_out[2217];
    assign layer4_out[286] = ~layer3_out[5671];
    assign layer4_out[287] = layer3_out[4739];
    assign layer4_out[288] = ~(layer3_out[1277] & layer3_out[1278]);
    assign layer4_out[289] = layer3_out[18];
    assign layer4_out[290] = layer3_out[2976] ^ layer3_out[2977];
    assign layer4_out[291] = ~(layer3_out[7404] ^ layer3_out[7405]);
    assign layer4_out[292] = layer3_out[7576] & ~layer3_out[7577];
    assign layer4_out[293] = ~layer3_out[3017] | layer3_out[3018];
    assign layer4_out[294] = ~layer3_out[1861];
    assign layer4_out[295] = layer3_out[5898];
    assign layer4_out[296] = ~layer3_out[781];
    assign layer4_out[297] = ~(layer3_out[7318] | layer3_out[7319]);
    assign layer4_out[298] = ~layer3_out[1664] | layer3_out[1665];
    assign layer4_out[299] = ~layer3_out[1342];
    assign layer4_out[300] = ~layer3_out[373] | layer3_out[374];
    assign layer4_out[301] = layer3_out[2705];
    assign layer4_out[302] = ~layer3_out[3227];
    assign layer4_out[303] = ~(layer3_out[6786] ^ layer3_out[6787]);
    assign layer4_out[304] = ~layer3_out[6536];
    assign layer4_out[305] = layer3_out[3907];
    assign layer4_out[306] = layer3_out[4436] ^ layer3_out[4437];
    assign layer4_out[307] = layer3_out[2650] | layer3_out[2651];
    assign layer4_out[308] = ~(layer3_out[4331] | layer3_out[4332]);
    assign layer4_out[309] = ~layer3_out[2348];
    assign layer4_out[310] = layer3_out[6537] & ~layer3_out[6536];
    assign layer4_out[311] = 1'b0;
    assign layer4_out[312] = layer3_out[5831] & layer3_out[5832];
    assign layer4_out[313] = ~(layer3_out[578] ^ layer3_out[579]);
    assign layer4_out[314] = layer3_out[3065];
    assign layer4_out[315] = ~(layer3_out[409] | layer3_out[410]);
    assign layer4_out[316] = ~layer3_out[6271];
    assign layer4_out[317] = ~(layer3_out[4831] & layer3_out[4832]);
    assign layer4_out[318] = layer3_out[717] & ~layer3_out[716];
    assign layer4_out[319] = ~layer3_out[344];
    assign layer4_out[320] = layer3_out[7394] & layer3_out[7395];
    assign layer4_out[321] = layer3_out[3748] & layer3_out[3749];
    assign layer4_out[322] = layer3_out[1526];
    assign layer4_out[323] = ~layer3_out[4480];
    assign layer4_out[324] = ~layer3_out[1540] | layer3_out[1539];
    assign layer4_out[325] = 1'b1;
    assign layer4_out[326] = layer3_out[6228] | layer3_out[6229];
    assign layer4_out[327] = layer3_out[1721];
    assign layer4_out[328] = ~(layer3_out[6630] ^ layer3_out[6631]);
    assign layer4_out[329] = ~(layer3_out[7117] ^ layer3_out[7118]);
    assign layer4_out[330] = ~layer3_out[3097];
    assign layer4_out[331] = layer3_out[4698];
    assign layer4_out[332] = layer3_out[941] ^ layer3_out[942];
    assign layer4_out[333] = layer3_out[4860] ^ layer3_out[4861];
    assign layer4_out[334] = ~(layer3_out[2051] | layer3_out[2052]);
    assign layer4_out[335] = ~layer3_out[2070];
    assign layer4_out[336] = ~(layer3_out[1135] & layer3_out[1136]);
    assign layer4_out[337] = layer3_out[6706];
    assign layer4_out[338] = layer3_out[5192];
    assign layer4_out[339] = ~layer3_out[4202] | layer3_out[4201];
    assign layer4_out[340] = ~layer3_out[6619];
    assign layer4_out[341] = ~layer3_out[7651] | layer3_out[7650];
    assign layer4_out[342] = layer3_out[5487] & layer3_out[5488];
    assign layer4_out[343] = layer3_out[5988] ^ layer3_out[5989];
    assign layer4_out[344] = ~(layer3_out[3122] & layer3_out[3123]);
    assign layer4_out[345] = layer3_out[4338] ^ layer3_out[4339];
    assign layer4_out[346] = ~(layer3_out[335] | layer3_out[336]);
    assign layer4_out[347] = layer3_out[4631] ^ layer3_out[4632];
    assign layer4_out[348] = layer3_out[1822];
    assign layer4_out[349] = layer3_out[2142];
    assign layer4_out[350] = layer3_out[426];
    assign layer4_out[351] = layer3_out[7743] & ~layer3_out[7744];
    assign layer4_out[352] = layer3_out[4199] ^ layer3_out[4200];
    assign layer4_out[353] = layer3_out[5032] ^ layer3_out[5033];
    assign layer4_out[354] = ~layer3_out[4003];
    assign layer4_out[355] = layer3_out[7595];
    assign layer4_out[356] = layer3_out[488] & ~layer3_out[487];
    assign layer4_out[357] = layer3_out[6031] & layer3_out[6032];
    assign layer4_out[358] = ~(layer3_out[6689] ^ layer3_out[6690]);
    assign layer4_out[359] = layer3_out[6219];
    assign layer4_out[360] = layer3_out[7824] & ~layer3_out[7825];
    assign layer4_out[361] = ~layer3_out[1070] | layer3_out[1071];
    assign layer4_out[362] = layer3_out[5471] | layer3_out[5472];
    assign layer4_out[363] = layer3_out[273] & layer3_out[274];
    assign layer4_out[364] = layer3_out[2989] | layer3_out[2990];
    assign layer4_out[365] = ~layer3_out[2972];
    assign layer4_out[366] = layer3_out[6904] ^ layer3_out[6905];
    assign layer4_out[367] = layer3_out[1155] & ~layer3_out[1156];
    assign layer4_out[368] = ~layer3_out[6902] | layer3_out[6901];
    assign layer4_out[369] = layer3_out[5101] ^ layer3_out[5102];
    assign layer4_out[370] = ~layer3_out[4930];
    assign layer4_out[371] = layer3_out[4380] & ~layer3_out[4381];
    assign layer4_out[372] = ~(layer3_out[6066] ^ layer3_out[6067]);
    assign layer4_out[373] = ~(layer3_out[1007] ^ layer3_out[1008]);
    assign layer4_out[374] = ~layer3_out[5515];
    assign layer4_out[375] = layer3_out[2471] & layer3_out[2472];
    assign layer4_out[376] = layer3_out[6022];
    assign layer4_out[377] = ~layer3_out[6967];
    assign layer4_out[378] = layer3_out[6910] ^ layer3_out[6911];
    assign layer4_out[379] = layer3_out[2531] & ~layer3_out[2532];
    assign layer4_out[380] = ~(layer3_out[2489] ^ layer3_out[2490]);
    assign layer4_out[381] = layer3_out[4443] & layer3_out[4444];
    assign layer4_out[382] = ~layer3_out[4341];
    assign layer4_out[383] = layer3_out[6860] ^ layer3_out[6861];
    assign layer4_out[384] = layer3_out[609] & ~layer3_out[610];
    assign layer4_out[385] = ~layer3_out[4220];
    assign layer4_out[386] = layer3_out[7963];
    assign layer4_out[387] = layer3_out[7054] & ~layer3_out[7053];
    assign layer4_out[388] = ~(layer3_out[1356] ^ layer3_out[1357]);
    assign layer4_out[389] = ~(layer3_out[938] | layer3_out[939]);
    assign layer4_out[390] = ~(layer3_out[2212] & layer3_out[2213]);
    assign layer4_out[391] = ~(layer3_out[6821] & layer3_out[6822]);
    assign layer4_out[392] = layer3_out[6516];
    assign layer4_out[393] = layer3_out[6669];
    assign layer4_out[394] = layer3_out[5701];
    assign layer4_out[395] = ~(layer3_out[3551] ^ layer3_out[3552]);
    assign layer4_out[396] = layer3_out[6254] & layer3_out[6255];
    assign layer4_out[397] = ~layer3_out[4306];
    assign layer4_out[398] = layer3_out[7364] ^ layer3_out[7365];
    assign layer4_out[399] = layer3_out[1934];
    assign layer4_out[400] = ~layer3_out[625] | layer3_out[626];
    assign layer4_out[401] = layer3_out[1672] ^ layer3_out[1673];
    assign layer4_out[402] = ~layer3_out[2685];
    assign layer4_out[403] = layer3_out[4636] & ~layer3_out[4635];
    assign layer4_out[404] = layer3_out[5743] & ~layer3_out[5744];
    assign layer4_out[405] = ~layer3_out[5274] | layer3_out[5273];
    assign layer4_out[406] = layer3_out[3052];
    assign layer4_out[407] = layer3_out[2635];
    assign layer4_out[408] = ~layer3_out[5851];
    assign layer4_out[409] = layer3_out[4481];
    assign layer4_out[410] = ~layer3_out[1274];
    assign layer4_out[411] = ~layer3_out[6534];
    assign layer4_out[412] = ~layer3_out[899] | layer3_out[898];
    assign layer4_out[413] = layer3_out[7038] | layer3_out[7039];
    assign layer4_out[414] = ~layer3_out[4874];
    assign layer4_out[415] = layer3_out[5244] ^ layer3_out[5245];
    assign layer4_out[416] = layer3_out[6059] | layer3_out[6060];
    assign layer4_out[417] = layer3_out[4859];
    assign layer4_out[418] = ~(layer3_out[2389] & layer3_out[2390]);
    assign layer4_out[419] = layer3_out[1953];
    assign layer4_out[420] = ~layer3_out[5693];
    assign layer4_out[421] = layer3_out[4498];
    assign layer4_out[422] = ~layer3_out[1769] | layer3_out[1768];
    assign layer4_out[423] = ~(layer3_out[349] ^ layer3_out[350]);
    assign layer4_out[424] = layer3_out[6187];
    assign layer4_out[425] = layer3_out[1981] & layer3_out[1982];
    assign layer4_out[426] = ~layer3_out[1556] | layer3_out[1555];
    assign layer4_out[427] = layer3_out[2309] ^ layer3_out[2310];
    assign layer4_out[428] = ~layer3_out[5931];
    assign layer4_out[429] = layer3_out[3057] & layer3_out[3058];
    assign layer4_out[430] = layer3_out[6349] | layer3_out[6350];
    assign layer4_out[431] = layer3_out[1058];
    assign layer4_out[432] = layer3_out[6368] & ~layer3_out[6369];
    assign layer4_out[433] = ~layer3_out[2072];
    assign layer4_out[434] = ~(layer3_out[1604] ^ layer3_out[1605]);
    assign layer4_out[435] = layer3_out[7389] ^ layer3_out[7390];
    assign layer4_out[436] = ~(layer3_out[7587] | layer3_out[7588]);
    assign layer4_out[437] = layer3_out[6818];
    assign layer4_out[438] = ~(layer3_out[1471] | layer3_out[1472]);
    assign layer4_out[439] = ~(layer3_out[2658] ^ layer3_out[2659]);
    assign layer4_out[440] = layer3_out[2059];
    assign layer4_out[441] = ~layer3_out[7395];
    assign layer4_out[442] = layer3_out[373];
    assign layer4_out[443] = layer3_out[4567] & ~layer3_out[4566];
    assign layer4_out[444] = layer3_out[3536];
    assign layer4_out[445] = layer3_out[5396] & ~layer3_out[5395];
    assign layer4_out[446] = layer3_out[975] & ~layer3_out[974];
    assign layer4_out[447] = layer3_out[5272] & ~layer3_out[5271];
    assign layer4_out[448] = ~(layer3_out[1958] | layer3_out[1959]);
    assign layer4_out[449] = layer3_out[2569];
    assign layer4_out[450] = ~(layer3_out[6121] | layer3_out[6122]);
    assign layer4_out[451] = layer3_out[7798];
    assign layer4_out[452] = layer3_out[5015] ^ layer3_out[5016];
    assign layer4_out[453] = layer3_out[1907] & ~layer3_out[1906];
    assign layer4_out[454] = layer3_out[4015] & layer3_out[4016];
    assign layer4_out[455] = layer3_out[4370];
    assign layer4_out[456] = ~layer3_out[4933];
    assign layer4_out[457] = ~layer3_out[7298];
    assign layer4_out[458] = layer3_out[7726];
    assign layer4_out[459] = layer3_out[3706];
    assign layer4_out[460] = layer3_out[2643];
    assign layer4_out[461] = layer3_out[2206];
    assign layer4_out[462] = layer3_out[6042] & ~layer3_out[6041];
    assign layer4_out[463] = layer3_out[5752];
    assign layer4_out[464] = layer3_out[6717];
    assign layer4_out[465] = layer3_out[7734];
    assign layer4_out[466] = ~layer3_out[7957] | layer3_out[7956];
    assign layer4_out[467] = ~(layer3_out[5914] & layer3_out[5915]);
    assign layer4_out[468] = layer3_out[2537] & ~layer3_out[2536];
    assign layer4_out[469] = layer3_out[4073] ^ layer3_out[4074];
    assign layer4_out[470] = ~layer3_out[41];
    assign layer4_out[471] = layer3_out[7116] & layer3_out[7117];
    assign layer4_out[472] = layer3_out[3887] ^ layer3_out[3888];
    assign layer4_out[473] = ~(layer3_out[7937] ^ layer3_out[7938]);
    assign layer4_out[474] = layer3_out[3907];
    assign layer4_out[475] = layer3_out[1091];
    assign layer4_out[476] = ~layer3_out[3076];
    assign layer4_out[477] = layer3_out[204] & ~layer3_out[203];
    assign layer4_out[478] = ~layer3_out[628];
    assign layer4_out[479] = ~(layer3_out[207] & layer3_out[208]);
    assign layer4_out[480] = layer3_out[6197] & ~layer3_out[6196];
    assign layer4_out[481] = layer3_out[4648];
    assign layer4_out[482] = ~layer3_out[1393] | layer3_out[1392];
    assign layer4_out[483] = ~(layer3_out[5427] | layer3_out[5428]);
    assign layer4_out[484] = layer3_out[4169] & ~layer3_out[4170];
    assign layer4_out[485] = ~layer3_out[5467] | layer3_out[5468];
    assign layer4_out[486] = layer3_out[1112];
    assign layer4_out[487] = ~(layer3_out[7885] ^ layer3_out[7886]);
    assign layer4_out[488] = ~layer3_out[7942];
    assign layer4_out[489] = ~layer3_out[422] | layer3_out[421];
    assign layer4_out[490] = layer3_out[6185] & ~layer3_out[6184];
    assign layer4_out[491] = ~layer3_out[4599] | layer3_out[4600];
    assign layer4_out[492] = layer3_out[7074];
    assign layer4_out[493] = layer3_out[1411];
    assign layer4_out[494] = 1'b0;
    assign layer4_out[495] = layer3_out[5291];
    assign layer4_out[496] = layer3_out[3859];
    assign layer4_out[497] = layer3_out[5216] & layer3_out[5217];
    assign layer4_out[498] = layer3_out[4683] & ~layer3_out[4684];
    assign layer4_out[499] = layer3_out[5856] ^ layer3_out[5857];
    assign layer4_out[500] = layer3_out[6774];
    assign layer4_out[501] = layer3_out[5655];
    assign layer4_out[502] = ~layer3_out[223] | layer3_out[224];
    assign layer4_out[503] = ~layer3_out[6471];
    assign layer4_out[504] = 1'b0;
    assign layer4_out[505] = layer3_out[4986] ^ layer3_out[4987];
    assign layer4_out[506] = ~(layer3_out[7021] ^ layer3_out[7022]);
    assign layer4_out[507] = layer3_out[3869];
    assign layer4_out[508] = ~(layer3_out[3001] & layer3_out[3002]);
    assign layer4_out[509] = ~layer3_out[6841] | layer3_out[6842];
    assign layer4_out[510] = ~layer3_out[4506];
    assign layer4_out[511] = ~layer3_out[5663] | layer3_out[5664];
    assign layer4_out[512] = layer3_out[4179] & layer3_out[4180];
    assign layer4_out[513] = ~(layer3_out[6130] & layer3_out[6131]);
    assign layer4_out[514] = ~layer3_out[1719] | layer3_out[1720];
    assign layer4_out[515] = ~layer3_out[5607];
    assign layer4_out[516] = layer3_out[2056];
    assign layer4_out[517] = layer3_out[6523] ^ layer3_out[6524];
    assign layer4_out[518] = layer3_out[2784] ^ layer3_out[2785];
    assign layer4_out[519] = ~layer3_out[4574] | layer3_out[4575];
    assign layer4_out[520] = layer3_out[5925];
    assign layer4_out[521] = layer3_out[5666] ^ layer3_out[5667];
    assign layer4_out[522] = ~(layer3_out[924] | layer3_out[925]);
    assign layer4_out[523] = layer3_out[6518];
    assign layer4_out[524] = ~layer3_out[7506];
    assign layer4_out[525] = layer3_out[7477];
    assign layer4_out[526] = ~layer3_out[5457];
    assign layer4_out[527] = ~layer3_out[841] | layer3_out[842];
    assign layer4_out[528] = ~layer3_out[743];
    assign layer4_out[529] = ~layer3_out[1413];
    assign layer4_out[530] = ~(layer3_out[4412] ^ layer3_out[4413]);
    assign layer4_out[531] = layer3_out[1903];
    assign layer4_out[532] = ~layer3_out[3326];
    assign layer4_out[533] = layer3_out[4450];
    assign layer4_out[534] = ~(layer3_out[4359] ^ layer3_out[4360]);
    assign layer4_out[535] = layer3_out[6443];
    assign layer4_out[536] = ~layer3_out[5103];
    assign layer4_out[537] = ~(layer3_out[1347] & layer3_out[1348]);
    assign layer4_out[538] = layer3_out[807] ^ layer3_out[808];
    assign layer4_out[539] = ~layer3_out[176] | layer3_out[177];
    assign layer4_out[540] = ~(layer3_out[6975] ^ layer3_out[6976]);
    assign layer4_out[541] = layer3_out[2787] & ~layer3_out[2786];
    assign layer4_out[542] = layer3_out[5165] & ~layer3_out[5164];
    assign layer4_out[543] = ~layer3_out[5628];
    assign layer4_out[544] = ~layer3_out[6355];
    assign layer4_out[545] = ~layer3_out[3680];
    assign layer4_out[546] = ~(layer3_out[956] & layer3_out[957]);
    assign layer4_out[547] = ~(layer3_out[4391] ^ layer3_out[4392]);
    assign layer4_out[548] = layer3_out[142];
    assign layer4_out[549] = ~layer3_out[6985] | layer3_out[6986];
    assign layer4_out[550] = ~(layer3_out[912] ^ layer3_out[913]);
    assign layer4_out[551] = layer3_out[3008];
    assign layer4_out[552] = ~layer3_out[6351];
    assign layer4_out[553] = ~layer3_out[2816];
    assign layer4_out[554] = layer3_out[7269] & layer3_out[7270];
    assign layer4_out[555] = ~(layer3_out[610] | layer3_out[611]);
    assign layer4_out[556] = layer3_out[6234];
    assign layer4_out[557] = layer3_out[3034];
    assign layer4_out[558] = ~(layer3_out[6411] ^ layer3_out[6412]);
    assign layer4_out[559] = ~layer3_out[1220] | layer3_out[1219];
    assign layer4_out[560] = layer3_out[5453];
    assign layer4_out[561] = layer3_out[6186] | layer3_out[6187];
    assign layer4_out[562] = ~layer3_out[3295];
    assign layer4_out[563] = layer3_out[5329] & ~layer3_out[5330];
    assign layer4_out[564] = ~(layer3_out[1728] ^ layer3_out[1729]);
    assign layer4_out[565] = ~(layer3_out[5916] | layer3_out[5917]);
    assign layer4_out[566] = ~layer3_out[4754] | layer3_out[4753];
    assign layer4_out[567] = ~layer3_out[3321];
    assign layer4_out[568] = ~(layer3_out[5617] | layer3_out[5618]);
    assign layer4_out[569] = ~layer3_out[960];
    assign layer4_out[570] = layer3_out[2369] & ~layer3_out[2368];
    assign layer4_out[571] = layer3_out[5608] ^ layer3_out[5609];
    assign layer4_out[572] = ~(layer3_out[873] ^ layer3_out[874]);
    assign layer4_out[573] = layer3_out[2609] ^ layer3_out[2610];
    assign layer4_out[574] = layer3_out[4103] ^ layer3_out[4104];
    assign layer4_out[575] = ~(layer3_out[2360] ^ layer3_out[2361]);
    assign layer4_out[576] = layer3_out[6374];
    assign layer4_out[577] = 1'b0;
    assign layer4_out[578] = ~(layer3_out[3892] | layer3_out[3893]);
    assign layer4_out[579] = ~layer3_out[6790];
    assign layer4_out[580] = ~layer3_out[2981];
    assign layer4_out[581] = ~layer3_out[6216];
    assign layer4_out[582] = layer3_out[7934] ^ layer3_out[7935];
    assign layer4_out[583] = ~layer3_out[1998];
    assign layer4_out[584] = ~(layer3_out[7694] | layer3_out[7695]);
    assign layer4_out[585] = layer3_out[2134];
    assign layer4_out[586] = ~layer3_out[3793];
    assign layer4_out[587] = ~layer3_out[3274] | layer3_out[3275];
    assign layer4_out[588] = layer3_out[3054] & ~layer3_out[3053];
    assign layer4_out[589] = layer3_out[1433] ^ layer3_out[1434];
    assign layer4_out[590] = layer3_out[4442];
    assign layer4_out[591] = layer3_out[3028] & layer3_out[3029];
    assign layer4_out[592] = ~layer3_out[3806];
    assign layer4_out[593] = layer3_out[7068] | layer3_out[7069];
    assign layer4_out[594] = layer3_out[5205] ^ layer3_out[5206];
    assign layer4_out[595] = layer3_out[4730] & ~layer3_out[4731];
    assign layer4_out[596] = ~layer3_out[6859] | layer3_out[6858];
    assign layer4_out[597] = ~(layer3_out[7728] ^ layer3_out[7729]);
    assign layer4_out[598] = ~(layer3_out[458] | layer3_out[459]);
    assign layer4_out[599] = ~(layer3_out[7836] | layer3_out[7837]);
    assign layer4_out[600] = ~layer3_out[1634] | layer3_out[1635];
    assign layer4_out[601] = ~layer3_out[2493];
    assign layer4_out[602] = ~(layer3_out[360] ^ layer3_out[361]);
    assign layer4_out[603] = 1'b1;
    assign layer4_out[604] = layer3_out[7409] ^ layer3_out[7410];
    assign layer4_out[605] = ~layer3_out[3640];
    assign layer4_out[606] = ~layer3_out[7729];
    assign layer4_out[607] = layer3_out[6936] & ~layer3_out[6935];
    assign layer4_out[608] = layer3_out[5495] ^ layer3_out[5496];
    assign layer4_out[609] = layer3_out[6749];
    assign layer4_out[610] = layer3_out[7961];
    assign layer4_out[611] = layer3_out[5962];
    assign layer4_out[612] = ~layer3_out[3495];
    assign layer4_out[613] = layer3_out[4848];
    assign layer4_out[614] = ~(layer3_out[381] ^ layer3_out[382]);
    assign layer4_out[615] = ~layer3_out[6816] | layer3_out[6817];
    assign layer4_out[616] = layer3_out[5840];
    assign layer4_out[617] = ~(layer3_out[4588] ^ layer3_out[4589]);
    assign layer4_out[618] = layer3_out[4947];
    assign layer4_out[619] = ~layer3_out[5948];
    assign layer4_out[620] = ~(layer3_out[3345] | layer3_out[3346]);
    assign layer4_out[621] = ~layer3_out[958] | layer3_out[959];
    assign layer4_out[622] = layer3_out[2344];
    assign layer4_out[623] = ~(layer3_out[1122] | layer3_out[1123]);
    assign layer4_out[624] = ~layer3_out[7049];
    assign layer4_out[625] = 1'b1;
    assign layer4_out[626] = ~layer3_out[5517] | layer3_out[5516];
    assign layer4_out[627] = layer3_out[570] & ~layer3_out[571];
    assign layer4_out[628] = layer3_out[6855] ^ layer3_out[6856];
    assign layer4_out[629] = ~layer3_out[6912];
    assign layer4_out[630] = layer3_out[3911];
    assign layer4_out[631] = layer3_out[177] ^ layer3_out[178];
    assign layer4_out[632] = ~(layer3_out[1367] | layer3_out[1368]);
    assign layer4_out[633] = ~(layer3_out[931] & layer3_out[932]);
    assign layer4_out[634] = layer3_out[4990];
    assign layer4_out[635] = layer3_out[6806] ^ layer3_out[6807];
    assign layer4_out[636] = layer3_out[1847];
    assign layer4_out[637] = ~layer3_out[1404] | layer3_out[1403];
    assign layer4_out[638] = layer3_out[6880];
    assign layer4_out[639] = ~(layer3_out[4610] & layer3_out[4611]);
    assign layer4_out[640] = layer3_out[7433] | layer3_out[7434];
    assign layer4_out[641] = ~(layer3_out[1133] & layer3_out[1134]);
    assign layer4_out[642] = layer3_out[7397] & layer3_out[7398];
    assign layer4_out[643] = layer3_out[1904];
    assign layer4_out[644] = ~(layer3_out[4078] ^ layer3_out[4079]);
    assign layer4_out[645] = ~layer3_out[7035] | layer3_out[7036];
    assign layer4_out[646] = layer3_out[5777];
    assign layer4_out[647] = ~(layer3_out[4868] ^ layer3_out[4869]);
    assign layer4_out[648] = ~(layer3_out[4795] | layer3_out[4796]);
    assign layer4_out[649] = ~layer3_out[1774];
    assign layer4_out[650] = layer3_out[2146] & layer3_out[2147];
    assign layer4_out[651] = layer3_out[4097];
    assign layer4_out[652] = layer3_out[1031];
    assign layer4_out[653] = ~layer3_out[2978];
    assign layer4_out[654] = layer3_out[5237];
    assign layer4_out[655] = ~layer3_out[2156];
    assign layer4_out[656] = ~(layer3_out[5504] | layer3_out[5505]);
    assign layer4_out[657] = layer3_out[4845] & ~layer3_out[4846];
    assign layer4_out[658] = layer3_out[2100] & ~layer3_out[2101];
    assign layer4_out[659] = ~layer3_out[5002] | layer3_out[5003];
    assign layer4_out[660] = ~(layer3_out[7641] ^ layer3_out[7642]);
    assign layer4_out[661] = layer3_out[1844] & ~layer3_out[1843];
    assign layer4_out[662] = layer3_out[1109] ^ layer3_out[1110];
    assign layer4_out[663] = layer3_out[3739] ^ layer3_out[3740];
    assign layer4_out[664] = layer3_out[6299] | layer3_out[6300];
    assign layer4_out[665] = layer3_out[1770] | layer3_out[1771];
    assign layer4_out[666] = layer3_out[345];
    assign layer4_out[667] = layer3_out[6462] ^ layer3_out[6463];
    assign layer4_out[668] = ~layer3_out[4561];
    assign layer4_out[669] = layer3_out[5291];
    assign layer4_out[670] = ~(layer3_out[3963] ^ layer3_out[3964]);
    assign layer4_out[671] = layer3_out[6091] & layer3_out[6092];
    assign layer4_out[672] = layer3_out[3094];
    assign layer4_out[673] = layer3_out[1725] ^ layer3_out[1726];
    assign layer4_out[674] = 1'b0;
    assign layer4_out[675] = layer3_out[784] & layer3_out[785];
    assign layer4_out[676] = layer3_out[3645];
    assign layer4_out[677] = layer3_out[7380] ^ layer3_out[7381];
    assign layer4_out[678] = ~layer3_out[6632] | layer3_out[6631];
    assign layer4_out[679] = ~layer3_out[689];
    assign layer4_out[680] = layer3_out[2526] & ~layer3_out[2525];
    assign layer4_out[681] = ~layer3_out[2852];
    assign layer4_out[682] = ~layer3_out[2239];
    assign layer4_out[683] = layer3_out[1472] ^ layer3_out[1473];
    assign layer4_out[684] = layer3_out[2415];
    assign layer4_out[685] = ~layer3_out[5415];
    assign layer4_out[686] = layer3_out[2278] & layer3_out[2279];
    assign layer4_out[687] = ~(layer3_out[1668] ^ layer3_out[1669]);
    assign layer4_out[688] = layer3_out[7507] | layer3_out[7508];
    assign layer4_out[689] = layer3_out[7029];
    assign layer4_out[690] = ~layer3_out[448];
    assign layer4_out[691] = layer3_out[1310] & ~layer3_out[1311];
    assign layer4_out[692] = ~layer3_out[2374];
    assign layer4_out[693] = layer3_out[2034] & ~layer3_out[2033];
    assign layer4_out[694] = layer3_out[7263];
    assign layer4_out[695] = ~layer3_out[4031];
    assign layer4_out[696] = ~layer3_out[3824];
    assign layer4_out[697] = ~(layer3_out[7435] ^ layer3_out[7436]);
    assign layer4_out[698] = ~(layer3_out[6419] | layer3_out[6420]);
    assign layer4_out[699] = layer3_out[6508] | layer3_out[6509];
    assign layer4_out[700] = layer3_out[7066];
    assign layer4_out[701] = ~layer3_out[7399] | layer3_out[7398];
    assign layer4_out[702] = layer3_out[3439] & layer3_out[3440];
    assign layer4_out[703] = layer3_out[6865];
    assign layer4_out[704] = layer3_out[7557];
    assign layer4_out[705] = ~layer3_out[7913] | layer3_out[7912];
    assign layer4_out[706] = layer3_out[7031] & ~layer3_out[7032];
    assign layer4_out[707] = ~(layer3_out[2084] | layer3_out[2085]);
    assign layer4_out[708] = layer3_out[1743] & ~layer3_out[1744];
    assign layer4_out[709] = ~layer3_out[5132];
    assign layer4_out[710] = layer3_out[2282] & ~layer3_out[2283];
    assign layer4_out[711] = ~layer3_out[419] | layer3_out[420];
    assign layer4_out[712] = layer3_out[1005] | layer3_out[1006];
    assign layer4_out[713] = ~layer3_out[4394];
    assign layer4_out[714] = layer3_out[4288] & ~layer3_out[4287];
    assign layer4_out[715] = layer3_out[2876];
    assign layer4_out[716] = ~layer3_out[4825] | layer3_out[4826];
    assign layer4_out[717] = layer3_out[6617] & layer3_out[6618];
    assign layer4_out[718] = ~layer3_out[5616];
    assign layer4_out[719] = layer3_out[4416] & layer3_out[4417];
    assign layer4_out[720] = layer3_out[5181];
    assign layer4_out[721] = layer3_out[3840];
    assign layer4_out[722] = ~layer3_out[460] | layer3_out[459];
    assign layer4_out[723] = ~(layer3_out[1832] ^ layer3_out[1833]);
    assign layer4_out[724] = layer3_out[4085] ^ layer3_out[4086];
    assign layer4_out[725] = ~layer3_out[1900];
    assign layer4_out[726] = layer3_out[1206];
    assign layer4_out[727] = ~layer3_out[5238] | layer3_out[5237];
    assign layer4_out[728] = layer3_out[3182] | layer3_out[3183];
    assign layer4_out[729] = ~layer3_out[68];
    assign layer4_out[730] = layer3_out[7010];
    assign layer4_out[731] = ~layer3_out[4928];
    assign layer4_out[732] = ~(layer3_out[6251] | layer3_out[6252]);
    assign layer4_out[733] = ~layer3_out[6455] | layer3_out[6454];
    assign layer4_out[734] = layer3_out[7134] & layer3_out[7135];
    assign layer4_out[735] = ~layer3_out[6161];
    assign layer4_out[736] = layer3_out[4680] ^ layer3_out[4681];
    assign layer4_out[737] = layer3_out[3855];
    assign layer4_out[738] = layer3_out[4966] ^ layer3_out[4967];
    assign layer4_out[739] = layer3_out[7508] ^ layer3_out[7509];
    assign layer4_out[740] = layer3_out[5989];
    assign layer4_out[741] = layer3_out[738] & layer3_out[739];
    assign layer4_out[742] = ~layer3_out[3526];
    assign layer4_out[743] = ~(layer3_out[7350] | layer3_out[7351]);
    assign layer4_out[744] = layer3_out[2268];
    assign layer4_out[745] = layer3_out[3966];
    assign layer4_out[746] = layer3_out[5117] & layer3_out[5118];
    assign layer4_out[747] = layer3_out[4910] ^ layer3_out[4911];
    assign layer4_out[748] = layer3_out[4806];
    assign layer4_out[749] = layer3_out[5588] & ~layer3_out[5589];
    assign layer4_out[750] = ~layer3_out[7231];
    assign layer4_out[751] = ~layer3_out[5689] | layer3_out[5688];
    assign layer4_out[752] = ~layer3_out[3882];
    assign layer4_out[753] = layer3_out[778];
    assign layer4_out[754] = ~layer3_out[683] | layer3_out[684];
    assign layer4_out[755] = layer3_out[4529];
    assign layer4_out[756] = layer3_out[6074] & ~layer3_out[6075];
    assign layer4_out[757] = layer3_out[2515] | layer3_out[2516];
    assign layer4_out[758] = ~layer3_out[398] | layer3_out[397];
    assign layer4_out[759] = layer3_out[4622] ^ layer3_out[4623];
    assign layer4_out[760] = ~layer3_out[7147] | layer3_out[7148];
    assign layer4_out[761] = layer3_out[915] & layer3_out[916];
    assign layer4_out[762] = layer3_out[1793] & ~layer3_out[1792];
    assign layer4_out[763] = layer3_out[7315] & layer3_out[7316];
    assign layer4_out[764] = layer3_out[3620];
    assign layer4_out[765] = layer3_out[7491] & ~layer3_out[7492];
    assign layer4_out[766] = ~layer3_out[1867] | layer3_out[1866];
    assign layer4_out[767] = layer3_out[3960];
    assign layer4_out[768] = layer3_out[2359] ^ layer3_out[2360];
    assign layer4_out[769] = layer3_out[6786];
    assign layer4_out[770] = ~layer3_out[287];
    assign layer4_out[771] = ~layer3_out[7966] | layer3_out[7967];
    assign layer4_out[772] = layer3_out[1230];
    assign layer4_out[773] = ~(layer3_out[2889] | layer3_out[2890]);
    assign layer4_out[774] = ~layer3_out[4932];
    assign layer4_out[775] = ~(layer3_out[7149] ^ layer3_out[7150]);
    assign layer4_out[776] = ~layer3_out[2126];
    assign layer4_out[777] = ~layer3_out[7571];
    assign layer4_out[778] = layer3_out[338] & layer3_out[339];
    assign layer4_out[779] = ~(layer3_out[6601] ^ layer3_out[6602]);
    assign layer4_out[780] = layer3_out[4250] & layer3_out[4251];
    assign layer4_out[781] = layer3_out[5612];
    assign layer4_out[782] = ~layer3_out[851];
    assign layer4_out[783] = layer3_out[5072] & ~layer3_out[5071];
    assign layer4_out[784] = layer3_out[6216] & layer3_out[6217];
    assign layer4_out[785] = layer3_out[7383] & layer3_out[7384];
    assign layer4_out[786] = layer3_out[6376] & ~layer3_out[6375];
    assign layer4_out[787] = ~layer3_out[6714];
    assign layer4_out[788] = ~(layer3_out[2932] & layer3_out[2933]);
    assign layer4_out[789] = ~layer3_out[6075];
    assign layer4_out[790] = ~layer3_out[7582];
    assign layer4_out[791] = layer3_out[68];
    assign layer4_out[792] = layer3_out[7566] & ~layer3_out[7565];
    assign layer4_out[793] = layer3_out[5194] & ~layer3_out[5195];
    assign layer4_out[794] = layer3_out[4106];
    assign layer4_out[795] = ~layer3_out[3836] | layer3_out[3835];
    assign layer4_out[796] = ~layer3_out[2942] | layer3_out[2941];
    assign layer4_out[797] = ~layer3_out[2354];
    assign layer4_out[798] = layer3_out[2464];
    assign layer4_out[799] = layer3_out[6699];
    assign layer4_out[800] = ~(layer3_out[4044] ^ layer3_out[4045]);
    assign layer4_out[801] = ~layer3_out[5034] | layer3_out[5033];
    assign layer4_out[802] = ~(layer3_out[2204] ^ layer3_out[2205]);
    assign layer4_out[803] = ~layer3_out[3757] | layer3_out[3758];
    assign layer4_out[804] = layer3_out[5056];
    assign layer4_out[805] = ~(layer3_out[5475] ^ layer3_out[5476]);
    assign layer4_out[806] = layer3_out[1891] ^ layer3_out[1892];
    assign layer4_out[807] = ~layer3_out[2023] | layer3_out[2022];
    assign layer4_out[808] = layer3_out[6122];
    assign layer4_out[809] = layer3_out[6486];
    assign layer4_out[810] = layer3_out[7087] ^ layer3_out[7088];
    assign layer4_out[811] = ~(layer3_out[1484] ^ layer3_out[1485]);
    assign layer4_out[812] = ~layer3_out[3428];
    assign layer4_out[813] = layer3_out[6352];
    assign layer4_out[814] = layer3_out[2851] & ~layer3_out[2850];
    assign layer4_out[815] = layer3_out[2904] ^ layer3_out[2905];
    assign layer4_out[816] = ~layer3_out[7210] | layer3_out[7211];
    assign layer4_out[817] = layer3_out[887] ^ layer3_out[888];
    assign layer4_out[818] = layer3_out[2255] & ~layer3_out[2254];
    assign layer4_out[819] = layer3_out[7410] | layer3_out[7411];
    assign layer4_out[820] = ~layer3_out[6142];
    assign layer4_out[821] = ~(layer3_out[3765] | layer3_out[3766]);
    assign layer4_out[822] = ~layer3_out[3489];
    assign layer4_out[823] = layer3_out[4692] & ~layer3_out[4693];
    assign layer4_out[824] = layer3_out[706] & layer3_out[707];
    assign layer4_out[825] = ~(layer3_out[1756] | layer3_out[1757]);
    assign layer4_out[826] = 1'b0;
    assign layer4_out[827] = ~(layer3_out[2714] | layer3_out[2715]);
    assign layer4_out[828] = layer3_out[3808];
    assign layer4_out[829] = ~layer3_out[6363];
    assign layer4_out[830] = ~(layer3_out[639] ^ layer3_out[640]);
    assign layer4_out[831] = ~layer3_out[808];
    assign layer4_out[832] = layer3_out[5869] ^ layer3_out[5870];
    assign layer4_out[833] = ~layer3_out[2936];
    assign layer4_out[834] = layer3_out[7973];
    assign layer4_out[835] = layer3_out[7235];
    assign layer4_out[836] = layer3_out[1];
    assign layer4_out[837] = ~layer3_out[492];
    assign layer4_out[838] = layer3_out[3699];
    assign layer4_out[839] = ~layer3_out[5175];
    assign layer4_out[840] = layer3_out[60] & layer3_out[61];
    assign layer4_out[841] = layer3_out[1625];
    assign layer4_out[842] = ~(layer3_out[855] | layer3_out[856]);
    assign layer4_out[843] = layer3_out[1487] & ~layer3_out[1486];
    assign layer4_out[844] = layer3_out[2668];
    assign layer4_out[845] = layer3_out[6169] | layer3_out[6170];
    assign layer4_out[846] = ~layer3_out[7218];
    assign layer4_out[847] = ~layer3_out[4432] | layer3_out[4431];
    assign layer4_out[848] = layer3_out[352];
    assign layer4_out[849] = layer3_out[3323];
    assign layer4_out[850] = layer3_out[1302] ^ layer3_out[1303];
    assign layer4_out[851] = ~(layer3_out[2276] ^ layer3_out[2277]);
    assign layer4_out[852] = layer3_out[2886] | layer3_out[2887];
    assign layer4_out[853] = layer3_out[8];
    assign layer4_out[854] = ~layer3_out[3453];
    assign layer4_out[855] = ~(layer3_out[0] ^ layer3_out[2]);
    assign layer4_out[856] = layer3_out[1105] | layer3_out[1106];
    assign layer4_out[857] = layer3_out[2753];
    assign layer4_out[858] = layer3_out[4068];
    assign layer4_out[859] = ~layer3_out[5634];
    assign layer4_out[860] = ~(layer3_out[2419] & layer3_out[2420]);
    assign layer4_out[861] = layer3_out[7746] | layer3_out[7747];
    assign layer4_out[862] = ~layer3_out[7324];
    assign layer4_out[863] = ~layer3_out[447];
    assign layer4_out[864] = layer3_out[6624];
    assign layer4_out[865] = layer3_out[6612];
    assign layer4_out[866] = layer3_out[6955] & ~layer3_out[6954];
    assign layer4_out[867] = layer3_out[1567] ^ layer3_out[1568];
    assign layer4_out[868] = ~(layer3_out[5829] ^ layer3_out[5830]);
    assign layer4_out[869] = ~layer3_out[6567] | layer3_out[6568];
    assign layer4_out[870] = ~(layer3_out[5351] & layer3_out[5352]);
    assign layer4_out[871] = layer3_out[5882] & ~layer3_out[5883];
    assign layer4_out[872] = layer3_out[4613];
    assign layer4_out[873] = layer3_out[6928];
    assign layer4_out[874] = layer3_out[1966];
    assign layer4_out[875] = layer3_out[6380];
    assign layer4_out[876] = layer3_out[1464] & ~layer3_out[1465];
    assign layer4_out[877] = layer3_out[1512];
    assign layer4_out[878] = layer3_out[5038];
    assign layer4_out[879] = ~layer3_out[512] | layer3_out[513];
    assign layer4_out[880] = ~layer3_out[2698];
    assign layer4_out[881] = ~(layer3_out[6356] ^ layer3_out[6357]);
    assign layer4_out[882] = ~layer3_out[3034];
    assign layer4_out[883] = layer3_out[7530];
    assign layer4_out[884] = ~(layer3_out[701] | layer3_out[702]);
    assign layer4_out[885] = layer3_out[6446];
    assign layer4_out[886] = ~(layer3_out[4092] ^ layer3_out[4093]);
    assign layer4_out[887] = layer3_out[1028] & ~layer3_out[1029];
    assign layer4_out[888] = layer3_out[6867] ^ layer3_out[6868];
    assign layer4_out[889] = layer3_out[7839];
    assign layer4_out[890] = layer3_out[6052];
    assign layer4_out[891] = ~layer3_out[4011];
    assign layer4_out[892] = layer3_out[1506];
    assign layer4_out[893] = ~layer3_out[3635] | layer3_out[3636];
    assign layer4_out[894] = layer3_out[6674];
    assign layer4_out[895] = ~layer3_out[2131];
    assign layer4_out[896] = ~layer3_out[2301];
    assign layer4_out[897] = ~layer3_out[5226];
    assign layer4_out[898] = ~layer3_out[1380];
    assign layer4_out[899] = ~(layer3_out[3402] | layer3_out[3403]);
    assign layer4_out[900] = layer3_out[3220];
    assign layer4_out[901] = ~(layer3_out[7514] ^ layer3_out[7515]);
    assign layer4_out[902] = layer3_out[264] & ~layer3_out[265];
    assign layer4_out[903] = layer3_out[1827];
    assign layer4_out[904] = layer3_out[3918] & ~layer3_out[3919];
    assign layer4_out[905] = ~(layer3_out[4578] | layer3_out[4579]);
    assign layer4_out[906] = ~(layer3_out[821] | layer3_out[822]);
    assign layer4_out[907] = ~(layer3_out[1838] | layer3_out[1839]);
    assign layer4_out[908] = layer3_out[4110];
    assign layer4_out[909] = layer3_out[3212] ^ layer3_out[3213];
    assign layer4_out[910] = ~layer3_out[3530];
    assign layer4_out[911] = ~layer3_out[7620];
    assign layer4_out[912] = layer3_out[6163];
    assign layer4_out[913] = ~layer3_out[3145];
    assign layer4_out[914] = ~layer3_out[6994];
    assign layer4_out[915] = ~layer3_out[5537];
    assign layer4_out[916] = layer3_out[7679];
    assign layer4_out[917] = ~layer3_out[877];
    assign layer4_out[918] = ~layer3_out[3024] | layer3_out[3025];
    assign layer4_out[919] = ~layer3_out[4876];
    assign layer4_out[920] = layer3_out[121];
    assign layer4_out[921] = ~layer3_out[3792];
    assign layer4_out[922] = ~(layer3_out[6410] | layer3_out[6411]);
    assign layer4_out[923] = layer3_out[7684] | layer3_out[7685];
    assign layer4_out[924] = layer3_out[3781] & layer3_out[3782];
    assign layer4_out[925] = layer3_out[2514];
    assign layer4_out[926] = ~(layer3_out[2436] & layer3_out[2437]);
    assign layer4_out[927] = ~(layer3_out[4822] ^ layer3_out[4823]);
    assign layer4_out[928] = layer3_out[4526] ^ layer3_out[4527];
    assign layer4_out[929] = ~layer3_out[6843];
    assign layer4_out[930] = layer3_out[4368] | layer3_out[4369];
    assign layer4_out[931] = ~layer3_out[6378];
    assign layer4_out[932] = ~layer3_out[3282];
    assign layer4_out[933] = layer3_out[7232] & ~layer3_out[7231];
    assign layer4_out[934] = layer3_out[4818] | layer3_out[4819];
    assign layer4_out[935] = layer3_out[6872] ^ layer3_out[6873];
    assign layer4_out[936] = layer3_out[5953];
    assign layer4_out[937] = layer3_out[2047] & ~layer3_out[2048];
    assign layer4_out[938] = layer3_out[6179] | layer3_out[6180];
    assign layer4_out[939] = layer3_out[3970] | layer3_out[3971];
    assign layer4_out[940] = layer3_out[7490];
    assign layer4_out[941] = ~layer3_out[4077] | layer3_out[4078];
    assign layer4_out[942] = ~layer3_out[1013];
    assign layer4_out[943] = ~layer3_out[370];
    assign layer4_out[944] = layer3_out[5905] | layer3_out[5906];
    assign layer4_out[945] = ~layer3_out[1090];
    assign layer4_out[946] = layer3_out[2838] & ~layer3_out[2837];
    assign layer4_out[947] = ~(layer3_out[3088] & layer3_out[3089]);
    assign layer4_out[948] = ~layer3_out[2027] | layer3_out[2026];
    assign layer4_out[949] = ~layer3_out[422];
    assign layer4_out[950] = ~layer3_out[2624];
    assign layer4_out[951] = ~layer3_out[5289];
    assign layer4_out[952] = ~layer3_out[5424] | layer3_out[5423];
    assign layer4_out[953] = layer3_out[5569] ^ layer3_out[5570];
    assign layer4_out[954] = layer3_out[7440] | layer3_out[7441];
    assign layer4_out[955] = ~layer3_out[4299];
    assign layer4_out[956] = layer3_out[1082] ^ layer3_out[1083];
    assign layer4_out[957] = layer3_out[870] ^ layer3_out[871];
    assign layer4_out[958] = ~layer3_out[2250];
    assign layer4_out[959] = layer3_out[7246] & ~layer3_out[7247];
    assign layer4_out[960] = layer3_out[4445] ^ layer3_out[4446];
    assign layer4_out[961] = ~(layer3_out[276] & layer3_out[277]);
    assign layer4_out[962] = ~layer3_out[6497];
    assign layer4_out[963] = layer3_out[564] ^ layer3_out[565];
    assign layer4_out[964] = layer3_out[3674] & ~layer3_out[3675];
    assign layer4_out[965] = layer3_out[1728];
    assign layer4_out[966] = ~layer3_out[3920];
    assign layer4_out[967] = ~(layer3_out[4773] ^ layer3_out[4774]);
    assign layer4_out[968] = layer3_out[3718];
    assign layer4_out[969] = ~(layer3_out[3512] & layer3_out[3513]);
    assign layer4_out[970] = ~(layer3_out[4665] ^ layer3_out[4666]);
    assign layer4_out[971] = layer3_out[5964];
    assign layer4_out[972] = ~layer3_out[5853];
    assign layer4_out[973] = ~(layer3_out[3728] & layer3_out[3729]);
    assign layer4_out[974] = layer3_out[1874] & ~layer3_out[1875];
    assign layer4_out[975] = ~layer3_out[6017];
    assign layer4_out[976] = layer3_out[6533] | layer3_out[6534];
    assign layer4_out[977] = layer3_out[249];
    assign layer4_out[978] = layer3_out[5293] | layer3_out[5294];
    assign layer4_out[979] = layer3_out[2855] & ~layer3_out[2854];
    assign layer4_out[980] = layer3_out[1246] ^ layer3_out[1247];
    assign layer4_out[981] = ~layer3_out[1915];
    assign layer4_out[982] = layer3_out[749] & ~layer3_out[748];
    assign layer4_out[983] = layer3_out[334] & ~layer3_out[335];
    assign layer4_out[984] = ~layer3_out[5668];
    assign layer4_out[985] = ~layer3_out[6476];
    assign layer4_out[986] = ~(layer3_out[3880] & layer3_out[3881]);
    assign layer4_out[987] = ~layer3_out[1406] | layer3_out[1405];
    assign layer4_out[988] = layer3_out[2252] & layer3_out[2253];
    assign layer4_out[989] = ~(layer3_out[3243] & layer3_out[3244]);
    assign layer4_out[990] = layer3_out[6798];
    assign layer4_out[991] = ~layer3_out[2404] | layer3_out[2405];
    assign layer4_out[992] = layer3_out[4792];
    assign layer4_out[993] = ~layer3_out[4539] | layer3_out[4538];
    assign layer4_out[994] = ~layer3_out[3236];
    assign layer4_out[995] = ~(layer3_out[5085] ^ layer3_out[5086]);
    assign layer4_out[996] = layer3_out[7207] & layer3_out[7208];
    assign layer4_out[997] = ~layer3_out[5422] | layer3_out[5421];
    assign layer4_out[998] = layer3_out[1049] | layer3_out[1050];
    assign layer4_out[999] = ~layer3_out[3547] | layer3_out[3546];
    assign layer4_out[1000] = layer3_out[2292];
    assign layer4_out[1001] = layer3_out[148] & ~layer3_out[147];
    assign layer4_out[1002] = ~layer3_out[1830];
    assign layer4_out[1003] = ~layer3_out[6118];
    assign layer4_out[1004] = ~layer3_out[2261];
    assign layer4_out[1005] = layer3_out[4586] & ~layer3_out[4587];
    assign layer4_out[1006] = layer3_out[5168] ^ layer3_out[5169];
    assign layer4_out[1007] = layer3_out[3462] | layer3_out[3463];
    assign layer4_out[1008] = layer3_out[6922];
    assign layer4_out[1009] = ~(layer3_out[5899] | layer3_out[5900]);
    assign layer4_out[1010] = layer3_out[582];
    assign layer4_out[1011] = layer3_out[6913];
    assign layer4_out[1012] = ~layer3_out[7203];
    assign layer4_out[1013] = ~layer3_out[5655];
    assign layer4_out[1014] = ~layer3_out[7706] | layer3_out[7707];
    assign layer4_out[1015] = layer3_out[5167] ^ layer3_out[5168];
    assign layer4_out[1016] = layer3_out[6226];
    assign layer4_out[1017] = layer3_out[6805];
    assign layer4_out[1018] = layer3_out[652];
    assign layer4_out[1019] = ~layer3_out[6977];
    assign layer4_out[1020] = ~(layer3_out[5702] ^ layer3_out[5703]);
    assign layer4_out[1021] = layer3_out[433] ^ layer3_out[434];
    assign layer4_out[1022] = layer3_out[3741] ^ layer3_out[3742];
    assign layer4_out[1023] = layer3_out[2502];
    assign layer4_out[1024] = ~layer3_out[4440];
    assign layer4_out[1025] = ~layer3_out[4660];
    assign layer4_out[1026] = layer3_out[5190];
    assign layer4_out[1027] = layer3_out[188] ^ layer3_out[189];
    assign layer4_out[1028] = ~layer3_out[1144];
    assign layer4_out[1029] = layer3_out[2321] & layer3_out[2322];
    assign layer4_out[1030] = ~(layer3_out[7024] ^ layer3_out[7025]);
    assign layer4_out[1031] = layer3_out[815];
    assign layer4_out[1032] = ~(layer3_out[4661] ^ layer3_out[4662]);
    assign layer4_out[1033] = ~layer3_out[2888];
    assign layer4_out[1034] = ~layer3_out[3790];
    assign layer4_out[1035] = ~layer3_out[261];
    assign layer4_out[1036] = ~layer3_out[474];
    assign layer4_out[1037] = layer3_out[6032];
    assign layer4_out[1038] = ~layer3_out[1640] | layer3_out[1641];
    assign layer4_out[1039] = layer3_out[1373];
    assign layer4_out[1040] = ~(layer3_out[3922] ^ layer3_out[3923]);
    assign layer4_out[1041] = ~layer3_out[3993];
    assign layer4_out[1042] = ~layer3_out[2688];
    assign layer4_out[1043] = layer3_out[1033];
    assign layer4_out[1044] = layer3_out[2785];
    assign layer4_out[1045] = ~layer3_out[7810] | layer3_out[7811];
    assign layer4_out[1046] = ~layer3_out[6232];
    assign layer4_out[1047] = ~layer3_out[2355] | layer3_out[2354];
    assign layer4_out[1048] = ~layer3_out[7585] | layer3_out[7586];
    assign layer4_out[1049] = layer3_out[1490] & ~layer3_out[1489];
    assign layer4_out[1050] = ~layer3_out[5769] | layer3_out[5770];
    assign layer4_out[1051] = ~layer3_out[2450];
    assign layer4_out[1052] = layer3_out[1818] & layer3_out[1819];
    assign layer4_out[1053] = ~(layer3_out[387] ^ layer3_out[388]);
    assign layer4_out[1054] = ~layer3_out[2782];
    assign layer4_out[1055] = ~layer3_out[6688];
    assign layer4_out[1056] = ~(layer3_out[336] & layer3_out[337]);
    assign layer4_out[1057] = layer3_out[7438] & layer3_out[7439];
    assign layer4_out[1058] = ~layer3_out[3911];
    assign layer4_out[1059] = layer3_out[5701] & layer3_out[5702];
    assign layer4_out[1060] = ~layer3_out[7771];
    assign layer4_out[1061] = layer3_out[4035] & ~layer3_out[4034];
    assign layer4_out[1062] = layer3_out[2964] & ~layer3_out[2965];
    assign layer4_out[1063] = layer3_out[175] | layer3_out[176];
    assign layer4_out[1064] = ~layer3_out[7217];
    assign layer4_out[1065] = ~(layer3_out[86] & layer3_out[87]);
    assign layer4_out[1066] = layer3_out[4127] & ~layer3_out[4128];
    assign layer4_out[1067] = layer3_out[4184] & layer3_out[4185];
    assign layer4_out[1068] = ~layer3_out[5954];
    assign layer4_out[1069] = layer3_out[6322];
    assign layer4_out[1070] = ~(layer3_out[1061] ^ layer3_out[1062]);
    assign layer4_out[1071] = layer3_out[5357] ^ layer3_out[5358];
    assign layer4_out[1072] = layer3_out[1207];
    assign layer4_out[1073] = ~layer3_out[5719];
    assign layer4_out[1074] = ~layer3_out[1019];
    assign layer4_out[1075] = ~(layer3_out[4516] | layer3_out[4517]);
    assign layer4_out[1076] = ~layer3_out[6370];
    assign layer4_out[1077] = ~layer3_out[4241];
    assign layer4_out[1078] = layer3_out[6305];
    assign layer4_out[1079] = ~layer3_out[6649] | layer3_out[6648];
    assign layer4_out[1080] = layer3_out[1249];
    assign layer4_out[1081] = layer3_out[7996] & ~layer3_out[7997];
    assign layer4_out[1082] = layer3_out[2834] & ~layer3_out[2833];
    assign layer4_out[1083] = layer3_out[5090];
    assign layer4_out[1084] = ~layer3_out[273] | layer3_out[272];
    assign layer4_out[1085] = ~(layer3_out[1638] | layer3_out[1639]);
    assign layer4_out[1086] = ~layer3_out[7146];
    assign layer4_out[1087] = ~(layer3_out[6780] ^ layer3_out[6781]);
    assign layer4_out[1088] = ~layer3_out[4585];
    assign layer4_out[1089] = layer3_out[3458];
    assign layer4_out[1090] = ~layer3_out[7271];
    assign layer4_out[1091] = ~layer3_out[3623];
    assign layer4_out[1092] = 1'b1;
    assign layer4_out[1093] = layer3_out[4498] ^ layer3_out[4499];
    assign layer4_out[1094] = layer3_out[522] & layer3_out[523];
    assign layer4_out[1095] = layer3_out[666] & ~layer3_out[665];
    assign layer4_out[1096] = layer3_out[5886];
    assign layer4_out[1097] = ~(layer3_out[6649] ^ layer3_out[6650]);
    assign layer4_out[1098] = layer3_out[6401] & ~layer3_out[6402];
    assign layer4_out[1099] = ~(layer3_out[7833] ^ layer3_out[7834]);
    assign layer4_out[1100] = ~layer3_out[1046];
    assign layer4_out[1101] = layer3_out[6693] ^ layer3_out[6694];
    assign layer4_out[1102] = ~(layer3_out[4472] ^ layer3_out[4473]);
    assign layer4_out[1103] = layer3_out[6993] | layer3_out[6994];
    assign layer4_out[1104] = ~layer3_out[4625] | layer3_out[4626];
    assign layer4_out[1105] = layer3_out[4253] ^ layer3_out[4254];
    assign layer4_out[1106] = layer3_out[5098] ^ layer3_out[5099];
    assign layer4_out[1107] = layer3_out[1737] & ~layer3_out[1736];
    assign layer4_out[1108] = layer3_out[4403] & ~layer3_out[4404];
    assign layer4_out[1109] = layer3_out[4863] ^ layer3_out[4864];
    assign layer4_out[1110] = ~layer3_out[5031];
    assign layer4_out[1111] = layer3_out[5105];
    assign layer4_out[1112] = ~layer3_out[2863];
    assign layer4_out[1113] = ~(layer3_out[4934] ^ layer3_out[4935]);
    assign layer4_out[1114] = ~(layer3_out[7522] & layer3_out[7523]);
    assign layer4_out[1115] = ~layer3_out[1694];
    assign layer4_out[1116] = layer3_out[4518] & ~layer3_out[4519];
    assign layer4_out[1117] = ~layer3_out[3528] | layer3_out[3529];
    assign layer4_out[1118] = ~(layer3_out[4405] & layer3_out[4406]);
    assign layer4_out[1119] = layer3_out[2291];
    assign layer4_out[1120] = layer3_out[622] | layer3_out[623];
    assign layer4_out[1121] = layer3_out[5778] | layer3_out[5779];
    assign layer4_out[1122] = layer3_out[174] ^ layer3_out[175];
    assign layer4_out[1123] = layer3_out[437] | layer3_out[438];
    assign layer4_out[1124] = layer3_out[6708];
    assign layer4_out[1125] = layer3_out[245] ^ layer3_out[246];
    assign layer4_out[1126] = ~(layer3_out[248] & layer3_out[249]);
    assign layer4_out[1127] = ~layer3_out[1528];
    assign layer4_out[1128] = ~(layer3_out[6768] ^ layer3_out[6769]);
    assign layer4_out[1129] = layer3_out[1903] | layer3_out[1904];
    assign layer4_out[1130] = layer3_out[5831];
    assign layer4_out[1131] = ~layer3_out[4318] | layer3_out[4319];
    assign layer4_out[1132] = ~layer3_out[4648];
    assign layer4_out[1133] = ~(layer3_out[2129] | layer3_out[2130]);
    assign layer4_out[1134] = ~layer3_out[6298] | layer3_out[6299];
    assign layer4_out[1135] = ~(layer3_out[2381] | layer3_out[2382]);
    assign layer4_out[1136] = ~(layer3_out[2587] & layer3_out[2588]);
    assign layer4_out[1137] = ~(layer3_out[1264] ^ layer3_out[1265]);
    assign layer4_out[1138] = layer3_out[6524];
    assign layer4_out[1139] = ~layer3_out[794];
    assign layer4_out[1140] = ~(layer3_out[5575] ^ layer3_out[5576]);
    assign layer4_out[1141] = ~layer3_out[5643];
    assign layer4_out[1142] = layer3_out[5795];
    assign layer4_out[1143] = layer3_out[3010] & ~layer3_out[3009];
    assign layer4_out[1144] = layer3_out[7564] | layer3_out[7565];
    assign layer4_out[1145] = ~layer3_out[4163];
    assign layer4_out[1146] = layer3_out[752];
    assign layer4_out[1147] = ~layer3_out[270] | layer3_out[269];
    assign layer4_out[1148] = layer3_out[6797];
    assign layer4_out[1149] = ~layer3_out[7312] | layer3_out[7313];
    assign layer4_out[1150] = ~(layer3_out[105] & layer3_out[106]);
    assign layer4_out[1151] = layer3_out[1497];
    assign layer4_out[1152] = ~layer3_out[4490] | layer3_out[4489];
    assign layer4_out[1153] = layer3_out[838] & ~layer3_out[839];
    assign layer4_out[1154] = ~layer3_out[7110];
    assign layer4_out[1155] = ~(layer3_out[4915] & layer3_out[4916]);
    assign layer4_out[1156] = ~(layer3_out[3936] ^ layer3_out[3937]);
    assign layer4_out[1157] = ~layer3_out[6678] | layer3_out[6679];
    assign layer4_out[1158] = layer3_out[6810] ^ layer3_out[6811];
    assign layer4_out[1159] = layer3_out[6457];
    assign layer4_out[1160] = layer3_out[4161];
    assign layer4_out[1161] = layer3_out[377];
    assign layer4_out[1162] = layer3_out[199] & ~layer3_out[198];
    assign layer4_out[1163] = layer3_out[7113] ^ layer3_out[7114];
    assign layer4_out[1164] = ~(layer3_out[7490] ^ layer3_out[7491]);
    assign layer4_out[1165] = ~(layer3_out[2407] | layer3_out[2408]);
    assign layer4_out[1166] = layer3_out[6155] ^ layer3_out[6156];
    assign layer4_out[1167] = layer3_out[3532] | layer3_out[3533];
    assign layer4_out[1168] = layer3_out[113] & ~layer3_out[114];
    assign layer4_out[1169] = layer3_out[4057];
    assign layer4_out[1170] = ~(layer3_out[5023] ^ layer3_out[5024]);
    assign layer4_out[1171] = layer3_out[661] & ~layer3_out[662];
    assign layer4_out[1172] = layer3_out[5626] & layer3_out[5627];
    assign layer4_out[1173] = layer3_out[6359];
    assign layer4_out[1174] = ~layer3_out[1234];
    assign layer4_out[1175] = layer3_out[6024] & layer3_out[6025];
    assign layer4_out[1176] = layer3_out[2342] & ~layer3_out[2341];
    assign layer4_out[1177] = ~(layer3_out[5365] | layer3_out[5366]);
    assign layer4_out[1178] = layer3_out[4284];
    assign layer4_out[1179] = layer3_out[5910];
    assign layer4_out[1180] = layer3_out[2605];
    assign layer4_out[1181] = layer3_out[3312];
    assign layer4_out[1182] = ~(layer3_out[5292] & layer3_out[5293]);
    assign layer4_out[1183] = layer3_out[3745];
    assign layer4_out[1184] = ~(layer3_out[5716] | layer3_out[5717]);
    assign layer4_out[1185] = ~layer3_out[2118] | layer3_out[2119];
    assign layer4_out[1186] = layer3_out[4322] ^ layer3_out[4323];
    assign layer4_out[1187] = layer3_out[5636] & ~layer3_out[5637];
    assign layer4_out[1188] = layer3_out[2091] ^ layer3_out[2092];
    assign layer4_out[1189] = ~layer3_out[2849] | layer3_out[2850];
    assign layer4_out[1190] = layer3_out[138] & ~layer3_out[139];
    assign layer4_out[1191] = ~layer3_out[2136] | layer3_out[2135];
    assign layer4_out[1192] = ~layer3_out[596] | layer3_out[597];
    assign layer4_out[1193] = ~(layer3_out[2243] ^ layer3_out[2244]);
    assign layer4_out[1194] = layer3_out[7092] & ~layer3_out[7091];
    assign layer4_out[1195] = ~(layer3_out[2322] & layer3_out[2323]);
    assign layer4_out[1196] = ~(layer3_out[5909] & layer3_out[5910]);
    assign layer4_out[1197] = ~layer3_out[919];
    assign layer4_out[1198] = ~layer3_out[5392] | layer3_out[5391];
    assign layer4_out[1199] = ~layer3_out[636] | layer3_out[637];
    assign layer4_out[1200] = ~layer3_out[6886];
    assign layer4_out[1201] = layer3_out[7431] & layer3_out[7432];
    assign layer4_out[1202] = layer3_out[2591] & layer3_out[2592];
    assign layer4_out[1203] = ~layer3_out[4851];
    assign layer4_out[1204] = layer3_out[6525] | layer3_out[6526];
    assign layer4_out[1205] = layer3_out[5281];
    assign layer4_out[1206] = layer3_out[1378] ^ layer3_out[1379];
    assign layer4_out[1207] = ~layer3_out[3485] | layer3_out[3484];
    assign layer4_out[1208] = ~layer3_out[4491] | layer3_out[4492];
    assign layer4_out[1209] = ~(layer3_out[7022] ^ layer3_out[7023]);
    assign layer4_out[1210] = layer3_out[5567];
    assign layer4_out[1211] = layer3_out[5795];
    assign layer4_out[1212] = ~layer3_out[4042];
    assign layer4_out[1213] = ~layer3_out[4804];
    assign layer4_out[1214] = layer3_out[137];
    assign layer4_out[1215] = layer3_out[7704];
    assign layer4_out[1216] = layer3_out[6671] & ~layer3_out[6672];
    assign layer4_out[1217] = layer3_out[2073] | layer3_out[2074];
    assign layer4_out[1218] = ~layer3_out[6896];
    assign layer4_out[1219] = ~(layer3_out[5284] ^ layer3_out[5285]);
    assign layer4_out[1220] = ~(layer3_out[7274] ^ layer3_out[7275]);
    assign layer4_out[1221] = ~layer3_out[2421];
    assign layer4_out[1222] = ~(layer3_out[3301] & layer3_out[3302]);
    assign layer4_out[1223] = layer3_out[4079] & layer3_out[4080];
    assign layer4_out[1224] = ~(layer3_out[3870] ^ layer3_out[3871]);
    assign layer4_out[1225] = ~layer3_out[6391];
    assign layer4_out[1226] = ~layer3_out[6657];
    assign layer4_out[1227] = ~layer3_out[1161];
    assign layer4_out[1228] = layer3_out[2198];
    assign layer4_out[1229] = ~(layer3_out[4404] | layer3_out[4405]);
    assign layer4_out[1230] = layer3_out[2374] ^ layer3_out[2375];
    assign layer4_out[1231] = ~layer3_out[7899] | layer3_out[7900];
    assign layer4_out[1232] = layer3_out[981] | layer3_out[982];
    assign layer4_out[1233] = ~(layer3_out[4984] ^ layer3_out[4985]);
    assign layer4_out[1234] = ~layer3_out[5812];
    assign layer4_out[1235] = layer3_out[527] ^ layer3_out[528];
    assign layer4_out[1236] = ~layer3_out[303];
    assign layer4_out[1237] = layer3_out[3140];
    assign layer4_out[1238] = layer3_out[839] ^ layer3_out[840];
    assign layer4_out[1239] = ~(layer3_out[3108] & layer3_out[3109]);
    assign layer4_out[1240] = ~(layer3_out[3376] & layer3_out[3377]);
    assign layer4_out[1241] = layer3_out[715];
    assign layer4_out[1242] = ~layer3_out[1353];
    assign layer4_out[1243] = ~layer3_out[6565] | layer3_out[6566];
    assign layer4_out[1244] = layer3_out[4764] ^ layer3_out[4765];
    assign layer4_out[1245] = layer3_out[1353] ^ layer3_out[1354];
    assign layer4_out[1246] = layer3_out[368];
    assign layer4_out[1247] = layer3_out[4462];
    assign layer4_out[1248] = ~layer3_out[7580];
    assign layer4_out[1249] = layer3_out[5068];
    assign layer4_out[1250] = ~layer3_out[3176];
    assign layer4_out[1251] = ~(layer3_out[1411] ^ layer3_out[1412]);
    assign layer4_out[1252] = ~layer3_out[4175];
    assign layer4_out[1253] = layer3_out[2164];
    assign layer4_out[1254] = ~layer3_out[1528];
    assign layer4_out[1255] = ~(layer3_out[4901] | layer3_out[4902]);
    assign layer4_out[1256] = layer3_out[7752] | layer3_out[7753];
    assign layer4_out[1257] = layer3_out[234] ^ layer3_out[235];
    assign layer4_out[1258] = layer3_out[424];
    assign layer4_out[1259] = ~layer3_out[2028] | layer3_out[2029];
    assign layer4_out[1260] = layer3_out[2400] & layer3_out[2401];
    assign layer4_out[1261] = layer3_out[2533] ^ layer3_out[2534];
    assign layer4_out[1262] = ~layer3_out[6745];
    assign layer4_out[1263] = ~layer3_out[2902];
    assign layer4_out[1264] = layer3_out[1111];
    assign layer4_out[1265] = ~(layer3_out[5169] & layer3_out[5170]);
    assign layer4_out[1266] = ~layer3_out[7303];
    assign layer4_out[1267] = ~(layer3_out[6881] ^ layer3_out[6882]);
    assign layer4_out[1268] = layer3_out[3417] & ~layer3_out[3416];
    assign layer4_out[1269] = ~layer3_out[5308] | layer3_out[5309];
    assign layer4_out[1270] = ~(layer3_out[6398] ^ layer3_out[6399]);
    assign layer4_out[1271] = ~layer3_out[3613];
    assign layer4_out[1272] = layer3_out[1217] ^ layer3_out[1218];
    assign layer4_out[1273] = layer3_out[6313];
    assign layer4_out[1274] = ~layer3_out[5592] | layer3_out[5591];
    assign layer4_out[1275] = ~(layer3_out[1950] | layer3_out[1951]);
    assign layer4_out[1276] = layer3_out[2936];
    assign layer4_out[1277] = layer3_out[6852] | layer3_out[6853];
    assign layer4_out[1278] = ~layer3_out[7543];
    assign layer4_out[1279] = layer3_out[3789] & ~layer3_out[3788];
    assign layer4_out[1280] = layer3_out[3602];
    assign layer4_out[1281] = ~(layer3_out[2294] ^ layer3_out[2295]);
    assign layer4_out[1282] = layer3_out[6129] | layer3_out[6130];
    assign layer4_out[1283] = ~layer3_out[3180];
    assign layer4_out[1284] = ~layer3_out[1616] | layer3_out[1615];
    assign layer4_out[1285] = layer3_out[72];
    assign layer4_out[1286] = layer3_out[1983];
    assign layer4_out[1287] = ~layer3_out[1210];
    assign layer4_out[1288] = ~(layer3_out[2070] & layer3_out[2071]);
    assign layer4_out[1289] = 1'b0;
    assign layer4_out[1290] = layer3_out[1202];
    assign layer4_out[1291] = layer3_out[5510] ^ layer3_out[5511];
    assign layer4_out[1292] = layer3_out[5333];
    assign layer4_out[1293] = layer3_out[2061] & layer3_out[2062];
    assign layer4_out[1294] = ~layer3_out[2722];
    assign layer4_out[1295] = ~(layer3_out[6111] ^ layer3_out[6112]);
    assign layer4_out[1296] = layer3_out[5388];
    assign layer4_out[1297] = layer3_out[2961] & layer3_out[2962];
    assign layer4_out[1298] = layer3_out[147];
    assign layer4_out[1299] = ~(layer3_out[2911] | layer3_out[2912]);
    assign layer4_out[1300] = layer3_out[302] | layer3_out[303];
    assign layer4_out[1301] = ~(layer3_out[5206] ^ layer3_out[5207]);
    assign layer4_out[1302] = layer3_out[4953] | layer3_out[4954];
    assign layer4_out[1303] = layer3_out[4852] | layer3_out[4853];
    assign layer4_out[1304] = ~(layer3_out[6682] & layer3_out[6683]);
    assign layer4_out[1305] = layer3_out[615];
    assign layer4_out[1306] = ~layer3_out[4571];
    assign layer4_out[1307] = ~(layer3_out[7198] | layer3_out[7199]);
    assign layer4_out[1308] = ~(layer3_out[7328] | layer3_out[7329]);
    assign layer4_out[1309] = layer3_out[2464] & ~layer3_out[2465];
    assign layer4_out[1310] = ~layer3_out[4604] | layer3_out[4605];
    assign layer4_out[1311] = ~layer3_out[6086];
    assign layer4_out[1312] = ~(layer3_out[653] & layer3_out[654]);
    assign layer4_out[1313] = ~(layer3_out[6106] ^ layer3_out[6107]);
    assign layer4_out[1314] = ~layer3_out[4040];
    assign layer4_out[1315] = layer3_out[6774] | layer3_out[6775];
    assign layer4_out[1316] = layer3_out[3708] & layer3_out[3709];
    assign layer4_out[1317] = ~(layer3_out[3803] | layer3_out[3804]);
    assign layer4_out[1318] = ~layer3_out[1212] | layer3_out[1211];
    assign layer4_out[1319] = layer3_out[7162] ^ layer3_out[7163];
    assign layer4_out[1320] = ~layer3_out[6113];
    assign layer4_out[1321] = ~(layer3_out[4757] | layer3_out[4758]);
    assign layer4_out[1322] = ~layer3_out[6115];
    assign layer4_out[1323] = layer3_out[5640] & ~layer3_out[5641];
    assign layer4_out[1324] = layer3_out[7904] & layer3_out[7905];
    assign layer4_out[1325] = ~layer3_out[1464] | layer3_out[1463];
    assign layer4_out[1326] = layer3_out[3111] ^ layer3_out[3112];
    assign layer4_out[1327] = ~layer3_out[6278];
    assign layer4_out[1328] = layer3_out[6321];
    assign layer4_out[1329] = layer3_out[7748] | layer3_out[7749];
    assign layer4_out[1330] = ~layer3_out[5096];
    assign layer4_out[1331] = layer3_out[6722] ^ layer3_out[6723];
    assign layer4_out[1332] = layer3_out[2694] ^ layer3_out[2695];
    assign layer4_out[1333] = ~layer3_out[1793] | layer3_out[1794];
    assign layer4_out[1334] = ~(layer3_out[5332] & layer3_out[5333]);
    assign layer4_out[1335] = ~layer3_out[6010] | layer3_out[6011];
    assign layer4_out[1336] = layer3_out[7342] & ~layer3_out[7343];
    assign layer4_out[1337] = layer3_out[7093] ^ layer3_out[7094];
    assign layer4_out[1338] = layer3_out[1297] & ~layer3_out[1296];
    assign layer4_out[1339] = ~layer3_out[1944];
    assign layer4_out[1340] = layer3_out[1585];
    assign layer4_out[1341] = 1'b1;
    assign layer4_out[1342] = ~layer3_out[1877];
    assign layer4_out[1343] = layer3_out[6641] ^ layer3_out[6642];
    assign layer4_out[1344] = layer3_out[7737];
    assign layer4_out[1345] = layer3_out[5843] | layer3_out[5844];
    assign layer4_out[1346] = layer3_out[5745];
    assign layer4_out[1347] = layer3_out[7444] & layer3_out[7445];
    assign layer4_out[1348] = ~(layer3_out[4710] ^ layer3_out[4711]);
    assign layer4_out[1349] = ~layer3_out[962];
    assign layer4_out[1350] = layer3_out[4273] ^ layer3_out[4274];
    assign layer4_out[1351] = ~layer3_out[2377] | layer3_out[2376];
    assign layer4_out[1352] = layer3_out[5894];
    assign layer4_out[1353] = ~layer3_out[126];
    assign layer4_out[1354] = ~layer3_out[7742] | layer3_out[7741];
    assign layer4_out[1355] = layer3_out[2342] | layer3_out[2343];
    assign layer4_out[1356] = ~layer3_out[3582] | layer3_out[3583];
    assign layer4_out[1357] = ~layer3_out[5639] | layer3_out[5640];
    assign layer4_out[1358] = ~layer3_out[3460] | layer3_out[3459];
    assign layer4_out[1359] = layer3_out[896];
    assign layer4_out[1360] = ~(layer3_out[6869] ^ layer3_out[6870]);
    assign layer4_out[1361] = layer3_out[3037] & ~layer3_out[3036];
    assign layer4_out[1362] = layer3_out[5432] | layer3_out[5433];
    assign layer4_out[1363] = ~layer3_out[3799] | layer3_out[3798];
    assign layer4_out[1364] = ~(layer3_out[6737] & layer3_out[6738]);
    assign layer4_out[1365] = ~(layer3_out[3407] ^ layer3_out[3408]);
    assign layer4_out[1366] = layer3_out[7335] & layer3_out[7336];
    assign layer4_out[1367] = ~layer3_out[5614] | layer3_out[5613];
    assign layer4_out[1368] = ~layer3_out[3876];
    assign layer4_out[1369] = layer3_out[5790] & layer3_out[5791];
    assign layer4_out[1370] = ~layer3_out[4077] | layer3_out[4076];
    assign layer4_out[1371] = ~(layer3_out[785] & layer3_out[786]);
    assign layer4_out[1372] = layer3_out[2899];
    assign layer4_out[1373] = ~layer3_out[7416];
    assign layer4_out[1374] = ~layer3_out[7391] | layer3_out[7392];
    assign layer4_out[1375] = ~layer3_out[550];
    assign layer4_out[1376] = ~layer3_out[7960];
    assign layer4_out[1377] = ~layer3_out[2339];
    assign layer4_out[1378] = layer3_out[7488];
    assign layer4_out[1379] = layer3_out[5114];
    assign layer4_out[1380] = layer3_out[7894] ^ layer3_out[7895];
    assign layer4_out[1381] = layer3_out[2622];
    assign layer4_out[1382] = ~layer3_out[6749] | layer3_out[6748];
    assign layer4_out[1383] = ~(layer3_out[575] ^ layer3_out[576]);
    assign layer4_out[1384] = ~layer3_out[2549] | layer3_out[2548];
    assign layer4_out[1385] = layer3_out[362] & ~layer3_out[361];
    assign layer4_out[1386] = ~layer3_out[1104];
    assign layer4_out[1387] = ~(layer3_out[5104] & layer3_out[5105]);
    assign layer4_out[1388] = ~layer3_out[7251] | layer3_out[7252];
    assign layer4_out[1389] = layer3_out[4346];
    assign layer4_out[1390] = layer3_out[3267];
    assign layer4_out[1391] = layer3_out[3163] ^ layer3_out[3164];
    assign layer4_out[1392] = layer3_out[7486] & ~layer3_out[7487];
    assign layer4_out[1393] = ~layer3_out[1287];
    assign layer4_out[1394] = ~(layer3_out[6402] ^ layer3_out[6403]);
    assign layer4_out[1395] = layer3_out[427] & layer3_out[428];
    assign layer4_out[1396] = ~(layer3_out[3273] ^ layer3_out[3274]);
    assign layer4_out[1397] = layer3_out[2873] & ~layer3_out[2872];
    assign layer4_out[1398] = ~layer3_out[4867] | layer3_out[4868];
    assign layer4_out[1399] = ~layer3_out[798] | layer3_out[799];
    assign layer4_out[1400] = layer3_out[3842] ^ layer3_out[3843];
    assign layer4_out[1401] = layer3_out[2028];
    assign layer4_out[1402] = layer3_out[6238];
    assign layer4_out[1403] = ~(layer3_out[29] ^ layer3_out[30]);
    assign layer4_out[1404] = ~(layer3_out[2382] ^ layer3_out[2383]);
    assign layer4_out[1405] = ~(layer3_out[5378] & layer3_out[5379]);
    assign layer4_out[1406] = ~layer3_out[1830];
    assign layer4_out[1407] = layer3_out[2373] & ~layer3_out[2372];
    assign layer4_out[1408] = ~layer3_out[671];
    assign layer4_out[1409] = layer3_out[1180] ^ layer3_out[1181];
    assign layer4_out[1410] = ~layer3_out[7307];
    assign layer4_out[1411] = layer3_out[4824] ^ layer3_out[4825];
    assign layer4_out[1412] = ~(layer3_out[858] & layer3_out[859]);
    assign layer4_out[1413] = layer3_out[7599];
    assign layer4_out[1414] = ~(layer3_out[1152] & layer3_out[1153]);
    assign layer4_out[1415] = ~(layer3_out[316] | layer3_out[317]);
    assign layer4_out[1416] = ~(layer3_out[5994] ^ layer3_out[5995]);
    assign layer4_out[1417] = layer3_out[5155] & ~layer3_out[5156];
    assign layer4_out[1418] = ~layer3_out[725];
    assign layer4_out[1419] = ~layer3_out[749];
    assign layer4_out[1420] = layer3_out[3944] & layer3_out[3945];
    assign layer4_out[1421] = ~layer3_out[4232] | layer3_out[4231];
    assign layer4_out[1422] = layer3_out[379];
    assign layer4_out[1423] = ~layer3_out[1131] | layer3_out[1130];
    assign layer4_out[1424] = ~(layer3_out[2825] | layer3_out[2826]);
    assign layer4_out[1425] = layer3_out[542];
    assign layer4_out[1426] = ~layer3_out[890];
    assign layer4_out[1427] = layer3_out[1060];
    assign layer4_out[1428] = ~layer3_out[4171];
    assign layer4_out[1429] = ~layer3_out[3360];
    assign layer4_out[1430] = ~layer3_out[294];
    assign layer4_out[1431] = layer3_out[194] | layer3_out[195];
    assign layer4_out[1432] = layer3_out[4880] | layer3_out[4881];
    assign layer4_out[1433] = ~layer3_out[7937];
    assign layer4_out[1434] = layer3_out[1119];
    assign layer4_out[1435] = ~(layer3_out[5844] | layer3_out[5845]);
    assign layer4_out[1436] = ~(layer3_out[2078] & layer3_out[2079]);
    assign layer4_out[1437] = ~layer3_out[5406];
    assign layer4_out[1438] = layer3_out[7321] & layer3_out[7322];
    assign layer4_out[1439] = ~(layer3_out[894] ^ layer3_out[895]);
    assign layer4_out[1440] = layer3_out[4324];
    assign layer4_out[1441] = ~layer3_out[81] | layer3_out[80];
    assign layer4_out[1442] = ~layer3_out[6594];
    assign layer4_out[1443] = layer3_out[6923] | layer3_out[6924];
    assign layer4_out[1444] = layer3_out[4967] ^ layer3_out[4968];
    assign layer4_out[1445] = layer3_out[7111] ^ layer3_out[7112];
    assign layer4_out[1446] = ~(layer3_out[4533] ^ layer3_out[4534]);
    assign layer4_out[1447] = 1'b1;
    assign layer4_out[1448] = ~layer3_out[7291];
    assign layer4_out[1449] = ~layer3_out[3084] | layer3_out[3083];
    assign layer4_out[1450] = layer3_out[243];
    assign layer4_out[1451] = ~(layer3_out[6883] ^ layer3_out[6884]);
    assign layer4_out[1452] = ~(layer3_out[663] & layer3_out[664]);
    assign layer4_out[1453] = ~(layer3_out[2902] | layer3_out[2903]);
    assign layer4_out[1454] = layer3_out[116] & ~layer3_out[115];
    assign layer4_out[1455] = layer3_out[498] & ~layer3_out[499];
    assign layer4_out[1456] = ~layer3_out[1091];
    assign layer4_out[1457] = layer3_out[181] ^ layer3_out[182];
    assign layer4_out[1458] = layer3_out[5297];
    assign layer4_out[1459] = ~(layer3_out[7831] & layer3_out[7832]);
    assign layer4_out[1460] = ~layer3_out[3289];
    assign layer4_out[1461] = layer3_out[2121];
    assign layer4_out[1462] = ~(layer3_out[1120] ^ layer3_out[1121]);
    assign layer4_out[1463] = layer3_out[5189];
    assign layer4_out[1464] = layer3_out[5518];
    assign layer4_out[1465] = layer3_out[574] & ~layer3_out[573];
    assign layer4_out[1466] = ~layer3_out[3065];
    assign layer4_out[1467] = layer3_out[5136];
    assign layer4_out[1468] = layer3_out[924];
    assign layer4_out[1469] = layer3_out[5294];
    assign layer4_out[1470] = ~layer3_out[3579];
    assign layer4_out[1471] = layer3_out[6725] & ~layer3_out[6726];
    assign layer4_out[1472] = ~layer3_out[7666] | layer3_out[7667];
    assign layer4_out[1473] = ~(layer3_out[3811] | layer3_out[3812]);
    assign layer4_out[1474] = layer3_out[2046];
    assign layer4_out[1475] = ~(layer3_out[4033] | layer3_out[4034]);
    assign layer4_out[1476] = layer3_out[3239] | layer3_out[3240];
    assign layer4_out[1477] = ~(layer3_out[980] & layer3_out[981]);
    assign layer4_out[1478] = layer3_out[5326] & ~layer3_out[5327];
    assign layer4_out[1479] = ~(layer3_out[3125] & layer3_out[3126]);
    assign layer4_out[1480] = ~(layer3_out[3186] | layer3_out[3187]);
    assign layer4_out[1481] = ~layer3_out[4918] | layer3_out[4919];
    assign layer4_out[1482] = ~(layer3_out[814] & layer3_out[815]);
    assign layer4_out[1483] = ~layer3_out[6192];
    assign layer4_out[1484] = ~layer3_out[3134];
    assign layer4_out[1485] = ~(layer3_out[3560] & layer3_out[3561]);
    assign layer4_out[1486] = layer3_out[5374] & ~layer3_out[5375];
    assign layer4_out[1487] = ~layer3_out[4965] | layer3_out[4964];
    assign layer4_out[1488] = layer3_out[4471];
    assign layer4_out[1489] = ~(layer3_out[2928] ^ layer3_out[2929]);
    assign layer4_out[1490] = ~(layer3_out[5430] ^ layer3_out[5431]);
    assign layer4_out[1491] = ~layer3_out[5605] | layer3_out[5606];
    assign layer4_out[1492] = layer3_out[7120] ^ layer3_out[7121];
    assign layer4_out[1493] = layer3_out[1577];
    assign layer4_out[1494] = ~(layer3_out[2648] & layer3_out[2649]);
    assign layer4_out[1495] = ~(layer3_out[2275] | layer3_out[2276]);
    assign layer4_out[1496] = ~(layer3_out[1281] ^ layer3_out[1282]);
    assign layer4_out[1497] = ~(layer3_out[7081] & layer3_out[7082]);
    assign layer4_out[1498] = layer3_out[2011];
    assign layer4_out[1499] = ~layer3_out[3252];
    assign layer4_out[1500] = layer3_out[6210] & ~layer3_out[6209];
    assign layer4_out[1501] = layer3_out[6021];
    assign layer4_out[1502] = layer3_out[5982] & layer3_out[5983];
    assign layer4_out[1503] = layer3_out[340];
    assign layer4_out[1504] = layer3_out[6366] & ~layer3_out[6367];
    assign layer4_out[1505] = layer3_out[6128];
    assign layer4_out[1506] = layer3_out[7847] ^ layer3_out[7848];
    assign layer4_out[1507] = ~(layer3_out[6049] | layer3_out[6050]);
    assign layer4_out[1508] = layer3_out[2712];
    assign layer4_out[1509] = ~layer3_out[2263];
    assign layer4_out[1510] = ~layer3_out[5577];
    assign layer4_out[1511] = layer3_out[1964] & ~layer3_out[1965];
    assign layer4_out[1512] = layer3_out[4777] ^ layer3_out[4778];
    assign layer4_out[1513] = layer3_out[7002] & layer3_out[7003];
    assign layer4_out[1514] = layer3_out[2414];
    assign layer4_out[1515] = ~layer3_out[3944] | layer3_out[3943];
    assign layer4_out[1516] = layer3_out[6055] & ~layer3_out[6056];
    assign layer4_out[1517] = ~(layer3_out[3346] | layer3_out[3347]);
    assign layer4_out[1518] = ~layer3_out[1763] | layer3_out[1762];
    assign layer4_out[1519] = layer3_out[1999] ^ layer3_out[2000];
    assign layer4_out[1520] = ~layer3_out[729];
    assign layer4_out[1521] = layer3_out[6670] ^ layer3_out[6671];
    assign layer4_out[1522] = layer3_out[7837] ^ layer3_out[7838];
    assign layer4_out[1523] = 1'b1;
    assign layer4_out[1524] = layer3_out[6114];
    assign layer4_out[1525] = ~(layer3_out[562] ^ layer3_out[563]);
    assign layer4_out[1526] = ~layer3_out[5363] | layer3_out[5364];
    assign layer4_out[1527] = ~layer3_out[3423];
    assign layer4_out[1528] = ~(layer3_out[3956] & layer3_out[3957]);
    assign layer4_out[1529] = layer3_out[4685] | layer3_out[4686];
    assign layer4_out[1530] = ~(layer3_out[2120] & layer3_out[2121]);
    assign layer4_out[1531] = ~(layer3_out[2820] | layer3_out[2821]);
    assign layer4_out[1532] = layer3_out[5537] & layer3_out[5538];
    assign layer4_out[1533] = layer3_out[7798];
    assign layer4_out[1534] = layer3_out[6355] | layer3_out[6356];
    assign layer4_out[1535] = layer3_out[4727];
    assign layer4_out[1536] = layer3_out[4147] ^ layer3_out[4148];
    assign layer4_out[1537] = layer3_out[1441] | layer3_out[1442];
    assign layer4_out[1538] = layer3_out[7122] ^ layer3_out[7123];
    assign layer4_out[1539] = ~(layer3_out[6333] & layer3_out[6334]);
    assign layer4_out[1540] = layer3_out[1661] ^ layer3_out[1662];
    assign layer4_out[1541] = 1'b0;
    assign layer4_out[1542] = layer3_out[6559];
    assign layer4_out[1543] = layer3_out[2326];
    assign layer4_out[1544] = ~layer3_out[6148];
    assign layer4_out[1545] = ~layer3_out[5712];
    assign layer4_out[1546] = ~(layer3_out[4877] ^ layer3_out[4878]);
    assign layer4_out[1547] = layer3_out[4558];
    assign layer4_out[1548] = layer3_out[1426];
    assign layer4_out[1549] = layer3_out[7477] ^ layer3_out[7478];
    assign layer4_out[1550] = ~layer3_out[4012];
    assign layer4_out[1551] = ~layer3_out[5177];
    assign layer4_out[1552] = layer3_out[7938] ^ layer3_out[7939];
    assign layer4_out[1553] = layer3_out[2319];
    assign layer4_out[1554] = layer3_out[7675];
    assign layer4_out[1555] = ~(layer3_out[2586] ^ layer3_out[2587]);
    assign layer4_out[1556] = layer3_out[5864] | layer3_out[5865];
    assign layer4_out[1557] = layer3_out[3902] & ~layer3_out[3903];
    assign layer4_out[1558] = ~layer3_out[3650];
    assign layer4_out[1559] = ~layer3_out[7864];
    assign layer4_out[1560] = ~(layer3_out[2424] ^ layer3_out[2425]);
    assign layer4_out[1561] = ~layer3_out[4920];
    assign layer4_out[1562] = ~(layer3_out[2915] ^ layer3_out[2916]);
    assign layer4_out[1563] = ~layer3_out[3150] | layer3_out[3149];
    assign layer4_out[1564] = ~layer3_out[4071];
    assign layer4_out[1565] = layer3_out[3494] ^ layer3_out[3495];
    assign layer4_out[1566] = layer3_out[7185];
    assign layer4_out[1567] = layer3_out[6246];
    assign layer4_out[1568] = layer3_out[6244];
    assign layer4_out[1569] = layer3_out[1899];
    assign layer4_out[1570] = ~layer3_out[4355];
    assign layer4_out[1571] = ~layer3_out[3592];
    assign layer4_out[1572] = layer3_out[151] & layer3_out[152];
    assign layer4_out[1573] = ~(layer3_out[817] & layer3_out[818]);
    assign layer4_out[1574] = layer3_out[3651];
    assign layer4_out[1575] = layer3_out[49];
    assign layer4_out[1576] = layer3_out[1724] ^ layer3_out[1725];
    assign layer4_out[1577] = layer3_out[3388] | layer3_out[3389];
    assign layer4_out[1578] = layer3_out[6808];
    assign layer4_out[1579] = layer3_out[628];
    assign layer4_out[1580] = ~layer3_out[2430] | layer3_out[2429];
    assign layer4_out[1581] = layer3_out[2968];
    assign layer4_out[1582] = layer3_out[4064];
    assign layer4_out[1583] = ~layer3_out[502];
    assign layer4_out[1584] = layer3_out[1555] & ~layer3_out[1554];
    assign layer4_out[1585] = ~layer3_out[4114] | layer3_out[4113];
    assign layer4_out[1586] = ~(layer3_out[2089] | layer3_out[2090]);
    assign layer4_out[1587] = layer3_out[1652];
    assign layer4_out[1588] = ~(layer3_out[1465] | layer3_out[1466]);
    assign layer4_out[1589] = layer3_out[4355];
    assign layer4_out[1590] = layer3_out[4297] ^ layer3_out[4298];
    assign layer4_out[1591] = ~layer3_out[2025];
    assign layer4_out[1592] = ~layer3_out[3036];
    assign layer4_out[1593] = layer3_out[4855] & ~layer3_out[4856];
    assign layer4_out[1594] = ~(layer3_out[1492] ^ layer3_out[1493]);
    assign layer4_out[1595] = ~layer3_out[5028];
    assign layer4_out[1596] = layer3_out[2375] & layer3_out[2376];
    assign layer4_out[1597] = layer3_out[5208] & layer3_out[5209];
    assign layer4_out[1598] = ~layer3_out[1665] | layer3_out[1666];
    assign layer4_out[1599] = ~(layer3_out[4389] ^ layer3_out[4390]);
    assign layer4_out[1600] = ~layer3_out[7420];
    assign layer4_out[1601] = layer3_out[5793];
    assign layer4_out[1602] = layer3_out[2172] | layer3_out[2173];
    assign layer4_out[1603] = layer3_out[1833] ^ layer3_out[1834];
    assign layer4_out[1604] = layer3_out[4053] ^ layer3_out[4054];
    assign layer4_out[1605] = ~layer3_out[58] | layer3_out[57];
    assign layer4_out[1606] = ~layer3_out[6687];
    assign layer4_out[1607] = layer3_out[602] & ~layer3_out[603];
    assign layer4_out[1608] = layer3_out[3984];
    assign layer4_out[1609] = ~(layer3_out[2527] ^ layer3_out[2528]);
    assign layer4_out[1610] = ~(layer3_out[2023] ^ layer3_out[2024]);
    assign layer4_out[1611] = ~layer3_out[6720];
    assign layer4_out[1612] = layer3_out[6831] & layer3_out[6832];
    assign layer4_out[1613] = ~layer3_out[1218];
    assign layer4_out[1614] = ~layer3_out[7593] | layer3_out[7594];
    assign layer4_out[1615] = ~layer3_out[383];
    assign layer4_out[1616] = ~layer3_out[359] | layer3_out[358];
    assign layer4_out[1617] = layer3_out[7443];
    assign layer4_out[1618] = layer3_out[5310] & ~layer3_out[5311];
    assign layer4_out[1619] = layer3_out[2044];
    assign layer4_out[1620] = layer3_out[736];
    assign layer4_out[1621] = layer3_out[2043] & ~layer3_out[2042];
    assign layer4_out[1622] = ~layer3_out[6528] | layer3_out[6529];
    assign layer4_out[1623] = ~layer3_out[2585] | layer3_out[2586];
    assign layer4_out[1624] = layer3_out[3092] ^ layer3_out[3093];
    assign layer4_out[1625] = ~layer3_out[3995] | layer3_out[3996];
    assign layer4_out[1626] = layer3_out[1735] | layer3_out[1736];
    assign layer4_out[1627] = ~(layer3_out[4750] & layer3_out[4751]);
    assign layer4_out[1628] = layer3_out[3395];
    assign layer4_out[1629] = layer3_out[2817] & ~layer3_out[2816];
    assign layer4_out[1630] = layer3_out[5546];
    assign layer4_out[1631] = layer3_out[3469];
    assign layer4_out[1632] = ~layer3_out[6521] | layer3_out[6522];
    assign layer4_out[1633] = ~layer3_out[3783];
    assign layer4_out[1634] = ~layer3_out[5218] | layer3_out[5219];
    assign layer4_out[1635] = ~(layer3_out[4476] ^ layer3_out[4477]);
    assign layer4_out[1636] = layer3_out[4636] | layer3_out[4637];
    assign layer4_out[1637] = layer3_out[3930] ^ layer3_out[3931];
    assign layer4_out[1638] = ~layer3_out[2012] | layer3_out[2013];
    assign layer4_out[1639] = layer3_out[5074];
    assign layer4_out[1640] = ~(layer3_out[4854] & layer3_out[4855]);
    assign layer4_out[1641] = layer3_out[2277] & layer3_out[2278];
    assign layer4_out[1642] = ~layer3_out[625] | layer3_out[624];
    assign layer4_out[1643] = ~layer3_out[3900];
    assign layer4_out[1644] = layer3_out[5185] & ~layer3_out[5184];
    assign layer4_out[1645] = layer3_out[3541];
    assign layer4_out[1646] = layer3_out[832] & ~layer3_out[831];
    assign layer4_out[1647] = ~layer3_out[2313];
    assign layer4_out[1648] = layer3_out[7352] & layer3_out[7353];
    assign layer4_out[1649] = ~layer3_out[1761];
    assign layer4_out[1650] = ~layer3_out[5495] | layer3_out[5494];
    assign layer4_out[1651] = ~layer3_out[1475];
    assign layer4_out[1652] = layer3_out[7319];
    assign layer4_out[1653] = ~(layer3_out[129] ^ layer3_out[130]);
    assign layer4_out[1654] = ~(layer3_out[5535] ^ layer3_out[5536]);
    assign layer4_out[1655] = layer3_out[4666];
    assign layer4_out[1656] = layer3_out[4787] & ~layer3_out[4788];
    assign layer4_out[1657] = ~layer3_out[533];
    assign layer4_out[1658] = ~(layer3_out[3442] & layer3_out[3443]);
    assign layer4_out[1659] = layer3_out[1469];
    assign layer4_out[1660] = layer3_out[6560] & ~layer3_out[6559];
    assign layer4_out[1661] = ~(layer3_out[633] & layer3_out[634]);
    assign layer4_out[1662] = ~layer3_out[1657];
    assign layer4_out[1663] = ~(layer3_out[6878] ^ layer3_out[6879]);
    assign layer4_out[1664] = layer3_out[5364] & ~layer3_out[5365];
    assign layer4_out[1665] = layer3_out[5708];
    assign layer4_out[1666] = layer3_out[4242];
    assign layer4_out[1667] = layer3_out[1446] & ~layer3_out[1447];
    assign layer4_out[1668] = ~(layer3_out[3723] | layer3_out[3724]);
    assign layer4_out[1669] = layer3_out[2018];
    assign layer4_out[1670] = ~layer3_out[893] | layer3_out[892];
    assign layer4_out[1671] = layer3_out[1028] & ~layer3_out[1027];
    assign layer4_out[1672] = ~layer3_out[2517];
    assign layer4_out[1673] = ~(layer3_out[3901] & layer3_out[3902]);
    assign layer4_out[1674] = ~layer3_out[3816];
    assign layer4_out[1675] = ~layer3_out[929];
    assign layer4_out[1676] = ~layer3_out[301];
    assign layer4_out[1677] = ~(layer3_out[649] | layer3_out[650]);
    assign layer4_out[1678] = ~(layer3_out[762] | layer3_out[763]);
    assign layer4_out[1679] = ~(layer3_out[6337] | layer3_out[6338]);
    assign layer4_out[1680] = ~layer3_out[2031];
    assign layer4_out[1681] = layer3_out[6621] & ~layer3_out[6622];
    assign layer4_out[1682] = layer3_out[3827] ^ layer3_out[3828];
    assign layer4_out[1683] = ~layer3_out[1714];
    assign layer4_out[1684] = ~layer3_out[3737];
    assign layer4_out[1685] = ~(layer3_out[537] ^ layer3_out[538]);
    assign layer4_out[1686] = ~layer3_out[4467];
    assign layer4_out[1687] = ~layer3_out[7352];
    assign layer4_out[1688] = ~(layer3_out[6477] ^ layer3_out[6478]);
    assign layer4_out[1689] = layer3_out[5917];
    assign layer4_out[1690] = layer3_out[872] & ~layer3_out[871];
    assign layer4_out[1691] = layer3_out[7772] & layer3_out[7773];
    assign layer4_out[1692] = ~(layer3_out[3634] & layer3_out[3635]);
    assign layer4_out[1693] = layer3_out[73] & ~layer3_out[74];
    assign layer4_out[1694] = layer3_out[5318] & layer3_out[5319];
    assign layer4_out[1695] = ~layer3_out[6412] | layer3_out[6413];
    assign layer4_out[1696] = ~(layer3_out[327] | layer3_out[328]);
    assign layer4_out[1697] = ~(layer3_out[3921] ^ layer3_out[3922]);
    assign layer4_out[1698] = ~(layer3_out[4121] & layer3_out[4122]);
    assign layer4_out[1699] = ~layer3_out[3753];
    assign layer4_out[1700] = layer3_out[2460] & ~layer3_out[2461];
    assign layer4_out[1701] = layer3_out[3711] & ~layer3_out[3712];
    assign layer4_out[1702] = ~(layer3_out[3767] & layer3_out[3768]);
    assign layer4_out[1703] = ~(layer3_out[3690] & layer3_out[3691]);
    assign layer4_out[1704] = layer3_out[4365];
    assign layer4_out[1705] = ~layer3_out[2046];
    assign layer4_out[1706] = 1'b0;
    assign layer4_out[1707] = ~layer3_out[1787] | layer3_out[1786];
    assign layer4_out[1708] = ~layer3_out[4310];
    assign layer4_out[1709] = ~layer3_out[4218] | layer3_out[4217];
    assign layer4_out[1710] = ~layer3_out[3755];
    assign layer4_out[1711] = layer3_out[7858];
    assign layer4_out[1712] = ~(layer3_out[7441] | layer3_out[7442]);
    assign layer4_out[1713] = ~layer3_out[7687];
    assign layer4_out[1714] = layer3_out[7961];
    assign layer4_out[1715] = layer3_out[7456] & ~layer3_out[7457];
    assign layer4_out[1716] = ~(layer3_out[1013] ^ layer3_out[1014]);
    assign layer4_out[1717] = layer3_out[4066] & layer3_out[4067];
    assign layer4_out[1718] = ~(layer3_out[2601] & layer3_out[2602]);
    assign layer4_out[1719] = ~layer3_out[4988];
    assign layer4_out[1720] = ~(layer3_out[5075] & layer3_out[5076]);
    assign layer4_out[1721] = layer3_out[3463] ^ layer3_out[3464];
    assign layer4_out[1722] = 1'b0;
    assign layer4_out[1723] = layer3_out[3059] ^ layer3_out[3060];
    assign layer4_out[1724] = ~(layer3_out[6099] ^ layer3_out[6100]);
    assign layer4_out[1725] = ~layer3_out[6734];
    assign layer4_out[1726] = ~layer3_out[6286] | layer3_out[6285];
    assign layer4_out[1727] = layer3_out[1660];
    assign layer4_out[1728] = ~layer3_out[2231];
    assign layer4_out[1729] = layer3_out[3367];
    assign layer4_out[1730] = layer3_out[1603];
    assign layer4_out[1731] = layer3_out[1362] & ~layer3_out[1361];
    assign layer4_out[1732] = layer3_out[3897] ^ layer3_out[3898];
    assign layer4_out[1733] = layer3_out[6192] ^ layer3_out[6193];
    assign layer4_out[1734] = ~layer3_out[3738] | layer3_out[3737];
    assign layer4_out[1735] = ~(layer3_out[3566] | layer3_out[3567]);
    assign layer4_out[1736] = ~layer3_out[3028];
    assign layer4_out[1737] = ~layer3_out[7605];
    assign layer4_out[1738] = layer3_out[259] & layer3_out[260];
    assign layer4_out[1739] = ~(layer3_out[2041] ^ layer3_out[2042]);
    assign layer4_out[1740] = ~layer3_out[5748] | layer3_out[5749];
    assign layer4_out[1741] = layer3_out[1001] ^ layer3_out[1002];
    assign layer4_out[1742] = ~layer3_out[3286] | layer3_out[3287];
    assign layer4_out[1743] = ~layer3_out[2858];
    assign layer4_out[1744] = 1'b1;
    assign layer4_out[1745] = layer3_out[7535];
    assign layer4_out[1746] = layer3_out[2624];
    assign layer4_out[1747] = ~layer3_out[5620];
    assign layer4_out[1748] = layer3_out[5502];
    assign layer4_out[1749] = ~layer3_out[7809];
    assign layer4_out[1750] = layer3_out[2995] & layer3_out[2996];
    assign layer4_out[1751] = ~(layer3_out[4650] | layer3_out[4651]);
    assign layer4_out[1752] = layer3_out[3853];
    assign layer4_out[1753] = ~layer3_out[568];
    assign layer4_out[1754] = ~layer3_out[2480];
    assign layer4_out[1755] = layer3_out[911] & ~layer3_out[912];
    assign layer4_out[1756] = ~(layer3_out[1574] ^ layer3_out[1575]);
    assign layer4_out[1757] = layer3_out[1552] ^ layer3_out[1553];
    assign layer4_out[1758] = ~layer3_out[7828];
    assign layer4_out[1759] = ~layer3_out[6736];
    assign layer4_out[1760] = ~(layer3_out[6400] ^ layer3_out[6401]);
    assign layer4_out[1761] = layer3_out[3721];
    assign layer4_out[1762] = ~layer3_out[7106];
    assign layer4_out[1763] = ~layer3_out[2272];
    assign layer4_out[1764] = layer3_out[6756];
    assign layer4_out[1765] = ~(layer3_out[6791] & layer3_out[6792]);
    assign layer4_out[1766] = layer3_out[1753];
    assign layer4_out[1767] = layer3_out[4005];
    assign layer4_out[1768] = layer3_out[1521] ^ layer3_out[1522];
    assign layer4_out[1769] = ~(layer3_out[7365] | layer3_out[7366]);
    assign layer4_out[1770] = ~layer3_out[6430] | layer3_out[6429];
    assign layer4_out[1771] = ~(layer3_out[4688] ^ layer3_out[4689]);
    assign layer4_out[1772] = ~layer3_out[5497] | layer3_out[5496];
    assign layer4_out[1773] = ~layer3_out[4114] | layer3_out[4115];
    assign layer4_out[1774] = ~layer3_out[1570];
    assign layer4_out[1775] = ~(layer3_out[7645] & layer3_out[7646]);
    assign layer4_out[1776] = ~layer3_out[5827];
    assign layer4_out[1777] = ~(layer3_out[6961] | layer3_out[6962]);
    assign layer4_out[1778] = layer3_out[4087];
    assign layer4_out[1779] = 1'b0;
    assign layer4_out[1780] = layer3_out[6625];
    assign layer4_out[1781] = ~layer3_out[1491];
    assign layer4_out[1782] = layer3_out[4638] & layer3_out[4639];
    assign layer4_out[1783] = ~(layer3_out[6280] ^ layer3_out[6281]);
    assign layer4_out[1784] = layer3_out[7716];
    assign layer4_out[1785] = layer3_out[228];
    assign layer4_out[1786] = ~(layer3_out[1470] & layer3_out[1471]);
    assign layer4_out[1787] = ~(layer3_out[1365] & layer3_out[1366]);
    assign layer4_out[1788] = layer3_out[1697] ^ layer3_out[1698];
    assign layer4_out[1789] = ~layer3_out[6464];
    assign layer4_out[1790] = ~layer3_out[2519];
    assign layer4_out[1791] = layer3_out[6054] & ~layer3_out[6053];
    assign layer4_out[1792] = layer3_out[553] ^ layer3_out[554];
    assign layer4_out[1793] = layer3_out[2818] & layer3_out[2819];
    assign layer4_out[1794] = layer3_out[6717] ^ layer3_out[6718];
    assign layer4_out[1795] = layer3_out[1850];
    assign layer4_out[1796] = ~(layer3_out[2269] ^ layer3_out[2270]);
    assign layer4_out[1797] = ~layer3_out[7247];
    assign layer4_out[1798] = ~layer3_out[6872];
    assign layer4_out[1799] = layer3_out[622];
    assign layer4_out[1800] = ~layer3_out[6136];
    assign layer4_out[1801] = ~layer3_out[4523] | layer3_out[4522];
    assign layer4_out[1802] = layer3_out[3752];
    assign layer4_out[1803] = layer3_out[6497];
    assign layer4_out[1804] = ~layer3_out[6703];
    assign layer4_out[1805] = layer3_out[2638] & ~layer3_out[2639];
    assign layer4_out[1806] = layer3_out[5185] | layer3_out[5186];
    assign layer4_out[1807] = layer3_out[353] ^ layer3_out[354];
    assign layer4_out[1808] = ~layer3_out[4737];
    assign layer4_out[1809] = layer3_out[6116] & ~layer3_out[6117];
    assign layer4_out[1810] = layer3_out[7169] | layer3_out[7170];
    assign layer4_out[1811] = layer3_out[676];
    assign layer4_out[1812] = ~layer3_out[7738];
    assign layer4_out[1813] = layer3_out[5540] ^ layer3_out[5541];
    assign layer4_out[1814] = ~layer3_out[4173];
    assign layer4_out[1815] = ~layer3_out[7787] | layer3_out[7786];
    assign layer4_out[1816] = layer3_out[6329];
    assign layer4_out[1817] = layer3_out[1297] & layer3_out[1298];
    assign layer4_out[1818] = ~layer3_out[7095];
    assign layer4_out[1819] = layer3_out[4447];
    assign layer4_out[1820] = ~layer3_out[2202] | layer3_out[2203];
    assign layer4_out[1821] = layer3_out[2311] ^ layer3_out[2312];
    assign layer4_out[1822] = ~layer3_out[7927];
    assign layer4_out[1823] = ~layer3_out[1365] | layer3_out[1364];
    assign layer4_out[1824] = ~layer3_out[5704] | layer3_out[5705];
    assign layer4_out[1825] = ~(layer3_out[6245] | layer3_out[6246]);
    assign layer4_out[1826] = layer3_out[7931] & ~layer3_out[7932];
    assign layer4_out[1827] = layer3_out[7849] | layer3_out[7850];
    assign layer4_out[1828] = ~(layer3_out[2208] | layer3_out[2209]);
    assign layer4_out[1829] = layer3_out[89];
    assign layer4_out[1830] = layer3_out[3743] | layer3_out[3744];
    assign layer4_out[1831] = layer3_out[5438] | layer3_out[5439];
    assign layer4_out[1832] = ~layer3_out[5693] | layer3_out[5692];
    assign layer4_out[1833] = layer3_out[7284] ^ layer3_out[7285];
    assign layer4_out[1834] = layer3_out[1127];
    assign layer4_out[1835] = 1'b0;
    assign layer4_out[1836] = ~(layer3_out[2158] ^ layer3_out[2159]);
    assign layer4_out[1837] = layer3_out[6510] & layer3_out[6511];
    assign layer4_out[1838] = layer3_out[6669];
    assign layer4_out[1839] = layer3_out[3292] & ~layer3_out[3293];
    assign layer4_out[1840] = ~layer3_out[368] | layer3_out[369];
    assign layer4_out[1841] = layer3_out[3985];
    assign layer4_out[1842] = ~layer3_out[5525];
    assign layer4_out[1843] = ~layer3_out[5418] | layer3_out[5419];
    assign layer4_out[1844] = ~layer3_out[5335];
    assign layer4_out[1845] = layer3_out[1077];
    assign layer4_out[1846] = layer3_out[7447] | layer3_out[7448];
    assign layer4_out[1847] = layer3_out[1960] | layer3_out[1961];
    assign layer4_out[1848] = layer3_out[1502] & ~layer3_out[1503];
    assign layer4_out[1849] = layer3_out[7019];
    assign layer4_out[1850] = ~layer3_out[7439];
    assign layer4_out[1851] = layer3_out[7856];
    assign layer4_out[1852] = layer3_out[2755];
    assign layer4_out[1853] = ~(layer3_out[4245] | layer3_out[4246]);
    assign layer4_out[1854] = layer3_out[3021] & ~layer3_out[3020];
    assign layer4_out[1855] = layer3_out[3026] & layer3_out[3027];
    assign layer4_out[1856] = layer3_out[2384];
    assign layer4_out[1857] = ~layer3_out[4700];
    assign layer4_out[1858] = layer3_out[7153];
    assign layer4_out[1859] = layer3_out[6275];
    assign layer4_out[1860] = layer3_out[5854];
    assign layer4_out[1861] = ~(layer3_out[5330] | layer3_out[5331]);
    assign layer4_out[1862] = layer3_out[1222];
    assign layer4_out[1863] = ~layer3_out[490];
    assign layer4_out[1864] = ~(layer3_out[2064] | layer3_out[2065]);
    assign layer4_out[1865] = ~(layer3_out[3126] ^ layer3_out[3127]);
    assign layer4_out[1866] = layer3_out[3518];
    assign layer4_out[1867] = layer3_out[7631] ^ layer3_out[7632];
    assign layer4_out[1868] = layer3_out[824];
    assign layer4_out[1869] = ~(layer3_out[1428] | layer3_out[1429]);
    assign layer4_out[1870] = layer3_out[3335] ^ layer3_out[3336];
    assign layer4_out[1871] = ~layer3_out[5945];
    assign layer4_out[1872] = layer3_out[4343];
    assign layer4_out[1873] = ~layer3_out[4142] | layer3_out[4143];
    assign layer4_out[1874] = ~layer3_out[1628] | layer3_out[1629];
    assign layer4_out[1875] = ~layer3_out[2662];
    assign layer4_out[1876] = ~layer3_out[2432];
    assign layer4_out[1877] = ~(layer3_out[2830] ^ layer3_out[2831]);
    assign layer4_out[1878] = ~layer3_out[4584] | layer3_out[4585];
    assign layer4_out[1879] = ~layer3_out[7553];
    assign layer4_out[1880] = ~layer3_out[4751] | layer3_out[4752];
    assign layer4_out[1881] = layer3_out[1783] & ~layer3_out[1784];
    assign layer4_out[1882] = ~layer3_out[4194] | layer3_out[4195];
    assign layer4_out[1883] = layer3_out[1123] ^ layer3_out[1124];
    assign layer4_out[1884] = layer3_out[3438];
    assign layer4_out[1885] = ~layer3_out[5101] | layer3_out[5100];
    assign layer4_out[1886] = layer3_out[2378];
    assign layer4_out[1887] = layer3_out[1339];
    assign layer4_out[1888] = ~(layer3_out[4454] & layer3_out[4455]);
    assign layer4_out[1889] = 1'b1;
    assign layer4_out[1890] = layer3_out[2946];
    assign layer4_out[1891] = 1'b0;
    assign layer4_out[1892] = layer3_out[937];
    assign layer4_out[1893] = ~layer3_out[2727];
    assign layer4_out[1894] = 1'b1;
    assign layer4_out[1895] = ~layer3_out[4830];
    assign layer4_out[1896] = ~layer3_out[3435];
    assign layer4_out[1897] = ~(layer3_out[6213] ^ layer3_out[6214]);
    assign layer4_out[1898] = layer3_out[5764] & ~layer3_out[5765];
    assign layer4_out[1899] = layer3_out[103] & ~layer3_out[102];
    assign layer4_out[1900] = layer3_out[4549] ^ layer3_out[4550];
    assign layer4_out[1901] = layer3_out[3446];
    assign layer4_out[1902] = layer3_out[6583];
    assign layer4_out[1903] = ~layer3_out[6964];
    assign layer4_out[1904] = layer3_out[4964];
    assign layer4_out[1905] = layer3_out[835];
    assign layer4_out[1906] = layer3_out[5488] | layer3_out[5489];
    assign layer4_out[1907] = layer3_out[6808] ^ layer3_out[6809];
    assign layer4_out[1908] = layer3_out[5985];
    assign layer4_out[1909] = ~layer3_out[7084];
    assign layer4_out[1910] = layer3_out[7408] | layer3_out[7409];
    assign layer4_out[1911] = layer3_out[4557];
    assign layer4_out[1912] = ~layer3_out[3629];
    assign layer4_out[1913] = ~layer3_out[6070] | layer3_out[6069];
    assign layer4_out[1914] = 1'b0;
    assign layer4_out[1915] = ~(layer3_out[6143] & layer3_out[6144]);
    assign layer4_out[1916] = layer3_out[3263];
    assign layer4_out[1917] = layer3_out[4319] & layer3_out[4320];
    assign layer4_out[1918] = layer3_out[1682];
    assign layer4_out[1919] = layer3_out[2974];
    assign layer4_out[1920] = ~layer3_out[7715];
    assign layer4_out[1921] = layer3_out[5560];
    assign layer4_out[1922] = layer3_out[4784] ^ layer3_out[4785];
    assign layer4_out[1923] = ~layer3_out[4835];
    assign layer4_out[1924] = ~layer3_out[2723];
    assign layer4_out[1925] = layer3_out[631];
    assign layer4_out[1926] = ~layer3_out[2993] | layer3_out[2994];
    assign layer4_out[1927] = layer3_out[7299] ^ layer3_out[7300];
    assign layer4_out[1928] = ~layer3_out[1543];
    assign layer4_out[1929] = layer3_out[6738] & ~layer3_out[6739];
    assign layer4_out[1930] = ~(layer3_out[969] ^ layer3_out[970]);
    assign layer4_out[1931] = layer3_out[6581] ^ layer3_out[6582];
    assign layer4_out[1932] = layer3_out[5930] | layer3_out[5931];
    assign layer4_out[1933] = layer3_out[540] & ~layer3_out[541];
    assign layer4_out[1934] = ~(layer3_out[169] & layer3_out[170]);
    assign layer4_out[1935] = layer3_out[6203];
    assign layer4_out[1936] = layer3_out[3674];
    assign layer4_out[1937] = layer3_out[6449];
    assign layer4_out[1938] = layer3_out[5157] & ~layer3_out[5156];
    assign layer4_out[1939] = ~(layer3_out[1938] ^ layer3_out[1939]);
    assign layer4_out[1940] = ~layer3_out[3373];
    assign layer4_out[1941] = layer3_out[6445] ^ layer3_out[6446];
    assign layer4_out[1942] = ~layer3_out[5601];
    assign layer4_out[1943] = layer3_out[3261];
    assign layer4_out[1944] = layer3_out[7754];
    assign layer4_out[1945] = layer3_out[4619];
    assign layer4_out[1946] = layer3_out[902];
    assign layer4_out[1947] = ~layer3_out[6383];
    assign layer4_out[1948] = ~layer3_out[1440];
    assign layer4_out[1949] = ~layer3_out[5300] | layer3_out[5301];
    assign layer4_out[1950] = ~layer3_out[3464];
    assign layer4_out[1951] = 1'b0;
    assign layer4_out[1952] = ~(layer3_out[5036] ^ layer3_out[5037]);
    assign layer4_out[1953] = ~layer3_out[6557];
    assign layer4_out[1954] = ~(layer3_out[3663] & layer3_out[3664]);
    assign layer4_out[1955] = ~(layer3_out[5880] ^ layer3_out[5881]);
    assign layer4_out[1956] = ~layer3_out[5695];
    assign layer4_out[1957] = ~layer3_out[5277];
    assign layer4_out[1958] = ~layer3_out[1592] | layer3_out[1593];
    assign layer4_out[1959] = ~layer3_out[7130];
    assign layer4_out[1960] = layer3_out[7857] & ~layer3_out[7858];
    assign layer4_out[1961] = ~layer3_out[3084];
    assign layer4_out[1962] = ~(layer3_out[6079] ^ layer3_out[6080]);
    assign layer4_out[1963] = ~(layer3_out[4024] ^ layer3_out[4025]);
    assign layer4_out[1964] = layer3_out[4496];
    assign layer4_out[1965] = layer3_out[3086] | layer3_out[3087];
    assign layer4_out[1966] = layer3_out[2752] ^ layer3_out[2753];
    assign layer4_out[1967] = ~layer3_out[7524];
    assign layer4_out[1968] = ~layer3_out[6026];
    assign layer4_out[1969] = layer3_out[6935];
    assign layer4_out[1970] = layer3_out[7155];
    assign layer4_out[1971] = ~(layer3_out[4663] ^ layer3_out[4664]);
    assign layer4_out[1972] = ~(layer3_out[1778] | layer3_out[1779]);
    assign layer4_out[1973] = ~layer3_out[5194];
    assign layer4_out[1974] = layer3_out[2777] ^ layer3_out[2778];
    assign layer4_out[1975] = layer3_out[7933];
    assign layer4_out[1976] = layer3_out[7861] & ~layer3_out[7860];
    assign layer4_out[1977] = ~layer3_out[1063] | layer3_out[1064];
    assign layer4_out[1978] = layer3_out[1532];
    assign layer4_out[1979] = layer3_out[1287];
    assign layer4_out[1980] = ~layer3_out[2111];
    assign layer4_out[1981] = layer3_out[3769] ^ layer3_out[3770];
    assign layer4_out[1982] = ~layer3_out[31];
    assign layer4_out[1983] = ~layer3_out[7211] | layer3_out[7212];
    assign layer4_out[1984] = layer3_out[2985] & layer3_out[2986];
    assign layer4_out[1985] = layer3_out[1170] ^ layer3_out[1171];
    assign layer4_out[1986] = layer3_out[5807] ^ layer3_out[5808];
    assign layer4_out[1987] = ~layer3_out[7287];
    assign layer4_out[1988] = layer3_out[6173];
    assign layer4_out[1989] = ~layer3_out[7674];
    assign layer4_out[1990] = layer3_out[4249] & ~layer3_out[4248];
    assign layer4_out[1991] = ~layer3_out[955];
    assign layer4_out[1992] = ~layer3_out[267];
    assign layer4_out[1993] = layer3_out[3446];
    assign layer4_out[1994] = layer3_out[2881];
    assign layer4_out[1995] = ~(layer3_out[1817] & layer3_out[1818]);
    assign layer4_out[1996] = ~layer3_out[2637];
    assign layer4_out[1997] = layer3_out[617] | layer3_out[618];
    assign layer4_out[1998] = ~(layer3_out[3903] | layer3_out[3904]);
    assign layer4_out[1999] = layer3_out[2021];
    assign layer4_out[2000] = layer3_out[6967] | layer3_out[6968];
    assign layer4_out[2001] = layer3_out[5611];
    assign layer4_out[2002] = layer3_out[1003] ^ layer3_out[1004];
    assign layer4_out[2003] = ~layer3_out[2406];
    assign layer4_out[2004] = ~(layer3_out[1282] ^ layer3_out[1283]);
    assign layer4_out[2005] = layer3_out[6310] & ~layer3_out[6309];
    assign layer4_out[2006] = ~(layer3_out[1968] & layer3_out[1969]);
    assign layer4_out[2007] = layer3_out[7119] ^ layer3_out[7120];
    assign layer4_out[2008] = ~layer3_out[7424];
    assign layer4_out[2009] = layer3_out[1424];
    assign layer4_out[2010] = layer3_out[1541] ^ layer3_out[1542];
    assign layer4_out[2011] = ~(layer3_out[1231] & layer3_out[1232]);
    assign layer4_out[2012] = ~layer3_out[348] | layer3_out[349];
    assign layer4_out[2013] = ~layer3_out[2140];
    assign layer4_out[2014] = layer3_out[2860] | layer3_out[2861];
    assign layer4_out[2015] = ~layer3_out[1015] | layer3_out[1016];
    assign layer4_out[2016] = ~(layer3_out[4141] | layer3_out[4142]);
    assign layer4_out[2017] = layer3_out[7357] ^ layer3_out[7358];
    assign layer4_out[2018] = layer3_out[1671] ^ layer3_out[1672];
    assign layer4_out[2019] = layer3_out[1437] & ~layer3_out[1438];
    assign layer4_out[2020] = ~layer3_out[7445] | layer3_out[7446];
    assign layer4_out[2021] = layer3_out[2139] & layer3_out[2140];
    assign layer4_out[2022] = layer3_out[6879];
    assign layer4_out[2023] = ~(layer3_out[2728] | layer3_out[2729]);
    assign layer4_out[2024] = ~layer3_out[4511];
    assign layer4_out[2025] = ~layer3_out[5376];
    assign layer4_out[2026] = layer3_out[3013];
    assign layer4_out[2027] = layer3_out[2701] ^ layer3_out[2702];
    assign layer4_out[2028] = ~(layer3_out[7192] & layer3_out[7193]);
    assign layer4_out[2029] = ~layer3_out[6672];
    assign layer4_out[2030] = layer3_out[612] ^ layer3_out[613];
    assign layer4_out[2031] = layer3_out[6646];
    assign layer4_out[2032] = ~layer3_out[2491] | layer3_out[2492];
    assign layer4_out[2033] = layer3_out[7541] & ~layer3_out[7542];
    assign layer4_out[2034] = ~(layer3_out[120] ^ layer3_out[121]);
    assign layer4_out[2035] = ~layer3_out[589];
    assign layer4_out[2036] = layer3_out[4743] & ~layer3_out[4742];
    assign layer4_out[2037] = layer3_out[994];
    assign layer4_out[2038] = ~layer3_out[7888];
    assign layer4_out[2039] = 1'b0;
    assign layer4_out[2040] = ~layer3_out[4862] | layer3_out[4863];
    assign layer4_out[2041] = 1'b0;
    assign layer4_out[2042] = ~(layer3_out[2097] ^ layer3_out[2098]);
    assign layer4_out[2043] = layer3_out[2747];
    assign layer4_out[2044] = layer3_out[7046] & layer3_out[7047];
    assign layer4_out[2045] = layer3_out[3130] | layer3_out[3131];
    assign layer4_out[2046] = ~(layer3_out[3627] | layer3_out[3628]);
    assign layer4_out[2047] = layer3_out[4982] & ~layer3_out[4983];
    assign layer4_out[2048] = layer3_out[3192];
    assign layer4_out[2049] = layer3_out[2803] | layer3_out[2804];
    assign layer4_out[2050] = ~layer3_out[4216] | layer3_out[4217];
    assign layer4_out[2051] = ~(layer3_out[2919] ^ layer3_out[2920]);
    assign layer4_out[2052] = layer3_out[4003] ^ layer3_out[4004];
    assign layer4_out[2053] = ~layer3_out[1859];
    assign layer4_out[2054] = ~(layer3_out[2903] | layer3_out[2904]);
    assign layer4_out[2055] = ~layer3_out[5650] | layer3_out[5651];
    assign layer4_out[2056] = ~layer3_out[1716] | layer3_out[1717];
    assign layer4_out[2057] = layer3_out[3209] ^ layer3_out[3210];
    assign layer4_out[2058] = layer3_out[772];
    assign layer4_out[2059] = ~layer3_out[2387];
    assign layer4_out[2060] = layer3_out[3259] & ~layer3_out[3258];
    assign layer4_out[2061] = layer3_out[3134];
    assign layer4_out[2062] = layer3_out[5784] & ~layer3_out[5785];
    assign layer4_out[2063] = ~layer3_out[7869];
    assign layer4_out[2064] = ~(layer3_out[3828] & layer3_out[3829]);
    assign layer4_out[2065] = layer3_out[4321] & ~layer3_out[4322];
    assign layer4_out[2066] = layer3_out[1754] | layer3_out[1755];
    assign layer4_out[2067] = ~(layer3_out[6336] ^ layer3_out[6337]);
    assign layer4_out[2068] = layer3_out[6048];
    assign layer4_out[2069] = layer3_out[623];
    assign layer4_out[2070] = layer3_out[5009] & ~layer3_out[5010];
    assign layer4_out[2071] = layer3_out[4134] & layer3_out[4135];
    assign layer4_out[2072] = layer3_out[3569] & layer3_out[3570];
    assign layer4_out[2073] = layer3_out[1400];
    assign layer4_out[2074] = layer3_out[3241];
    assign layer4_out[2075] = layer3_out[7055];
    assign layer4_out[2076] = ~layer3_out[5686];
    assign layer4_out[2077] = ~(layer3_out[112] | layer3_out[113]);
    assign layer4_out[2078] = layer3_out[3032] & ~layer3_out[3033];
    assign layer4_out[2079] = 1'b0;
    assign layer4_out[2080] = layer3_out[6365] ^ layer3_out[6366];
    assign layer4_out[2081] = ~layer3_out[1557] | layer3_out[1556];
    assign layer4_out[2082] = ~(layer3_out[2614] & layer3_out[2615]);
    assign layer4_out[2083] = ~(layer3_out[760] ^ layer3_out[761]);
    assign layer4_out[2084] = layer3_out[1887] & layer3_out[1888];
    assign layer4_out[2085] = layer3_out[4641];
    assign layer4_out[2086] = ~(layer3_out[2616] ^ layer3_out[2617]);
    assign layer4_out[2087] = layer3_out[6864] & ~layer3_out[6865];
    assign layer4_out[2088] = ~(layer3_out[6572] ^ layer3_out[6573]);
    assign layer4_out[2089] = layer3_out[7526] ^ layer3_out[7527];
    assign layer4_out[2090] = ~layer3_out[6848];
    assign layer4_out[2091] = layer3_out[5912] & layer3_out[5913];
    assign layer4_out[2092] = layer3_out[4278];
    assign layer4_out[2093] = layer3_out[3130] & ~layer3_out[3129];
    assign layer4_out[2094] = layer3_out[4864] & ~layer3_out[4865];
    assign layer4_out[2095] = layer3_out[7009];
    assign layer4_out[2096] = layer3_out[7401];
    assign layer4_out[2097] = layer3_out[37];
    assign layer4_out[2098] = layer3_out[4124] | layer3_out[4125];
    assign layer4_out[2099] = ~layer3_out[127];
    assign layer4_out[2100] = layer3_out[89] & ~layer3_out[88];
    assign layer4_out[2101] = ~layer3_out[7344] | layer3_out[7343];
    assign layer4_out[2102] = layer3_out[4207] ^ layer3_out[4208];
    assign layer4_out[2103] = ~layer3_out[3271];
    assign layer4_out[2104] = ~(layer3_out[1800] ^ layer3_out[1801]);
    assign layer4_out[2105] = ~(layer3_out[3476] & layer3_out[3477]);
    assign layer4_out[2106] = ~layer3_out[2196] | layer3_out[2195];
    assign layer4_out[2107] = layer3_out[4353];
    assign layer4_out[2108] = ~layer3_out[2196];
    assign layer4_out[2109] = layer3_out[7229] ^ layer3_out[7230];
    assign layer4_out[2110] = ~layer3_out[6340] | layer3_out[6341];
    assign layer4_out[2111] = layer3_out[2933] ^ layer3_out[2934];
    assign layer4_out[2112] = layer3_out[4606] | layer3_out[4607];
    assign layer4_out[2113] = layer3_out[6250] ^ layer3_out[6251];
    assign layer4_out[2114] = ~(layer3_out[1283] ^ layer3_out[1284]);
    assign layer4_out[2115] = layer3_out[1526] & ~layer3_out[1527];
    assign layer4_out[2116] = layer3_out[6795] ^ layer3_out[6796];
    assign layer4_out[2117] = ~layer3_out[1030];
    assign layer4_out[2118] = layer3_out[7378] ^ layer3_out[7379];
    assign layer4_out[2119] = ~layer3_out[2422] | layer3_out[2423];
    assign layer4_out[2120] = ~layer3_out[4882];
    assign layer4_out[2121] = layer3_out[3259];
    assign layer4_out[2122] = ~layer3_out[7350] | layer3_out[7349];
    assign layer4_out[2123] = layer3_out[6297];
    assign layer4_out[2124] = ~layer3_out[7265];
    assign layer4_out[2125] = ~layer3_out[4478];
    assign layer4_out[2126] = layer3_out[7307] & layer3_out[7308];
    assign layer4_out[2127] = ~(layer3_out[4371] ^ layer3_out[4372]);
    assign layer4_out[2128] = ~layer3_out[3460];
    assign layer4_out[2129] = layer3_out[6424] ^ layer3_out[6425];
    assign layer4_out[2130] = ~layer3_out[2717] | layer3_out[2718];
    assign layer4_out[2131] = ~(layer3_out[7346] | layer3_out[7347]);
    assign layer4_out[2132] = ~layer3_out[2148];
    assign layer4_out[2133] = layer3_out[103];
    assign layer4_out[2134] = ~layer3_out[1734];
    assign layer4_out[2135] = layer3_out[1108];
    assign layer4_out[2136] = ~(layer3_out[583] & layer3_out[584]);
    assign layer4_out[2137] = layer3_out[5464];
    assign layer4_out[2138] = layer3_out[4519] | layer3_out[4520];
    assign layer4_out[2139] = ~layer3_out[7597] | layer3_out[7596];
    assign layer4_out[2140] = ~layer3_out[7071];
    assign layer4_out[2141] = ~layer3_out[1477];
    assign layer4_out[2142] = layer3_out[5047];
    assign layer4_out[2143] = ~layer3_out[47];
    assign layer4_out[2144] = ~(layer3_out[6597] ^ layer3_out[6598]);
    assign layer4_out[2145] = ~(layer3_out[4045] ^ layer3_out[4046]);
    assign layer4_out[2146] = ~(layer3_out[3564] ^ layer3_out[3565]);
    assign layer4_out[2147] = ~layer3_out[6031] | layer3_out[6030];
    assign layer4_out[2148] = ~layer3_out[2504] | layer3_out[2505];
    assign layer4_out[2149] = ~layer3_out[7805] | layer3_out[7806];
    assign layer4_out[2150] = layer3_out[796] & ~layer3_out[797];
    assign layer4_out[2151] = layer3_out[4453];
    assign layer4_out[2152] = ~layer3_out[4120];
    assign layer4_out[2153] = ~(layer3_out[2385] | layer3_out[2386]);
    assign layer4_out[2154] = ~layer3_out[6604];
    assign layer4_out[2155] = ~layer3_out[1225];
    assign layer4_out[2156] = ~(layer3_out[1259] | layer3_out[1260]);
    assign layer4_out[2157] = layer3_out[5574];
    assign layer4_out[2158] = ~layer3_out[5242];
    assign layer4_out[2159] = layer3_out[1822] | layer3_out[1823];
    assign layer4_out[2160] = layer3_out[4993];
    assign layer4_out[2161] = ~layer3_out[566];
    assign layer4_out[2162] = ~(layer3_out[4972] & layer3_out[4973]);
    assign layer4_out[2163] = layer3_out[5578];
    assign layer4_out[2164] = ~layer3_out[4237] | layer3_out[4236];
    assign layer4_out[2165] = ~layer3_out[704];
    assign layer4_out[2166] = layer3_out[5998];
    assign layer4_out[2167] = layer3_out[2584];
    assign layer4_out[2168] = layer3_out[2337] ^ layer3_out[2338];
    assign layer4_out[2169] = layer3_out[3386] | layer3_out[3387];
    assign layer4_out[2170] = layer3_out[3985];
    assign layer4_out[2171] = ~(layer3_out[4965] & layer3_out[4966]);
    assign layer4_out[2172] = ~(layer3_out[5731] ^ layer3_out[5732]);
    assign layer4_out[2173] = layer3_out[2660];
    assign layer4_out[2174] = ~(layer3_out[3688] ^ layer3_out[3689]);
    assign layer4_out[2175] = layer3_out[4711] & layer3_out[4712];
    assign layer4_out[2176] = ~layer3_out[6719] | layer3_out[6718];
    assign layer4_out[2177] = layer3_out[4626] ^ layer3_out[4627];
    assign layer4_out[2178] = layer3_out[1185] ^ layer3_out[1186];
    assign layer4_out[2179] = layer3_out[7177] & ~layer3_out[7178];
    assign layer4_out[2180] = ~(layer3_out[1755] ^ layer3_out[1756]);
    assign layer4_out[2181] = layer3_out[2367] ^ layer3_out[2368];
    assign layer4_out[2182] = layer3_out[7428] | layer3_out[7429];
    assign layer4_out[2183] = ~layer3_out[2620];
    assign layer4_out[2184] = layer3_out[6235];
    assign layer4_out[2185] = layer3_out[5063];
    assign layer4_out[2186] = ~(layer3_out[3588] | layer3_out[3589]);
    assign layer4_out[2187] = ~layer3_out[2015];
    assign layer4_out[2188] = ~layer3_out[674] | layer3_out[673];
    assign layer4_out[2189] = layer3_out[940] & layer3_out[941];
    assign layer4_out[2190] = layer3_out[4962] ^ layer3_out[4963];
    assign layer4_out[2191] = ~(layer3_out[7848] | layer3_out[7849]);
    assign layer4_out[2192] = ~layer3_out[1655] | layer3_out[1656];
    assign layer4_out[2193] = ~layer3_out[4989] | layer3_out[4988];
    assign layer4_out[2194] = layer3_out[2206];
    assign layer4_out[2195] = layer3_out[6443] | layer3_out[6444];
    assign layer4_out[2196] = ~layer3_out[3703];
    assign layer4_out[2197] = layer3_out[6972] ^ layer3_out[6973];
    assign layer4_out[2198] = layer3_out[1788] ^ layer3_out[1789];
    assign layer4_out[2199] = ~layer3_out[6362] | layer3_out[6361];
    assign layer4_out[2200] = ~layer3_out[3030] | layer3_out[3031];
    assign layer4_out[2201] = layer3_out[5159] & ~layer3_out[5160];
    assign layer4_out[2202] = ~layer3_out[5491] | layer3_out[5492];
    assign layer4_out[2203] = ~layer3_out[2417] | layer3_out[2418];
    assign layer4_out[2204] = layer3_out[1738] & ~layer3_out[1737];
    assign layer4_out[2205] = ~layer3_out[5680];
    assign layer4_out[2206] = layer3_out[123] & layer3_out[124];
    assign layer4_out[2207] = layer3_out[3394];
    assign layer4_out[2208] = ~layer3_out[3216] | layer3_out[3217];
    assign layer4_out[2209] = ~layer3_out[6909] | layer3_out[6910];
    assign layer4_out[2210] = layer3_out[3225] & ~layer3_out[3224];
    assign layer4_out[2211] = ~layer3_out[31];
    assign layer4_out[2212] = ~layer3_out[4026];
    assign layer4_out[2213] = layer3_out[7670] | layer3_out[7671];
    assign layer4_out[2214] = layer3_out[4171];
    assign layer4_out[2215] = layer3_out[5000] | layer3_out[5001];
    assign layer4_out[2216] = layer3_out[6089] ^ layer3_out[6090];
    assign layer4_out[2217] = ~layer3_out[1883] | layer3_out[1882];
    assign layer4_out[2218] = layer3_out[7509] ^ layer3_out[7510];
    assign layer4_out[2219] = layer3_out[2926];
    assign layer4_out[2220] = ~(layer3_out[5452] ^ layer3_out[5453]);
    assign layer4_out[2221] = layer3_out[1782] & ~layer3_out[1783];
    assign layer4_out[2222] = ~layer3_out[2365] | layer3_out[2366];
    assign layer4_out[2223] = ~layer3_out[3946];
    assign layer4_out[2224] = ~layer3_out[486];
    assign layer4_out[2225] = ~layer3_out[3351];
    assign layer4_out[2226] = ~(layer3_out[208] & layer3_out[209]);
    assign layer4_out[2227] = layer3_out[3760];
    assign layer4_out[2228] = layer3_out[2564];
    assign layer4_out[2229] = ~layer3_out[6119];
    assign layer4_out[2230] = layer3_out[402] & ~layer3_out[403];
    assign layer4_out[2231] = layer3_out[7386] & ~layer3_out[7387];
    assign layer4_out[2232] = layer3_out[7922] ^ layer3_out[7923];
    assign layer4_out[2233] = ~(layer3_out[488] & layer3_out[489]);
    assign layer4_out[2234] = ~(layer3_out[5935] | layer3_out[5936]);
    assign layer4_out[2235] = layer3_out[3888] ^ layer3_out[3889];
    assign layer4_out[2236] = layer3_out[183] & ~layer3_out[182];
    assign layer4_out[2237] = layer3_out[3770] ^ layer3_out[3771];
    assign layer4_out[2238] = layer3_out[3548];
    assign layer4_out[2239] = ~(layer3_out[2593] | layer3_out[2594]);
    assign layer4_out[2240] = layer3_out[6302] & layer3_out[6303];
    assign layer4_out[2241] = layer3_out[3624] & ~layer3_out[3625];
    assign layer4_out[2242] = ~layer3_out[3974] | layer3_out[3975];
    assign layer4_out[2243] = layer3_out[2304] & ~layer3_out[2305];
    assign layer4_out[2244] = layer3_out[4794];
    assign layer4_out[2245] = layer3_out[7223] & ~layer3_out[7224];
    assign layer4_out[2246] = ~layer3_out[7723] | layer3_out[7722];
    assign layer4_out[2247] = ~layer3_out[3995] | layer3_out[3994];
    assign layer4_out[2248] = ~layer3_out[52];
    assign layer4_out[2249] = ~layer3_out[3831] | layer3_out[3830];
    assign layer4_out[2250] = ~layer3_out[7073] | layer3_out[7074];
    assign layer4_out[2251] = ~layer3_out[938] | layer3_out[937];
    assign layer4_out[2252] = ~(layer3_out[7204] ^ layer3_out[7205]);
    assign layer4_out[2253] = ~(layer3_out[5616] ^ layer3_out[5617]);
    assign layer4_out[2254] = layer3_out[4919] | layer3_out[4920];
    assign layer4_out[2255] = layer3_out[4722] | layer3_out[4723];
    assign layer4_out[2256] = layer3_out[6292];
    assign layer4_out[2257] = layer3_out[5909];
    assign layer4_out[2258] = layer3_out[4725] | layer3_out[4726];
    assign layer4_out[2259] = layer3_out[3772] & ~layer3_out[3771];
    assign layer4_out[2260] = layer3_out[7083];
    assign layer4_out[2261] = layer3_out[3706];
    assign layer4_out[2262] = layer3_out[7647];
    assign layer4_out[2263] = ~layer3_out[4572] | layer3_out[4573];
    assign layer4_out[2264] = layer3_out[6329];
    assign layer4_out[2265] = layer3_out[7286] & ~layer3_out[7285];
    assign layer4_out[2266] = ~(layer3_out[4020] & layer3_out[4021]);
    assign layer4_out[2267] = ~layer3_out[3153];
    assign layer4_out[2268] = layer3_out[2176];
    assign layer4_out[2269] = layer3_out[4018] | layer3_out[4019];
    assign layer4_out[2270] = layer3_out[5978];
    assign layer4_out[2271] = layer3_out[4735] & ~layer3_out[4734];
    assign layer4_out[2272] = 1'b1;
    assign layer4_out[2273] = ~(layer3_out[6397] | layer3_out[6398]);
    assign layer4_out[2274] = ~(layer3_out[3677] | layer3_out[3678]);
    assign layer4_out[2275] = layer3_out[5870] & ~layer3_out[5871];
    assign layer4_out[2276] = ~layer3_out[4627];
    assign layer4_out[2277] = ~layer3_out[3576];
    assign layer4_out[2278] = layer3_out[4548] | layer3_out[4549];
    assign layer4_out[2279] = ~layer3_out[3653];
    assign layer4_out[2280] = ~(layer3_out[7276] & layer3_out[7277]);
    assign layer4_out[2281] = ~layer3_out[3472];
    assign layer4_out[2282] = layer3_out[3101];
    assign layer4_out[2283] = layer3_out[4311];
    assign layer4_out[2284] = ~layer3_out[5484] | layer3_out[5485];
    assign layer4_out[2285] = ~layer3_out[7575] | layer3_out[7574];
    assign layer4_out[2286] = ~(layer3_out[5876] ^ layer3_out[5877]);
    assign layer4_out[2287] = layer3_out[7539] ^ layer3_out[7540];
    assign layer4_out[2288] = layer3_out[3833] & ~layer3_out[3832];
    assign layer4_out[2289] = layer3_out[1568] & ~layer3_out[1569];
    assign layer4_out[2290] = layer3_out[2059];
    assign layer4_out[2291] = layer3_out[5229] ^ layer3_out[5230];
    assign layer4_out[2292] = ~layer3_out[7268];
    assign layer4_out[2293] = ~layer3_out[7281] | layer3_out[7280];
    assign layer4_out[2294] = layer3_out[2154] & ~layer3_out[2155];
    assign layer4_out[2295] = layer3_out[7981];
    assign layer4_out[2296] = layer3_out[4349] ^ layer3_out[4350];
    assign layer4_out[2297] = layer3_out[3971] ^ layer3_out[3972];
    assign layer4_out[2298] = ~layer3_out[6139];
    assign layer4_out[2299] = layer3_out[4835] & ~layer3_out[4836];
    assign layer4_out[2300] = ~layer3_out[1462] | layer3_out[1463];
    assign layer4_out[2301] = layer3_out[6261];
    assign layer4_out[2302] = layer3_out[431] ^ layer3_out[432];
    assign layer4_out[2303] = ~layer3_out[6074];
    assign layer4_out[2304] = layer3_out[3486] ^ layer3_out[3487];
    assign layer4_out[2305] = layer3_out[7403];
    assign layer4_out[2306] = ~layer3_out[1598];
    assign layer4_out[2307] = layer3_out[7692] | layer3_out[7693];
    assign layer4_out[2308] = layer3_out[2808];
    assign layer4_out[2309] = layer3_out[1409] ^ layer3_out[1410];
    assign layer4_out[2310] = ~layer3_out[6042] | layer3_out[6043];
    assign layer4_out[2311] = ~layer3_out[1115];
    assign layer4_out[2312] = ~(layer3_out[2274] & layer3_out[2275]);
    assign layer4_out[2313] = ~layer3_out[4596];
    assign layer4_out[2314] = ~layer3_out[2826];
    assign layer4_out[2315] = ~(layer3_out[7778] ^ layer3_out[7779]);
    assign layer4_out[2316] = ~layer3_out[484];
    assign layer4_out[2317] = layer3_out[5013] & ~layer3_out[5014];
    assign layer4_out[2318] = ~(layer3_out[6131] & layer3_out[6132]);
    assign layer4_out[2319] = ~layer3_out[4632] | layer3_out[4633];
    assign layer4_out[2320] = 1'b1;
    assign layer4_out[2321] = layer3_out[7066] & layer3_out[7067];
    assign layer4_out[2322] = ~layer3_out[866];
    assign layer4_out[2323] = layer3_out[3874] ^ layer3_out[3875];
    assign layer4_out[2324] = ~layer3_out[5558];
    assign layer4_out[2325] = ~layer3_out[7585] | layer3_out[7584];
    assign layer4_out[2326] = ~layer3_out[2264] | layer3_out[2265];
    assign layer4_out[2327] = layer3_out[7921];
    assign layer4_out[2328] = layer3_out[1872] | layer3_out[1873];
    assign layer4_out[2329] = layer3_out[7612] ^ layer3_out[7613];
    assign layer4_out[2330] = ~layer3_out[2487] | layer3_out[2486];
    assign layer4_out[2331] = ~(layer3_out[1675] ^ layer3_out[1676]);
    assign layer4_out[2332] = ~layer3_out[2725];
    assign layer4_out[2333] = ~layer3_out[240];
    assign layer4_out[2334] = ~layer3_out[6550];
    assign layer4_out[2335] = layer3_out[999] & ~layer3_out[1000];
    assign layer4_out[2336] = ~layer3_out[5776];
    assign layer4_out[2337] = layer3_out[5547] ^ layer3_out[5548];
    assign layer4_out[2338] = ~layer3_out[7640] | layer3_out[7639];
    assign layer4_out[2339] = ~(layer3_out[2798] ^ layer3_out[2799]);
    assign layer4_out[2340] = layer3_out[21];
    assign layer4_out[2341] = layer3_out[6950] & ~layer3_out[6951];
    assign layer4_out[2342] = layer3_out[6667] & ~layer3_out[6668];
    assign layer4_out[2343] = layer3_out[3614];
    assign layer4_out[2344] = ~(layer3_out[2308] | layer3_out[2309]);
    assign layer4_out[2345] = layer3_out[5559] & ~layer3_out[5558];
    assign layer4_out[2346] = ~layer3_out[7197] | layer3_out[7196];
    assign layer4_out[2347] = layer3_out[1451] | layer3_out[1452];
    assign layer4_out[2348] = layer3_out[2655] | layer3_out[2656];
    assign layer4_out[2349] = ~layer3_out[7373] | layer3_out[7374];
    assign layer4_out[2350] = 1'b0;
    assign layer4_out[2351] = ~(layer3_out[3356] ^ layer3_out[3357]);
    assign layer4_out[2352] = layer3_out[9] ^ layer3_out[10];
    assign layer4_out[2353] = layer3_out[2478];
    assign layer4_out[2354] = layer3_out[1976] & ~layer3_out[1975];
    assign layer4_out[2355] = layer3_out[1858];
    assign layer4_out[2356] = ~(layer3_out[5858] ^ layer3_out[5859]);
    assign layer4_out[2357] = layer3_out[4247] ^ layer3_out[4248];
    assign layer4_out[2358] = ~(layer3_out[4143] ^ layer3_out[4144]);
    assign layer4_out[2359] = layer3_out[6006] | layer3_out[6007];
    assign layer4_out[2360] = layer3_out[6653] ^ layer3_out[6654];
    assign layer4_out[2361] = ~layer3_out[678];
    assign layer4_out[2362] = layer3_out[165] & ~layer3_out[166];
    assign layer4_out[2363] = ~(layer3_out[7969] ^ layer3_out[7970]);
    assign layer4_out[2364] = ~layer3_out[4137];
    assign layer4_out[2365] = layer3_out[868];
    assign layer4_out[2366] = layer3_out[675] & layer3_out[676];
    assign layer4_out[2367] = layer3_out[167] & layer3_out[168];
    assign layer4_out[2368] = layer3_out[1098];
    assign layer4_out[2369] = ~(layer3_out[5419] & layer3_out[5420]);
    assign layer4_out[2370] = layer3_out[6727];
    assign layer4_out[2371] = ~layer3_out[4625];
    assign layer4_out[2372] = ~layer3_out[3969] | layer3_out[3970];
    assign layer4_out[2373] = ~layer3_out[6544];
    assign layer4_out[2374] = layer3_out[366] & ~layer3_out[365];
    assign layer4_out[2375] = layer3_out[2495] ^ layer3_out[2496];
    assign layer4_out[2376] = layer3_out[7897];
    assign layer4_out[2377] = layer3_out[6959];
    assign layer4_out[2378] = ~layer3_out[6982];
    assign layer4_out[2379] = layer3_out[1079] ^ layer3_out[1080];
    assign layer4_out[2380] = layer3_out[3467];
    assign layer4_out[2381] = ~(layer3_out[4105] ^ layer3_out[4106]);
    assign layer4_out[2382] = ~layer3_out[659];
    assign layer4_out[2383] = layer3_out[3825] & layer3_out[3826];
    assign layer4_out[2384] = ~layer3_out[7101];
    assign layer4_out[2385] = ~(layer3_out[4951] | layer3_out[4952]);
    assign layer4_out[2386] = layer3_out[5754];
    assign layer4_out[2387] = ~layer3_out[2828] | layer3_out[2827];
    assign layer4_out[2388] = ~layer3_out[705] | layer3_out[704];
    assign layer4_out[2389] = layer3_out[6512] & ~layer3_out[6511];
    assign layer4_out[2390] = layer3_out[2153];
    assign layer4_out[2391] = ~layer3_out[4778];
    assign layer4_out[2392] = ~(layer3_out[6138] | layer3_out[6139]);
    assign layer4_out[2393] = layer3_out[2738] & ~layer3_out[2739];
    assign layer4_out[2394] = layer3_out[2530] & ~layer3_out[2529];
    assign layer4_out[2395] = layer3_out[2566];
    assign layer4_out[2396] = layer3_out[6499];
    assign layer4_out[2397] = ~layer3_out[7843];
    assign layer4_out[2398] = ~layer3_out[2603];
    assign layer4_out[2399] = ~(layer3_out[1124] ^ layer3_out[1125]);
    assign layer4_out[2400] = ~layer3_out[4872] | layer3_out[4873];
    assign layer4_out[2401] = layer3_out[2813];
    assign layer4_out[2402] = layer3_out[4438] ^ layer3_out[4439];
    assign layer4_out[2403] = layer3_out[6330] ^ layer3_out[6331];
    assign layer4_out[2404] = layer3_out[4265] & layer3_out[4266];
    assign layer4_out[2405] = layer3_out[3153];
    assign layer4_out[2406] = ~layer3_out[252] | layer3_out[251];
    assign layer4_out[2407] = ~(layer3_out[3381] | layer3_out[3382]);
    assign layer4_out[2408] = layer3_out[2191] & ~layer3_out[2190];
    assign layer4_out[2409] = ~(layer3_out[7143] | layer3_out[7144]);
    assign layer4_out[2410] = ~layer3_out[4489];
    assign layer4_out[2411] = ~layer3_out[5192];
    assign layer4_out[2412] = ~layer3_out[4309] | layer3_out[4308];
    assign layer4_out[2413] = layer3_out[1824] & ~layer3_out[1823];
    assign layer4_out[2414] = ~layer3_out[1597];
    assign layer4_out[2415] = ~(layer3_out[5052] & layer3_out[5053]);
    assign layer4_out[2416] = ~(layer3_out[1701] ^ layer3_out[1702]);
    assign layer4_out[2417] = layer3_out[6777] ^ layer3_out[6778];
    assign layer4_out[2418] = layer3_out[7188] & ~layer3_out[7187];
    assign layer4_out[2419] = layer3_out[293] ^ layer3_out[294];
    assign layer4_out[2420] = ~(layer3_out[1080] | layer3_out[1081]);
    assign layer4_out[2421] = ~layer3_out[5199] | layer3_out[5198];
    assign layer4_out[2422] = ~layer3_out[7668];
    assign layer4_out[2423] = layer3_out[6839] | layer3_out[6840];
    assign layer4_out[2424] = ~(layer3_out[1632] | layer3_out[1633]);
    assign layer4_out[2425] = layer3_out[4878] & ~layer3_out[4879];
    assign layer4_out[2426] = ~layer3_out[914] | layer3_out[915];
    assign layer4_out[2427] = ~layer3_out[7098];
    assign layer4_out[2428] = layer3_out[4512] & layer3_out[4513];
    assign layer4_out[2429] = layer3_out[3957] & ~layer3_out[3958];
    assign layer4_out[2430] = ~layer3_out[2456] | layer3_out[2457];
    assign layer4_out[2431] = ~layer3_out[1162];
    assign layer4_out[2432] = layer3_out[2343] ^ layer3_out[2344];
    assign layer4_out[2433] = layer3_out[6503] & ~layer3_out[6502];
    assign layer4_out[2434] = ~layer3_out[4278];
    assign layer4_out[2435] = layer3_out[3928];
    assign layer4_out[2436] = ~layer3_out[2483];
    assign layer4_out[2437] = layer3_out[655];
    assign layer4_out[2438] = layer3_out[5331] ^ layer3_out[5332];
    assign layer4_out[2439] = ~(layer3_out[584] ^ layer3_out[585]);
    assign layer4_out[2440] = ~layer3_out[1546];
    assign layer4_out[2441] = ~(layer3_out[256] | layer3_out[257]);
    assign layer4_out[2442] = ~layer3_out[1200] | layer3_out[1199];
    assign layer4_out[2443] = ~(layer3_out[751] | layer3_out[752]);
    assign layer4_out[2444] = ~layer3_out[7483];
    assign layer4_out[2445] = layer3_out[5203] & ~layer3_out[5204];
    assign layer4_out[2446] = ~(layer3_out[463] ^ layer3_out[464]);
    assign layer4_out[2447] = layer3_out[6936] ^ layer3_out[6937];
    assign layer4_out[2448] = ~layer3_out[7722];
    assign layer4_out[2449] = 1'b0;
    assign layer4_out[2450] = ~layer3_out[3655] | layer3_out[3654];
    assign layer4_out[2451] = layer3_out[3562] & ~layer3_out[3563];
    assign layer4_out[2452] = layer3_out[300] ^ layer3_out[301];
    assign layer4_out[2453] = ~layer3_out[279];
    assign layer4_out[2454] = ~layer3_out[5025];
    assign layer4_out[2455] = layer3_out[5952];
    assign layer4_out[2456] = ~(layer3_out[1256] | layer3_out[1257]);
    assign layer4_out[2457] = ~layer3_out[6480];
    assign layer4_out[2458] = ~layer3_out[79];
    assign layer4_out[2459] = layer3_out[7732] | layer3_out[7733];
    assign layer4_out[2460] = ~(layer3_out[2388] ^ layer3_out[2389]);
    assign layer4_out[2461] = ~(layer3_out[5828] ^ layer3_out[5829]);
    assign layer4_out[2462] = ~layer3_out[6169] | layer3_out[6168];
    assign layer4_out[2463] = ~layer3_out[1685] | layer3_out[1686];
    assign layer4_out[2464] = ~(layer3_out[4237] | layer3_out[4238]);
    assign layer4_out[2465] = layer3_out[3942] | layer3_out[3943];
    assign layer4_out[2466] = layer3_out[5434] & layer3_out[5435];
    assign layer4_out[2467] = layer3_out[4908] & ~layer3_out[4907];
    assign layer4_out[2468] = layer3_out[6147] ^ layer3_out[6148];
    assign layer4_out[2469] = ~layer3_out[5447] | layer3_out[5446];
    assign layer4_out[2470] = layer3_out[2066] & ~layer3_out[2067];
    assign layer4_out[2471] = layer3_out[4395];
    assign layer4_out[2472] = layer3_out[1462];
    assign layer4_out[2473] = ~layer3_out[5210];
    assign layer4_out[2474] = ~layer3_out[7255] | layer3_out[7256];
    assign layer4_out[2475] = layer3_out[2113];
    assign layer4_out[2476] = layer3_out[768] & ~layer3_out[767];
    assign layer4_out[2477] = ~layer3_out[2327] | layer3_out[2328];
    assign layer4_out[2478] = ~(layer3_out[1868] ^ layer3_out[1869]);
    assign layer4_out[2479] = layer3_out[5745] ^ layer3_out[5746];
    assign layer4_out[2480] = layer3_out[2771];
    assign layer4_out[2481] = ~layer3_out[4940];
    assign layer4_out[2482] = ~(layer3_out[1132] & layer3_out[1133]);
    assign layer4_out[2483] = ~(layer3_out[5082] | layer3_out[5083]);
    assign layer4_out[2484] = layer3_out[5469];
    assign layer4_out[2485] = ~layer3_out[5490] | layer3_out[5489];
    assign layer4_out[2486] = ~layer3_out[2932];
    assign layer4_out[2487] = layer3_out[3653];
    assign layer4_out[2488] = layer3_out[1281];
    assign layer4_out[2489] = ~(layer3_out[5118] & layer3_out[5119]);
    assign layer4_out[2490] = ~(layer3_out[736] ^ layer3_out[737]);
    assign layer4_out[2491] = ~layer3_out[1191];
    assign layer4_out[2492] = layer3_out[396];
    assign layer4_out[2493] = ~layer3_out[4598];
    assign layer4_out[2494] = layer3_out[2236] ^ layer3_out[2237];
    assign layer4_out[2495] = layer3_out[863] ^ layer3_out[864];
    assign layer4_out[2496] = ~(layer3_out[4732] ^ layer3_out[4733]);
    assign layer4_out[2497] = ~layer3_out[6288];
    assign layer4_out[2498] = ~layer3_out[2668];
    assign layer4_out[2499] = layer3_out[5490] ^ layer3_out[5491];
    assign layer4_out[2500] = ~layer3_out[4348];
    assign layer4_out[2501] = ~layer3_out[155];
    assign layer4_out[2502] = layer3_out[405] ^ layer3_out[406];
    assign layer4_out[2503] = ~(layer3_out[5520] | layer3_out[5521]);
    assign layer4_out[2504] = ~layer3_out[1260];
    assign layer4_out[2505] = ~layer3_out[3206];
    assign layer4_out[2506] = layer3_out[7011] | layer3_out[7012];
    assign layer4_out[2507] = ~(layer3_out[1935] | layer3_out[1936]);
    assign layer4_out[2508] = layer3_out[217];
    assign layer4_out[2509] = ~layer3_out[1912];
    assign layer4_out[2510] = layer3_out[7017];
    assign layer4_out[2511] = layer3_out[607];
    assign layer4_out[2512] = ~(layer3_out[7911] ^ layer3_out[7912]);
    assign layer4_out[2513] = layer3_out[1358];
    assign layer4_out[2514] = ~(layer3_out[5672] ^ layer3_out[5673]);
    assign layer4_out[2515] = ~(layer3_out[2470] & layer3_out[2471]);
    assign layer4_out[2516] = ~layer3_out[7172] | layer3_out[7171];
    assign layer4_out[2517] = ~(layer3_out[1730] & layer3_out[1731]);
    assign layer4_out[2518] = ~(layer3_out[2687] | layer3_out[2688]);
    assign layer4_out[2519] = layer3_out[5324] & ~layer3_out[5323];
    assign layer4_out[2520] = ~layer3_out[2998] | layer3_out[2997];
    assign layer4_out[2521] = ~(layer3_out[723] & layer3_out[724]);
    assign layer4_out[2522] = ~layer3_out[3455];
    assign layer4_out[2523] = ~(layer3_out[1454] ^ layer3_out[1455]);
    assign layer4_out[2524] = ~(layer3_out[5965] | layer3_out[5966]);
    assign layer4_out[2525] = ~layer3_out[2400] | layer3_out[2399];
    assign layer4_out[2526] = layer3_out[2652];
    assign layer4_out[2527] = ~layer3_out[2506];
    assign layer4_out[2528] = ~layer3_out[819] | layer3_out[818];
    assign layer4_out[2529] = layer3_out[5529];
    assign layer4_out[2530] = layer3_out[5857] & layer3_out[5858];
    assign layer4_out[2531] = 1'b0;
    assign layer4_out[2532] = layer3_out[3573] & layer3_out[3574];
    assign layer4_out[2533] = ~layer3_out[7146];
    assign layer4_out[2534] = layer3_out[5070] | layer3_out[5071];
    assign layer4_out[2535] = layer3_out[6255] ^ layer3_out[6256];
    assign layer4_out[2536] = ~(layer3_out[6259] ^ layer3_out[6260]);
    assign layer4_out[2537] = ~layer3_out[1988];
    assign layer4_out[2538] = layer3_out[5012] | layer3_out[5013];
    assign layer4_out[2539] = ~(layer3_out[3260] ^ layer3_out[3261]);
    assign layer4_out[2540] = layer3_out[4942] ^ layer3_out[4943];
    assign layer4_out[2541] = ~(layer3_out[3665] ^ layer3_out[3666]);
    assign layer4_out[2542] = layer3_out[1030];
    assign layer4_out[2543] = ~layer3_out[6645];
    assign layer4_out[2544] = layer3_out[5515];
    assign layer4_out[2545] = ~(layer3_out[6614] | layer3_out[6615]);
    assign layer4_out[2546] = ~(layer3_out[2371] ^ layer3_out[2372]);
    assign layer4_out[2547] = ~layer3_out[7780] | layer3_out[7781];
    assign layer4_out[2548] = ~layer3_out[7964];
    assign layer4_out[2549] = ~layer3_out[2003] | layer3_out[2002];
    assign layer4_out[2550] = layer3_out[3668] & layer3_out[3669];
    assign layer4_out[2551] = ~(layer3_out[7862] ^ layer3_out[7863]);
    assign layer4_out[2552] = layer3_out[7118] & layer3_out[7119];
    assign layer4_out[2553] = layer3_out[773];
    assign layer4_out[2554] = layer3_out[825];
    assign layer4_out[2555] = ~layer3_out[155];
    assign layer4_out[2556] = ~(layer3_out[7815] & layer3_out[7816]);
    assign layer4_out[2557] = layer3_out[787];
    assign layer4_out[2558] = layer3_out[4256];
    assign layer4_out[2559] = ~layer3_out[7015];
    assign layer4_out[2560] = layer3_out[3693] ^ layer3_out[3694];
    assign layer4_out[2561] = layer3_out[1361] & ~layer3_out[1360];
    assign layer4_out[2562] = ~layer3_out[5815];
    assign layer4_out[2563] = layer3_out[6812] & ~layer3_out[6813];
    assign layer4_out[2564] = layer3_out[4276] ^ layer3_out[4277];
    assign layer4_out[2565] = ~layer3_out[7369];
    assign layer4_out[2566] = ~(layer3_out[4869] & layer3_out[4870]);
    assign layer4_out[2567] = layer3_out[2788] | layer3_out[2789];
    assign layer4_out[2568] = layer3_out[6108] ^ layer3_out[6109];
    assign layer4_out[2569] = ~layer3_out[4242];
    assign layer4_out[2570] = ~(layer3_out[1825] & layer3_out[1826]);
    assign layer4_out[2571] = ~layer3_out[7194];
    assign layer4_out[2572] = layer3_out[7609] & ~layer3_out[7608];
    assign layer4_out[2573] = ~layer3_out[4449];
    assign layer4_out[2574] = layer3_out[413];
    assign layer4_out[2575] = ~layer3_out[3321];
    assign layer4_out[2576] = ~layer3_out[3620] | layer3_out[3619];
    assign layer4_out[2577] = ~layer3_out[4019];
    assign layer4_out[2578] = layer3_out[3778];
    assign layer4_out[2579] = ~layer3_out[5407];
    assign layer4_out[2580] = layer3_out[5622] ^ layer3_out[5623];
    assign layer4_out[2581] = 1'b0;
    assign layer4_out[2582] = ~(layer3_out[6126] ^ layer3_out[6127]);
    assign layer4_out[2583] = ~layer3_out[5345] | layer3_out[5344];
    assign layer4_out[2584] = ~layer3_out[4990];
    assign layer4_out[2585] = ~layer3_out[6121] | layer3_out[6120];
    assign layer4_out[2586] = ~layer3_out[6109];
    assign layer4_out[2587] = ~(layer3_out[2492] ^ layer3_out[2493]);
    assign layer4_out[2588] = layer3_out[162];
    assign layer4_out[2589] = layer3_out[5924] & ~layer3_out[5925];
    assign layer4_out[2590] = ~layer3_out[1234];
    assign layer4_out[2591] = ~layer3_out[3659];
    assign layer4_out[2592] = ~layer3_out[770];
    assign layer4_out[2593] = ~layer3_out[5903];
    assign layer4_out[2594] = layer3_out[5059];
    assign layer4_out[2595] = ~layer3_out[5264];
    assign layer4_out[2596] = ~layer3_out[1483];
    assign layer4_out[2597] = ~layer3_out[1239];
    assign layer4_out[2598] = ~(layer3_out[7948] ^ layer3_out[7949]);
    assign layer4_out[2599] = ~(layer3_out[1102] ^ layer3_out[1103]);
    assign layer4_out[2600] = layer3_out[3419];
    assign layer4_out[2601] = layer3_out[3561] & layer3_out[3562];
    assign layer4_out[2602] = ~(layer3_out[4693] | layer3_out[4694]);
    assign layer4_out[2603] = layer3_out[792] ^ layer3_out[793];
    assign layer4_out[2604] = ~(layer3_out[6396] ^ layer3_out[6397]);
    assign layer4_out[2605] = 1'b0;
    assign layer4_out[2606] = ~(layer3_out[5212] ^ layer3_out[5213]);
    assign layer4_out[2607] = ~layer3_out[6633];
    assign layer4_out[2608] = layer3_out[2189] & layer3_out[2190];
    assign layer4_out[2609] = ~layer3_out[2177];
    assign layer4_out[2610] = ~layer3_out[7305] | layer3_out[7304];
    assign layer4_out[2611] = layer3_out[6944];
    assign layer4_out[2612] = ~layer3_out[5130];
    assign layer4_out[2613] = ~layer3_out[7598] | layer3_out[7599];
    assign layer4_out[2614] = layer3_out[3058] & layer3_out[3059];
    assign layer4_out[2615] = ~layer3_out[6953] | layer3_out[6952];
    assign layer4_out[2616] = ~layer3_out[6932] | layer3_out[6931];
    assign layer4_out[2617] = layer3_out[7993];
    assign layer4_out[2618] = ~layer3_out[5972] | layer3_out[5973];
    assign layer4_out[2619] = layer3_out[282] & layer3_out[283];
    assign layer4_out[2620] = layer3_out[5538] ^ layer3_out[5539];
    assign layer4_out[2621] = layer3_out[1884];
    assign layer4_out[2622] = layer3_out[3289] & ~layer3_out[3290];
    assign layer4_out[2623] = ~layer3_out[6854];
    assign layer4_out[2624] = ~layer3_out[837];
    assign layer4_out[2625] = layer3_out[3632] ^ layer3_out[3633];
    assign layer4_out[2626] = ~layer3_out[7981];
    assign layer4_out[2627] = layer3_out[5222] & ~layer3_out[5223];
    assign layer4_out[2628] = layer3_out[3909];
    assign layer4_out[2629] = ~layer3_out[350];
    assign layer4_out[2630] = layer3_out[467] & ~layer3_out[468];
    assign layer4_out[2631] = layer3_out[2952] ^ layer3_out[2953];
    assign layer4_out[2632] = layer3_out[7677];
    assign layer4_out[2633] = ~(layer3_out[5915] ^ layer3_out[5916]);
    assign layer4_out[2634] = ~layer3_out[7733];
    assign layer4_out[2635] = ~layer3_out[968];
    assign layer4_out[2636] = layer3_out[2115] & ~layer3_out[2114];
    assign layer4_out[2637] = layer3_out[6644];
    assign layer4_out[2638] = layer3_out[1468] & ~layer3_out[1467];
    assign layer4_out[2639] = layer3_out[2341];
    assign layer4_out[2640] = layer3_out[2700] & layer3_out[2701];
    assign layer4_out[2641] = ~layer3_out[3121];
    assign layer4_out[2642] = layer3_out[7742] & layer3_out[7743];
    assign layer4_out[2643] = ~layer3_out[4822];
    assign layer4_out[2644] = ~(layer3_out[2074] ^ layer3_out[2075]);
    assign layer4_out[2645] = ~layer3_out[4095];
    assign layer4_out[2646] = layer3_out[3879] | layer3_out[3880];
    assign layer4_out[2647] = layer3_out[1429] | layer3_out[1430];
    assign layer4_out[2648] = layer3_out[5058] & ~layer3_out[5059];
    assign layer4_out[2649] = layer3_out[3938];
    assign layer4_out[2650] = layer3_out[3501] ^ layer3_out[3502];
    assign layer4_out[2651] = layer3_out[4099] & ~layer3_out[4100];
    assign layer4_out[2652] = ~(layer3_out[6836] & layer3_out[6837]);
    assign layer4_out[2653] = ~layer3_out[4883] | layer3_out[4882];
    assign layer4_out[2654] = layer3_out[1349] & ~layer3_out[1348];
    assign layer4_out[2655] = ~layer3_out[7719];
    assign layer4_out[2656] = ~(layer3_out[6698] ^ layer3_out[6699]);
    assign layer4_out[2657] = layer3_out[5803] & layer3_out[5804];
    assign layer4_out[2658] = layer3_out[2517] | layer3_out[2518];
    assign layer4_out[2659] = layer3_out[7121] & layer3_out[7122];
    assign layer4_out[2660] = ~layer3_out[561] | layer3_out[560];
    assign layer4_out[2661] = ~(layer3_out[3367] | layer3_out[3368]);
    assign layer4_out[2662] = ~(layer3_out[5040] | layer3_out[5041]);
    assign layer4_out[2663] = ~layer3_out[874] | layer3_out[875];
    assign layer4_out[2664] = layer3_out[6828] & ~layer3_out[6827];
    assign layer4_out[2665] = ~(layer3_out[2874] ^ layer3_out[2875]);
    assign layer4_out[2666] = ~layer3_out[399];
    assign layer4_out[2667] = ~layer3_out[7889];
    assign layer4_out[2668] = ~(layer3_out[5278] ^ layer3_out[5279]);
    assign layer4_out[2669] = layer3_out[384] & ~layer3_out[385];
    assign layer4_out[2670] = layer3_out[7356];
    assign layer4_out[2671] = layer3_out[5166] & layer3_out[5167];
    assign layer4_out[2672] = layer3_out[187] | layer3_out[188];
    assign layer4_out[2673] = layer3_out[3405];
    assign layer4_out[2674] = ~(layer3_out[6207] & layer3_out[6208]);
    assign layer4_out[2675] = ~layer3_out[4088] | layer3_out[4089];
    assign layer4_out[2676] = layer3_out[132] ^ layer3_out[133];
    assign layer4_out[2677] = layer3_out[1953] & layer3_out[1954];
    assign layer4_out[2678] = layer3_out[6650] & ~layer3_out[6651];
    assign layer4_out[2679] = layer3_out[7156] ^ layer3_out[7157];
    assign layer4_out[2680] = ~layer3_out[7326];
    assign layer4_out[2681] = ~layer3_out[4895];
    assign layer4_out[2682] = ~layer3_out[3977];
    assign layer4_out[2683] = layer3_out[3490] ^ layer3_out[3491];
    assign layer4_out[2684] = ~(layer3_out[4300] ^ layer3_out[4301]);
    assign layer4_out[2685] = ~(layer3_out[4386] & layer3_out[4387]);
    assign layer4_out[2686] = ~layer3_out[3194] | layer3_out[3193];
    assign layer4_out[2687] = ~layer3_out[3568];
    assign layer4_out[2688] = layer3_out[2631];
    assign layer4_out[2689] = layer3_out[1244];
    assign layer4_out[2690] = ~(layer3_out[1078] ^ layer3_out[1079]);
    assign layer4_out[2691] = ~(layer3_out[1835] ^ layer3_out[1836]);
    assign layer4_out[2692] = layer3_out[3745];
    assign layer4_out[2693] = ~layer3_out[7774];
    assign layer4_out[2694] = ~layer3_out[991];
    assign layer4_out[2695] = layer3_out[5867];
    assign layer4_out[2696] = layer3_out[110];
    assign layer4_out[2697] = layer3_out[1911];
    assign layer4_out[2698] = ~layer3_out[2589];
    assign layer4_out[2699] = layer3_out[1838] & ~layer3_out[1837];
    assign layer4_out[2700] = layer3_out[5951];
    assign layer4_out[2701] = layer3_out[3773];
    assign layer4_out[2702] = ~layer3_out[2579];
    assign layer4_out[2703] = ~layer3_out[4471] | layer3_out[4472];
    assign layer4_out[2704] = layer3_out[6762];
    assign layer4_out[2705] = ~(layer3_out[746] ^ layer3_out[747]);
    assign layer4_out[2706] = layer3_out[7859];
    assign layer4_out[2707] = layer3_out[1629];
    assign layer4_out[2708] = layer3_out[3807] | layer3_out[3808];
    assign layer4_out[2709] = ~layer3_out[431];
    assign layer4_out[2710] = layer3_out[5934];
    assign layer4_out[2711] = layer3_out[7466] | layer3_out[7467];
    assign layer4_out[2712] = layer3_out[5492];
    assign layer4_out[2713] = layer3_out[1189];
    assign layer4_out[2714] = layer3_out[2862] & layer3_out[2863];
    assign layer4_out[2715] = ~layer3_out[5445];
    assign layer4_out[2716] = ~(layer3_out[3822] & layer3_out[3823]);
    assign layer4_out[2717] = ~layer3_out[1713];
    assign layer4_out[2718] = layer3_out[1734] & ~layer3_out[1733];
    assign layer4_out[2719] = 1'b0;
    assign layer4_out[2720] = ~layer3_out[6594];
    assign layer4_out[2721] = ~(layer3_out[5010] ^ layer3_out[5011]);
    assign layer4_out[2722] = ~layer3_out[4270];
    assign layer4_out[2723] = ~layer3_out[5937];
    assign layer4_out[2724] = ~layer3_out[4905];
    assign layer4_out[2725] = layer3_out[4275] | layer3_out[4276];
    assign layer4_out[2726] = ~layer3_out[4317];
    assign layer4_out[2727] = layer3_out[1078] & ~layer3_out[1077];
    assign layer4_out[2728] = layer3_out[6560];
    assign layer4_out[2729] = ~(layer3_out[691] & layer3_out[692]);
    assign layer4_out[2730] = ~(layer3_out[2953] & layer3_out[2954]);
    assign layer4_out[2731] = layer3_out[7312];
    assign layer4_out[2732] = layer3_out[5178] & ~layer3_out[5179];
    assign layer4_out[2733] = ~layer3_out[1301];
    assign layer4_out[2734] = ~layer3_out[482];
    assign layer4_out[2735] = ~(layer3_out[4158] | layer3_out[4159]);
    assign layer4_out[2736] = ~(layer3_out[1867] ^ layer3_out[1868]);
    assign layer4_out[2737] = ~layer3_out[5412] | layer3_out[5411];
    assign layer4_out[2738] = ~layer3_out[5549];
    assign layer4_out[2739] = layer3_out[6676];
    assign layer4_out[2740] = layer3_out[3477] & layer3_out[3478];
    assign layer4_out[2741] = ~layer3_out[7194];
    assign layer4_out[2742] = ~(layer3_out[6282] & layer3_out[6283]);
    assign layer4_out[2743] = layer3_out[3948] ^ layer3_out[3949];
    assign layer4_out[2744] = layer3_out[4291] & layer3_out[4292];
    assign layer4_out[2745] = ~layer3_out[7076] | layer3_out[7077];
    assign layer4_out[2746] = layer3_out[6367] & ~layer3_out[6368];
    assign layer4_out[2747] = ~(layer3_out[5204] ^ layer3_out[5205]);
    assign layer4_out[2748] = ~(layer3_out[5634] | layer3_out[5635]);
    assign layer4_out[2749] = layer3_out[4210] & ~layer3_out[4209];
    assign layer4_out[2750] = ~layer3_out[3437];
    assign layer4_out[2751] = layer3_out[2897];
    assign layer4_out[2752] = ~layer3_out[3814] | layer3_out[3815];
    assign layer4_out[2753] = layer3_out[3353] & ~layer3_out[3354];
    assign layer4_out[2754] = ~(layer3_out[5350] | layer3_out[5351]);
    assign layer4_out[2755] = layer3_out[6428];
    assign layer4_out[2756] = layer3_out[4082] ^ layer3_out[4083];
    assign layer4_out[2757] = layer3_out[7300];
    assign layer4_out[2758] = layer3_out[1669] ^ layer3_out[1670];
    assign layer4_out[2759] = layer3_out[2079];
    assign layer4_out[2760] = ~(layer3_out[2164] ^ layer3_out[2165]);
    assign layer4_out[2761] = ~layer3_out[400];
    assign layer4_out[2762] = layer3_out[7005];
    assign layer4_out[2763] = ~layer3_out[4827];
    assign layer4_out[2764] = ~(layer3_out[4837] | layer3_out[4838]);
    assign layer4_out[2765] = layer3_out[3885] & ~layer3_out[3884];
    assign layer4_out[2766] = layer3_out[2310] ^ layer3_out[2311];
    assign layer4_out[2767] = ~layer3_out[6214];
    assign layer4_out[2768] = layer3_out[828];
    assign layer4_out[2769] = layer3_out[4126];
    assign layer4_out[2770] = ~(layer3_out[3531] ^ layer3_out[3532]);
    assign layer4_out[2771] = layer3_out[6201];
    assign layer4_out[2772] = layer3_out[6982] & layer3_out[6983];
    assign layer4_out[2773] = layer3_out[7238] ^ layer3_out[7239];
    assign layer4_out[2774] = ~(layer3_out[7001] | layer3_out[7002]);
    assign layer4_out[2775] = layer3_out[1459];
    assign layer4_out[2776] = layer3_out[1722] & layer3_out[1723];
    assign layer4_out[2777] = layer3_out[6455];
    assign layer4_out[2778] = layer3_out[4956] | layer3_out[4957];
    assign layer4_out[2779] = ~layer3_out[744] | layer3_out[743];
    assign layer4_out[2780] = ~(layer3_out[3724] | layer3_out[3725]);
    assign layer4_out[2781] = ~(layer3_out[224] ^ layer3_out[225]);
    assign layer4_out[2782] = ~layer3_out[6458];
    assign layer4_out[2783] = layer3_out[2647] & layer3_out[2648];
    assign layer4_out[2784] = layer3_out[119];
    assign layer4_out[2785] = ~layer3_out[6334] | layer3_out[6335];
    assign layer4_out[2786] = layer3_out[6804] & ~layer3_out[6803];
    assign layer4_out[2787] = ~layer3_out[6877];
    assign layer4_out[2788] = layer3_out[1095] | layer3_out[1096];
    assign layer4_out[2789] = ~(layer3_out[2950] ^ layer3_out[2951]);
    assign layer4_out[2790] = layer3_out[5556];
    assign layer4_out[2791] = ~layer3_out[3682];
    assign layer4_out[2792] = layer3_out[6816];
    assign layer4_out[2793] = layer3_out[6014] & ~layer3_out[6013];
    assign layer4_out[2794] = layer3_out[6374] ^ layer3_out[6375];
    assign layer4_out[2795] = ~(layer3_out[7170] | layer3_out[7171]);
    assign layer4_out[2796] = ~(layer3_out[606] ^ layer3_out[607]);
    assign layer4_out[2797] = layer3_out[2443];
    assign layer4_out[2798] = ~(layer3_out[5080] ^ layer3_out[5081]);
    assign layer4_out[2799] = layer3_out[2544] | layer3_out[2545];
    assign layer4_out[2800] = layer3_out[5604];
    assign layer4_out[2801] = ~(layer3_out[504] ^ layer3_out[505]);
    assign layer4_out[2802] = layer3_out[594];
    assign layer4_out[2803] = ~layer3_out[4010] | layer3_out[4009];
    assign layer4_out[2804] = ~layer3_out[6766];
    assign layer4_out[2805] = layer3_out[7314] ^ layer3_out[7315];
    assign layer4_out[2806] = layer3_out[7200];
    assign layer4_out[2807] = ~(layer3_out[7176] | layer3_out[7177]);
    assign layer4_out[2808] = layer3_out[949];
    assign layer4_out[2809] = layer3_out[69] ^ layer3_out[70];
    assign layer4_out[2810] = ~layer3_out[4748];
    assign layer4_out[2811] = ~layer3_out[1643];
    assign layer4_out[2812] = layer3_out[3005] & ~layer3_out[3004];
    assign layer4_out[2813] = layer3_out[909] & ~layer3_out[910];
    assign layer4_out[2814] = layer3_out[4724] ^ layer3_out[4725];
    assign layer4_out[2815] = ~layer3_out[553];
    assign layer4_out[2816] = ~(layer3_out[1775] & layer3_out[1776]);
    assign layer4_out[2817] = layer3_out[2184] | layer3_out[2185];
    assign layer4_out[2818] = layer3_out[4705] & ~layer3_out[4706];
    assign layer4_out[2819] = ~(layer3_out[6920] & layer3_out[6921]);
    assign layer4_out[2820] = ~(layer3_out[1478] ^ layer3_out[1479]);
    assign layer4_out[2821] = layer3_out[1327] & ~layer3_out[1326];
    assign layer4_out[2822] = layer3_out[3715];
    assign layer4_out[2823] = layer3_out[7822] ^ layer3_out[7823];
    assign layer4_out[2824] = layer3_out[5763] & ~layer3_out[5762];
    assign layer4_out[2825] = layer3_out[4564];
    assign layer4_out[2826] = ~(layer3_out[5030] | layer3_out[5031]);
    assign layer4_out[2827] = layer3_out[6505];
    assign layer4_out[2828] = layer3_out[6731];
    assign layer4_out[2829] = layer3_out[2102] ^ layer3_out[2103];
    assign layer4_out[2830] = layer3_out[3118];
    assign layer4_out[2831] = ~layer3_out[6014] | layer3_out[6015];
    assign layer4_out[2832] = ~(layer3_out[4846] & layer3_out[4847]);
    assign layer4_out[2833] = ~layer3_out[7458] | layer3_out[7459];
    assign layer4_out[2834] = ~layer3_out[3665] | layer3_out[3664];
    assign layer4_out[2835] = layer3_out[891] & ~layer3_out[890];
    assign layer4_out[2836] = ~(layer3_out[7865] | layer3_out[7866]);
    assign layer4_out[2837] = ~layer3_out[3735] | layer3_out[3736];
    assign layer4_out[2838] = ~(layer3_out[1019] | layer3_out[1020]);
    assign layer4_out[2839] = ~layer3_out[667];
    assign layer4_out[2840] = ~(layer3_out[6888] ^ layer3_out[6889]);
    assign layer4_out[2841] = layer3_out[7951] ^ layer3_out[7952];
    assign layer4_out[2842] = ~(layer3_out[7502] ^ layer3_out[7503]);
    assign layer4_out[2843] = ~layer3_out[1790] | layer3_out[1791];
    assign layer4_out[2844] = layer3_out[7545] & ~layer3_out[7544];
    assign layer4_out[2845] = layer3_out[2233] & ~layer3_out[2232];
    assign layer4_out[2846] = ~layer3_out[381];
    assign layer4_out[2847] = ~(layer3_out[1408] & layer3_out[1409]);
    assign layer4_out[2848] = layer3_out[3449];
    assign layer4_out[2849] = layer3_out[2858] ^ layer3_out[2859];
    assign layer4_out[2850] = ~layer3_out[5833] | layer3_out[5832];
    assign layer4_out[2851] = layer3_out[1798] ^ layer3_out[1799];
    assign layer4_out[2852] = layer3_out[54] | layer3_out[55];
    assign layer4_out[2853] = ~(layer3_out[5327] ^ layer3_out[5328]);
    assign layer4_out[2854] = layer3_out[7949];
    assign layer4_out[2855] = ~layer3_out[242] | layer3_out[241];
    assign layer4_out[2856] = ~(layer3_out[2242] & layer3_out[2243]);
    assign layer4_out[2857] = ~layer3_out[442];
    assign layer4_out[2858] = ~layer3_out[2606];
    assign layer4_out[2859] = layer3_out[7243] & ~layer3_out[7244];
    assign layer4_out[2860] = ~layer3_out[6754] | layer3_out[6755];
    assign layer4_out[2861] = layer3_out[2038] & ~layer3_out[2039];
    assign layer4_out[2862] = ~layer3_out[7488] | layer3_out[7487];
    assign layer4_out[2863] = layer3_out[7039];
    assign layer4_out[2864] = layer3_out[6918];
    assign layer4_out[2865] = ~layer3_out[1388];
    assign layer4_out[2866] = layer3_out[7614] & ~layer3_out[7613];
    assign layer4_out[2867] = ~layer3_out[1015] | layer3_out[1014];
    assign layer4_out[2868] = ~(layer3_out[5802] | layer3_out[5803]);
    assign layer4_out[2869] = ~layer3_out[1318] | layer3_out[1317];
    assign layer4_out[2870] = ~layer3_out[6765] | layer3_out[6766];
    assign layer4_out[2871] = layer3_out[2323] ^ layer3_out[2324];
    assign layer4_out[2872] = layer3_out[5872];
    assign layer4_out[2873] = layer3_out[6829];
    assign layer4_out[2874] = ~layer3_out[5502];
    assign layer4_out[2875] = layer3_out[5443] & layer3_out[5444];
    assign layer4_out[2876] = layer3_out[6489] ^ layer3_out[6490];
    assign layer4_out[2877] = ~(layer3_out[3178] | layer3_out[3179]);
    assign layer4_out[2878] = ~layer3_out[1705];
    assign layer4_out[2879] = ~layer3_out[3048] | layer3_out[3047];
    assign layer4_out[2880] = ~layer3_out[7152];
    assign layer4_out[2881] = ~layer3_out[6311];
    assign layer4_out[2882] = layer3_out[7768];
    assign layer4_out[2883] = layer3_out[5732] ^ layer3_out[5733];
    assign layer4_out[2884] = ~(layer3_out[7800] ^ layer3_out[7801]);
    assign layer4_out[2885] = layer3_out[2689];
    assign layer4_out[2886] = ~layer3_out[4209];
    assign layer4_out[2887] = layer3_out[6084] ^ layer3_out[6085];
    assign layer4_out[2888] = layer3_out[2149] & ~layer3_out[2150];
    assign layer4_out[2889] = ~(layer3_out[3542] ^ layer3_out[3543]);
    assign layer4_out[2890] = ~layer3_out[212];
    assign layer4_out[2891] = layer3_out[2148] & ~layer3_out[2147];
    assign layer4_out[2892] = ~layer3_out[1623] | layer3_out[1622];
    assign layer4_out[2893] = ~layer3_out[4956] | layer3_out[4955];
    assign layer4_out[2894] = ~(layer3_out[6372] ^ layer3_out[6373]);
    assign layer4_out[2895] = ~layer3_out[173];
    assign layer4_out[2896] = ~layer3_out[1799];
    assign layer4_out[2897] = ~layer3_out[1749];
    assign layer4_out[2898] = layer3_out[6066] & ~layer3_out[6065];
    assign layer4_out[2899] = layer3_out[3327];
    assign layer4_out[2900] = ~(layer3_out[383] | layer3_out[384]);
    assign layer4_out[2901] = layer3_out[1802] ^ layer3_out[1803];
    assign layer4_out[2902] = ~layer3_out[4772];
    assign layer4_out[2903] = ~(layer3_out[4948] ^ layer3_out[4949]);
    assign layer4_out[2904] = layer3_out[5735] & layer3_out[5736];
    assign layer4_out[2905] = ~layer3_out[3415];
    assign layer4_out[2906] = ~(layer3_out[7052] & layer3_out[7053]);
    assign layer4_out[2907] = ~layer3_out[1319];
    assign layer4_out[2908] = layer3_out[2509] & ~layer3_out[2510];
    assign layer4_out[2909] = layer3_out[1519];
    assign layer4_out[2910] = ~(layer3_out[5251] ^ layer3_out[5252]);
    assign layer4_out[2911] = ~layer3_out[1624];
    assign layer4_out[2912] = ~(layer3_out[4432] ^ layer3_out[4433]);
    assign layer4_out[2913] = ~(layer3_out[6062] | layer3_out[6063]);
    assign layer4_out[2914] = layer3_out[6181] ^ layer3_out[6182];
    assign layer4_out[2915] = layer3_out[321] | layer3_out[322];
    assign layer4_out[2916] = layer3_out[19] & ~layer3_out[20];
    assign layer4_out[2917] = ~layer3_out[3905];
    assign layer4_out[2918] = ~layer3_out[377];
    assign layer4_out[2919] = layer3_out[7272];
    assign layer4_out[2920] = ~layer3_out[1938];
    assign layer4_out[2921] = ~(layer3_out[6005] | layer3_out[6006]);
    assign layer4_out[2922] = layer3_out[7427];
    assign layer4_out[2923] = ~(layer3_out[5586] ^ layer3_out[5587]);
    assign layer4_out[2924] = ~(layer3_out[1242] ^ layer3_out[1243]);
    assign layer4_out[2925] = layer3_out[2019];
    assign layer4_out[2926] = ~layer3_out[567] | layer3_out[568];
    assign layer4_out[2927] = layer3_out[7946];
    assign layer4_out[2928] = layer3_out[3550] & ~layer3_out[3551];
    assign layer4_out[2929] = ~(layer3_out[2773] ^ layer3_out[2774]);
    assign layer4_out[2930] = layer3_out[2301] ^ layer3_out[2302];
    assign layer4_out[2931] = layer3_out[220] | layer3_out[221];
    assign layer4_out[2932] = ~layer3_out[5261];
    assign layer4_out[2933] = layer3_out[6918] & ~layer3_out[6919];
    assign layer4_out[2934] = layer3_out[3536];
    assign layer4_out[2935] = layer3_out[4857];
    assign layer4_out[2936] = layer3_out[4600] | layer3_out[4601];
    assign layer4_out[2937] = layer3_out[4812];
    assign layer4_out[2938] = ~(layer3_out[1424] ^ layer3_out[1425]);
    assign layer4_out[2939] = layer3_out[6743];
    assign layer4_out[2940] = layer3_out[2970] & ~layer3_out[2969];
    assign layer4_out[2941] = ~layer3_out[3282];
    assign layer4_out[2942] = ~layer3_out[1092];
    assign layer4_out[2943] = ~layer3_out[4386] | layer3_out[4385];
    assign layer4_out[2944] = ~layer3_out[7670];
    assign layer4_out[2945] = layer3_out[7153];
    assign layer4_out[2946] = layer3_out[2561] ^ layer3_out[2562];
    assign layer4_out[2947] = layer3_out[7575] | layer3_out[7576];
    assign layer4_out[2948] = 1'b1;
    assign layer4_out[2949] = ~(layer3_out[5707] ^ layer3_out[5708]);
    assign layer4_out[2950] = layer3_out[1415] & ~layer3_out[1414];
    assign layer4_out[2951] = layer3_out[2111];
    assign layer4_out[2952] = layer3_out[3170];
    assign layer4_out[2953] = ~layer3_out[1990];
    assign layer4_out[2954] = layer3_out[2686];
    assign layer4_out[2955] = ~layer3_out[659];
    assign layer4_out[2956] = ~(layer3_out[6854] & layer3_out[6855]);
    assign layer4_out[2957] = ~layer3_out[7181];
    assign layer4_out[2958] = layer3_out[5730] & ~layer3_out[5731];
    assign layer4_out[2959] = layer3_out[6999] | layer3_out[7000];
    assign layer4_out[2960] = ~(layer3_out[4655] & layer3_out[4656]);
    assign layer4_out[2961] = ~layer3_out[2363];
    assign layer4_out[2962] = layer3_out[911];
    assign layer4_out[2963] = ~layer3_out[2871];
    assign layer4_out[2964] = 1'b1;
    assign layer4_out[2965] = layer3_out[6023];
    assign layer4_out[2966] = ~(layer3_out[5183] | layer3_out[5184]);
    assign layer4_out[2967] = layer3_out[3809] ^ layer3_out[3810];
    assign layer4_out[2968] = ~layer3_out[3244];
    assign layer4_out[2969] = ~layer3_out[7604] | layer3_out[7605];
    assign layer4_out[2970] = ~layer3_out[7274] | layer3_out[7273];
    assign layer4_out[2971] = layer3_out[478] ^ layer3_out[479];
    assign layer4_out[2972] = ~layer3_out[1608] | layer3_out[1607];
    assign layer4_out[2973] = ~(layer3_out[4104] ^ layer3_out[4105]);
    assign layer4_out[2974] = ~layer3_out[5322];
    assign layer4_out[2975] = layer3_out[7989] ^ layer3_out[7990];
    assign layer4_out[2976] = ~(layer3_out[1505] & layer3_out[1506]);
    assign layer4_out[2977] = layer3_out[3710] & ~layer3_out[3711];
    assign layer4_out[2978] = ~layer3_out[6991];
    assign layer4_out[2979] = ~(layer3_out[4945] & layer3_out[4946]);
    assign layer4_out[2980] = ~layer3_out[1976] | layer3_out[1977];
    assign layer4_out[2981] = layer3_out[6002] ^ layer3_out[6003];
    assign layer4_out[2982] = layer3_out[7682];
    assign layer4_out[2983] = ~layer3_out[6253];
    assign layer4_out[2984] = layer3_out[4760];
    assign layer4_out[2985] = layer3_out[2431];
    assign layer4_out[2986] = layer3_out[7469] & ~layer3_out[7468];
    assign layer4_out[2987] = ~(layer3_out[5420] & layer3_out[5421]);
    assign layer4_out[2988] = ~layer3_out[4082] | layer3_out[4081];
    assign layer4_out[2989] = layer3_out[5400];
    assign layer4_out[2990] = layer3_out[6610] ^ layer3_out[6611];
    assign layer4_out[2991] = ~layer3_out[6953];
    assign layer4_out[2992] = ~layer3_out[3466];
    assign layer4_out[2993] = layer3_out[2710];
    assign layer4_out[2994] = ~layer3_out[1380];
    assign layer4_out[2995] = layer3_out[4888];
    assign layer4_out[2996] = ~(layer3_out[1862] & layer3_out[1863]);
    assign layer4_out[2997] = ~(layer3_out[5913] ^ layer3_out[5914]);
    assign layer4_out[2998] = ~layer3_out[1573];
    assign layer4_out[2999] = layer3_out[4070] ^ layer3_out[4071];
    assign layer4_out[3000] = ~layer3_out[4615] | layer3_out[4614];
    assign layer4_out[3001] = layer3_out[7479];
    assign layer4_out[3002] = layer3_out[7050] ^ layer3_out[7051];
    assign layer4_out[3003] = ~layer3_out[3127] | layer3_out[3128];
    assign layer4_out[3004] = ~layer3_out[2335];
    assign layer4_out[3005] = layer3_out[6729] ^ layer3_out[6730];
    assign layer4_out[3006] = layer3_out[4057] ^ layer3_out[4058];
    assign layer4_out[3007] = layer3_out[759] & ~layer3_out[758];
    assign layer4_out[3008] = layer3_out[4210] ^ layer3_out[4211];
    assign layer4_out[3009] = ~(layer3_out[2480] ^ layer3_out[2481]);
    assign layer4_out[3010] = layer3_out[5978];
    assign layer4_out[3011] = layer3_out[1359] | layer3_out[1360];
    assign layer4_out[3012] = layer3_out[3290] ^ layer3_out[3291];
    assign layer4_out[3013] = ~(layer3_out[2550] ^ layer3_out[2551]);
    assign layer4_out[3014] = layer3_out[1369] & ~layer3_out[1370];
    assign layer4_out[3015] = layer3_out[1875];
    assign layer4_out[3016] = ~layer3_out[4746];
    assign layer4_out[3017] = layer3_out[6837];
    assign layer4_out[3018] = layer3_out[2441];
    assign layer4_out[3019] = ~layer3_out[5393];
    assign layer4_out[3020] = ~layer3_out[3371];
    assign layer4_out[3021] = ~layer3_out[4524];
    assign layer4_out[3022] = ~(layer3_out[3254] ^ layer3_out[3255]);
    assign layer4_out[3023] = 1'b1;
    assign layer4_out[3024] = ~layer3_out[5284];
    assign layer4_out[3025] = layer3_out[4768];
    assign layer4_out[3026] = layer3_out[1748];
    assign layer4_out[3027] = ~(layer3_out[6937] | layer3_out[6938]);
    assign layer4_out[3028] = layer3_out[3171] ^ layer3_out[3172];
    assign layer4_out[3029] = ~(layer3_out[6588] | layer3_out[6589]);
    assign layer4_out[3030] = layer3_out[2926];
    assign layer4_out[3031] = layer3_out[2570] ^ layer3_out[2571];
    assign layer4_out[3032] = layer3_out[2052] ^ layer3_out[2053];
    assign layer4_out[3033] = ~(layer3_out[4973] ^ layer3_out[4974]);
    assign layer4_out[3034] = ~layer3_out[161];
    assign layer4_out[3035] = ~layer3_out[7770];
    assign layer4_out[3036] = ~layer3_out[6205];
    assign layer4_out[3037] = layer3_out[2984] ^ layer3_out[2985];
    assign layer4_out[3038] = ~(layer3_out[2003] | layer3_out[2004]);
    assign layer4_out[3039] = layer3_out[7209] | layer3_out[7210];
    assign layer4_out[3040] = layer3_out[34] ^ layer3_out[35];
    assign layer4_out[3041] = layer3_out[117] | layer3_out[118];
    assign layer4_out[3042] = ~layer3_out[902] | layer3_out[901];
    assign layer4_out[3043] = layer3_out[7633] | layer3_out[7634];
    assign layer4_out[3044] = layer3_out[2512];
    assign layer4_out[3045] = ~layer3_out[1894];
    assign layer4_out[3046] = layer3_out[1443] & ~layer3_out[1444];
    assign layer4_out[3047] = ~layer3_out[5561] | layer3_out[5560];
    assign layer4_out[3048] = layer3_out[4755] & ~layer3_out[4754];
    assign layer4_out[3049] = layer3_out[4596];
    assign layer4_out[3050] = layer3_out[7288] ^ layer3_out[7289];
    assign layer4_out[3051] = layer3_out[1623] ^ layer3_out[1624];
    assign layer4_out[3052] = ~layer3_out[7701];
    assign layer4_out[3053] = layer3_out[2490];
    assign layer4_out[3054] = layer3_out[5258];
    assign layer4_out[3055] = ~layer3_out[4836];
    assign layer4_out[3056] = ~(layer3_out[5808] | layer3_out[5809]);
    assign layer4_out[3057] = layer3_out[3238] ^ layer3_out[3239];
    assign layer4_out[3058] = layer3_out[5055] | layer3_out[5056];
    assign layer4_out[3059] = layer3_out[4689] | layer3_out[4690];
    assign layer4_out[3060] = ~layer3_out[1890];
    assign layer4_out[3061] = layer3_out[7725] | layer3_out[7726];
    assign layer4_out[3062] = layer3_out[1178] | layer3_out[1179];
    assign layer4_out[3063] = ~layer3_out[4922];
    assign layer4_out[3064] = ~layer3_out[1878];
    assign layer4_out[3065] = ~layer3_out[7318];
    assign layer4_out[3066] = layer3_out[5264] ^ layer3_out[5265];
    assign layer4_out[3067] = ~layer3_out[2550];
    assign layer4_out[3068] = ~layer3_out[3120];
    assign layer4_out[3069] = layer3_out[4205] ^ layer3_out[4206];
    assign layer4_out[3070] = layer3_out[4400];
    assign layer4_out[3071] = layer3_out[5478] & layer3_out[5479];
    assign layer4_out[3072] = layer3_out[4983] & layer3_out[4984];
    assign layer4_out[3073] = layer3_out[5337];
    assign layer4_out[3074] = layer3_out[4720];
    assign layer4_out[3075] = ~layer3_out[2181];
    assign layer4_out[3076] = layer3_out[7925] & ~layer3_out[7926];
    assign layer4_out[3077] = ~(layer3_out[6327] ^ layer3_out[6328]);
    assign layer4_out[3078] = ~layer3_out[7165] | layer3_out[7166];
    assign layer4_out[3079] = layer3_out[2473] & ~layer3_out[2474];
    assign layer4_out[3080] = ~layer3_out[6483] | layer3_out[6484];
    assign layer4_out[3081] = layer3_out[1372] ^ layer3_out[1373];
    assign layer4_out[3082] = layer3_out[4877];
    assign layer4_out[3083] = ~(layer3_out[6876] & layer3_out[6877]);
    assign layer4_out[3084] = layer3_out[4891] & ~layer3_out[4890];
    assign layer4_out[3085] = layer3_out[6828] ^ layer3_out[6829];
    assign layer4_out[3086] = layer3_out[7080] ^ layer3_out[7081];
    assign layer4_out[3087] = layer3_out[3386];
    assign layer4_out[3088] = ~layer3_out[7062];
    assign layer4_out[3089] = ~layer3_out[5780] | layer3_out[5779];
    assign layer4_out[3090] = layer3_out[5023];
    assign layer4_out[3091] = layer3_out[5053];
    assign layer4_out[3092] = ~layer3_out[2269];
    assign layer4_out[3093] = layer3_out[2582] ^ layer3_out[2583];
    assign layer4_out[3094] = ~layer3_out[274] | layer3_out[275];
    assign layer4_out[3095] = layer3_out[4244] & layer3_out[4245];
    assign layer4_out[3096] = ~layer3_out[3];
    assign layer4_out[3097] = ~layer3_out[14] | layer3_out[15];
    assign layer4_out[3098] = layer3_out[5635] & layer3_out[5636];
    assign layer4_out[3099] = ~layer3_out[3941];
    assign layer4_out[3100] = ~(layer3_out[4889] & layer3_out[4890]);
    assign layer4_out[3101] = layer3_out[6418];
    assign layer4_out[3102] = ~layer3_out[7020];
    assign layer4_out[3103] = ~(layer3_out[3886] ^ layer3_out[3887]);
    assign layer4_out[3104] = layer3_out[4333];
    assign layer4_out[3105] = ~(layer3_out[3854] | layer3_out[3855]);
    assign layer4_out[3106] = layer3_out[5986] ^ layer3_out[5987];
    assign layer4_out[3107] = layer3_out[4294];
    assign layer4_out[3108] = layer3_out[6473];
    assign layer4_out[3109] = ~layer3_out[4748];
    assign layer4_out[3110] = ~layer3_out[587];
    assign layer4_out[3111] = ~layer3_out[5780];
    assign layer4_out[3112] = layer3_out[5340] & ~layer3_out[5339];
    assign layer4_out[3113] = ~(layer3_out[2177] ^ layer3_out[2178]);
    assign layer4_out[3114] = layer3_out[433] & ~layer3_out[432];
    assign layer4_out[3115] = layer3_out[5190] & layer3_out[5191];
    assign layer4_out[3116] = layer3_out[502] | layer3_out[503];
    assign layer4_out[3117] = ~layer3_out[4900];
    assign layer4_out[3118] = ~layer3_out[4098] | layer3_out[4099];
    assign layer4_out[3119] = ~layer3_out[2797];
    assign layer4_out[3120] = ~(layer3_out[1842] ^ layer3_out[1843]);
    assign layer4_out[3121] = ~layer3_out[7562] | layer3_out[7563];
    assign layer4_out[3122] = ~layer3_out[2618];
    assign layer4_out[3123] = layer3_out[1764] | layer3_out[1765];
    assign layer4_out[3124] = layer3_out[776];
    assign layer4_out[3125] = ~layer3_out[713];
    assign layer4_out[3126] = layer3_out[1892] ^ layer3_out[1893];
    assign layer4_out[3127] = 1'b1;
    assign layer4_out[3128] = ~(layer3_out[5927] ^ layer3_out[5928]);
    assign layer4_out[3129] = ~layer3_out[4937] | layer3_out[4938];
    assign layer4_out[3130] = ~(layer3_out[2248] ^ layer3_out[2249]);
    assign layer4_out[3131] = ~layer3_out[5970];
    assign layer4_out[3132] = layer3_out[7228] & ~layer3_out[7229];
    assign layer4_out[3133] = ~layer3_out[1515] | layer3_out[1514];
    assign layer4_out[3134] = layer3_out[5818] ^ layer3_out[5819];
    assign layer4_out[3135] = layer3_out[5513] & ~layer3_out[5514];
    assign layer4_out[3136] = ~(layer3_out[4286] ^ layer3_out[4287]);
    assign layer4_out[3137] = layer3_out[7698] & layer3_out[7699];
    assign layer4_out[3138] = layer3_out[5942];
    assign layer4_out[3139] = layer3_out[1980] & ~layer3_out[1979];
    assign layer4_out[3140] = layer3_out[4888];
    assign layer4_out[3141] = ~layer3_out[3678];
    assign layer4_out[3142] = layer3_out[7061] & ~layer3_out[7062];
    assign layer4_out[3143] = ~(layer3_out[3818] | layer3_out[3819]);
    assign layer4_out[3144] = ~(layer3_out[6969] ^ layer3_out[6970]);
    assign layer4_out[3145] = ~layer3_out[2150];
    assign layer4_out[3146] = layer3_out[6656];
    assign layer4_out[3147] = layer3_out[801] & ~layer3_out[800];
    assign layer4_out[3148] = layer3_out[3147];
    assign layer4_out[3149] = ~(layer3_out[333] | layer3_out[334]);
    assign layer4_out[3150] = ~layer3_out[481] | layer3_out[480];
    assign layer4_out[3151] = ~(layer3_out[761] & layer3_out[762]);
    assign layer4_out[3152] = ~(layer3_out[5410] | layer3_out[5411]);
    assign layer4_out[3153] = layer3_out[2999] & layer3_out[3000];
    assign layer4_out[3154] = layer3_out[2682] & ~layer3_out[2681];
    assign layer4_out[3155] = layer3_out[1951] & layer3_out[1952];
    assign layer4_out[3156] = ~(layer3_out[144] ^ layer3_out[145]);
    assign layer4_out[3157] = layer3_out[1571] & ~layer3_out[1572];
    assign layer4_out[3158] = layer3_out[5463] & ~layer3_out[5462];
    assign layer4_out[3159] = ~layer3_out[1466] | layer3_out[1467];
    assign layer4_out[3160] = ~layer3_out[1088];
    assign layer4_out[3161] = layer3_out[3475];
    assign layer4_out[3162] = ~layer3_out[4069] | layer3_out[4070];
    assign layer4_out[3163] = layer3_out[80];
    assign layer4_out[3164] = ~layer3_out[6291] | layer3_out[6290];
    assign layer4_out[3165] = layer3_out[511] | layer3_out[512];
    assign layer4_out[3166] = layer3_out[832] ^ layer3_out[833];
    assign layer4_out[3167] = ~(layer3_out[7971] ^ layer3_out[7972]);
    assign layer4_out[3168] = ~(layer3_out[3191] ^ layer3_out[3192]);
    assign layer4_out[3169] = layer3_out[627];
    assign layer4_out[3170] = layer3_out[6039] & ~layer3_out[6040];
    assign layer4_out[3171] = ~(layer3_out[268] ^ layer3_out[269]);
    assign layer4_out[3172] = layer3_out[2134] ^ layer3_out[2135];
    assign layer4_out[3173] = ~layer3_out[4188];
    assign layer4_out[3174] = layer3_out[601];
    assign layer4_out[3175] = ~layer3_out[4590] | layer3_out[4589];
    assign layer4_out[3176] = ~layer3_out[2665];
    assign layer4_out[3177] = layer3_out[1995] & ~layer3_out[1996];
    assign layer4_out[3178] = layer3_out[1862] & ~layer3_out[1861];
    assign layer4_out[3179] = ~layer3_out[7820];
    assign layer4_out[3180] = layer3_out[5543];
    assign layer4_out[3181] = ~layer3_out[1330];
    assign layer4_out[3182] = layer3_out[6283] & layer3_out[6284];
    assign layer4_out[3183] = ~layer3_out[1212];
    assign layer4_out[3184] = layer3_out[4611];
    assign layer4_out[3185] = layer3_out[391] & layer3_out[392];
    assign layer4_out[3186] = layer3_out[1631] & ~layer3_out[1630];
    assign layer4_out[3187] = layer3_out[5799];
    assign layer4_out[3188] = layer3_out[528] | layer3_out[529];
    assign layer4_out[3189] = ~(layer3_out[2912] | layer3_out[2913]);
    assign layer4_out[3190] = ~layer3_out[48];
    assign layer4_out[3191] = ~(layer3_out[329] ^ layer3_out[330]);
    assign layer4_out[3192] = layer3_out[1269];
    assign layer4_out[3193] = layer3_out[312];
    assign layer4_out[3194] = ~layer3_out[5286] | layer3_out[5287];
    assign layer4_out[3195] = ~layer3_out[6938];
    assign layer4_out[3196] = ~(layer3_out[5705] ^ layer3_out[5706]);
    assign layer4_out[3197] = ~layer3_out[1355];
    assign layer4_out[3198] = ~layer3_out[7157];
    assign layer4_out[3199] = layer3_out[4155] & layer3_out[4156];
    assign layer4_out[3200] = ~layer3_out[6136];
    assign layer4_out[3201] = layer3_out[6008] ^ layer3_out[6009];
    assign layer4_out[3202] = layer3_out[5594] ^ layer3_out[5595];
    assign layer4_out[3203] = 1'b1;
    assign layer4_out[3204] = layer3_out[7142] ^ layer3_out[7143];
    assign layer4_out[3205] = layer3_out[4456];
    assign layer4_out[3206] = layer3_out[7215];
    assign layer4_out[3207] = ~(layer3_out[7060] & layer3_out[7061]);
    assign layer4_out[3208] = layer3_out[4718] ^ layer3_out[4719];
    assign layer4_out[3209] = ~layer3_out[3152] | layer3_out[3151];
    assign layer4_out[3210] = layer3_out[6315] | layer3_out[6316];
    assign layer4_out[3211] = layer3_out[5122];
    assign layer4_out[3212] = ~(layer3_out[7326] & layer3_out[7327]);
    assign layer4_out[3213] = ~layer3_out[2646];
    assign layer4_out[3214] = ~(layer3_out[1127] | layer3_out[1128]);
    assign layer4_out[3215] = ~layer3_out[7739];
    assign layer4_out[3216] = layer3_out[1558] & ~layer3_out[1559];
    assign layer4_out[3217] = layer3_out[6564];
    assign layer4_out[3218] = layer3_out[3493] | layer3_out[3494];
    assign layer4_out[3219] = layer3_out[4951];
    assign layer4_out[3220] = ~(layer3_out[7781] & layer3_out[7782]);
    assign layer4_out[3221] = layer3_out[3913] & layer3_out[3914];
    assign layer4_out[3222] = ~(layer3_out[3530] ^ layer3_out[3531]);
    assign layer4_out[3223] = ~layer3_out[4604];
    assign layer4_out[3224] = layer3_out[2783];
    assign layer4_out[3225] = ~layer3_out[2879];
    assign layer4_out[3226] = layer3_out[1649];
    assign layer4_out[3227] = layer3_out[4337] ^ layer3_out[4338];
    assign layer4_out[3228] = layer3_out[6338] & ~layer3_out[6339];
    assign layer4_out[3229] = ~(layer3_out[5063] ^ layer3_out[5064]);
    assign layer4_out[3230] = layer3_out[7237] & layer3_out[7238];
    assign layer4_out[3231] = ~(layer3_out[4239] ^ layer3_out[4240]);
    assign layer4_out[3232] = ~layer3_out[994];
    assign layer4_out[3233] = layer3_out[6794] ^ layer3_out[6795];
    assign layer4_out[3234] = ~layer3_out[6267];
    assign layer4_out[3235] = layer3_out[4858];
    assign layer4_out[3236] = 1'b1;
    assign layer4_out[3237] = layer3_out[5220] ^ layer3_out[5221];
    assign layer4_out[3238] = ~layer3_out[3849];
    assign layer4_out[3239] = layer3_out[457] & ~layer3_out[456];
    assign layer4_out[3240] = layer3_out[7106] | layer3_out[7107];
    assign layer4_out[3241] = layer3_out[6506] & ~layer3_out[6507];
    assign layer4_out[3242] = ~(layer3_out[7407] ^ layer3_out[7408]);
    assign layer4_out[3243] = layer3_out[1828] & ~layer3_out[1829];
    assign layer4_out[3244] = layer3_out[7794] ^ layer3_out[7795];
    assign layer4_out[3245] = layer3_out[5067] & ~layer3_out[5066];
    assign layer4_out[3246] = ~layer3_out[7310];
    assign layer4_out[3247] = ~layer3_out[7195];
    assign layer4_out[3248] = layer3_out[4381] & ~layer3_out[4382];
    assign layer4_out[3249] = ~(layer3_out[3444] & layer3_out[3445]);
    assign layer4_out[3250] = ~(layer3_out[4350] & layer3_out[4351]);
    assign layer4_out[3251] = layer3_out[3255];
    assign layer4_out[3252] = ~layer3_out[3612];
    assign layer4_out[3253] = layer3_out[440] | layer3_out[441];
    assign layer4_out[3254] = layer3_out[991] & ~layer3_out[990];
    assign layer4_out[3255] = ~layer3_out[1376];
    assign layer4_out[3256] = layer3_out[291] & ~layer3_out[290];
    assign layer4_out[3257] = layer3_out[2890] | layer3_out[2891];
    assign layer4_out[3258] = layer3_out[1594] ^ layer3_out[1595];
    assign layer4_out[3259] = ~layer3_out[1889];
    assign layer4_out[3260] = layer3_out[834];
    assign layer4_out[3261] = ~layer3_out[1294];
    assign layer4_out[3262] = ~layer3_out[955];
    assign layer4_out[3263] = ~(layer3_out[2330] & layer3_out[2331]);
    assign layer4_out[3264] = layer3_out[7851];
    assign layer4_out[3265] = ~layer3_out[5158];
    assign layer4_out[3266] = ~(layer3_out[5213] ^ layer3_out[5214]);
    assign layer4_out[3267] = layer3_out[3589] ^ layer3_out[3590];
    assign layer4_out[3268] = layer3_out[7881];
    assign layer4_out[3269] = layer3_out[951];
    assign layer4_out[3270] = ~layer3_out[4521] | layer3_out[4520];
    assign layer4_out[3271] = layer3_out[4036] & layer3_out[4037];
    assign layer4_out[3272] = layer3_out[2467];
    assign layer4_out[3273] = ~layer3_out[1073];
    assign layer4_out[3274] = layer3_out[2475] & ~layer3_out[2474];
    assign layer4_out[3275] = ~(layer3_out[6957] & layer3_out[6958]);
    assign layer4_out[3276] = layer3_out[3139];
    assign layer4_out[3277] = layer3_out[4686] ^ layer3_out[4687];
    assign layer4_out[3278] = layer3_out[4252] ^ layer3_out[4253];
    assign layer4_out[3279] = ~layer3_out[4122];
    assign layer4_out[3280] = layer3_out[2006];
    assign layer4_out[3281] = ~layer3_out[3247] | layer3_out[3248];
    assign layer4_out[3282] = layer3_out[7257];
    assign layer4_out[3283] = layer3_out[4602] ^ layer3_out[4603];
    assign layer4_out[3284] = layer3_out[156] & layer3_out[157];
    assign layer4_out[3285] = layer3_out[637] & ~layer3_out[638];
    assign layer4_out[3286] = ~layer3_out[3811];
    assign layer4_out[3287] = layer3_out[7461];
    assign layer4_out[3288] = layer3_out[1710] & layer3_out[1711];
    assign layer4_out[3289] = layer3_out[3204];
    assign layer4_out[3290] = layer3_out[1159] & ~layer3_out[1160];
    assign layer4_out[3291] = layer3_out[3838] & ~layer3_out[3837];
    assign layer4_out[3292] = layer3_out[7257] & ~layer3_out[7258];
    assign layer4_out[3293] = ~layer3_out[6730] | layer3_out[6731];
    assign layer4_out[3294] = layer3_out[1786];
    assign layer4_out[3295] = ~(layer3_out[4980] | layer3_out[4981]);
    assign layer4_out[3296] = ~layer3_out[2733];
    assign layer4_out[3297] = layer3_out[5806] & ~layer3_out[5807];
    assign layer4_out[3298] = ~layer3_out[4554];
    assign layer4_out[3299] = layer3_out[5472];
    assign layer4_out[3300] = ~(layer3_out[133] | layer3_out[134]);
    assign layer4_out[3301] = layer3_out[1400] ^ layer3_out[1401];
    assign layer4_out[3302] = ~layer3_out[7662] | layer3_out[7661];
    assign layer4_out[3303] = layer3_out[255] & ~layer3_out[254];
    assign layer4_out[3304] = layer3_out[7864];
    assign layer4_out[3305] = layer3_out[2732];
    assign layer4_out[3306] = layer3_out[1970] & layer3_out[1971];
    assign layer4_out[3307] = layer3_out[2067] & ~layer3_out[2068];
    assign layer4_out[3308] = ~layer3_out[6648] | layer3_out[6647];
    assign layer4_out[3309] = layer3_out[5298] | layer3_out[5299];
    assign layer4_out[3310] = ~layer3_out[5996];
    assign layer4_out[3311] = layer3_out[5144] ^ layer3_out[5145];
    assign layer4_out[3312] = layer3_out[6956];
    assign layer4_out[3313] = ~(layer3_out[2906] | layer3_out[2907]);
    assign layer4_out[3314] = layer3_out[7330];
    assign layer4_out[3315] = ~(layer3_out[3725] ^ layer3_out[3726]);
    assign layer4_out[3316] = layer3_out[5661] | layer3_out[5662];
    assign layer4_out[3317] = ~layer3_out[852] | layer3_out[853];
    assign layer4_out[3318] = layer3_out[1117] & ~layer3_out[1116];
    assign layer4_out[3319] = ~layer3_out[7094] | layer3_out[7095];
    assign layer4_out[3320] = ~layer3_out[3792];
    assign layer4_out[3321] = layer3_out[4558] & ~layer3_out[4559];
    assign layer4_out[3322] = layer3_out[7725];
    assign layer4_out[3323] = ~layer3_out[5210] | layer3_out[5209];
    assign layer4_out[3324] = ~(layer3_out[5919] ^ layer3_out[5920]);
    assign layer4_out[3325] = ~(layer3_out[5320] & layer3_out[5321]);
    assign layer4_out[3326] = ~layer3_out[7803];
    assign layer4_out[3327] = ~layer3_out[4102] | layer3_out[4103];
    assign layer4_out[3328] = layer3_out[1746] | layer3_out[1747];
    assign layer4_out[3329] = layer3_out[5375];
    assign layer4_out[3330] = layer3_out[5624];
    assign layer4_out[3331] = ~layer3_out[1606] | layer3_out[1605];
    assign layer4_out[3332] = ~layer3_out[418];
    assign layer4_out[3333] = layer3_out[4993];
    assign layer4_out[3334] = layer3_out[4859] | layer3_out[4860];
    assign layer4_out[3335] = ~layer3_out[3672] | layer3_out[3671];
    assign layer4_out[3336] = ~(layer3_out[3951] ^ layer3_out[3952]);
    assign layer4_out[3337] = layer3_out[42] | layer3_out[43];
    assign layer4_out[3338] = layer3_out[1579];
    assign layer4_out[3339] = layer3_out[4424];
    assign layer4_out[3340] = ~layer3_out[6716] | layer3_out[6715];
    assign layer4_out[3341] = ~layer3_out[1312];
    assign layer4_out[3342] = layer3_out[1187] & ~layer3_out[1188];
    assign layer4_out[3343] = ~layer3_out[4756] | layer3_out[4755];
    assign layer4_out[3344] = ~layer3_out[3931] | layer3_out[3932];
    assign layer4_out[3345] = layer3_out[4491];
    assign layer4_out[3346] = layer3_out[3777] & ~layer3_out[3776];
    assign layer4_out[3347] = layer3_out[7672] | layer3_out[7673];
    assign layer4_out[3348] = ~layer3_out[3062] | layer3_out[3063];
    assign layer4_out[3349] = ~layer3_out[5449];
    assign layer4_out[3350] = layer3_out[6834] | layer3_out[6835];
    assign layer4_out[3351] = layer3_out[7529];
    assign layer4_out[3352] = layer3_out[2049] & layer3_out[2050];
    assign layer4_out[3353] = layer3_out[3947];
    assign layer4_out[3354] = layer3_out[1335];
    assign layer4_out[3355] = ~(layer3_out[3310] ^ layer3_out[3311]);
    assign layer4_out[3356] = layer3_out[1853] & layer3_out[1854];
    assign layer4_out[3357] = ~layer3_out[3456];
    assign layer4_out[3358] = layer3_out[2799] & layer3_out[2800];
    assign layer4_out[3359] = ~layer3_out[1816];
    assign layer4_out[3360] = layer3_out[3731] | layer3_out[3732];
    assign layer4_out[3361] = layer3_out[7916];
    assign layer4_out[3362] = layer3_out[5563] | layer3_out[5564];
    assign layer4_out[3363] = layer3_out[2393] ^ layer3_out[2394];
    assign layer4_out[3364] = layer3_out[7757] & ~layer3_out[7758];
    assign layer4_out[3365] = ~(layer3_out[7297] ^ layer3_out[7298]);
    assign layer4_out[3366] = 1'b0;
    assign layer4_out[3367] = ~layer3_out[6153] | layer3_out[6152];
    assign layer4_out[3368] = ~(layer3_out[2072] | layer3_out[2073]);
    assign layer4_out[3369] = layer3_out[2747] | layer3_out[2748];
    assign layer4_out[3370] = ~(layer3_out[3473] ^ layer3_out[3474]);
    assign layer4_out[3371] = layer3_out[1523] ^ layer3_out[1524];
    assign layer4_out[3372] = ~layer3_out[5135];
    assign layer4_out[3373] = ~layer3_out[446];
    assign layer4_out[3374] = layer3_out[4388] & layer3_out[4389];
    assign layer4_out[3375] = layer3_out[6278] & ~layer3_out[6279];
    assign layer4_out[3376] = ~(layer3_out[3966] & layer3_out[3967]);
    assign layer4_out[3377] = ~layer3_out[6458];
    assign layer4_out[3378] = ~(layer3_out[1631] | layer3_out[1632]);
    assign layer4_out[3379] = ~layer3_out[2812];
    assign layer4_out[3380] = ~layer3_out[3978];
    assign layer4_out[3381] = ~layer3_out[2273];
    assign layer4_out[3382] = ~layer3_out[263];
    assign layer4_out[3383] = layer3_out[7569];
    assign layer4_out[3384] = ~(layer3_out[2223] & layer3_out[2224]);
    assign layer4_out[3385] = ~layer3_out[6921];
    assign layer4_out[3386] = layer3_out[2737] | layer3_out[2738];
    assign layer4_out[3387] = layer3_out[3383];
    assign layer4_out[3388] = ~layer3_out[1275] | layer3_out[1276];
    assign layer4_out[3389] = layer3_out[7653] & ~layer3_out[7652];
    assign layer4_out[3390] = ~layer3_out[2843] | layer3_out[2842];
    assign layer4_out[3391] = ~layer3_out[3799];
    assign layer4_out[3392] = ~layer3_out[985] | layer3_out[986];
    assign layer4_out[3393] = layer3_out[6821];
    assign layer4_out[3394] = ~layer3_out[7375];
    assign layer4_out[3395] = ~(layer3_out[2503] & layer3_out[2504]);
    assign layer4_out[3396] = ~layer3_out[4678] | layer3_out[4679];
    assign layer4_out[3397] = ~(layer3_out[5433] & layer3_out[5434]);
    assign layer4_out[3398] = layer3_out[2616] & ~layer3_out[2615];
    assign layer4_out[3399] = layer3_out[5579] ^ layer3_out[5580];
    assign layer4_out[3400] = layer3_out[3226] & ~layer3_out[3227];
    assign layer4_out[3401] = ~layer3_out[5057];
    assign layer4_out[3402] = ~layer3_out[5836];
    assign layer4_out[3403] = layer3_out[6951];
    assign layer4_out[3404] = layer3_out[6629] | layer3_out[6630];
    assign layer4_out[3405] = ~layer3_out[4642] | layer3_out[4643];
    assign layer4_out[3406] = ~layer3_out[3528];
    assign layer4_out[3407] = ~layer3_out[1739] | layer3_out[1738];
    assign layer4_out[3408] = ~layer3_out[771] | layer3_out[770];
    assign layer4_out[3409] = layer3_out[4833];
    assign layer4_out[3410] = layer3_out[3605] & ~layer3_out[3606];
    assign layer4_out[3411] = ~(layer3_out[6945] ^ layer3_out[6946]);
    assign layer4_out[3412] = ~(layer3_out[7854] ^ layer3_out[7855]);
    assign layer4_out[3413] = layer3_out[4383] & layer3_out[4384];
    assign layer4_out[3414] = layer3_out[3091] ^ layer3_out[3092];
    assign layer4_out[3415] = ~(layer3_out[6208] ^ layer3_out[6209]);
    assign layer4_out[3416] = ~(layer3_out[4052] ^ layer3_out[4053]);
    assign layer4_out[3417] = layer3_out[479] | layer3_out[480];
    assign layer4_out[3418] = ~layer3_out[4707] | layer3_out[4706];
    assign layer4_out[3419] = layer3_out[3751];
    assign layer4_out[3420] = layer3_out[6772];
    assign layer4_out[3421] = ~(layer3_out[4615] ^ layer3_out[4616]);
    assign layer4_out[3422] = layer3_out[6284] & layer3_out[6285];
    assign layer4_out[3423] = ~layer3_out[4732] | layer3_out[4731];
    assign layer4_out[3424] = ~(layer3_out[457] ^ layer3_out[458]);
    assign layer4_out[3425] = layer3_out[5743];
    assign layer4_out[3426] = layer3_out[5750] ^ layer3_out[5751];
    assign layer4_out[3427] = ~layer3_out[7777];
    assign layer4_out[3428] = ~layer3_out[5061];
    assign layer4_out[3429] = ~(layer3_out[7583] ^ layer3_out[7584]);
    assign layer4_out[3430] = 1'b0;
    assign layer4_out[3431] = layer3_out[5892];
    assign layer4_out[3432] = ~layer3_out[2207];
    assign layer4_out[3433] = layer3_out[6799];
    assign layer4_out[3434] = layer3_out[5449];
    assign layer4_out[3435] = layer3_out[5848] & ~layer3_out[5847];
    assign layer4_out[3436] = ~layer3_out[1147];
    assign layer4_out[3437] = layer3_out[6225] ^ layer3_out[6226];
    assign layer4_out[3438] = ~(layer3_out[429] ^ layer3_out[430]);
    assign layer4_out[3439] = ~(layer3_out[6517] ^ layer3_out[6518]);
    assign layer4_out[3440] = ~(layer3_out[3322] | layer3_out[3323]);
    assign layer4_out[3441] = layer3_out[6258];
    assign layer4_out[3442] = layer3_out[374] & ~layer3_out[375];
    assign layer4_out[3443] = layer3_out[7506] | layer3_out[7507];
    assign layer4_out[3444] = ~(layer3_out[6223] & layer3_out[6224]);
    assign layer4_out[3445] = layer3_out[7246] & ~layer3_out[7245];
    assign layer4_out[3446] = ~layer3_out[3873];
    assign layer4_out[3447] = ~(layer3_out[6194] | layer3_out[6195]);
    assign layer4_out[3448] = ~layer3_out[3196];
    assign layer4_out[3449] = layer3_out[6291];
    assign layer4_out[3450] = layer3_out[820];
    assign layer4_out[3451] = ~layer3_out[4605];
    assign layer4_out[3452] = ~(layer3_out[4892] | layer3_out[4893]);
    assign layer4_out[3453] = layer3_out[950];
    assign layer4_out[3454] = layer3_out[3525];
    assign layer4_out[3455] = layer3_out[3049] & ~layer3_out[3050];
    assign layer4_out[3456] = ~layer3_out[5569] | layer3_out[5568];
    assign layer4_out[3457] = ~(layer3_out[6289] | layer3_out[6290]);
    assign layer4_out[3458] = layer3_out[6286] ^ layer3_out[6287];
    assign layer4_out[3459] = layer3_out[3580];
    assign layer4_out[3460] = ~layer3_out[7389];
    assign layer4_out[3461] = ~layer3_out[186];
    assign layer4_out[3462] = ~layer3_out[6150];
    assign layer4_out[3463] = ~(layer3_out[4601] & layer3_out[4602]);
    assign layer4_out[3464] = layer3_out[1175] & ~layer3_out[1174];
    assign layer4_out[3465] = ~layer3_out[3660];
    assign layer4_out[3466] = ~(layer3_out[5319] | layer3_out[5320]);
    assign layer4_out[3467] = layer3_out[6176];
    assign layer4_out[3468] = layer3_out[2920] ^ layer3_out[2921];
    assign layer4_out[3469] = layer3_out[5518];
    assign layer4_out[3470] = ~layer3_out[6762] | layer3_out[6761];
    assign layer4_out[3471] = layer3_out[5493];
    assign layer4_out[3472] = ~layer3_out[5153];
    assign layer4_out[3473] = ~(layer3_out[21] ^ layer3_out[22]);
    assign layer4_out[3474] = ~layer3_out[4637];
    assign layer4_out[3475] = layer3_out[362] & layer3_out[363];
    assign layer4_out[3476] = ~(layer3_out[7567] ^ layer3_out[7568]);
    assign layer4_out[3477] = ~layer3_out[5138];
    assign layer4_out[3478] = layer3_out[829];
    assign layer4_out[3479] = ~layer3_out[2856] | layer3_out[2857];
    assign layer4_out[3480] = layer3_out[3836];
    assign layer4_out[3481] = layer3_out[685] & ~layer3_out[684];
    assign layer4_out[3482] = ~(layer3_out[2756] | layer3_out[2757]);
    assign layer4_out[3483] = layer3_out[5926];
    assign layer4_out[3484] = layer3_out[3597];
    assign layer4_out[3485] = ~(layer3_out[4058] ^ layer3_out[4059]);
    assign layer4_out[3486] = ~layer3_out[4073] | layer3_out[4072];
    assign layer4_out[3487] = ~(layer3_out[3779] ^ layer3_out[3780]);
    assign layer4_out[3488] = ~layer3_out[7453] | layer3_out[7454];
    assign layer4_out[3489] = layer3_out[7693] ^ layer3_out[7694];
    assign layer4_out[3490] = ~layer3_out[3850] | layer3_out[3851];
    assign layer4_out[3491] = layer3_out[5202] & ~layer3_out[5201];
    assign layer4_out[3492] = layer3_out[1962];
    assign layer4_out[3493] = layer3_out[7950];
    assign layer4_out[3494] = ~layer3_out[7557];
    assign layer4_out[3495] = layer3_out[979];
    assign layer4_out[3496] = ~(layer3_out[3481] ^ layer3_out[3482]);
    assign layer4_out[3497] = layer3_out[4866] & ~layer3_out[4865];
    assign layer4_out[3498] = ~layer3_out[3334];
    assign layer4_out[3499] = ~(layer3_out[5584] ^ layer3_out[5585]);
    assign layer4_out[3500] = layer3_out[5862];
    assign layer4_out[3501] = ~layer3_out[2911];
    assign layer4_out[3502] = layer3_out[652] ^ layer3_out[653];
    assign layer4_out[3503] = ~(layer3_out[7967] ^ layer3_out[7968]);
    assign layer4_out[3504] = layer3_out[1677] & ~layer3_out[1678];
    assign layer4_out[3505] = ~layer3_out[263];
    assign layer4_out[3506] = layer3_out[6909];
    assign layer4_out[3507] = layer3_out[2249];
    assign layer4_out[3508] = ~layer3_out[6377];
    assign layer4_out[3509] = layer3_out[5814];
    assign layer4_out[3510] = layer3_out[3158] & layer3_out[3159];
    assign layer4_out[3511] = ~(layer3_out[280] | layer3_out[281]);
    assign layer4_out[3512] = layer3_out[3838] ^ layer3_out[3839];
    assign layer4_out[3513] = layer3_out[1787] ^ layer3_out[1788];
    assign layer4_out[3514] = layer3_out[940] & ~layer3_out[939];
    assign layer4_out[3515] = ~(layer3_out[4065] ^ layer3_out[4066]);
    assign layer4_out[3516] = ~layer3_out[4935] | layer3_out[4936];
    assign layer4_out[3517] = ~(layer3_out[5842] & layer3_out[5843]);
    assign layer4_out[3518] = ~layer3_out[6232];
    assign layer4_out[3519] = layer3_out[7242] & layer3_out[7243];
    assign layer4_out[3520] = layer3_out[2123];
    assign layer4_out[3521] = ~(layer3_out[2409] & layer3_out[2410]);
    assign layer4_out[3522] = ~layer3_out[314];
    assign layer4_out[3523] = layer3_out[6748] & ~layer3_out[6747];
    assign layer4_out[3524] = ~layer3_out[107];
    assign layer4_out[3525] = layer3_out[2017] & ~layer3_out[2018];
    assign layer4_out[3526] = layer3_out[159];
    assign layer4_out[3527] = ~layer3_out[389];
    assign layer4_out[3528] = layer3_out[7976] ^ layer3_out[7977];
    assign layer4_out[3529] = layer3_out[615] | layer3_out[616];
    assign layer4_out[3530] = ~(layer3_out[4543] & layer3_out[4544]);
    assign layer4_out[3531] = ~(layer3_out[6707] | layer3_out[6708]);
    assign layer4_out[3532] = layer3_out[6606];
    assign layer4_out[3533] = ~layer3_out[586] | layer3_out[585];
    assign layer4_out[3534] = layer3_out[6104];
    assign layer4_out[3535] = layer3_out[1041] & layer3_out[1042];
    assign layer4_out[3536] = layer3_out[2696];
    assign layer4_out[3537] = ~layer3_out[5939];
    assign layer4_out[3538] = layer3_out[5106] ^ layer3_out[5107];
    assign layer4_out[3539] = ~(layer3_out[2104] & layer3_out[2105]);
    assign layer4_out[3540] = ~(layer3_out[3221] & layer3_out[3222]);
    assign layer4_out[3541] = layer3_out[5665] ^ layer3_out[5666];
    assign layer4_out[3542] = layer3_out[6231] & ~layer3_out[6230];
    assign layer4_out[3543] = layer3_out[2403];
    assign layer4_out[3544] = layer3_out[3418];
    assign layer4_out[3545] = ~(layer3_out[7687] | layer3_out[7688]);
    assign layer4_out[3546] = layer3_out[5121] & ~layer3_out[5120];
    assign layer4_out[3547] = ~layer3_out[313];
    assign layer4_out[3548] = layer3_out[271];
    assign layer4_out[3549] = layer3_out[6137];
    assign layer4_out[3550] = layer3_out[6469];
    assign layer4_out[3551] = ~layer3_out[6693];
    assign layer4_out[3552] = 1'b0;
    assign layer4_out[3553] = ~layer3_out[6782];
    assign layer4_out[3554] = ~(layer3_out[1901] & layer3_out[1902]);
    assign layer4_out[3555] = ~layer3_out[4776] | layer3_out[4775];
    assign layer4_out[3556] = ~layer3_out[2832];
    assign layer4_out[3557] = ~layer3_out[131] | layer3_out[130];
    assign layer4_out[3558] = layer3_out[2162] & layer3_out[2163];
    assign layer4_out[3559] = ~(layer3_out[3722] | layer3_out[3723]);
    assign layer4_out[3560] = ~layer3_out[4746];
    assign layer4_out[3561] = ~layer3_out[572] | layer3_out[573];
    assign layer4_out[3562] = layer3_out[2435] & ~layer3_out[2436];
    assign layer4_out[3563] = ~(layer3_out[6712] ^ layer3_out[6713]);
    assign layer4_out[3564] = layer3_out[6263] | layer3_out[6264];
    assign layer4_out[3565] = layer3_out[1864] & ~layer3_out[1865];
    assign layer4_out[3566] = ~(layer3_out[3215] ^ layer3_out[3216]);
    assign layer4_out[3567] = ~layer3_out[6947] | layer3_out[6948];
    assign layer4_out[3568] = layer3_out[6407] | layer3_out[6408];
    assign layer4_out[3569] = ~(layer3_out[3119] | layer3_out[3120]);
    assign layer4_out[3570] = ~(layer3_out[6081] ^ layer3_out[6082]);
    assign layer4_out[3571] = ~layer3_out[5791] | layer3_out[5792];
    assign layer4_out[3572] = layer3_out[3202];
    assign layer4_out[3573] = ~layer3_out[4928];
    assign layer4_out[3574] = layer3_out[253] & ~layer3_out[252];
    assign layer4_out[3575] = ~layer3_out[3337];
    assign layer4_out[3576] = ~layer3_out[5672];
    assign layer4_out[3577] = ~layer3_out[4119];
    assign layer4_out[3578] = ~(layer3_out[7578] ^ layer3_out[7579]);
    assign layer4_out[3579] = ~layer3_out[7543];
    assign layer4_out[3580] = layer3_out[153];
    assign layer4_out[3581] = ~layer3_out[5942];
    assign layer4_out[3582] = ~layer3_out[1512];
    assign layer4_out[3583] = layer3_out[876];
    assign layer4_out[3584] = ~layer3_out[7190];
    assign layer4_out[3585] = ~layer3_out[1340];
    assign layer4_out[3586] = layer3_out[3375];
    assign layer4_out[3587] = layer3_out[7369];
    assign layer4_out[3588] = ~(layer3_out[7213] ^ layer3_out[7214]);
    assign layer4_out[3589] = ~(layer3_out[6620] | layer3_out[6621]);
    assign layer4_out[3590] = layer3_out[5163] & ~layer3_out[5164];
    assign layer4_out[3591] = ~layer3_out[3231];
    assign layer4_out[3592] = layer3_out[1138] | layer3_out[1139];
    assign layer4_out[3593] = layer3_out[1359];
    assign layer4_out[3594] = ~(layer3_out[6316] & layer3_out[6317]);
    assign layer4_out[3595] = ~layer3_out[1648];
    assign layer4_out[3596] = layer3_out[3315] ^ layer3_out[3316];
    assign layer4_out[3597] = ~(layer3_out[265] | layer3_out[266]);
    assign layer4_out[3598] = layer3_out[7624] & ~layer3_out[7623];
    assign layer4_out[3599] = layer3_out[3726] & layer3_out[3727];
    assign layer4_out[3600] = layer3_out[5038] & ~layer3_out[5037];
    assign layer4_out[3601] = layer3_out[509];
    assign layer4_out[3602] = ~layer3_out[4547];
    assign layer4_out[3603] = layer3_out[14] & ~layer3_out[13];
    assign layer4_out[3604] = ~(layer3_out[1024] & layer3_out[1025]);
    assign layer4_out[3605] = layer3_out[4001];
    assign layer4_out[3606] = ~layer3_out[7294] | layer3_out[7295];
    assign layer4_out[3607] = layer3_out[3581] | layer3_out[3582];
    assign layer4_out[3608] = layer3_out[7800];
    assign layer4_out[3609] = layer3_out[5825];
    assign layer4_out[3610] = ~layer3_out[5259];
    assign layer4_out[3611] = layer3_out[5207];
    assign layer4_out[3612] = layer3_out[844] & ~layer3_out[843];
    assign layer4_out[3613] = layer3_out[4146] & layer3_out[4147];
    assign layer4_out[3614] = 1'b1;
    assign layer4_out[3615] = ~(layer3_out[3148] ^ layer3_out[3149]);
    assign layer4_out[3616] = ~layer3_out[5892];
    assign layer4_out[3617] = layer3_out[5729];
    assign layer4_out[3618] = layer3_out[6331];
    assign layer4_out[3619] = layer3_out[5040];
    assign layer4_out[3620] = ~layer3_out[4046] | layer3_out[4047];
    assign layer4_out[3621] = layer3_out[291] ^ layer3_out[292];
    assign layer4_out[3622] = layer3_out[5397] ^ layer3_out[5398];
    assign layer4_out[3623] = ~layer3_out[1986] | layer3_out[1985];
    assign layer4_out[3624] = layer3_out[4313];
    assign layer4_out[3625] = ~layer3_out[3718] | layer3_out[3717];
    assign layer4_out[3626] = ~layer3_out[4960] | layer3_out[4959];
    assign layer4_out[3627] = ~layer3_out[3468];
    assign layer4_out[3628] = layer3_out[7647];
    assign layer4_out[3629] = layer3_out[1691] & ~layer3_out[1690];
    assign layer4_out[3630] = ~layer3_out[7227];
    assign layer4_out[3631] = ~(layer3_out[1228] | layer3_out[1229]);
    assign layer4_out[3632] = layer3_out[2417];
    assign layer4_out[3633] = ~layer3_out[4266] | layer3_out[4267];
    assign layer4_out[3634] = ~layer3_out[1675];
    assign layer4_out[3635] = layer3_out[562];
    assign layer4_out[3636] = ~(layer3_out[7844] & layer3_out[7845]);
    assign layer4_out[3637] = ~layer3_out[7309];
    assign layer4_out[3638] = layer3_out[1967];
    assign layer4_out[3639] = layer3_out[5424] ^ layer3_out[5425];
    assign layer4_out[3640] = layer3_out[4833];
    assign layer4_out[3641] = layer3_out[4817];
    assign layer4_out[3642] = layer3_out[395] & layer3_out[396];
    assign layer4_out[3643] = ~layer3_out[4483] | layer3_out[4482];
    assign layer4_out[3644] = layer3_out[7766] ^ layer3_out[7767];
    assign layer4_out[3645] = ~(layer3_out[5131] | layer3_out[5132]);
    assign layer4_out[3646] = layer3_out[5422] & layer3_out[5423];
    assign layer4_out[3647] = layer3_out[190] & layer3_out[191];
    assign layer4_out[3648] = layer3_out[3833];
    assign layer4_out[3649] = ~(layer3_out[4924] & layer3_out[4925]);
    assign layer4_out[3650] = ~layer3_out[2349];
    assign layer4_out[3651] = ~layer3_out[524];
    assign layer4_out[3652] = ~layer3_out[4799];
    assign layer4_out[3653] = ~layer3_out[1796] | layer3_out[1797];
    assign layer4_out[3654] = ~(layer3_out[2094] | layer3_out[2095]);
    assign layer4_out[3655] = layer3_out[3109];
    assign layer4_out[3656] = layer3_out[678];
    assign layer4_out[3657] = ~layer3_out[1055];
    assign layer4_out[3658] = ~layer3_out[3044];
    assign layer4_out[3659] = ~(layer3_out[7356] | layer3_out[7357]);
    assign layer4_out[3660] = ~(layer3_out[1707] | layer3_out[1708]);
    assign layer4_out[3661] = layer3_out[7953] ^ layer3_out[7954];
    assign layer4_out[3662] = layer3_out[1254] ^ layer3_out[1255];
    assign layer4_out[3663] = layer3_out[7322] ^ layer3_out[7323];
    assign layer4_out[3664] = ~(layer3_out[5897] ^ layer3_out[5898]);
    assign layer4_out[3665] = ~layer3_out[6893];
    assign layer4_out[3666] = layer3_out[6496];
    assign layer4_out[3667] = layer3_out[5724] ^ layer3_out[5725];
    assign layer4_out[3668] = ~(layer3_out[6308] & layer3_out[6309]);
    assign layer4_out[3669] = ~(layer3_out[4043] ^ layer3_out[4044]);
    assign layer4_out[3670] = layer3_out[2081] & layer3_out[2082];
    assign layer4_out[3671] = layer3_out[3141];
    assign layer4_out[3672] = layer3_out[2757] & ~layer3_out[2758];
    assign layer4_out[3673] = layer3_out[4712] & layer3_out[4713];
    assign layer4_out[3674] = ~layer3_out[1923];
    assign layer4_out[3675] = ~(layer3_out[2032] | layer3_out[2033]);
    assign layer4_out[3676] = ~layer3_out[4283];
    assign layer4_out[3677] = layer3_out[5438] & ~layer3_out[5437];
    assign layer4_out[3678] = ~(layer3_out[2992] & layer3_out[2993]);
    assign layer4_out[3679] = 1'b1;
    assign layer4_out[3680] = ~layer3_out[3082] | layer3_out[3081];
    assign layer4_out[3681] = layer3_out[7975];
    assign layer4_out[3682] = ~(layer3_out[1608] & layer3_out[1609]);
    assign layer4_out[3683] = layer3_out[385] ^ layer3_out[386];
    assign layer4_out[3684] = layer3_out[4871];
    assign layer4_out[3685] = layer3_out[74] | layer3_out[75];
    assign layer4_out[3686] = ~layer3_out[5532];
    assign layer4_out[3687] = ~layer3_out[3358] | layer3_out[3359];
    assign layer4_out[3688] = ~(layer3_out[4884] ^ layer3_out[4885]);
    assign layer4_out[3689] = layer3_out[4401];
    assign layer4_out[3690] = layer3_out[1777];
    assign layer4_out[3691] = layer3_out[2399];
    assign layer4_out[3692] = ~layer3_out[620] | layer3_out[619];
    assign layer4_out[3693] = layer3_out[2795] & ~layer3_out[2794];
    assign layer4_out[3694] = ~(layer3_out[2563] ^ layer3_out[2564]);
    assign layer4_out[3695] = layer3_out[3318] & ~layer3_out[3317];
    assign layer4_out[3696] = layer3_out[863];
    assign layer4_out[3697] = layer3_out[3306] ^ layer3_out[3307];
    assign layer4_out[3698] = ~layer3_out[6570];
    assign layer4_out[3699] = ~layer3_out[1890] | layer3_out[1891];
    assign layer4_out[3700] = layer3_out[6695] ^ layer3_out[6696];
    assign layer4_out[3701] = layer3_out[2509];
    assign layer4_out[3702] = ~layer3_out[3787];
    assign layer4_out[3703] = ~(layer3_out[6849] | layer3_out[6850]);
    assign layer4_out[3704] = ~layer3_out[6038];
    assign layer4_out[3705] = layer3_out[5648];
    assign layer4_out[3706] = layer3_out[3585];
    assign layer4_out[3707] = ~layer3_out[406];
    assign layer4_out[3708] = ~layer3_out[4707];
    assign layer4_out[3709] = ~layer3_out[7420];
    assign layer4_out[3710] = ~(layer3_out[5390] ^ layer3_out[5391]);
    assign layer4_out[3711] = ~(layer3_out[2087] ^ layer3_out[2088]);
    assign layer4_out[3712] = ~layer3_out[1688];
    assign layer4_out[3713] = ~layer3_out[7468];
    assign layer4_out[3714] = ~layer3_out[7886];
    assign layer4_out[3715] = layer3_out[217] | layer3_out[218];
    assign layer4_out[3716] = ~layer3_out[6791];
    assign layer4_out[3717] = layer3_out[5653] ^ layer3_out[5654];
    assign layer4_out[3718] = layer3_out[7222];
    assign layer4_out[3719] = layer3_out[1582] & layer3_out[1583];
    assign layer4_out[3720] = layer3_out[1881] & layer3_out[1882];
    assign layer4_out[3721] = ~layer3_out[6072] | layer3_out[6071];
    assign layer4_out[3722] = layer3_out[7175];
    assign layer4_out[3723] = ~layer3_out[5247];
    assign layer4_out[3724] = layer3_out[7622] | layer3_out[7623];
    assign layer4_out[3725] = layer3_out[4912];
    assign layer4_out[3726] = layer3_out[3607];
    assign layer4_out[3727] = layer3_out[4591];
    assign layer4_out[3728] = ~layer3_out[3693];
    assign layer4_out[3729] = layer3_out[4576] & ~layer3_out[4575];
    assign layer4_out[3730] = layer3_out[7713];
    assign layer4_out[3731] = layer3_out[5714] | layer3_out[5715];
    assign layer4_out[3732] = ~(layer3_out[5894] | layer3_out[5895]);
    assign layer4_out[3733] = ~(layer3_out[2577] ^ layer3_out[2578]);
    assign layer4_out[3734] = layer3_out[3829] & layer3_out[3830];
    assign layer4_out[3735] = layer3_out[7671] | layer3_out[7672];
    assign layer4_out[3736] = ~(layer3_out[4097] ^ layer3_out[4098]);
    assign layer4_out[3737] = layer3_out[5301] & layer3_out[5302];
    assign layer4_out[3738] = 1'b1;
    assign layer4_out[3739] = layer3_out[983] | layer3_out[984];
    assign layer4_out[3740] = layer3_out[5148] | layer3_out[5149];
    assign layer4_out[3741] = layer3_out[6569];
    assign layer4_out[3742] = layer3_out[129];
    assign layer4_out[3743] = ~layer3_out[1601];
    assign layer4_out[3744] = layer3_out[5738] & ~layer3_out[5739];
    assign layer4_out[3745] = layer3_out[6805] ^ layer3_out[6806];
    assign layer4_out[3746] = layer3_out[4613] ^ layer3_out[4614];
    assign layer4_out[3747] = layer3_out[7769] | layer3_out[7770];
    assign layer4_out[3748] = layer3_out[6227] ^ layer3_out[6228];
    assign layer4_out[3749] = ~(layer3_out[6513] & layer3_out[6514]);
    assign layer4_out[3750] = ~layer3_out[7617] | layer3_out[7616];
    assign layer4_out[3751] = ~layer3_out[1197] | layer3_out[1198];
    assign layer4_out[3752] = layer3_out[3128] ^ layer3_out[3129];
    assign layer4_out[3753] = ~layer3_out[4440];
    assign layer4_out[3754] = ~(layer3_out[7413] ^ layer3_out[7414]);
    assign layer4_out[3755] = layer3_out[3853];
    assign layer4_out[3756] = layer3_out[6803];
    assign layer4_out[3757] = layer3_out[5020];
    assign layer4_out[3758] = ~layer3_out[3229];
    assign layer4_out[3759] = layer3_out[7105] & ~layer3_out[7104];
    assign layer4_out[3760] = ~(layer3_out[4022] ^ layer3_out[4023]);
    assign layer4_out[3761] = layer3_out[4268];
    assign layer4_out[3762] = ~layer3_out[6706] | layer3_out[6707];
    assign layer4_out[3763] = layer3_out[2396] & ~layer3_out[2395];
    assign layer4_out[3764] = layer3_out[4568];
    assign layer4_out[3765] = layer3_out[2307] ^ layer3_out[2308];
    assign layer4_out[3766] = ~layer3_out[3525];
    assign layer4_out[3767] = ~layer3_out[7704] | layer3_out[7705];
    assign layer4_out[3768] = layer3_out[756] ^ layer3_out[757];
    assign layer4_out[3769] = ~layer3_out[544];
    assign layer4_out[3770] = ~layer3_out[3087];
    assign layer4_out[3771] = layer3_out[4131];
    assign layer4_out[3772] = layer3_out[6102] | layer3_out[6103];
    assign layer4_out[3773] = ~layer3_out[2124];
    assign layer4_out[3774] = layer3_out[1798];
    assign layer4_out[3775] = layer3_out[3926];
    assign layer4_out[3776] = ~layer3_out[1940];
    assign layer4_out[3777] = layer3_out[4316];
    assign layer4_out[3778] = ~layer3_out[7116];
    assign layer4_out[3779] = layer3_out[6222] & ~layer3_out[6223];
    assign layer4_out[3780] = ~layer3_out[4435] | layer3_out[4434];
    assign layer4_out[3781] = layer3_out[5154] & ~layer3_out[5155];
    assign layer4_out[3782] = ~layer3_out[2778] | layer3_out[2779];
    assign layer4_out[3783] = ~(layer3_out[7313] ^ layer3_out[7314]);
    assign layer4_out[3784] = layer3_out[6747] & ~layer3_out[6746];
    assign layer4_out[3785] = ~layer3_out[6659];
    assign layer4_out[3786] = layer3_out[6218] ^ layer3_out[6219];
    assign layer4_out[3787] = layer3_out[6661] & layer3_out[6662];
    assign layer4_out[3788] = ~layer3_out[7802];
    assign layer4_out[3789] = layer3_out[15] ^ layer3_out[16];
    assign layer4_out[3790] = ~(layer3_out[2691] | layer3_out[2692]);
    assign layer4_out[3791] = layer3_out[443] ^ layer3_out[444];
    assign layer4_out[3792] = layer3_out[3118] & ~layer3_out[3117];
    assign layer4_out[3793] = layer3_out[95] ^ layer3_out[96];
    assign layer4_out[3794] = ~(layer3_out[5243] & layer3_out[5244]);
    assign layer4_out[3795] = layer3_out[7254];
    assign layer4_out[3796] = layer3_out[707] & ~layer3_out[708];
    assign layer4_out[3797] = ~layer3_out[1928];
    assign layer4_out[3798] = layer3_out[6409] & layer3_out[6410];
    assign layer4_out[3799] = layer3_out[6460];
    assign layer4_out[3800] = layer3_out[277] ^ layer3_out[278];
    assign layer4_out[3801] = ~layer3_out[5232];
    assign layer4_out[3802] = ~layer3_out[5188];
    assign layer4_out[3803] = layer3_out[1885] & ~layer3_out[1886];
    assign layer4_out[3804] = ~(layer3_out[5116] | layer3_out[5117]);
    assign layer4_out[3805] = layer3_out[1635] ^ layer3_out[1636];
    assign layer4_out[3806] = ~layer3_out[3256];
    assign layer4_out[3807] = layer3_out[4054];
    assign layer4_out[3808] = layer3_out[1445] & layer3_out[1446];
    assign layer4_out[3809] = ~layer3_out[1402];
    assign layer4_out[3810] = ~(layer3_out[1657] & layer3_out[1658]);
    assign layer4_out[3811] = ~layer3_out[2533] | layer3_out[2532];
    assign layer4_out[3812] = ~(layer3_out[407] & layer3_out[408]);
    assign layer4_out[3813] = layer3_out[5437];
    assign layer4_out[3814] = ~(layer3_out[2086] ^ layer3_out[2087]);
    assign layer4_out[3815] = ~(layer3_out[508] ^ layer3_out[509]);
    assign layer4_out[3816] = layer3_out[2461] & ~layer3_out[2462];
    assign layer4_out[3817] = ~layer3_out[5349] | layer3_out[5350];
    assign layer4_out[3818] = layer3_out[6783];
    assign layer4_out[3819] = ~layer3_out[226];
    assign layer4_out[3820] = ~layer3_out[5025];
    assign layer4_out[3821] = layer3_out[6420] | layer3_out[6421];
    assign layer4_out[3822] = layer3_out[5090] & ~layer3_out[5091];
    assign layer4_out[3823] = ~layer3_out[1226];
    assign layer4_out[3824] = ~layer3_out[6947];
    assign layer4_out[3825] = ~(layer3_out[4565] ^ layer3_out[4566]);
    assign layer4_out[3826] = layer3_out[1766];
    assign layer4_out[3827] = ~layer3_out[6176];
    assign layer4_out[3828] = ~(layer3_out[1897] | layer3_out[1898]);
    assign layer4_out[3829] = ~(layer3_out[2200] ^ layer3_out[2201]);
    assign layer4_out[3830] = ~(layer3_out[235] ^ layer3_out[236]);
    assign layer4_out[3831] = layer3_out[1097] & ~layer3_out[1096];
    assign layer4_out[3832] = ~layer3_out[5069] | layer3_out[5070];
    assign layer4_out[3833] = ~layer3_out[6129];
    assign layer4_out[3834] = ~layer3_out[1578];
    assign layer4_out[3835] = layer3_out[7385] & ~layer3_out[7386];
    assign layer4_out[3836] = ~(layer3_out[6115] ^ layer3_out[6116]);
    assign layer4_out[3837] = ~layer3_out[4203] | layer3_out[4204];
    assign layer4_out[3838] = layer3_out[4029];
    assign layer4_out[3839] = layer3_out[807] & ~layer3_out[806];
    assign layer4_out[3840] = layer3_out[5179] | layer3_out[5180];
    assign layer4_out[3841] = ~(layer3_out[3919] ^ layer3_out[3920]);
    assign layer4_out[3842] = ~layer3_out[2866];
    assign layer4_out[3843] = ~layer3_out[4388];
    assign layer4_out[3844] = layer3_out[5911] | layer3_out[5912];
    assign layer4_out[3845] = layer3_out[4813];
    assign layer4_out[3846] = layer3_out[2501];
    assign layer4_out[3847] = ~(layer3_out[7454] ^ layer3_out[7455]);
    assign layer4_out[3848] = ~(layer3_out[1387] & layer3_out[1388]);
    assign layer4_out[3849] = ~layer3_out[5525] | layer3_out[5526];
    assign layer4_out[3850] = ~layer3_out[2499];
    assign layer4_out[3851] = ~layer3_out[4730];
    assign layer4_out[3852] = ~layer3_out[5718];
    assign layer4_out[3853] = ~(layer3_out[4339] ^ layer3_out[4340]);
    assign layer4_out[3854] = ~(layer3_out[2939] & layer3_out[2940]);
    assign layer4_out[3855] = layer3_out[921] & ~layer3_out[922];
    assign layer4_out[3856] = ~layer3_out[6924] | layer3_out[6925];
    assign layer4_out[3857] = ~(layer3_out[4913] & layer3_out[4914]);
    assign layer4_out[3858] = ~(layer3_out[3716] | layer3_out[3717]);
    assign layer4_out[3859] = ~layer3_out[7910];
    assign layer4_out[3860] = ~(layer3_out[4267] ^ layer3_out[4268]);
    assign layer4_out[3861] = ~layer3_out[3864];
    assign layer4_out[3862] = ~(layer3_out[7878] ^ layer3_out[7879]);
    assign layer4_out[3863] = ~(layer3_out[4815] ^ layer3_out[4816]);
    assign layer4_out[3864] = layer3_out[7832] & ~layer3_out[7833];
    assign layer4_out[3865] = layer3_out[2010];
    assign layer4_out[3866] = layer3_out[5932];
    assign layer4_out[3867] = ~(layer3_out[5940] | layer3_out[5941]);
    assign layer4_out[3868] = layer3_out[1336] | layer3_out[1337];
    assign layer4_out[3869] = layer3_out[5721] & ~layer3_out[5722];
    assign layer4_out[3870] = ~layer3_out[6124];
    assign layer4_out[3871] = layer3_out[4803];
    assign layer4_out[3872] = layer3_out[1325];
    assign layer4_out[3873] = layer3_out[7591] & ~layer3_out[7590];
    assign layer4_out[3874] = layer3_out[6364];
    assign layer4_out[3875] = layer3_out[418];
    assign layer4_out[3876] = layer3_out[7945] ^ layer3_out[7946];
    assign layer4_out[3877] = ~layer3_out[411];
    assign layer4_out[3878] = ~layer3_out[6171];
    assign layer4_out[3879] = layer3_out[168] & ~layer3_out[169];
    assign layer4_out[3880] = ~layer3_out[796] | layer3_out[795];
    assign layer4_out[3881] = ~layer3_out[5129];
    assign layer4_out[3882] = ~(layer3_out[6576] ^ layer3_out[6577]);
    assign layer4_out[3883] = ~(layer3_out[2108] & layer3_out[2109]);
    assign layer4_out[3884] = layer3_out[2524];
    assign layer4_out[3885] = ~layer3_out[2212] | layer3_out[2211];
    assign layer4_out[3886] = layer3_out[5874];
    assign layer4_out[3887] = ~layer3_out[7054];
    assign layer4_out[3888] = layer3_out[1877] & ~layer3_out[1878];
    assign layer4_out[3889] = layer3_out[2720];
    assign layer4_out[3890] = ~layer3_out[549] | layer3_out[548];
    assign layer4_out[3891] = ~(layer3_out[2938] | layer3_out[2939]);
    assign layer4_out[3892] = ~(layer3_out[1561] | layer3_out[1562]);
    assign layer4_out[3893] = layer3_out[6870] | layer3_out[6871];
    assign layer4_out[3894] = ~(layer3_out[2454] ^ layer3_out[2455]);
    assign layer4_out[3895] = ~layer3_out[342];
    assign layer4_out[3896] = layer3_out[7376];
    assign layer4_out[3897] = ~layer3_out[7086];
    assign layer4_out[3898] = layer3_out[285] ^ layer3_out[286];
    assign layer4_out[3899] = layer3_out[847] & ~layer3_out[848];
    assign layer4_out[3900] = layer3_out[2572];
    assign layer4_out[3901] = layer3_out[5018] | layer3_out[5019];
    assign layer4_out[3902] = ~layer3_out[4903] | layer3_out[4902];
    assign layer4_out[3903] = layer3_out[7259] ^ layer3_out[7260];
    assign layer4_out[3904] = layer3_out[1991] | layer3_out[1992];
    assign layer4_out[3905] = layer3_out[6581];
    assign layer4_out[3906] = layer3_out[455] & layer3_out[456];
    assign layer4_out[3907] = layer3_out[1941];
    assign layer4_out[3908] = ~(layer3_out[4537] & layer3_out[4538]);
    assign layer4_out[3909] = ~layer3_out[2641];
    assign layer4_out[3910] = ~layer3_out[298];
    assign layer4_out[3911] = layer3_out[2004];
    assign layer4_out[3912] = layer3_out[63];
    assign layer4_out[3913] = ~layer3_out[1185];
    assign layer4_out[3914] = layer3_out[7872] | layer3_out[7873];
    assign layer4_out[3915] = ~layer3_out[3912];
    assign layer4_out[3916] = ~layer3_out[3344];
    assign layer4_out[3917] = ~layer3_out[4095];
    assign layer4_out[3918] = layer3_out[6942] & ~layer3_out[6941];
    assign layer4_out[3919] = layer3_out[7493] ^ layer3_out[7494];
    assign layer4_out[3920] = layer3_out[4720] ^ layer3_out[4721];
    assign layer4_out[3921] = ~(layer3_out[1309] ^ layer3_out[1310]);
    assign layer4_out[3922] = layer3_out[563];
    assign layer4_out[3923] = ~layer3_out[2056];
    assign layer4_out[3924] = ~layer3_out[7573];
    assign layer4_out[3925] = ~layer3_out[6553];
    assign layer4_out[3926] = ~layer3_out[3085];
    assign layer4_out[3927] = layer3_out[6348];
    assign layer4_out[3928] = layer3_out[6273];
    assign layer4_out[3929] = ~(layer3_out[2447] & layer3_out[2448]);
    assign layer4_out[3930] = ~layer3_out[7640] | layer3_out[7641];
    assign layer4_out[3931] = layer3_out[6887] & ~layer3_out[6888];
    assign layer4_out[3932] = ~layer3_out[7895];
    assign layer4_out[3933] = ~(layer3_out[3303] ^ layer3_out[3304]);
    assign layer4_out[3934] = layer3_out[3396] & layer3_out[3397];
    assign layer4_out[3935] = ~layer3_out[1692];
    assign layer4_out[3936] = ~(layer3_out[4281] & layer3_out[4282]);
    assign layer4_out[3937] = ~layer3_out[186] | layer3_out[187];
    assign layer4_out[3938] = layer3_out[3859] & ~layer3_out[3860];
    assign layer4_out[3939] = layer3_out[6700];
    assign layer4_out[3940] = ~layer3_out[7040] | layer3_out[7041];
    assign layer4_out[3941] = ~layer3_out[6652];
    assign layer4_out[3942] = ~(layer3_out[6555] ^ layer3_out[6556]);
    assign layer4_out[3943] = layer3_out[4092];
    assign layer4_out[3944] = ~layer3_out[2541];
    assign layer4_out[3945] = ~layer3_out[4634] | layer3_out[4635];
    assign layer4_out[3946] = layer3_out[1808] ^ layer3_out[1809];
    assign layer4_out[3947] = ~layer3_out[6440];
    assign layer4_out[3948] = ~(layer3_out[1113] & layer3_out[1114]);
    assign layer4_out[3949] = ~(layer3_out[4373] ^ layer3_out[4374]);
    assign layer4_out[3950] = layer3_out[7968] ^ layer3_out[7969];
    assign layer4_out[3951] = ~(layer3_out[3795] ^ layer3_out[3796]);
    assign layer4_out[3952] = ~(layer3_out[3072] & layer3_out[3073]);
    assign layer4_out[3953] = ~(layer3_out[2598] & layer3_out[2599]);
    assign layer4_out[3954] = ~layer3_out[7502];
    assign layer4_out[3955] = layer3_out[5799];
    assign layer4_out[3956] = ~layer3_out[2553];
    assign layer4_out[3957] = ~layer3_out[1970];
    assign layer4_out[3958] = layer3_out[869];
    assign layer4_out[3959] = layer3_out[3079];
    assign layer4_out[3960] = ~layer3_out[2597];
    assign layer4_out[3961] = layer3_out[3187];
    assign layer4_out[3962] = layer3_out[1101];
    assign layer4_out[3963] = ~layer3_out[2335];
    assign layer4_out[3964] = layer3_out[167] & ~layer3_out[166];
    assign layer4_out[3965] = ~(layer3_out[1688] | layer3_out[1689]);
    assign layer4_out[3966] = layer3_out[1711];
    assign layer4_out[3967] = layer3_out[4100] & ~layer3_out[4101];
    assign layer4_out[3968] = layer3_out[7510] ^ layer3_out[7511];
    assign layer4_out[3969] = layer3_out[3950] & layer3_out[3951];
    assign layer4_out[3970] = ~layer3_out[3049] | layer3_out[3048];
    assign layer4_out[3971] = ~(layer3_out[1396] | layer3_out[1397]);
    assign layer4_out[3972] = ~(layer3_out[3694] | layer3_out[3695]);
    assign layer4_out[3973] = layer3_out[5962] & ~layer3_out[5961];
    assign layer4_out[3974] = layer3_out[1504];
    assign layer4_out[3975] = layer3_out[7327] ^ layer3_out[7328];
    assign layer4_out[3976] = ~layer3_out[4607];
    assign layer4_out[3977] = layer3_out[4257];
    assign layer4_out[3978] = layer3_out[3667];
    assign layer4_out[3979] = ~layer3_out[5197] | layer3_out[5198];
    assign layer4_out[3980] = layer3_out[4068];
    assign layer4_out[3981] = layer3_out[2248];
    assign layer4_out[3982] = layer3_out[2743] & ~layer3_out[2744];
    assign layer4_out[3983] = ~layer3_out[4884];
    assign layer4_out[3984] = ~(layer3_out[2137] | layer3_out[2138]);
    assign layer4_out[3985] = ~(layer3_out[4808] | layer3_out[4809]);
    assign layer4_out[3986] = ~layer3_out[220] | layer3_out[219];
    assign layer4_out[3987] = layer3_out[7589] & ~layer3_out[7590];
    assign layer4_out[3988] = ~layer3_out[2880];
    assign layer4_out[3989] = ~layer3_out[206];
    assign layer4_out[3990] = ~layer3_out[5699];
    assign layer4_out[3991] = layer3_out[1081];
    assign layer4_out[3992] = layer3_out[4484];
    assign layer4_out[3993] = ~layer3_out[5884] | layer3_out[5883];
    assign layer4_out[3994] = ~(layer3_out[4172] & layer3_out[4173]);
    assign layer4_out[3995] = ~(layer3_out[6732] & layer3_out[6733]);
    assign layer4_out[3996] = ~layer3_out[6596];
    assign layer4_out[3997] = layer3_out[2884] | layer3_out[2885];
    assign layer4_out[3998] = layer3_out[4229];
    assign layer4_out[3999] = ~layer3_out[5804];
    assign layer4_out[4000] = ~(layer3_out[7051] ^ layer3_out[7052]);
    assign layer4_out[4001] = ~layer3_out[613] | layer3_out[614];
    assign layer4_out[4002] = layer3_out[3423] ^ layer3_out[3424];
    assign layer4_out[4003] = ~(layer3_out[1537] ^ layer3_out[1538]);
    assign layer4_out[4004] = layer3_out[1268] ^ layer3_out[1269];
    assign layer4_out[4005] = ~layer3_out[2899];
    assign layer4_out[4006] = ~layer3_out[5849];
    assign layer4_out[4007] = ~layer3_out[5002];
    assign layer4_out[4008] = ~layer3_out[1232] | layer3_out[1233];
    assign layer4_out[4009] = layer3_out[7639];
    assign layer4_out[4010] = ~(layer3_out[2948] ^ layer3_out[2949]);
    assign layer4_out[4011] = layer3_out[6060] | layer3_out[6061];
    assign layer4_out[4012] = layer3_out[5509];
    assign layer4_out[4013] = layer3_out[230];
    assign layer4_out[4014] = ~layer3_out[6933];
    assign layer4_out[4015] = ~layer3_out[5937];
    assign layer4_out[4016] = ~layer3_out[5860];
    assign layer4_out[4017] = ~layer3_out[6270] | layer3_out[6269];
    assign layer4_out[4018] = layer3_out[1928] | layer3_out[1929];
    assign layer4_out[4019] = ~layer3_out[7630];
    assign layer4_out[4020] = layer3_out[7446] ^ layer3_out[7447];
    assign layer4_out[4021] = ~layer3_out[5710];
    assign layer4_out[4022] = ~layer3_out[5362];
    assign layer4_out[4023] = ~(layer3_out[4138] ^ layer3_out[4139]);
    assign layer4_out[4024] = ~layer3_out[5372] | layer3_out[5371];
    assign layer4_out[4025] = layer3_out[5321] ^ layer3_out[5322];
    assign layer4_out[4026] = layer3_out[638];
    assign layer4_out[4027] = layer3_out[706];
    assign layer4_out[4028] = ~layer3_out[2035];
    assign layer4_out[4029] = layer3_out[793] & layer3_out[794];
    assign layer4_out[4030] = ~layer3_out[6801] | layer3_out[6802];
    assign layer4_out[4031] = ~(layer3_out[3488] & layer3_out[3489]);
    assign layer4_out[4032] = layer3_out[3647] & layer3_out[3648];
    assign layer4_out[4033] = ~layer3_out[1157] | layer3_out[1158];
    assign layer4_out[4034] = ~(layer3_out[2225] & layer3_out[2226]);
    assign layer4_out[4035] = ~layer3_out[6461] | layer3_out[6462];
    assign layer4_out[4036] = layer3_out[6592];
    assign layer4_out[4037] = ~(layer3_out[4351] ^ layer3_out[4352]);
    assign layer4_out[4038] = layer3_out[530] & ~layer3_out[529];
    assign layer4_out[4039] = layer3_out[907];
    assign layer4_out[4040] = layer3_out[324] ^ layer3_out[325];
    assign layer4_out[4041] = layer3_out[5741];
    assign layer4_out[4042] = ~layer3_out[3078] | layer3_out[3077];
    assign layer4_out[4043] = ~(layer3_out[2453] ^ layer3_out[2454]);
    assign layer4_out[4044] = layer3_out[3073] ^ layer3_out[3074];
    assign layer4_out[4045] = ~(layer3_out[7521] & layer3_out[7522]);
    assign layer4_out[4046] = layer3_out[1268] & ~layer3_out[1267];
    assign layer4_out[4047] = ~(layer3_out[2199] ^ layer3_out[2200]);
    assign layer4_out[4048] = ~layer3_out[7664];
    assign layer4_out[4049] = layer3_out[5773] | layer3_out[5774];
    assign layer4_out[4050] = ~layer3_out[2487] | layer3_out[2488];
    assign layer4_out[4051] = ~(layer3_out[4135] ^ layer3_out[4136]);
    assign layer4_out[4052] = ~layer3_out[7829];
    assign layer4_out[4053] = ~(layer3_out[2165] ^ layer3_out[2166]);
    assign layer4_out[4054] = ~layer3_out[3317] | layer3_out[3316];
    assign layer4_out[4055] = layer3_out[6267] | layer3_out[6268];
    assign layer4_out[4056] = layer3_out[2255];
    assign layer4_out[4057] = ~layer3_out[1025] | layer3_out[1026];
    assign layer4_out[4058] = layer3_out[6825] ^ layer3_out[6826];
    assign layer4_out[4059] = layer3_out[4166];
    assign layer4_out[4060] = layer3_out[3667] | layer3_out[3668];
    assign layer4_out[4061] = layer3_out[1165];
    assign layer4_out[4062] = ~(layer3_out[5812] & layer3_out[5813]);
    assign layer4_out[4063] = ~layer3_out[2143];
    assign layer4_out[4064] = layer3_out[3436];
    assign layer4_out[4065] = 1'b0;
    assign layer4_out[4066] = layer3_out[845] & layer3_out[846];
    assign layer4_out[4067] = ~(layer3_out[1845] | layer3_out[1846]);
    assign layer4_out[4068] = ~(layer3_out[4908] & layer3_out[4909]);
    assign layer4_out[4069] = ~layer3_out[6676];
    assign layer4_out[4070] = layer3_out[1291] ^ layer3_out[1292];
    assign layer4_out[4071] = ~(layer3_out[7227] & layer3_out[7228]);
    assign layer4_out[4072] = ~layer3_out[6390];
    assign layer4_out[4073] = layer3_out[3041];
    assign layer4_out[4074] = ~layer3_out[3900];
    assign layer4_out[4075] = layer3_out[3143];
    assign layer4_out[4076] = ~layer3_out[5675];
    assign layer4_out[4077] = ~(layer3_out[3633] & layer3_out[3634]);
    assign layer4_out[4078] = ~(layer3_out[2944] ^ layer3_out[2945]);
    assign layer4_out[4079] = ~layer3_out[2790];
    assign layer4_out[4080] = layer3_out[7867] & ~layer3_out[7868];
    assign layer4_out[4081] = layer3_out[5991] ^ layer3_out[5992];
    assign layer4_out[4082] = layer3_out[3522] & ~layer3_out[3521];
    assign layer4_out[4083] = layer3_out[4227];
    assign layer4_out[4084] = 1'b1;
    assign layer4_out[4085] = layer3_out[1033] & ~layer3_out[1032];
    assign layer4_out[4086] = ~layer3_out[4879];
    assign layer4_out[4087] = layer3_out[461];
    assign layer4_out[4088] = ~layer3_out[7035];
    assign layer4_out[4089] = layer3_out[5730];
    assign layer4_out[4090] = ~layer3_out[4917];
    assign layer4_out[4091] = layer3_out[527] & ~layer3_out[526];
    assign layer4_out[4092] = layer3_out[2469] & ~layer3_out[2470];
    assign layer4_out[4093] = layer3_out[1227] | layer3_out[1228];
    assign layer4_out[4094] = layer3_out[1933];
    assign layer4_out[4095] = layer3_out[5368] & layer3_out[5369];
    assign layer4_out[4096] = ~layer3_out[4906];
    assign layer4_out[4097] = layer3_out[5756] & layer3_out[5757];
    assign layer4_out[4098] = layer3_out[2657];
    assign layer4_out[4099] = layer3_out[1085] | layer3_out[1086];
    assign layer4_out[4100] = layer3_out[1739];
    assign layer4_out[4101] = ~layer3_out[6391] | layer3_out[6392];
    assign layer4_out[4102] = ~layer3_out[7629];
    assign layer4_out[4103] = layer3_out[4772] & ~layer3_out[4771];
    assign layer4_out[4104] = ~layer3_out[2315] | layer3_out[2316];
    assign layer4_out[4105] = layer3_out[606] & ~layer3_out[605];
    assign layer4_out[4106] = layer3_out[7133] ^ layer3_out[7134];
    assign layer4_out[4107] = layer3_out[1175] ^ layer3_out[1176];
    assign layer4_out[4108] = ~layer3_out[1052];
    assign layer4_out[4109] = ~(layer3_out[3456] ^ layer3_out[3457]);
    assign layer4_out[4110] = layer3_out[4843];
    assign layer4_out[4111] = ~(layer3_out[7006] & layer3_out[7007]);
    assign layer4_out[4112] = layer3_out[4941];
    assign layer4_out[4113] = ~layer3_out[4848];
    assign layer4_out[4114] = layer3_out[7200] | layer3_out[7201];
    assign layer4_out[4115] = layer3_out[39] & ~layer3_out[40];
    assign layer4_out[4116] = layer3_out[3023] | layer3_out[3024];
    assign layer4_out[4117] = ~layer3_out[1136] | layer3_out[1137];
    assign layer4_out[4118] = ~(layer3_out[595] | layer3_out[596]);
    assign layer4_out[4119] = layer3_out[7360] & layer3_out[7361];
    assign layer4_out[4120] = layer3_out[6592] ^ layer3_out[6593];
    assign layer4_out[4121] = ~layer3_out[7265] | layer3_out[7264];
    assign layer4_out[4122] = layer3_out[2209];
    assign layer4_out[4123] = ~layer3_out[3716];
    assign layer4_out[4124] = ~layer3_out[4887];
    assign layer4_out[4125] = ~(layer3_out[6760] & layer3_out[6761]);
    assign layer4_out[4126] = ~layer3_out[2107] | layer3_out[2108];
    assign layer4_out[4127] = layer3_out[6505];
    assign layer4_out[4128] = ~(layer3_out[988] | layer3_out[989]);
    assign layer4_out[4129] = ~layer3_out[450];
    assign layer4_out[4130] = ~layer3_out[7208] | layer3_out[7209];
    assign layer4_out[4131] = layer3_out[5497] & layer3_out[5498];
    assign layer4_out[4132] = layer3_out[514];
    assign layer4_out[4133] = layer3_out[4327] ^ layer3_out[4328];
    assign layer4_out[4134] = ~(layer3_out[4021] | layer3_out[4022]);
    assign layer4_out[4135] = ~(layer3_out[5821] | layer3_out[5822]);
    assign layer4_out[4136] = layer3_out[7591] & ~layer3_out[7592];
    assign layer4_out[4137] = ~(layer3_out[6978] & layer3_out[6979]);
    assign layer4_out[4138] = layer3_out[1751];
    assign layer4_out[4139] = layer3_out[360];
    assign layer4_out[4140] = ~layer3_out[1717];
    assign layer4_out[4141] = layer3_out[6741];
    assign layer4_out[4142] = layer3_out[7515];
    assign layer4_out[4143] = ~layer3_out[1130];
    assign layer4_out[4144] = ~layer3_out[7160];
    assign layer4_out[4145] = layer3_out[3473];
    assign layer4_out[4146] = ~layer3_out[7033] | layer3_out[7034];
    assign layer4_out[4147] = ~layer3_out[3369];
    assign layer4_out[4148] = layer3_out[726] ^ layer3_out[727];
    assign layer4_out[4149] = layer3_out[1257] | layer3_out[1258];
    assign layer4_out[4150] = ~layer3_out[7907] | layer3_out[7906];
    assign layer4_out[4151] = layer3_out[2431];
    assign layer4_out[4152] = ~layer3_out[1036];
    assign layer4_out[4153] = ~layer3_out[3593];
    assign layer4_out[4154] = layer3_out[3286] & ~layer3_out[3285];
    assign layer4_out[4155] = ~(layer3_out[4260] | layer3_out[4261]);
    assign layer4_out[4156] = ~layer3_out[5093];
    assign layer4_out[4157] = layer3_out[5866];
    assign layer4_out[4158] = layer3_out[1978] & ~layer3_out[1977];
    assign layer4_out[4159] = 1'b1;
    assign layer4_out[4160] = layer3_out[3410];
    assign layer4_out[4161] = ~(layer3_out[2543] ^ layer3_out[2544]);
    assign layer4_out[4162] = layer3_out[2048] ^ layer3_out[2049];
    assign layer4_out[4163] = ~layer3_out[4485];
    assign layer4_out[4164] = layer3_out[1115];
    assign layer4_out[4165] = layer3_out[6343];
    assign layer4_out[4166] = layer3_out[5786];
    assign layer4_out[4167] = ~layer3_out[6340];
    assign layer4_out[4168] = layer3_out[7902];
    assign layer4_out[4169] = ~layer3_out[3513];
    assign layer4_out[4170] = ~layer3_out[7358];
    assign layer4_out[4171] = layer3_out[5468] & layer3_out[5469];
    assign layer4_out[4172] = ~layer3_out[6522] | layer3_out[6523];
    assign layer4_out[4173] = ~layer3_out[7723];
    assign layer4_out[4174] = ~layer3_out[5659];
    assign layer4_out[4175] = ~layer3_out[420] | layer3_out[421];
    assign layer4_out[4176] = ~layer3_out[860];
    assign layer4_out[4177] = layer3_out[7097];
    assign layer4_out[4178] = layer3_out[435] ^ layer3_out[436];
    assign layer4_out[4179] = layer3_out[7711];
    assign layer4_out[4180] = layer3_out[3291];
    assign layer4_out[4181] = layer3_out[719];
    assign layer4_out[4182] = ~layer3_out[7714];
    assign layer4_out[4183] = layer3_out[4413] ^ layer3_out[4414];
    assign layer4_out[4184] = ~layer3_out[3871] | layer3_out[3872];
    assign layer4_out[4185] = layer3_out[371] | layer3_out[372];
    assign layer4_out[4186] = layer3_out[3991] & ~layer3_out[3992];
    assign layer4_out[4187] = ~layer3_out[5938] | layer3_out[5939];
    assign layer4_out[4188] = ~layer3_out[437] | layer3_out[436];
    assign layer4_out[4189] = ~layer3_out[376];
    assign layer4_out[4190] = layer3_out[3852];
    assign layer4_out[4191] = ~layer3_out[3354];
    assign layer4_out[4192] = layer3_out[1763] & layer3_out[1764];
    assign layer4_out[4193] = ~layer3_out[4646];
    assign layer4_out[4194] = ~(layer3_out[7700] ^ layer3_out[7701]);
    assign layer4_out[4195] = ~layer3_out[4466];
    assign layer4_out[4196] = ~layer3_out[998] | layer3_out[997];
    assign layer4_out[4197] = layer3_out[782];
    assign layer4_out[4198] = layer3_out[6151] & ~layer3_out[6152];
    assign layer4_out[4199] = ~(layer3_out[6965] | layer3_out[6966]);
    assign layer4_out[4200] = ~(layer3_out[3264] & layer3_out[3265]);
    assign layer4_out[4201] = ~(layer3_out[1374] | layer3_out[1375]);
    assign layer4_out[4202] = ~(layer3_out[7205] | layer3_out[7206]);
    assign layer4_out[4203] = ~layer3_out[7412];
    assign layer4_out[4204] = layer3_out[5386];
    assign layer4_out[4205] = layer3_out[7854];
    assign layer4_out[4206] = ~layer3_out[1701];
    assign layer4_out[4207] = ~layer3_out[7633];
    assign layer4_out[4208] = ~layer3_out[3426];
    assign layer4_out[4209] = ~(layer3_out[1663] & layer3_out[1664]);
    assign layer4_out[4210] = ~layer3_out[756];
    assign layer4_out[4211] = ~(layer3_out[4515] ^ layer3_out[4516]);
    assign layer4_out[4212] = layer3_out[7037] & ~layer3_out[7036];
    assign layer4_out[4213] = layer3_out[2600] & layer3_out[2601];
    assign layer4_out[4214] = layer3_out[1261] ^ layer3_out[1262];
    assign layer4_out[4215] = ~layer3_out[2415];
    assign layer4_out[4216] = ~layer3_out[6703];
    assign layer4_out[4217] = ~(layer3_out[2712] & layer3_out[2713]);
    assign layer4_out[4218] = layer3_out[540];
    assign layer4_out[4219] = layer3_out[2498] | layer3_out[2499];
    assign layer4_out[4220] = layer3_out[5929] & layer3_out[5930];
    assign layer4_out[4221] = ~(layer3_out[1192] | layer3_out[1193]);
    assign layer4_out[4222] = ~layer3_out[4510];
    assign layer4_out[4223] = ~layer3_out[1007];
    assign layer4_out[4224] = ~layer3_out[63];
    assign layer4_out[4225] = layer3_out[33];
    assign layer4_out[4226] = layer3_out[2852];
    assign layer4_out[4227] = layer3_out[6789];
    assign layer4_out[4228] = ~(layer3_out[7545] & layer3_out[7546]);
    assign layer4_out[4229] = ~layer3_out[1011];
    assign layer4_out[4230] = layer3_out[1587];
    assign layer4_out[4231] = ~layer3_out[510];
    assign layer4_out[4232] = layer3_out[846] & ~layer3_out[847];
    assign layer4_out[4233] = ~(layer3_out[6415] & layer3_out[6416]);
    assign layer4_out[4234] = ~layer3_out[4244] | layer3_out[4243];
    assign layer4_out[4235] = layer3_out[1895] & ~layer3_out[1896];
    assign layer4_out[4236] = ~layer3_out[6575];
    assign layer4_out[4237] = layer3_out[1503] | layer3_out[1504];
    assign layer4_out[4238] = ~layer3_out[1148];
    assign layer4_out[4239] = ~layer3_out[5461];
    assign layer4_out[4240] = ~layer3_out[2013];
    assign layer4_out[4241] = layer3_out[1203];
    assign layer4_out[4242] = ~layer3_out[4410];
    assign layer4_out[4243] = layer3_out[5460];
    assign layer4_out[4244] = layer3_out[4493] & layer3_out[4494];
    assign layer4_out[4245] = ~layer3_out[6437] | layer3_out[6438];
    assign layer4_out[4246] = layer3_out[1216] & layer3_out[1217];
    assign layer4_out[4247] = ~(layer3_out[2333] | layer3_out[2334]);
    assign layer4_out[4248] = layer3_out[7412] & layer3_out[7413];
    assign layer4_out[4249] = layer3_out[3915] | layer3_out[3916];
    assign layer4_out[4250] = layer3_out[6190] | layer3_out[6191];
    assign layer4_out[4251] = layer3_out[2051] & ~layer3_out[2050];
    assign layer4_out[4252] = layer3_out[744] ^ layer3_out[745];
    assign layer4_out[4253] = layer3_out[2998];
    assign layer4_out[4254] = ~(layer3_out[4587] ^ layer3_out[4588]);
    assign layer4_out[4255] = ~layer3_out[2038];
    assign layer4_out[4256] = ~(layer3_out[7513] & layer3_out[7514]);
    assign layer4_out[4257] = layer3_out[83] ^ layer3_out[84];
    assign layer4_out[4258] = ~layer3_out[401] | layer3_out[402];
    assign layer4_out[4259] = ~layer3_out[5684] | layer3_out[5683];
    assign layer4_out[4260] = ~layer3_out[34];
    assign layer4_out[4261] = ~layer3_out[4850];
    assign layer4_out[4262] = layer3_out[4540] ^ layer3_out[4541];
    assign layer4_out[4263] = ~layer3_out[4540] | layer3_out[4539];
    assign layer4_out[4264] = ~layer3_out[1448];
    assign layer4_out[4265] = layer3_out[4361];
    assign layer4_out[4266] = layer3_out[4768] | layer3_out[4769];
    assign layer4_out[4267] = layer3_out[4653];
    assign layer4_out[4268] = layer3_out[2563];
    assign layer4_out[4269] = ~(layer3_out[7252] ^ layer3_out[7253]);
    assign layer4_out[4270] = ~(layer3_out[4435] | layer3_out[4436]);
    assign layer4_out[4271] = ~layer3_out[1575];
    assign layer4_out[4272] = ~layer3_out[4736];
    assign layer4_out[4273] = layer3_out[933] & layer3_out[934];
    assign layer4_out[4274] = layer3_out[7283];
    assign layer4_out[4275] = ~(layer3_out[6133] | layer3_out[6134]);
    assign layer4_out[4276] = ~(layer3_out[227] | layer3_out[228]);
    assign layer4_out[4277] = ~layer3_out[868];
    assign layer4_out[4278] = layer3_out[3600];
    assign layer4_out[4279] = layer3_out[1705] | layer3_out[1706];
    assign layer4_out[4280] = layer3_out[7586];
    assign layer4_out[4281] = layer3_out[577] & ~layer3_out[576];
    assign layer4_out[4282] = ~(layer3_out[2787] & layer3_out[2788]);
    assign layer4_out[4283] = ~(layer3_out[6478] ^ layer3_out[6479]);
    assign layer4_out[4284] = layer3_out[3549] ^ layer3_out[3550];
    assign layer4_out[4285] = layer3_out[2237] & ~layer3_out[2238];
    assign layer4_out[4286] = layer3_out[3499] | layer3_out[3500];
    assign layer4_out[4287] = ~layer3_out[4780] | layer3_out[4781];
    assign layer4_out[4288] = ~layer3_out[1304];
    assign layer4_out[4289] = ~(layer3_out[1083] ^ layer3_out[1084]);
    assign layer4_out[4290] = ~layer3_out[5359] | layer3_out[5360];
    assign layer4_out[4291] = layer3_out[6811] & layer3_out[6812];
    assign layer4_out[4292] = ~layer3_out[5268];
    assign layer4_out[4293] = layer3_out[6694];
    assign layer4_out[4294] = ~layer3_out[7126];
    assign layer4_out[4295] = layer3_out[370] & ~layer3_out[369];
    assign layer4_out[4296] = layer3_out[4800] | layer3_out[4801];
    assign layer4_out[4297] = ~(layer3_out[4817] ^ layer3_out[4818]);
    assign layer4_out[4298] = ~(layer3_out[7401] ^ layer3_out[7402]);
    assign layer4_out[4299] = ~layer3_out[4501] | layer3_out[4502];
    assign layer4_out[4300] = ~layer3_out[721];
    assign layer4_out[4301] = layer3_out[1914] & ~layer3_out[1913];
    assign layer4_out[4302] = ~layer3_out[2914] | layer3_out[2915];
    assign layer4_out[4303] = layer3_out[7092];
    assign layer4_out[4304] = ~layer3_out[2100];
    assign layer4_out[4305] = layer3_out[1559] ^ layer3_out[1560];
    assign layer4_out[4306] = ~layer3_out[85];
    assign layer4_out[4307] = layer3_out[1333] & ~layer3_out[1332];
    assign layer4_out[4308] = ~layer3_out[93];
    assign layer4_out[4309] = ~layer3_out[2566];
    assign layer4_out[4310] = ~layer3_out[3999];
    assign layer4_out[4311] = ~(layer3_out[6817] ^ layer3_out[6818]);
    assign layer4_out[4312] = ~layer3_out[1356];
    assign layer4_out[4313] = ~layer3_out[709];
    assign layer4_out[4314] = layer3_out[2599] | layer3_out[2600];
    assign layer4_out[4315] = ~(layer3_out[1243] | layer3_out[1244]);
    assign layer4_out[4316] = ~(layer3_out[5285] ^ layer3_out[5286]);
    assign layer4_out[4317] = ~layer3_out[2145];
    assign layer4_out[4318] = layer3_out[357];
    assign layer4_out[4319] = ~(layer3_out[7340] | layer3_out[7341]);
    assign layer4_out[4320] = ~layer3_out[4739];
    assign layer4_out[4321] = layer3_out[5607] ^ layer3_out[5608];
    assign layer4_out[4322] = layer3_out[1385] & layer3_out[1386];
    assign layer4_out[4323] = ~(layer3_out[3616] ^ layer3_out[3617]);
    assign layer4_out[4324] = ~layer3_out[7731] | layer3_out[7732];
    assign layer4_out[4325] = layer3_out[3251];
    assign layer4_out[4326] = ~layer3_out[6048];
    assign layer4_out[4327] = layer3_out[284] | layer3_out[285];
    assign layer4_out[4328] = layer3_out[7829] & layer3_out[7830];
    assign layer4_out[4329] = ~layer3_out[82] | layer3_out[83];
    assign layer4_out[4330] = layer3_out[5153];
    assign layer4_out[4331] = layer3_out[1290] & layer3_out[1291];
    assign layer4_out[4332] = layer3_out[1371] & ~layer3_out[1372];
    assign layer4_out[4333] = ~layer3_out[6595];
    assign layer4_out[4334] = layer3_out[879];
    assign layer4_out[4335] = layer3_out[450] & ~layer3_out[451];
    assign layer4_out[4336] = ~layer3_out[5750];
    assign layer4_out[4337] = layer3_out[5596] | layer3_out[5597];
    assign layer4_out[4338] = ~(layer3_out[5512] | layer3_out[5513]);
    assign layer4_out[4339] = layer3_out[4307] & ~layer3_out[4306];
    assign layer4_out[4340] = layer3_out[5603] & layer3_out[5604];
    assign layer4_out[4341] = 1'b0;
    assign layer4_out[4342] = ~(layer3_out[3360] | layer3_out[3361]);
    assign layer4_out[4343] = ~layer3_out[2883];
    assign layer4_out[4344] = ~layer3_out[2829];
    assign layer4_out[4345] = layer3_out[780] ^ layer3_out[781];
    assign layer4_out[4346] = ~layer3_out[2441];
    assign layer4_out[4347] = ~layer3_out[366];
    assign layer4_out[4348] = ~(layer3_out[7381] ^ layer3_out[7382]);
    assign layer4_out[4349] = 1'b1;
    assign layer4_out[4350] = ~layer3_out[1790];
    assign layer4_out[4351] = layer3_out[4995] | layer3_out[4996];
    assign layer4_out[4352] = ~layer3_out[5853] | layer3_out[5854];
    assign layer4_out[4353] = layer3_out[6728] | layer3_out[6729];
    assign layer4_out[4354] = layer3_out[7852];
    assign layer4_out[4355] = layer3_out[1134] ^ layer3_out[1135];
    assign layer4_out[4356] = ~(layer3_out[7898] ^ layer3_out[7899]);
    assign layer4_out[4357] = ~layer3_out[2379];
    assign layer4_out[4358] = layer3_out[4724] & ~layer3_out[4723];
    assign layer4_out[4359] = ~(layer3_out[7644] | layer3_out[7645]);
    assign layer4_out[4360] = ~layer3_out[3144];
    assign layer4_out[4361] = layer3_out[3461] ^ layer3_out[3462];
    assign layer4_out[4362] = ~layer3_out[6939] | layer3_out[6940];
    assign layer4_out[4363] = ~layer3_out[140];
    assign layer4_out[4364] = layer3_out[3517];
    assign layer4_out[4365] = ~(layer3_out[5884] ^ layer3_out[5885]);
    assign layer4_out[4366] = layer3_out[3522];
    assign layer4_out[4367] = ~layer3_out[5690];
    assign layer4_out[4368] = ~layer3_out[404];
    assign layer4_out[4369] = layer3_out[5582];
    assign layer4_out[4370] = ~layer3_out[2667];
    assign layer4_out[4371] = layer3_out[1532];
    assign layer4_out[4372] = ~(layer3_out[1859] & layer3_out[1860]);
    assign layer4_out[4373] = layer3_out[111] | layer3_out[112];
    assign layer4_out[4374] = ~layer3_out[5317] | layer3_out[5316];
    assign layer4_out[4375] = ~layer3_out[1280];
    assign layer4_out[4376] = layer3_out[3640] & ~layer3_out[3641];
    assign layer4_out[4377] = layer3_out[1530] | layer3_out[1531];
    assign layer4_out[4378] = ~layer3_out[6759];
    assign layer4_out[4379] = layer3_out[5463] & ~layer3_out[5464];
    assign layer4_out[4380] = ~(layer3_out[996] & layer3_out[997]);
    assign layer4_out[4381] = ~(layer3_out[4139] & layer3_out[4140]);
    assign layer4_out[4382] = 1'b0;
    assign layer4_out[4383] = layer3_out[879];
    assign layer4_out[4384] = layer3_out[5698] & ~layer3_out[5697];
    assign layer4_out[4385] = layer3_out[7908] & layer3_out[7909];
    assign layer4_out[4386] = ~layer3_out[5985];
    assign layer4_out[4387] = ~layer3_out[742];
    assign layer4_out[4388] = ~layer3_out[7710];
    assign layer4_out[4389] = ~layer3_out[6312];
    assign layer4_out[4390] = layer3_out[1985];
    assign layer4_out[4391] = layer3_out[1452] & ~layer3_out[1453];
    assign layer4_out[4392] = layer3_out[7958] & ~layer3_out[7957];
    assign layer4_out[4393] = ~layer3_out[3006] | layer3_out[3005];
    assign layer4_out[4394] = layer3_out[5079] & layer3_out[5080];
    assign layer4_out[4395] = layer3_out[5311];
    assign layer4_out[4396] = ~layer3_out[6388];
    assign layer4_out[4397] = ~layer3_out[5846] | layer3_out[5845];
    assign layer4_out[4398] = ~(layer3_out[1570] ^ layer3_out[1571]);
    assign layer4_out[4399] = 1'b0;
    assign layer4_out[4400] = layer3_out[5837] ^ layer3_out[5838];
    assign layer4_out[4401] = layer3_out[6844] ^ layer3_out[6845];
    assign layer4_out[4402] = 1'b0;
    assign layer4_out[4403] = ~layer3_out[2435] | layer3_out[2434];
    assign layer4_out[4404] = layer3_out[4885] | layer3_out[4886];
    assign layer4_out[4405] = ~(layer3_out[916] & layer3_out[917]);
    assign layer4_out[4406] = layer3_out[1920] ^ layer3_out[1921];
    assign layer4_out[4407] = ~layer3_out[5860];
    assign layer4_out[4408] = ~(layer3_out[4744] ^ layer3_out[4745]);
    assign layer4_out[4409] = ~layer3_out[660] | layer3_out[661];
    assign layer4_out[4410] = layer3_out[1008] ^ layer3_out[1009];
    assign layer4_out[4411] = layer3_out[2259];
    assign layer4_out[4412] = layer3_out[864] & ~layer3_out[865];
    assign layer4_out[4413] = ~(layer3_out[6724] & layer3_out[6725]);
    assign layer4_out[4414] = ~(layer3_out[4227] & layer3_out[4228]);
    assign layer4_out[4415] = layer3_out[2885] & ~layer3_out[2886];
    assign layer4_out[4416] = layer3_out[1534];
    assign layer4_out[4417] = ~layer3_out[471];
    assign layer4_out[4418] = ~layer3_out[1141];
    assign layer4_out[4419] = ~layer3_out[5765];
    assign layer4_out[4420] = ~(layer3_out[231] & layer3_out[232]);
    assign layer4_out[4421] = ~(layer3_out[2263] | layer3_out[2264]);
    assign layer4_out[4422] = layer3_out[4687] & ~layer3_out[4688];
    assign layer4_out[4423] = ~layer3_out[4090];
    assign layer4_out[4424] = 1'b0;
    assign layer4_out[4425] = ~layer3_out[5761];
    assign layer4_out[4426] = ~layer3_out[948];
    assign layer4_out[4427] = layer3_out[2053];
    assign layer4_out[4428] = ~layer3_out[693];
    assign layer4_out[4429] = 1'b0;
    assign layer4_out[4430] = layer3_out[6161];
    assign layer4_out[4431] = layer3_out[2875];
    assign layer4_out[4432] = layer3_out[3914];
    assign layer4_out[4433] = ~layer3_out[7561];
    assign layer4_out[4434] = layer3_out[5969] ^ layer3_out[5970];
    assign layer4_out[4435] = layer3_out[4272];
    assign layer4_out[4436] = layer3_out[7164];
    assign layer4_out[4437] = layer3_out[6956] & layer3_out[6957];
    assign layer4_out[4438] = layer3_out[247];
    assign layer4_out[4439] = ~layer3_out[1699];
    assign layer4_out[4440] = layer3_out[1139];
    assign layer4_out[4441] = ~layer3_out[7236];
    assign layer4_out[4442] = ~layer3_out[6404];
    assign layer4_out[4443] = ~(layer3_out[5539] ^ layer3_out[5540]);
    assign layer4_out[4444] = layer3_out[1646];
    assign layer4_out[4445] = layer3_out[1197];
    assign layer4_out[4446] = ~(layer3_out[2861] ^ layer3_out[2862]);
    assign layer4_out[4447] = ~layer3_out[674] | layer3_out[675];
    assign layer4_out[4448] = layer3_out[6874] & layer3_out[6875];
    assign layer4_out[4449] = ~layer3_out[7140] | layer3_out[7141];
    assign layer4_out[4450] = layer3_out[7921];
    assign layer4_out[4451] = layer3_out[5282];
    assign layer4_out[4452] = ~layer3_out[6100];
    assign layer4_out[4453] = ~layer3_out[7643] | layer3_out[7644];
    assign layer4_out[4454] = ~layer3_out[5695] | layer3_out[5696];
    assign layer4_out[4455] = ~(layer3_out[6452] ^ layer3_out[6453]);
    assign layer4_out[4456] = 1'b1;
    assign layer4_out[4457] = layer3_out[6838];
    assign layer4_out[4458] = ~(layer3_out[4958] | layer3_out[4959]);
    assign layer4_out[4459] = ~layer3_out[2156];
    assign layer4_out[4460] = ~layer3_out[3651];
    assign layer4_out[4461] = ~(layer3_out[7519] ^ layer3_out[7520]);
    assign layer4_out[4462] = layer3_out[1129];
    assign layer4_out[4463] = ~layer3_out[3099];
    assign layer4_out[4464] = ~(layer3_out[6775] | layer3_out[6776]);
    assign layer4_out[4465] = layer3_out[7719];
    assign layer4_out[4466] = ~layer3_out[6797];
    assign layer4_out[4467] = layer3_out[3917];
    assign layer4_out[4468] = ~layer3_out[3102];
    assign layer4_out[4469] = layer3_out[1214] | layer3_out[1215];
    assign layer4_out[4470] = layer3_out[6027];
    assign layer4_out[4471] = ~(layer3_out[5429] ^ layer3_out[5430]);
    assign layer4_out[4472] = ~(layer3_out[4457] | layer3_out[4458]);
    assign layer4_out[4473] = ~(layer3_out[7013] & layer3_out[7014]);
    assign layer4_out[4474] = layer3_out[257] ^ layer3_out[258];
    assign layer4_out[4475] = layer3_out[6893] & layer3_out[6894];
    assign layer4_out[4476] = ~(layer3_out[7773] & layer3_out[7774]);
    assign layer4_out[4477] = layer3_out[1125] & layer3_out[1126];
    assign layer4_out[4478] = layer3_out[486] & ~layer3_out[485];
    assign layer4_out[4479] = layer3_out[3254] & ~layer3_out[3253];
    assign layer4_out[4480] = layer3_out[5576];
    assign layer4_out[4481] = layer3_out[3385];
    assign layer4_out[4482] = ~layer3_out[2080] | layer3_out[2081];
    assign layer4_out[4483] = layer3_out[3847] ^ layer3_out[3848];
    assign layer4_out[4484] = ~layer3_out[4789] | layer3_out[4788];
    assign layer4_out[4485] = ~(layer3_out[7279] & layer3_out[7280]);
    assign layer4_out[4486] = layer3_out[3110];
    assign layer4_out[4487] = layer3_out[3604];
    assign layer4_out[4488] = ~(layer3_out[4594] & layer3_out[4595]);
    assign layer4_out[4489] = ~layer3_out[685];
    assign layer4_out[4490] = layer3_out[6045];
    assign layer4_out[4491] = ~layer3_out[891];
    assign layer4_out[4492] = ~(layer3_out[5341] & layer3_out[5342]);
    assign layer4_out[4493] = layer3_out[5276] | layer3_out[5277];
    assign layer4_out[4494] = ~layer3_out[3968];
    assign layer4_out[4495] = ~layer3_out[6164];
    assign layer4_out[4496] = ~layer3_out[1338] | layer3_out[1337];
    assign layer4_out[4497] = ~layer3_out[2380];
    assign layer4_out[4498] = layer3_out[7601];
    assign layer4_out[4499] = ~layer3_out[3064] | layer3_out[3063];
    assign layer4_out[4500] = layer3_out[295] & layer3_out[296];
    assign layer4_out[4501] = ~layer3_out[4153];
    assign layer4_out[4502] = layer3_out[118] & layer3_out[119];
    assign layer4_out[4503] = layer3_out[6607] ^ layer3_out[6608];
    assign layer4_out[4504] = layer3_out[7216] | layer3_out[7217];
    assign layer4_out[4505] = layer3_out[5887] & ~layer3_out[5888];
    assign layer4_out[4506] = ~layer3_out[1231];
    assign layer4_out[4507] = ~(layer3_out[4198] ^ layer3_out[4199]);
    assign layer4_out[4508] = ~layer3_out[2961] | layer3_out[2960];
    assign layer4_out[4509] = ~(layer3_out[3543] | layer3_out[3544]);
    assign layer4_out[4510] = layer3_out[5887];
    assign layer4_out[4511] = layer3_out[5398];
    assign layer4_out[4512] = ~layer3_out[5816];
    assign layer4_out[4513] = 1'b0;
    assign layer4_out[4514] = ~layer3_out[2524] | layer3_out[2525];
    assign layer4_out[4515] = ~(layer3_out[3483] ^ layer3_out[3484]);
    assign layer4_out[4516] = ~(layer3_out[7924] ^ layer3_out[7925]);
    assign layer4_out[4517] = layer3_out[5172] & layer3_out[5173];
    assign layer4_out[4518] = layer3_out[3775] ^ layer3_out[3776];
    assign layer4_out[4519] = layer3_out[180] ^ layer3_out[181];
    assign layer4_out[4520] = ~layer3_out[2315];
    assign layer4_out[4521] = layer3_out[3566] & ~layer3_out[3565];
    assign layer4_out[4522] = layer3_out[7906];
    assign layer4_out[4523] = layer3_out[4488];
    assign layer4_out[4524] = ~layer3_out[4051];
    assign layer4_out[4525] = ~layer3_out[3806];
    assign layer4_out[4526] = ~layer3_out[587] | layer3_out[586];
    assign layer4_out[4527] = ~layer3_out[5370] | layer3_out[5371];
    assign layer4_out[4528] = ~layer3_out[5416] | layer3_out[5417];
    assign layer4_out[4529] = ~(layer3_out[5402] & layer3_out[5403]);
    assign layer4_out[4530] = ~layer3_out[1767];
    assign layer4_out[4531] = layer3_out[1314] ^ layer3_out[1315];
    assign layer4_out[4532] = layer3_out[1344] | layer3_out[1345];
    assign layer4_out[4533] = layer3_out[1245] ^ layer3_out[1246];
    assign layer4_out[4534] = layer3_out[6778] & ~layer3_out[6779];
    assign layer4_out[4535] = ~layer3_out[87] | layer3_out[88];
    assign layer4_out[4536] = ~layer3_out[6494];
    assign layer4_out[4537] = layer3_out[3236];
    assign layer4_out[4538] = ~layer3_out[4212];
    assign layer4_out[4539] = ~(layer3_out[6900] | layer3_out[6901]);
    assign layer4_out[4540] = ~layer3_out[2092];
    assign layer4_out[4541] = layer3_out[2230];
    assign layer4_out[4542] = ~(layer3_out[3389] ^ layer3_out[3390]);
    assign layer4_out[4543] = layer3_out[783] & ~layer3_out[784];
    assign layer4_out[4544] = layer3_out[4699] & ~layer3_out[4698];
    assign layer4_out[4545] = layer3_out[45];
    assign layer4_out[4546] = layer3_out[1811];
    assign layer4_out[4547] = ~layer3_out[3787] | layer3_out[3788];
    assign layer4_out[4548] = ~layer3_out[2730];
    assign layer4_out[4549] = layer3_out[3613] & layer3_out[3614];
    assign layer4_out[4550] = layer3_out[6221] & ~layer3_out[6222];
    assign layer4_out[4551] = layer3_out[4526];
    assign layer4_out[4552] = layer3_out[2654] ^ layer3_out[2655];
    assign layer4_out[4553] = layer3_out[5861] & layer3_out[5862];
    assign layer4_out[4554] = layer3_out[5755] & ~layer3_out[5754];
    assign layer4_out[4555] = ~(layer3_out[7991] & layer3_out[7992]);
    assign layer4_out[4556] = layer3_out[6665] & ~layer3_out[6666];
    assign layer4_out[4557] = layer3_out[213] ^ layer3_out[214];
    assign layer4_out[4558] = layer3_out[2358];
    assign layer4_out[4559] = layer3_out[5551];
    assign layer4_out[4560] = ~layer3_out[3211] | layer3_out[3210];
    assign layer4_out[4561] = ~layer3_out[5652];
    assign layer4_out[4562] = ~layer3_out[6852];
    assign layer4_out[4563] = layer3_out[2663];
    assign layer4_out[4564] = ~layer3_out[3375] | layer3_out[3374];
    assign layer4_out[4565] = ~layer3_out[5083];
    assign layer4_out[4566] = layer3_out[2741] & ~layer3_out[2740];
    assign layer4_out[4567] = ~layer3_out[6712] | layer3_out[6711];
    assign layer4_out[4568] = layer3_out[13];
    assign layer4_out[4569] = layer3_out[2625] & layer3_out[2626];
    assign layer4_out[4570] = layer3_out[4344] & ~layer3_out[4345];
    assign layer4_out[4571] = layer3_out[5300];
    assign layer4_out[4572] = ~(layer3_out[4978] | layer3_out[4979]);
    assign layer4_out[4573] = ~layer3_out[3765];
    assign layer4_out[4574] = ~layer3_out[2463];
    assign layer4_out[4575] = ~layer3_out[5922];
    assign layer4_out[4576] = ~(layer3_out[3952] ^ layer3_out[3953]);
    assign layer4_out[4577] = layer3_out[3552] | layer3_out[3553];
    assign layer4_out[4578] = layer3_out[6348] & layer3_out[6349];
    assign layer4_out[4579] = layer3_out[4995];
    assign layer4_out[4580] = layer3_out[109] & ~layer3_out[108];
    assign layer4_out[4581] = layer3_out[7853];
    assign layer4_out[4582] = ~layer3_out[1037] | layer3_out[1038];
    assign layer4_out[4583] = layer3_out[4861] & layer3_out[4862];
    assign layer4_out[4584] = layer3_out[7902] & ~layer3_out[7901];
    assign layer4_out[4585] = layer3_out[2103];
    assign layer4_out[4586] = ~(layer3_out[7566] ^ layer3_out[7567]);
    assign layer4_out[4587] = ~(layer3_out[3268] | layer3_out[3269]);
    assign layer4_out[4588] = layer3_out[469];
    assign layer4_out[4589] = ~layer3_out[2132] | layer3_out[2131];
    assign layer4_out[4590] = ~layer3_out[164];
    assign layer4_out[4591] = ~layer3_out[3448] | layer3_out[3449];
    assign layer4_out[4592] = ~layer3_out[4673];
    assign layer4_out[4593] = layer3_out[2521];
    assign layer4_out[4594] = layer3_out[2629];
    assign layer4_out[4595] = ~(layer3_out[4658] | layer3_out[4659]);
    assign layer4_out[4596] = ~layer3_out[5599];
    assign layer4_out[4597] = layer3_out[1321];
    assign layer4_out[4598] = layer3_out[7705] ^ layer3_out[7706];
    assign layer4_out[4599] = ~(layer3_out[580] | layer3_out[581]);
    assign layer4_out[4600] = layer3_out[2458] | layer3_out[2459];
    assign layer4_out[4601] = ~layer3_out[3098] | layer3_out[3099];
    assign layer4_out[4602] = ~layer3_out[3642];
    assign layer4_out[4603] = layer3_out[4419];
    assign layer4_out[4604] = ~layer3_out[6471];
    assign layer4_out[4605] = ~layer3_out[6742];
    assign layer4_out[4606] = layer3_out[4644] & ~layer3_out[4645];
    assign layer4_out[4607] = ~layer3_out[5991];
    assign layer4_out[4608] = ~layer3_out[669] | layer3_out[668];
    assign layer4_out[4609] = layer3_out[2317] ^ layer3_out[2318];
    assign layer4_out[4610] = layer3_out[2273] & ~layer3_out[2274];
    assign layer4_out[4611] = layer3_out[3432];
    assign layer4_out[4612] = layer3_out[3673];
    assign layer4_out[4613] = ~layer3_out[6673];
    assign layer4_out[4614] = ~layer3_out[6975] | layer3_out[6974];
    assign layer4_out[4615] = layer3_out[4662] ^ layer3_out[4663];
    assign layer4_out[4616] = ~(layer3_out[7782] ^ layer3_out[7783]);
    assign layer4_out[4617] = layer3_out[1848] ^ layer3_out[1849];
    assign layer4_out[4618] = 1'b0;
    assign layer4_out[4619] = ~(layer3_out[1179] | layer3_out[1180]);
    assign layer4_out[4620] = ~(layer3_out[3347] | layer3_out[3348]);
    assign layer4_out[4621] = ~layer3_out[3661];
    assign layer4_out[4622] = ~layer3_out[4996];
    assign layer4_out[4623] = layer3_out[52] & layer3_out[53];
    assign layer4_out[4624] = layer3_out[258] | layer3_out[259];
    assign layer4_out[4625] = ~(layer3_out[2183] ^ layer3_out[2184]);
    assign layer4_out[4626] = layer3_out[5598];
    assign layer4_out[4627] = ~layer3_out[7777];
    assign layer4_out[4628] = ~layer3_out[5219];
    assign layer4_out[4629] = layer3_out[81] ^ layer3_out[82];
    assign layer4_out[4630] = layer3_out[1316];
    assign layer4_out[4631] = ~(layer3_out[2807] ^ layer3_out[2808]);
    assign layer4_out[4632] = ~(layer3_out[7520] & layer3_out[7521]);
    assign layer4_out[4633] = layer3_out[7014] | layer3_out[7015];
    assign layer4_out[4634] = ~(layer3_out[1989] & layer3_out[1990]);
    assign layer4_out[4635] = 1'b0;
    assign layer4_out[4636] = ~layer3_out[6530] | layer3_out[6531];
    assign layer4_out[4637] = ~(layer3_out[2001] ^ layer3_out[2002]);
    assign layer4_out[4638] = ~layer3_out[6220] | layer3_out[6221];
    assign layer4_out[4639] = ~(layer3_out[3246] & layer3_out[3247]);
    assign layer4_out[4640] = layer3_out[6234] ^ layer3_out[6235];
    assign layer4_out[4641] = layer3_out[1385];
    assign layer4_out[4642] = layer3_out[4503];
    assign layer4_out[4643] = layer3_out[1836] ^ layer3_out[1837];
    assign layer4_out[4644] = ~(layer3_out[3503] ^ layer3_out[3504]);
    assign layer4_out[4645] = ~layer3_out[2152] | layer3_out[2153];
    assign layer4_out[4646] = layer3_out[7124];
    assign layer4_out[4647] = layer3_out[452] & ~layer3_out[451];
    assign layer4_out[4648] = ~(layer3_out[1771] | layer3_out[1772]);
    assign layer4_out[4649] = ~layer3_out[1956];
    assign layer4_out[4650] = ~(layer3_out[7609] & layer3_out[7610]);
    assign layer4_out[4651] = ~layer3_out[3506];
    assign layer4_out[4652] = ~layer3_out[1272];
    assign layer4_out[4653] = ~(layer3_out[2859] | layer3_out[2860]);
    assign layer4_out[4654] = ~(layer3_out[4025] ^ layer3_out[4026]);
    assign layer4_out[4655] = ~layer3_out[3595];
    assign layer4_out[4656] = layer3_out[1075];
    assign layer4_out[4657] = layer3_out[5630] & layer3_out[5631];
    assign layer4_out[4658] = layer3_out[5329];
    assign layer4_out[4659] = layer3_out[2806];
    assign layer4_out[4660] = ~layer3_out[3276];
    assign layer4_out[4661] = layer3_out[1645];
    assign layer4_out[4662] = layer3_out[2127] & layer3_out[2128];
    assign layer4_out[4663] = ~layer3_out[7616];
    assign layer4_out[4664] = ~layer3_out[3420] | layer3_out[3421];
    assign layer4_out[4665] = ~(layer3_out[3537] | layer3_out[3538]);
    assign layer4_out[4666] = layer3_out[132];
    assign layer4_out[4667] = ~layer3_out[7564];
    assign layer4_out[4668] = ~layer3_out[1376];
    assign layer4_out[4669] = ~layer3_out[2595];
    assign layer4_out[4670] = layer3_out[6724];
    assign layer4_out[4671] = ~layer3_out[7339];
    assign layer4_out[4672] = layer3_out[2996];
    assign layer4_out[4673] = ~(layer3_out[1795] ^ layer3_out[1796]);
    assign layer4_out[4674] = ~(layer3_out[1695] ^ layer3_out[1696]);
    assign layer4_out[4675] = layer3_out[1278];
    assign layer4_out[4676] = layer3_out[298];
    assign layer4_out[4677] = ~layer3_out[4178];
    assign layer4_out[4678] = layer3_out[4292] & layer3_out[4293];
    assign layer4_out[4679] = ~(layer3_out[3862] ^ layer3_out[3863]);
    assign layer4_out[4680] = layer3_out[2608];
    assign layer4_out[4681] = layer3_out[6916] & layer3_out[6917];
    assign layer4_out[4682] = ~(layer3_out[2867] & layer3_out[2868]);
    assign layer4_out[4683] = ~layer3_out[5373] | layer3_out[5374];
    assign layer4_out[4684] = layer3_out[1750] | layer3_out[1751];
    assign layer4_out[4685] = layer3_out[5734];
    assign layer4_out[4686] = ~layer3_out[2693] | layer3_out[2692];
    assign layer4_out[4687] = layer3_out[5505];
    assign layer4_out[4688] = layer3_out[3557];
    assign layer4_out[4689] = ~layer3_out[1686];
    assign layer4_out[4690] = ~layer3_out[6155];
    assign layer4_out[4691] = layer3_out[4161] | layer3_out[4162];
    assign layer4_out[4692] = layer3_out[4215] & layer3_out[4216];
    assign layer4_out[4693] = ~(layer3_out[1972] & layer3_out[1973]);
    assign layer4_out[4694] = layer3_out[6544];
    assign layer4_out[4695] = ~layer3_out[2547];
    assign layer4_out[4696] = layer3_out[5625];
    assign layer4_out[4697] = layer3_out[6422] & ~layer3_out[6423];
    assign layer4_out[4698] = layer3_out[5343] ^ layer3_out[5344];
    assign layer4_out[4699] = ~layer3_out[6998] | layer3_out[6999];
    assign layer4_out[4700] = layer3_out[7414];
    assign layer4_out[4701] = ~(layer3_out[6248] ^ layer3_out[6249]);
    assign layer4_out[4702] = layer3_out[3939] ^ layer3_out[3940];
    assign layer4_out[4703] = ~layer3_out[7965];
    assign layer4_out[4704] = ~layer3_out[240] | layer3_out[241];
    assign layer4_out[4705] = ~layer3_out[4298] | layer3_out[4299];
    assign layer4_out[4706] = ~(layer3_out[5115] & layer3_out[5116]);
    assign layer4_out[4707] = layer3_out[2567] | layer3_out[2568];
    assign layer4_out[4708] = ~layer3_out[3865] | layer3_out[3866];
    assign layer4_out[4709] = layer3_out[6051] & ~layer3_out[6050];
    assign layer4_out[4710] = ~layer3_out[4176];
    assign layer4_out[4711] = ~(layer3_out[7405] ^ layer3_out[7406]);
    assign layer4_out[4712] = layer3_out[3223] & ~layer3_out[3224];
    assign layer4_out[4713] = layer3_out[6990];
    assign layer4_out[4714] = ~layer3_out[5386];
    assign layer4_out[4715] = ~layer3_out[7089];
    assign layer4_out[4716] = ~layer3_out[3801];
    assign layer4_out[4717] = ~layer3_out[338];
    assign layer4_out[4718] = ~(layer3_out[6180] | layer3_out[6181]);
    assign layer4_out[4719] = layer3_out[3426] ^ layer3_out[3427];
    assign layer4_out[4720] = layer3_out[6514];
    assign layer4_out[4721] = layer3_out[2592] & ~layer3_out[2593];
    assign layer4_out[4722] = ~layer3_out[1693];
    assign layer4_out[4723] = ~layer3_out[1209];
    assign layer4_out[4724] = ~layer3_out[4144];
    assign layer4_out[4725] = layer3_out[210] ^ layer3_out[211];
    assign layer4_out[4726] = 1'b1;
    assign layer4_out[4727] = layer3_out[6110] | layer3_out[6111];
    assign layer4_out[4728] = layer3_out[7057] ^ layer3_out[7058];
    assign layer4_out[4729] = layer3_out[2475] & layer3_out[2476];
    assign layer4_out[4730] = ~(layer3_out[2848] ^ layer3_out[2849]);
    assign layer4_out[4731] = ~layer3_out[7443];
    assign layer4_out[4732] = ~(layer3_out[2194] ^ layer3_out[2195]);
    assign layer4_out[4733] = ~(layer3_out[6449] | layer3_out[6450]);
    assign layer4_out[4734] = ~layer3_out[1271];
    assign layer4_out[4735] = layer3_out[816] & ~layer3_out[817];
    assign layer4_out[4736] = ~layer3_out[4362] | layer3_out[4361];
    assign layer4_out[4737] = layer3_out[7345] | layer3_out[7346];
    assign layer4_out[4738] = ~(layer3_out[1548] ^ layer3_out[1549]);
    assign layer4_out[4739] = layer3_out[2418] | layer3_out[2419];
    assign layer4_out[4740] = ~layer3_out[2740];
    assign layer4_out[4741] = layer3_out[5126] & layer3_out[5127];
    assign layer4_out[4742] = ~layer3_out[3198];
    assign layer4_out[4743] = layer3_out[3939] & ~layer3_out[3938];
    assign layer4_out[4744] = layer3_out[601] & ~layer3_out[602];
    assign layer4_out[4745] = ~(layer3_out[6624] ^ layer3_out[6625]);
    assign layer4_out[4746] = layer3_out[6126];
    assign layer4_out[4747] = layer3_out[4866] ^ layer3_out[4867];
    assign layer4_out[4748] = ~(layer3_out[2581] | layer3_out[2582]);
    assign layer4_out[4749] = layer3_out[5817] ^ layer3_out[5818];
    assign layer4_out[4750] = layer3_out[7750] & ~layer3_out[7749];
    assign layer4_out[4751] = ~(layer3_out[1538] & layer3_out[1539]);
    assign layer4_out[4752] = ~(layer3_out[4145] ^ layer3_out[4146]);
    assign layer4_out[4753] = layer3_out[1560];
    assign layer4_out[4754] = layer3_out[4810] & ~layer3_out[4811];
    assign layer4_out[4755] = ~layer3_out[579] | layer3_out[580];
    assign layer4_out[4756] = layer3_out[1342];
    assign layer4_out[4757] = ~layer3_out[1143];
    assign layer4_out[4758] = ~layer3_out[5474];
    assign layer4_out[4759] = layer3_out[1815];
    assign layer4_out[4760] = layer3_out[6546] & ~layer3_out[6547];
    assign layer4_out[4761] = ~layer3_out[2289];
    assign layer4_out[4762] = ~layer3_out[532] | layer3_out[531];
    assign layer4_out[4763] = ~layer3_out[5704];
    assign layer4_out[4764] = ~(layer3_out[4246] ^ layer3_out[4247]);
    assign layer4_out[4765] = ~layer3_out[7791];
    assign layer4_out[4766] = layer3_out[663];
    assign layer4_out[4767] = layer3_out[5337] & layer3_out[5338];
    assign layer4_out[4768] = layer3_out[2883] ^ layer3_out[2884];
    assign layer4_out[4769] = ~layer3_out[7431] | layer3_out[7430];
    assign layer4_out[4770] = ~layer3_out[7649];
    assign layer4_out[4771] = ~(layer3_out[225] ^ layer3_out[226]);
    assign layer4_out[4772] = layer3_out[6142];
    assign layer4_out[4773] = layer3_out[7384] & ~layer3_out[7385];
    assign layer4_out[4774] = ~layer3_out[1301] | layer3_out[1302];
    assign layer4_out[4775] = ~layer3_out[1742];
    assign layer4_out[4776] = layer3_out[2355] ^ layer3_out[2356];
    assign layer4_out[4777] = layer3_out[5960] & ~layer3_out[5961];
    assign layer4_out[4778] = layer3_out[4201];
    assign layer4_out[4779] = layer3_out[6491];
    assign layer4_out[4780] = ~layer3_out[4250] | layer3_out[4249];
    assign layer4_out[4781] = ~(layer3_out[4309] & layer3_out[4310]);
    assign layer4_out[4782] = ~layer3_out[5758];
    assign layer4_out[4783] = layer3_out[7339];
    assign layer4_out[4784] = ~layer3_out[7539] | layer3_out[7538];
    assign layer4_out[4785] = layer3_out[2438];
    assign layer4_out[4786] = ~layer3_out[3405];
    assign layer4_out[4787] = ~(layer3_out[3789] ^ layer3_out[3790]);
    assign layer4_out[4788] = layer3_out[7498];
    assign layer4_out[4789] = ~(layer3_out[1606] ^ layer3_out[1607]);
    assign layer4_out[4790] = ~(layer3_out[4568] ^ layer3_out[4569]);
    assign layer4_out[4791] = layer3_out[4111] & ~layer3_out[4110];
    assign layer4_out[4792] = layer3_out[6064];
    assign layer4_out[4793] = layer3_out[1940];
    assign layer4_out[4794] = layer3_out[1947] & ~layer3_out[1948];
    assign layer4_out[4795] = layer3_out[1578] & layer3_out[1579];
    assign layer4_out[4796] = layer3_out[3890];
    assign layer4_out[4797] = layer3_out[3997] ^ layer3_out[3998];
    assign layer4_out[4798] = ~(layer3_out[5223] ^ layer3_out[5224]);
    assign layer4_out[4799] = layer3_out[6862];
    assign layer4_out[4800] = ~layer3_out[4007] | layer3_out[4008];
    assign layer4_out[4801] = ~layer3_out[5723];
    assign layer4_out[4802] = layer3_out[4969];
    assign layer4_out[4803] = ~layer3_out[3677];
    assign layer4_out[4804] = ~layer3_out[7406] | layer3_out[7407];
    assign layer4_out[4805] = layer3_out[1112] ^ layer3_out[1113];
    assign layer4_out[4806] = ~(layer3_out[2656] | layer3_out[2657]);
    assign layer4_out[4807] = layer3_out[1437];
    assign layer4_out[4808] = ~layer3_out[5137] | layer3_out[5136];
    assign layer4_out[4809] = ~layer3_out[740];
    assign layer4_out[4810] = ~layer3_out[7842];
    assign layer4_out[4811] = layer3_out[3312];
    assign layer4_out[4812] = layer3_out[4682] & layer3_out[4683];
    assign layer4_out[4813] = ~layer3_out[6202];
    assign layer4_out[4814] = ~layer3_out[764] | layer3_out[763];
    assign layer4_out[4815] = ~(layer3_out[3935] ^ layer3_out[3936]);
    assign layer4_out[4816] = ~layer3_out[1239];
    assign layer4_out[4817] = ~layer3_out[6306];
    assign layer4_out[4818] = ~(layer3_out[1183] | layer3_out[1184]);
    assign layer4_out[4819] = layer3_out[2421] & layer3_out[2422];
    assign layer4_out[4820] = ~layer3_out[4998] | layer3_out[4997];
    assign layer4_out[4821] = ~(layer3_out[4649] ^ layer3_out[4650]);
    assign layer4_out[4822] = layer3_out[6273];
    assign layer4_out[4823] = layer3_out[1510] & layer3_out[1511];
    assign layer4_out[4824] = ~layer3_out[7220];
    assign layer4_out[4825] = ~layer3_out[2703];
    assign layer4_out[4826] = layer3_out[7715] & layer3_out[7716];
    assign layer4_out[4827] = layer3_out[7236];
    assign layer4_out[4828] = ~layer3_out[7155] | layer3_out[7154];
    assign layer4_out[4829] = ~layer3_out[3062] | layer3_out[3061];
    assign layer4_out[4830] = ~layer3_out[5787];
    assign layer4_out[4831] = layer3_out[3399];
    assign layer4_out[4832] = ~layer3_out[4797] | layer3_out[4798];
    assign layer4_out[4833] = layer3_out[4181];
    assign layer4_out[4834] = layer3_out[5260] & layer3_out[5261];
    assign layer4_out[4835] = ~layer3_out[452];
    assign layer4_out[4836] = layer3_out[1516] ^ layer3_out[1517];
    assign layer4_out[4837] = ~layer3_out[5373];
    assign layer4_out[4838] = ~layer3_out[230] | layer3_out[229];
    assign layer4_out[4839] = ~layer3_out[2992] | layer3_out[2991];
    assign layer4_out[4840] = ~layer3_out[7378] | layer3_out[7377];
    assign layer4_out[4841] = ~(layer3_out[618] | layer3_out[619]);
    assign layer4_out[4842] = layer3_out[2397];
    assign layer4_out[4843] = layer3_out[594] ^ layer3_out[595];
    assign layer4_out[4844] = ~layer3_out[5841];
    assign layer4_out[4845] = layer3_out[4186] ^ layer3_out[4187];
    assign layer4_out[4846] = ~layer3_out[4294];
    assign layer4_out[4847] = ~layer3_out[305];
    assign layer4_out[4848] = ~layer3_out[7958];
    assign layer4_out[4849] = layer3_out[6323] | layer3_out[6324];
    assign layer4_out[4850] = layer3_out[880] & layer3_out[881];
    assign layer4_out[4851] = ~(layer3_out[6035] | layer3_out[6036]);
    assign layer4_out[4852] = layer3_out[651] & ~layer3_out[650];
    assign layer4_out[4853] = 1'b1;
    assign layer4_out[4854] = layer3_out[3401] | layer3_out[3402];
    assign layer4_out[4855] = ~layer3_out[7790];
    assign layer4_out[4856] = ~layer3_out[29] | layer3_out[28];
    assign layer4_out[4857] = ~(layer3_out[571] ^ layer3_out[572]);
    assign layer4_out[4858] = ~(layer3_out[65] | layer3_out[66]);
    assign layer4_out[4859] = layer3_out[2802] & layer3_out[2803];
    assign layer4_out[4860] = ~layer3_out[820] | layer3_out[821];
    assign layer4_out[4861] = ~layer3_out[5819];
    assign layer4_out[4862] = layer3_out[5479];
    assign layer4_out[4863] = layer3_out[3993];
    assign layer4_out[4864] = layer3_out[4193];
    assign layer4_out[4865] = layer3_out[4660];
    assign layer4_out[4866] = ~layer3_out[4235] | layer3_out[4236];
    assign layer4_out[4867] = ~(layer3_out[970] & layer3_out[971]);
    assign layer4_out[4868] = layer3_out[1682];
    assign layer4_out[4869] = ~layer3_out[7079];
    assign layer4_out[4870] = ~layer3_out[6173] | layer3_out[6174];
    assign layer4_out[4871] = ~layer3_out[1921] | layer3_out[1922];
    assign layer4_out[4872] = layer3_out[4231];
    assign layer4_out[4873] = ~layer3_out[2318] | layer3_out[2319];
    assign layer4_out[4874] = layer3_out[6153] | layer3_out[6154];
    assign layer4_out[4875] = ~layer3_out[6914] | layer3_out[6915];
    assign layer4_out[4876] = ~(layer3_out[3046] | layer3_out[3047]);
    assign layer4_out[4877] = ~(layer3_out[5138] ^ layer3_out[5139]);
    assign layer4_out[4878] = ~layer3_out[5868];
    assign layer4_out[4879] = ~(layer3_out[6206] ^ layer3_out[6207]);
    assign layer4_out[4880] = layer3_out[1979];
    assign layer4_out[4881] = layer3_out[4151];
    assign layer4_out[4882] = layer3_out[5003] & ~layer3_out[5004];
    assign layer4_out[4883] = ~layer3_out[2967];
    assign layer4_out[4884] = layer3_out[3305] | layer3_out[3306];
    assign layer4_out[4885] = ~layer3_out[6857];
    assign layer4_out[4886] = ~(layer3_out[2571] | layer3_out[2572]);
    assign layer4_out[4887] = ~layer3_out[7248] | layer3_out[7249];
    assign layer4_out[4888] = layer3_out[4946] ^ layer3_out[4947];
    assign layer4_out[4889] = ~(layer3_out[6846] ^ layer3_out[6847]);
    assign layer4_out[4890] = ~layer3_out[1840] | layer3_out[1841];
    assign layer4_out[4891] = ~layer3_out[7697] | layer3_out[7696];
    assign layer4_out[4892] = layer3_out[4218];
    assign layer4_out[4893] = layer3_out[6529];
    assign layer4_out[4894] = ~layer3_out[6533] | layer3_out[6532];
    assign layer4_out[4895] = ~layer3_out[7898] | layer3_out[7897];
    assign layer4_out[4896] = layer3_out[4256] & ~layer3_out[4255];
    assign layer4_out[4897] = layer3_out[6488] ^ layer3_out[6489];
    assign layer4_out[4898] = layer3_out[7665] ^ layer3_out[7666];
    assign layer4_out[4899] = 1'b0;
    assign layer4_out[4900] = layer3_out[5826] & ~layer3_out[5827];
    assign layer4_out[4901] = layer3_out[5233] & ~layer3_out[5232];
    assign layer4_out[4902] = layer3_out[5050] & ~layer3_out[5051];
    assign layer4_out[4903] = ~layer3_out[2652];
    assign layer4_out[4904] = layer3_out[6384] ^ layer3_out[6385];
    assign layer4_out[4905] = layer3_out[5] & layer3_out[6];
    assign layer4_out[4906] = layer3_out[5436] & ~layer3_out[5435];
    assign layer4_out[4907] = layer3_out[550];
    assign layer4_out[4908] = layer3_out[247] | layer3_out[248];
    assign layer4_out[4909] = layer3_out[5088] & ~layer3_out[5087];
    assign layer4_out[4910] = layer3_out[5296] & ~layer3_out[5295];
    assign layer4_out[4911] = ~(layer3_out[5477] ^ layer3_out[5478]);
    assign layer4_out[4912] = layer3_out[1319];
    assign layer4_out[4913] = ~layer3_out[7071];
    assign layer4_out[4914] = ~(layer3_out[347] ^ layer3_out[348]);
    assign layer4_out[4915] = ~layer3_out[5216];
    assign layer4_out[4916] = layer3_out[2511] ^ layer3_out[2512];
    assign layer4_out[4917] = layer3_out[3891] ^ layer3_out[3892];
    assign layer4_out[4918] = ~layer3_out[856] | layer3_out[857];
    assign layer4_out[4919] = layer3_out[538] & layer3_out[539];
    assign layer4_out[4920] = ~layer3_out[4291];
    assign layer4_out[4921] = ~(layer3_out[1694] | layer3_out[1695]);
    assign layer4_out[4922] = ~(layer3_out[2113] & layer3_out[2114]);
    assign layer4_out[4923] = ~layer3_out[1417];
    assign layer4_out[4924] = layer3_out[3277] & ~layer3_out[3278];
    assign layer4_out[4925] = layer3_out[495];
    assign layer4_out[4926] = layer3_out[6467];
    assign layer4_out[4927] = ~(layer3_out[493] ^ layer3_out[494]);
    assign layer4_out[4928] = ~layer3_out[7337] | layer3_out[7338];
    assign layer4_out[4929] = layer3_out[6555];
    assign layer4_out[4930] = ~(layer3_out[7144] & layer3_out[7145]);
    assign layer4_out[4931] = ~layer3_out[5200];
    assign layer4_out[4932] = layer3_out[5369];
    assign layer4_out[4933] = layer3_out[2546] & ~layer3_out[2547];
    assign layer4_out[4934] = layer3_out[926] ^ layer3_out[927];
    assign layer4_out[4935] = layer3_out[3538] & layer3_out[3539];
    assign layer4_out[4936] = layer3_out[139] | layer3_out[140];
    assign layer4_out[4937] = ~layer3_out[1307];
    assign layer4_out[4938] = ~layer3_out[3644];
    assign layer4_out[4939] = ~layer3_out[1377];
    assign layer4_out[4940] = ~(layer3_out[7503] ^ layer3_out[7504]);
    assign layer4_out[4941] = ~(layer3_out[7642] & layer3_out[7643]);
    assign layer4_out[4942] = layer3_out[6441] | layer3_out[6442];
    assign layer4_out[4943] = layer3_out[6303];
    assign layer4_out[4944] = ~layer3_out[2194];
    assign layer4_out[4945] = ~layer3_out[7033];
    assign layer4_out[4946] = ~layer3_out[973];
    assign layer4_out[4947] = ~(layer3_out[6197] | layer3_out[6198]);
    assign layer4_out[4948] = layer3_out[3358];
    assign layer4_out[4949] = layer3_out[592] ^ layer3_out[593];
    assign layer4_out[4950] = layer3_out[4829];
    assign layer4_out[4951] = ~(layer3_out[4925] | layer3_out[4926]);
    assign layer4_out[4952] = layer3_out[2682];
    assign layer4_out[4953] = ~(layer3_out[2246] | layer3_out[2247]);
    assign layer4_out[4954] = ~(layer3_out[3514] & layer3_out[3515]);
    assign layer4_out[4955] = layer3_out[7494];
    assign layer4_out[4956] = layer3_out[2257] | layer3_out[2258];
    assign layer4_out[4957] = layer3_out[2201] & ~layer3_out[2202];
    assign layer4_out[4958] = ~(layer3_out[5645] ^ layer3_out[5646]);
    assign layer4_out[4959] = ~(layer3_out[4115] | layer3_out[4116]);
    assign layer4_out[4960] = layer3_out[7893] & layer3_out[7894];
    assign layer4_out[4961] = ~layer3_out[6841] | layer3_out[6840];
    assign layer4_out[4962] = layer3_out[1040];
    assign layer4_out[4963] = layer3_out[1298] ^ layer3_out[1299];
    assign layer4_out[4964] = ~(layer3_out[4390] ^ layer3_out[4391]);
    assign layer4_out[4965] = layer3_out[5476] & ~layer3_out[5477];
    assign layer4_out[4966] = ~(layer3_out[6403] ^ layer3_out[6404]);
    assign layer4_out[4967] = layer3_out[408] | layer3_out[409];
    assign layer4_out[4968] = 1'b1;
    assign layer4_out[4969] = layer3_out[3307] ^ layer3_out[3308];
    assign layer4_out[4970] = layer3_out[1643];
    assign layer4_out[4971] = ~layer3_out[6814] | layer3_out[6815];
    assign layer4_out[4972] = ~layer3_out[2321] | layer3_out[2320];
    assign layer4_out[4973] = ~(layer3_out[4030] & layer3_out[4031]);
    assign layer4_out[4974] = layer3_out[7621];
    assign layer4_out[4975] = layer3_out[5900];
    assign layer4_out[4976] = ~layer3_out[1043] | layer3_out[1044];
    assign layer4_out[4977] = layer3_out[4195] | layer3_out[4196];
    assign layer4_out[4978] = ~layer3_out[7045];
    assign layer4_out[4979] = ~(layer3_out[7990] ^ layer3_out[7991]);
    assign layer4_out[4980] = ~layer3_out[1930];
    assign layer4_out[4981] = ~layer3_out[343] | layer3_out[344];
    assign layer4_out[4982] = ~layer3_out[5234];
    assign layer4_out[4983] = ~(layer3_out[799] ^ layer3_out[800]);
    assign layer4_out[4984] = layer3_out[1284] ^ layer3_out[1285];
    assign layer4_out[4985] = ~layer3_out[3106] | layer3_out[3107];
    assign layer4_out[4986] = ~(layer3_out[5088] ^ layer3_out[5089]);
    assign layer4_out[4987] = layer3_out[3243];
    assign layer4_out[4988] = layer3_out[2639] & layer3_out[2640];
    assign layer4_out[4989] = ~(layer3_out[1086] ^ layer3_out[1087]);
    assign layer4_out[4990] = layer3_out[7971];
    assign layer4_out[4991] = layer3_out[4684] & layer3_out[4685];
    assign layer4_out[4992] = ~layer3_out[6961];
    assign layer4_out[4993] = ~layer3_out[3987];
    assign layer4_out[4994] = layer3_out[4903] & ~layer3_out[4904];
    assign layer4_out[4995] = layer3_out[2556] & ~layer3_out[2555];
    assign layer4_out[4996] = layer3_out[109] ^ layer3_out[110];
    assign layer4_out[4997] = layer3_out[3608] ^ layer3_out[3609];
    assign layer4_out[4998] = layer3_out[6174];
    assign layer4_out[4999] = layer3_out[7373];
    assign layer4_out[5000] = layer3_out[5326];
    assign layer4_out[5001] = ~(layer3_out[5174] | layer3_out[5175]);
    assign layer4_out[5002] = layer3_out[6058] ^ layer3_out[6059];
    assign layer4_out[5003] = ~layer3_out[4156];
    assign layer4_out[5004] = ~(layer3_out[514] ^ layer3_out[515]);
    assign layer4_out[5005] = ~(layer3_out[4801] ^ layer3_out[4802]);
    assign layer4_out[5006] = layer3_out[3294] & ~layer3_out[3295];
    assign layer4_out[5007] = layer3_out[759];
    assign layer4_out[5008] = ~layer3_out[1810];
    assign layer4_out[5009] = ~layer3_out[6431];
    assign layer4_out[5010] = ~(layer3_out[4429] | layer3_out[4430]);
    assign layer4_out[5011] = ~layer3_out[5772] | layer3_out[5771];
    assign layer4_out[5012] = ~(layer3_out[5262] | layer3_out[5263]);
    assign layer4_out[5013] = ~(layer3_out[3349] & layer3_out[3350]);
    assign layer4_out[5014] = ~(layer3_out[1678] & layer3_out[1679]);
    assign layer4_out[5015] = layer3_out[1499];
    assign layer4_out[5016] = 1'b0;
    assign layer4_out[5017] = layer3_out[7362];
    assign layer4_out[5018] = layer3_out[7735];
    assign layer4_out[5019] = ~layer3_out[5527];
    assign layer4_out[5020] = ~layer3_out[2590];
    assign layer4_out[5021] = layer3_out[964];
    assign layer4_out[5022] = ~layer3_out[5228] | layer3_out[5227];
    assign layer4_out[5023] = ~(layer3_out[7983] | layer3_out[7984]);
    assign layer4_out[5024] = ~layer3_out[7372];
    assign layer4_out[5025] = ~(layer3_out[2595] & layer3_out[2596]);
    assign layer4_out[5026] = ~layer3_out[2854] | layer3_out[2853];
    assign layer4_out[5027] = ~layer3_out[3044];
    assign layer4_out[5028] = layer3_out[6886];
    assign layer4_out[5029] = layer3_out[5866] ^ layer3_out[5867];
    assign layer4_out[5030] = ~layer3_out[1368];
    assign layer4_out[5031] = ~(layer3_out[3682] | layer3_out[3683]);
    assign layer4_out[5032] = ~layer3_out[320];
    assign layer4_out[5033] = layer3_out[4669];
    assign layer4_out[5034] = layer3_out[3433] | layer3_out[3434];
    assign layer4_out[5035] = layer3_out[6919] | layer3_out[6920];
    assign layer4_out[5036] = layer3_out[6710];
    assign layer4_out[5037] = layer3_out[6045];
    assign layer4_out[5038] = ~layer3_out[7825] | layer3_out[7826];
    assign layer4_out[5039] = layer3_out[710] & ~layer3_out[711];
    assign layer4_out[5040] = ~layer3_out[7114] | layer3_out[7115];
    assign layer4_out[5041] = ~(layer3_out[5377] ^ layer3_out[5378]);
    assign layer4_out[5042] = layer3_out[1104];
    assign layer4_out[5043] = layer3_out[5345] | layer3_out[5346];
    assign layer4_out[5044] = ~layer3_out[6949];
    assign layer4_out[5045] = ~(layer3_out[1266] & layer3_out[1267]);
    assign layer4_out[5046] = ~layer3_out[5482];
    assign layer4_out[5047] = ~(layer3_out[7636] ^ layer3_out[7637]);
    assign layer4_out[5048] = 1'b1;
    assign layer4_out[5049] = ~(layer3_out[2387] & layer3_out[2388]);
    assign layer4_out[5050] = layer3_out[2810];
    assign layer4_out[5051] = layer3_out[2096] | layer3_out[2097];
    assign layer4_out[5052] = ~(layer3_out[733] ^ layer3_out[734]);
    assign layer4_out[5053] = ~(layer3_out[2836] | layer3_out[2837]);
    assign layer4_out[5054] = layer3_out[1930];
    assign layer4_out[5055] = layer3_out[4774];
    assign layer4_out[5056] = ~layer3_out[7452];
    assign layer4_out[5057] = ~layer3_out[1869] | layer3_out[1870];
    assign layer4_out[5058] = layer3_out[4674] ^ layer3_out[4675];
    assign layer4_out[5059] = layer3_out[1496];
    assign layer4_out[5060] = ~layer3_out[6213] | layer3_out[6212];
    assign layer4_out[5061] = ~(layer3_out[1420] ^ layer3_out[1421]);
    assign layer4_out[5062] = ~layer3_out[3844];
    assign layer4_out[5063] = ~(layer3_out[4016] ^ layer3_out[4017]);
    assign layer4_out[5064] = layer3_out[1980] & layer3_out[1981];
    assign layer4_out[5065] = layer3_out[5562] & ~layer3_out[5561];
    assign layer4_out[5066] = ~layer3_out[6481];
    assign layer4_out[5067] = layer3_out[1370];
    assign layer4_out[5068] = ~(layer3_out[6896] ^ layer3_out[6897]);
    assign layer4_out[5069] = ~layer3_out[5060];
    assign layer4_out[5070] = ~(layer3_out[2119] ^ layer3_out[2120]);
    assign layer4_out[5071] = ~(layer3_out[7992] ^ layer3_out[7993]);
    assign layer4_out[5072] = ~(layer3_out[3272] ^ layer3_out[3273]);
    assign layer4_out[5073] = layer3_out[555];
    assign layer4_out[5074] = layer3_out[1524] & ~layer3_out[1525];
    assign layer4_out[5075] = ~(layer3_out[4296] & layer3_out[4297]);
    assign layer4_out[5076] = layer3_out[5098] & ~layer3_out[5097];
    assign layer4_out[5077] = layer3_out[3299];
    assign layer4_out[5078] = layer3_out[5839];
    assign layer4_out[5079] = layer3_out[6319];
    assign layer4_out[5080] = layer3_out[7283] & layer3_out[7284];
    assign layer4_out[5081] = ~(layer3_out[3079] | layer3_out[3080]);
    assign layer4_out[5082] = ~layer3_out[395];
    assign layer4_out[5083] = layer3_out[1871] | layer3_out[1872];
    assign layer4_out[5084] = ~(layer3_out[5788] ^ layer3_out[5789]);
    assign layer4_out[5085] = layer3_out[6096] & layer3_out[6097];
    assign layer4_out[5086] = ~layer3_out[6237];
    assign layer4_out[5087] = layer3_out[3452] & ~layer3_out[3453];
    assign layer4_out[5088] = layer3_out[7392] & ~layer3_out[7393];
    assign layer4_out[5089] = ~(layer3_out[2541] ^ layer3_out[2542]);
    assign layer4_out[5090] = layer3_out[1572] & ~layer3_out[1573];
    assign layer4_out[5091] = 1'b1;
    assign layer4_out[5092] = ~layer3_out[536];
    assign layer4_out[5093] = layer3_out[1659];
    assign layer4_out[5094] = layer3_out[4620] & layer3_out[4621];
    assign layer4_out[5095] = ~layer3_out[667];
    assign layer4_out[5096] = ~layer3_out[1596] | layer3_out[1595];
    assign layer4_out[5097] = layer3_out[6586] | layer3_out[6587];
    assign layer4_out[5098] = layer3_out[7345];
    assign layer4_out[5099] = layer3_out[1010] | layer3_out[1011];
    assign layer4_out[5100] = ~layer3_out[5890] | layer3_out[5891];
    assign layer4_out[5101] = layer3_out[27] & ~layer3_out[28];
    assign layer4_out[5102] = layer3_out[48] & ~layer3_out[47];
    assign layer4_out[5103] = layer3_out[196] ^ layer3_out[197];
    assign layer4_out[5104] = layer3_out[525];
    assign layer4_out[5105] = layer3_out[2574] ^ layer3_out[2575];
    assign layer4_out[5106] = layer3_out[6051];
    assign layer4_out[5107] = ~(layer3_out[3136] | layer3_out[3137]);
    assign layer4_out[5108] = ~(layer3_out[5565] & layer3_out[5566]);
    assign layer4_out[5109] = ~(layer3_out[6007] ^ layer3_out[6008]);
    assign layer4_out[5110] = ~(layer3_out[669] ^ layer3_out[670]);
    assign layer4_out[5111] = layer3_out[7930];
    assign layer4_out[5112] = layer3_out[3575];
    assign layer4_out[5113] = ~(layer3_out[4449] | layer3_out[4450]);
    assign layer4_out[5114] = ~layer3_out[5215];
    assign layer4_out[5115] = layer3_out[5761] ^ layer3_out[5762];
    assign layer4_out[5116] = layer3_out[1107];
    assign layer4_out[5117] = ~layer3_out[1912];
    assign layer4_out[5118] = ~(layer3_out[1182] & layer3_out[1183]);
    assign layer4_out[5119] = ~layer3_out[1480] | layer3_out[1479];
    assign layer4_out[5120] = layer3_out[798];
    assign layer4_out[5121] = layer3_out[6099];
    assign layer4_out[5122] = layer3_out[5451] | layer3_out[5452];
    assign layer4_out[5123] = layer3_out[4770] & ~layer3_out[4769];
    assign layer4_out[5124] = layer3_out[4130] & layer3_out[4131];
    assign layer4_out[5125] = ~(layer3_out[233] ^ layer3_out[234]);
    assign layer4_out[5126] = ~layer3_out[4617] | layer3_out[4618];
    assign layer4_out[5127] = ~layer3_out[2094];
    assign layer4_out[5128] = ~(layer3_out[2539] ^ layer3_out[2540]);
    assign layer4_out[5129] = ~layer3_out[3217];
    assign layer4_out[5130] = layer3_out[3469];
    assign layer4_out[5131] = ~(layer3_out[7496] & layer3_out[7497]);
    assign layer4_out[5132] = ~layer3_out[559];
    assign layer4_out[5133] = layer3_out[3895] & ~layer3_out[3894];
    assign layer4_out[5134] = layer3_out[2768] & layer3_out[2769];
    assign layer4_out[5135] = ~(layer3_out[1098] | layer3_out[1099]);
    assign layer4_out[5136] = layer3_out[3780] ^ layer3_out[3781];
    assign layer4_out[5137] = layer3_out[3841] & layer3_out[3842];
    assign layer4_out[5138] = layer3_out[5994] & ~layer3_out[5993];
    assign layer4_out[5139] = layer3_out[6300];
    assign layer4_out[5140] = ~(layer3_out[2661] ^ layer3_out[2662]);
    assign layer4_out[5141] = layer3_out[4899] & ~layer3_out[4900];
    assign layer4_out[5142] = ~layer3_out[6494];
    assign layer4_out[5143] = layer3_out[5852];
    assign layer4_out[5144] = layer3_out[657] ^ layer3_out[658];
    assign layer4_out[5145] = layer3_out[233] & ~layer3_out[232];
    assign layer4_out[5146] = layer3_out[6019] & ~layer3_out[6018];
    assign layer4_out[5147] = layer3_out[4552];
    assign layer4_out[5148] = ~layer3_out[2204];
    assign layer4_out[5149] = layer3_out[7279];
    assign layer4_out[5150] = layer3_out[5682] ^ layer3_out[5683];
    assign layer4_out[5151] = layer3_out[1955];
    assign layer4_out[5152] = layer3_out[3738];
    assign layer4_out[5153] = layer3_out[4569] ^ layer3_out[4570];
    assign layer4_out[5154] = ~layer3_out[1647] | layer3_out[1646];
    assign layer4_out[5155] = layer3_out[0] & layer3_out[1];
    assign layer4_out[5156] = layer3_out[6657] & ~layer3_out[6658];
    assign layer4_out[5157] = ~layer3_out[2011];
    assign layer4_out[5158] = ~layer3_out[5589];
    assign layer4_out[5159] = layer3_out[4760] ^ layer3_out[4761];
    assign layer4_out[5160] = ~layer3_out[2469] | layer3_out[2468];
    assign layer4_out[5161] = ~layer3_out[2691];
    assign layer4_out[5162] = layer3_out[1754];
    assign layer4_out[5163] = ~(layer3_out[1944] ^ layer3_out[1945]);
    assign layer4_out[5164] = layer3_out[2256] & ~layer3_out[2257];
    assign layer4_out[5165] = ~layer3_out[5276] | layer3_out[5275];
    assign layer4_out[5166] = ~layer3_out[5499] | layer3_out[5498];
    assign layer4_out[5167] = ~layer3_out[5790];
    assign layer4_out[5168] = ~(layer3_out[5775] & layer3_out[5776]);
    assign layer4_out[5169] = ~layer3_out[5401] | layer3_out[5402];
    assign layer4_out[5170] = ~(layer3_out[3213] & layer3_out[3214]);
    assign layer4_out[5171] = ~layer3_out[7363] | layer3_out[7364];
    assign layer4_out[5172] = ~(layer3_out[4954] | layer3_out[4955]);
    assign layer4_out[5173] = ~layer3_out[3684] | layer3_out[3683];
    assign layer4_out[5174] = ~layer3_out[2537] | layer3_out[2538];
    assign layer4_out[5175] = ~(layer3_out[6011] ^ layer3_out[6012]);
    assign layer4_out[5176] = ~layer3_out[4943];
    assign layer4_out[5177] = ~layer3_out[6503];
    assign layer4_out[5178] = layer3_out[7954] ^ layer3_out[7955];
    assign layer4_out[5179] = ~layer3_out[5143] | layer3_out[5142];
    assign layer4_out[5180] = ~(layer3_out[2444] ^ layer3_out[2445]);
    assign layer4_out[5181] = layer3_out[3785];
    assign layer4_out[5182] = layer3_out[1562];
    assign layer4_out[5183] = layer3_out[7293];
    assign layer4_out[5184] = ~(layer3_out[7047] ^ layer3_out[7048]);
    assign layer4_out[5185] = layer3_out[2589] ^ layer3_out[2590];
    assign layer4_out[5186] = ~layer3_out[5394];
    assign layer4_out[5187] = ~layer3_out[2825] | layer3_out[2824];
    assign layer4_out[5188] = ~layer3_out[7892];
    assign layer4_out[5189] = layer3_out[7994] & layer3_out[7995];
    assign layer4_out[5190] = ~layer3_out[5147] | layer3_out[5146];
    assign layer4_out[5191] = ~(layer3_out[4781] & layer3_out[4782]);
    assign layer4_out[5192] = ~(layer3_out[6527] ^ layer3_out[6528]);
    assign layer4_out[5193] = layer3_out[3380] & ~layer3_out[3379];
    assign layer4_out[5194] = layer3_out[6258];
    assign layer4_out[5195] = layer3_out[1622];
    assign layer4_out[5196] = layer3_out[1391] & layer3_out[1392];
    assign layer4_out[5197] = ~layer3_out[7759] | layer3_out[7760];
    assign layer4_out[5198] = layer3_out[100];
    assign layer4_out[5199] = layer3_out[1039] & layer3_out[1040];
    assign layer4_out[5200] = layer3_out[4063] ^ layer3_out[4064];
    assign layer4_out[5201] = ~layer3_out[4577] | layer3_out[4578];
    assign layer4_out[5202] = ~layer3_out[7206];
    assign layer4_out[5203] = layer3_out[1758] & ~layer3_out[1757];
    assign layer4_out[5204] = ~layer3_out[4582];
    assign layer4_out[5205] = layer3_out[6437] & ~layer3_out[6436];
    assign layer4_out[5206] = ~layer3_out[6469];
    assign layer4_out[5207] = ~layer3_out[7132] | layer3_out[7131];
    assign layer4_out[5208] = ~layer3_out[3577] | layer3_out[3578];
    assign layer4_out[5209] = ~(layer3_out[3975] | layer3_out[3976]);
    assign layer4_out[5210] = layer3_out[1483] & ~layer3_out[1482];
    assign layer4_out[5211] = layer3_out[5792] & ~layer3_out[5793];
    assign layer4_out[5212] = layer3_out[7883] & ~layer3_out[7884];
    assign layer4_out[5213] = ~layer3_out[4321];
    assign layer4_out[5214] = ~layer3_out[4336];
    assign layer4_out[5215] = ~layer3_out[5197];
    assign layer4_out[5216] = layer3_out[2795] ^ layer3_out[2796];
    assign layer4_out[5217] = layer3_out[6683];
    assign layer4_out[5218] = ~layer3_out[6103];
    assign layer4_out[5219] = layer3_out[4758] & ~layer3_out[4759];
    assign layer4_out[5220] = layer3_out[1343];
    assign layer4_out[5221] = ~layer3_out[2286];
    assign layer4_out[5222] = layer3_out[5157] ^ layer3_out[5158];
    assign layer4_out[5223] = ~layer3_out[7250];
    assign layer4_out[5224] = layer3_out[5504];
    assign layer4_out[5225] = ~(layer3_out[3237] ^ layer3_out[3238]);
    assign layer4_out[5226] = layer3_out[475] | layer3_out[476];
    assign layer4_out[5227] = layer3_out[6537] & ~layer3_out[6538];
    assign layer4_out[5228] = ~layer3_out[1022] | layer3_out[1023];
    assign layer4_out[5229] = layer3_out[6579];
    assign layer4_out[5230] = ~layer3_out[2427];
    assign layer4_out[5231] = layer3_out[6393];
    assign layer4_out[5232] = ~layer3_out[2975];
    assign layer4_out[5233] = layer3_out[6850];
    assign layer4_out[5234] = layer3_out[4264];
    assign layer4_out[5235] = ~(layer3_out[299] & layer3_out[300]);
    assign layer4_out[5236] = layer3_out[5733] ^ layer3_out[5734];
    assign layer4_out[5237] = layer3_out[1842] & ~layer3_out[1841];
    assign layer4_out[5238] = layer3_out[3474] & ~layer3_out[3475];
    assign layer4_out[5239] = layer3_out[6421];
    assign layer4_out[5240] = layer3_out[7484] & layer3_out[7485];
    assign layer4_out[5241] = layer3_out[1334];
    assign layer4_out[5242] = ~layer3_out[6091] | layer3_out[6090];
    assign layer4_out[5243] = layer3_out[3045] & ~layer3_out[3046];
    assign layer4_out[5244] = layer3_out[5522];
    assign layer4_out[5245] = ~layer3_out[2346];
    assign layer4_out[5246] = layer3_out[4059] & layer3_out[4060];
    assign layer4_out[5247] = layer3_out[4840] ^ layer3_out[4841];
    assign layer4_out[5248] = layer3_out[2868] | layer3_out[2869];
    assign layer4_out[5249] = ~layer3_out[2304];
    assign layer4_out[5250] = ~layer3_out[590];
    assign layer4_out[5251] = layer3_out[6666] ^ layer3_out[6667];
    assign layer4_out[5252] = layer3_out[3511];
    assign layer4_out[5253] = layer3_out[237];
    assign layer4_out[5254] = layer3_out[5553];
    assign layer4_out[5255] = ~layer3_out[1294];
    assign layer4_out[5256] = layer3_out[4770] ^ layer3_out[4771];
    assign layer4_out[5257] = ~layer3_out[2252] | layer3_out[2251];
    assign layer4_out[5258] = layer3_out[439] & ~layer3_out[438];
    assign layer4_out[5259] = ~(layer3_out[3554] ^ layer3_out[3555]);
    assign layer4_out[5260] = layer3_out[1508] & layer3_out[1509];
    assign layer4_out[5261] = layer3_out[2452] ^ layer3_out[2453];
    assign layer4_out[5262] = ~(layer3_out[5482] & layer3_out[5483]);
    assign layer4_out[5263] = ~layer3_out[4365];
    assign layer4_out[5264] = layer3_out[7612];
    assign layer4_out[5265] = layer3_out[5358] & layer3_out[5359];
    assign layer4_out[5266] = layer3_out[4211] & layer3_out[4212];
    assign layer4_out[5267] = layer3_out[7424] & ~layer3_out[7425];
    assign layer4_out[5268] = ~layer3_out[4713] | layer3_out[4714];
    assign layer4_out[5269] = layer3_out[3136];
    assign layer4_out[5270] = ~layer3_out[530];
    assign layer4_out[5271] = layer3_out[3169];
    assign layer4_out[5272] = ~layer3_out[6628];
    assign layer4_out[5273] = ~layer3_out[6779];
    assign layer4_out[5274] = ~(layer3_out[3961] ^ layer3_out[3962]);
    assign layer4_out[5275] = ~layer3_out[282];
    assign layer4_out[5276] = ~layer3_out[7745] | layer3_out[7744];
    assign layer4_out[5277] = layer3_out[3332] & layer3_out[3333];
    assign layer4_out[5278] = ~layer3_out[7427] | layer3_out[7426];
    assign layer4_out[5279] = ~layer3_out[6875];
    assign layer4_out[5280] = layer3_out[7549];
    assign layer4_out[5281] = layer3_out[2175];
    assign layer4_out[5282] = layer3_out[1304] & ~layer3_out[1303];
    assign layer4_out[5283] = layer3_out[7786];
    assign layer4_out[5284] = ~layer3_out[6426] | layer3_out[6425];
    assign layer4_out[5285] = ~(layer3_out[541] & layer3_out[542]);
    assign layer4_out[5286] = layer3_out[7821] ^ layer3_out[7822];
    assign layer4_out[5287] = layer3_out[1169] & ~layer3_out[1170];
    assign layer4_out[5288] = ~(layer3_out[153] & layer3_out[154]);
    assign layer4_out[5289] = ~layer3_out[1712];
    assign layer4_out[5290] = ~layer3_out[7254] | layer3_out[7255];
    assign layer4_out[5291] = layer3_out[6740];
    assign layer4_out[5292] = ~(layer3_out[3155] | layer3_out[3156]);
    assign layer4_out[5293] = 1'b1;
    assign layer4_out[5294] = ~layer3_out[4949];
    assign layer4_out[5295] = ~layer3_out[4383];
    assign layer4_out[5296] = layer3_out[1475];
    assign layer4_out[5297] = 1'b0;
    assign layer4_out[5298] = ~layer3_out[354] | layer3_out[355];
    assign layer4_out[5299] = ~layer3_out[6347];
    assign layer4_out[5300] = layer3_out[7324] ^ layer3_out[7325];
    assign layer4_out[5301] = 1'b1;
    assign layer4_out[5302] = layer3_out[3342] & layer3_out[3343];
    assign layer4_out[5303] = layer3_out[5670];
    assign layer4_out[5304] = ~(layer3_out[3933] ^ layer3_out[3934]);
    assign layer4_out[5305] = layer3_out[122] ^ layer3_out[123];
    assign layer4_out[5306] = layer3_out[2036];
    assign layer4_out[5307] = ~(layer3_out[6028] & layer3_out[6029]);
    assign layer4_out[5308] = layer3_out[2531];
    assign layer4_out[5309] = layer3_out[4408];
    assign layer4_out[5310] = ~layer3_out[4931];
    assign layer4_out[5311] = ~(layer3_out[4494] & layer3_out[4495]);
    assign layer4_out[5312] = layer3_out[3553] ^ layer3_out[3554];
    assign layer4_out[5313] = ~layer3_out[810];
    assign layer4_out[5314] = layer3_out[1362] ^ layer3_out[1363];
    assign layer4_out[5315] = ~layer3_out[2891] | layer3_out[2892];
    assign layer4_out[5316] = layer3_out[5760];
    assign layer4_out[5317] = layer3_out[779] & layer3_out[780];
    assign layer4_out[5318] = layer3_out[4074];
    assign layer4_out[5319] = ~layer3_out[6763];
    assign layer4_out[5320] = layer3_out[3279] | layer3_out[3280];
    assign layer4_out[5321] = layer3_out[672];
    assign layer4_out[5322] = ~layer3_out[5404];
    assign layer4_out[5323] = ~(layer3_out[3293] ^ layer3_out[3294]);
    assign layer4_out[5324] = ~layer3_out[7955];
    assign layer4_out[5325] = ~layer3_out[1340];
    assign layer4_out[5326] = ~layer3_out[5592] | layer3_out[5593];
    assign layer4_out[5327] = layer3_out[3735];
    assign layer4_out[5328] = layer3_out[6600];
    assign layer4_out[5329] = ~layer3_out[754];
    assign layer4_out[5330] = layer3_out[6727];
    assign layer4_out[5331] = ~layer3_out[1732];
    assign layer4_out[5332] = layer3_out[7099] ^ layer3_out[7100];
    assign layer4_out[5333] = ~layer3_out[4271];
    assign layer4_out[5334] = layer3_out[3802] & ~layer3_out[3803];
    assign layer4_out[5335] = layer3_out[923];
    assign layer4_out[5336] = ~layer3_out[1500];
    assign layer4_out[5337] = layer3_out[4366] | layer3_out[4367];
    assign layer4_out[5338] = ~layer3_out[7583];
    assign layer4_out[5339] = ~layer3_out[2897];
    assign layer4_out[5340] = ~(layer3_out[5324] & layer3_out[5325]);
    assign layer4_out[5341] = ~(layer3_out[1235] | layer3_out[1236]);
    assign layer4_out[5342] = ~layer3_out[1832];
    assign layer4_out[5343] = ~(layer3_out[5428] | layer3_out[5429]);
    assign layer4_out[5344] = ~layer3_out[1345] | layer3_out[1346];
    assign layer4_out[5345] = ~(layer3_out[7789] | layer3_out[7790]);
    assign layer4_out[5346] = ~layer3_out[1550];
    assign layer4_out[5347] = ~(layer3_out[1087] & layer3_out[1088]);
    assign layer4_out[5348] = layer3_out[7731];
    assign layer4_out[5349] = ~(layer3_out[5068] ^ layer3_out[5069]);
    assign layer4_out[5350] = layer3_out[5587] & layer3_out[5588];
    assign layer4_out[5351] = layer3_out[7947] ^ layer3_out[7948];
    assign layer4_out[5352] = ~layer3_out[1215];
    assign layer4_out[5353] = ~layer3_out[1094];
    assign layer4_out[5354] = ~layer3_out[4024] | layer3_out[4023];
    assign layer4_out[5355] = ~(layer3_out[7086] ^ layer3_out[7087]);
    assign layer4_out[5356] = ~(layer3_out[98] & layer3_out[99]);
    assign layer4_out[5357] = ~layer3_out[2000] | layer3_out[2001];
    assign layer4_out[5358] = layer3_out[4421] & ~layer3_out[4422];
    assign layer4_out[5359] = layer3_out[907] ^ layer3_out[908];
    assign layer4_out[5360] = ~layer3_out[7168] | layer3_out[7167];
    assign layer4_out[5361] = layer3_out[2166] ^ layer3_out[2167];
    assign layer4_out[5362] = layer3_out[7048] | layer3_out[7049];
    assign layer4_out[5363] = ~(layer3_out[3926] ^ layer3_out[3927]);
    assign layer4_out[5364] = layer3_out[5466];
    assign layer4_out[5365] = layer3_out[7665] & ~layer3_out[7664];
    assign layer4_out[5366] = layer3_out[6199] & ~layer3_out[6198];
    assign layer4_out[5367] = ~layer3_out[5685];
    assign layer4_out[5368] = ~layer3_out[1613];
    assign layer4_out[5369] = ~(layer3_out[2362] ^ layer3_out[2363]);
    assign layer4_out[5370] = ~layer3_out[2358];
    assign layer4_out[5371] = layer3_out[7835];
    assign layer4_out[5372] = ~(layer3_out[6598] ^ layer3_out[6599]);
    assign layer4_out[5373] = ~layer3_out[5279];
    assign layer4_out[5374] = 1'b1;
    assign layer4_out[5375] = layer3_out[7987] ^ layer3_out[7988];
    assign layer4_out[5376] = layer3_out[4644] & ~layer3_out[4643];
    assign layer4_out[5377] = layer3_out[331];
    assign layer4_out[5378] = ~layer3_out[1676];
    assign layer4_out[5379] = layer3_out[1879] ^ layer3_out[1880];
    assign layer4_out[5380] = ~layer3_out[3622];
    assign layer4_out[5381] = ~(layer3_out[5238] ^ layer3_out[5239]);
    assign layer4_out[5382] = layer3_out[1614] & ~layer3_out[1615];
    assign layer4_out[5383] = ~layer3_out[5610];
    assign layer4_out[5384] = ~(layer3_out[1564] & layer3_out[1565]);
    assign layer4_out[5385] = layer3_out[1473] & ~layer3_out[1474];
    assign layer4_out[5386] = layer3_out[2694];
    assign layer4_out[5387] = layer3_out[4325] | layer3_out[4326];
    assign layer4_out[5388] = ~layer3_out[194] | layer3_out[193];
    assign layer4_out[5389] = ~(layer3_out[7393] & layer3_out[7394]);
    assign layer4_out[5390] = layer3_out[4187] & layer3_out[4188];
    assign layer4_out[5391] = layer3_out[7426] & ~layer3_out[7425];
    assign layer4_out[5392] = layer3_out[3801] & ~layer3_out[3802];
    assign layer4_out[5393] = ~layer3_out[6019];
    assign layer4_out[5394] = layer3_out[1062] | layer3_out[1063];
    assign layer4_out[5395] = layer3_out[307] & ~layer3_out[306];
    assign layer4_out[5396] = layer3_out[4555] & ~layer3_out[4556];
    assign layer4_out[5397] = layer3_out[6601] & ~layer3_out[6600];
    assign layer4_out[5398] = layer3_out[4842] & layer3_out[4843];
    assign layer4_out[5399] = ~layer3_out[7527];
    assign layer4_out[5400] = ~layer3_out[3488] | layer3_out[3487];
    assign layer4_out[5401] = layer3_out[5820] & layer3_out[5821];
    assign layer4_out[5402] = layer3_out[1198] ^ layer3_out[1199];
    assign layer4_out[5403] = ~layer3_out[3631] | layer3_out[3630];
    assign layer4_out[5404] = ~(layer3_out[4703] & layer3_out[4704]);
    assign layer4_out[5405] = layer3_out[4696];
    assign layer4_out[5406] = ~layer3_out[7234];
    assign layer4_out[5407] = layer3_out[6150] & layer3_out[6151];
    assign layer4_out[5408] = layer3_out[6548];
    assign layer4_out[5409] = ~(layer3_out[3534] & layer3_out[3535]);
    assign layer4_out[5410] = layer3_out[3146] & layer3_out[3147];
    assign layer4_out[5411] = ~(layer3_out[1702] ^ layer3_out[1703]);
    assign layer4_out[5412] = ~layer3_out[3157];
    assign layer4_out[5413] = ~(layer3_out[6619] | layer3_out[6620]);
    assign layer4_out[5414] = layer3_out[5035];
    assign layer4_out[5415] = layer3_out[4129];
    assign layer4_out[5416] = layer3_out[4976];
    assign layer4_out[5417] = ~(layer3_out[3269] & layer3_out[3270]);
    assign layer4_out[5418] = ~(layer3_out[4702] ^ layer3_out[4703]);
    assign layer4_out[5419] = layer3_out[4346] | layer3_out[4347];
    assign layer4_out[5420] = ~(layer3_out[4111] ^ layer3_out[4112]);
    assign layer4_out[5421] = layer3_out[6447] | layer3_out[6448];
    assign layer4_out[5422] = ~layer3_out[1445] | layer3_out[1444];
    assign layer4_out[5423] = ~layer3_out[5170];
    assign layer4_out[5424] = ~(layer3_out[5509] & layer3_out[5510]);
    assign layer4_out[5425] = layer3_out[3500];
    assign layer4_out[5426] = layer3_out[3397];
    assign layer4_out[5427] = ~(layer3_out[524] ^ layer3_out[525]);
    assign layer4_out[5428] = ~layer3_out[5078] | layer3_out[5077];
    assign layer4_out[5429] = ~(layer3_out[3709] ^ layer3_out[3710]);
    assign layer4_out[5430] = layer3_out[713];
    assign layer4_out[5431] = ~layer3_out[4640] | layer3_out[4639];
    assign layer4_out[5432] = ~layer3_out[7225];
    assign layer4_out[5433] = ~(layer3_out[6015] | layer3_out[6016]);
    assign layer4_out[5434] = ~layer3_out[5810];
    assign layer4_out[5435] = ~(layer3_out[7680] ^ layer3_out[7681]);
    assign layer4_out[5436] = 1'b1;
    assign layer4_out[5437] = ~layer3_out[3205];
    assign layer4_out[5438] = layer3_out[1723] | layer3_out[1724];
    assign layer4_out[5439] = ~layer3_out[1398];
    assign layer4_out[5440] = layer3_out[6604];
    assign layer4_out[5441] = ~layer3_out[4830];
    assign layer4_out[5442] = ~(layer3_out[6224] & layer3_out[6225]);
    assign layer4_out[5443] = layer3_out[3443] & ~layer3_out[3444];
    assign layer4_out[5444] = layer3_out[178] ^ layer3_out[179];
    assign layer4_out[5445] = ~(layer3_out[7812] | layer3_out[7813]);
    assign layer4_out[5446] = layer3_out[2990] ^ layer3_out[2991];
    assign layer4_out[5447] = ~layer3_out[830];
    assign layer4_out[5448] = layer3_out[943];
    assign layer4_out[5449] = layer3_out[7135];
    assign layer4_out[5450] = layer3_out[3448];
    assign layer4_out[5451] = layer3_out[4226];
    assign layer4_out[5452] = layer3_out[2347];
    assign layer4_out[5453] = layer3_out[7139] & layer3_out[7140];
    assign layer4_out[5454] = layer3_out[6608] ^ layer3_out[6609];
    assign layer4_out[5455] = ~(layer3_out[5149] ^ layer3_out[5150]);
    assign layer4_out[5456] = ~layer3_out[2864] | layer3_out[2865];
    assign layer4_out[5457] = layer3_out[4592] & layer3_out[4593];
    assign layer4_out[5458] = layer3_out[3783] ^ layer3_out[3784];
    assign layer4_out[5459] = layer3_out[315] ^ layer3_out[316];
    assign layer4_out[5460] = ~layer3_out[3956] | layer3_out[3955];
    assign layer4_out[5461] = layer3_out[7067] & ~layer3_out[7068];
    assign layer4_out[5462] = ~(layer3_out[3502] ^ layer3_out[3503]);
    assign layer4_out[5463] = layer3_out[6576] & ~layer3_out[6575];
    assign layer4_out[5464] = ~layer3_out[3363];
    assign layer4_out[5465] = layer3_out[221] & layer3_out[222];
    assign layer4_out[5466] = layer3_out[1791];
    assign layer4_out[5467] = ~layer3_out[6501];
    assign layer4_out[5468] = ~layer3_out[1502];
    assign layer4_out[5469] = ~layer3_out[883];
    assign layer4_out[5470] = ~layer3_out[5018];
    assign layer4_out[5471] = ~layer3_out[4013] | layer3_out[4014];
    assign layer4_out[5472] = layer3_out[3452];
    assign layer4_out[5473] = layer3_out[4232] & ~layer3_out[4233];
    assign layer4_out[5474] = ~layer3_out[4427];
    assign layer4_out[5475] = layer3_out[4608] ^ layer3_out[4609];
    assign layer4_out[5476] = ~(layer3_out[7432] | layer3_out[7433]);
    assign layer4_out[5477] = ~(layer3_out[4463] & layer3_out[4464]);
    assign layer4_out[5478] = layer3_out[1813] | layer3_out[1814];
    assign layer4_out[5479] = layer3_out[7615] & ~layer3_out[7614];
    assign layer4_out[5480] = ~layer3_out[1137];
    assign layer4_out[5481] = layer3_out[664] ^ layer3_out[665];
    assign layer4_out[5482] = ~layer3_out[1557] | layer3_out[1558];
    assign layer4_out[5483] = layer3_out[643];
    assign layer4_out[5484] = layer3_out[7607];
    assign layer4_out[5485] = layer3_out[4897];
    assign layer4_out[5486] = ~layer3_out[5288];
    assign layer4_out[5487] = ~layer3_out[202];
    assign layer4_out[5488] = ~(layer3_out[551] ^ layer3_out[552]);
    assign layer4_out[5489] = ~layer3_out[1936] | layer3_out[1937];
    assign layer4_out[5490] = ~layer3_out[673];
    assign layer4_out[5491] = 1'b1;
    assign layer4_out[5492] = layer3_out[1581] ^ layer3_out[1582];
    assign layer4_out[5493] = layer3_out[3539] ^ layer3_out[3540];
    assign layer4_out[5494] = ~(layer3_out[340] ^ layer3_out[341]);
    assign layer4_out[5495] = ~(layer3_out[6063] ^ layer3_out[6064]);
    assign layer4_out[5496] = layer3_out[2918] & layer3_out[2919];
    assign layer4_out[5497] = layer3_out[719] ^ layer3_out[720];
    assign layer4_out[5498] = ~layer3_out[696];
    assign layer4_out[5499] = ~(layer3_out[4893] ^ layer3_out[4894]);
    assign layer4_out[5500] = ~layer3_out[4692];
    assign layer4_out[5501] = ~(layer3_out[1177] | layer3_out[1178]);
    assign layer4_out[5502] = ~(layer3_out[6416] | layer3_out[6417]);
    assign layer4_out[5503] = ~(layer3_out[7682] & layer3_out[7683]);
    assign layer4_out[5504] = layer3_out[1383];
    assign layer4_out[5505] = ~(layer3_out[5971] ^ layer3_out[5972]);
    assign layer4_out[5506] = layer3_out[4508] & ~layer3_out[4507];
    assign layer4_out[5507] = layer3_out[144];
    assign layer4_out[5508] = layer3_out[2804] ^ layer3_out[2805];
    assign layer4_out[5509] = ~layer3_out[3524];
    assign layer4_out[5510] = layer3_out[204] ^ layer3_out[205];
    assign layer4_out[5511] = ~(layer3_out[547] ^ layer3_out[548]);
    assign layer4_out[5512] = layer3_out[2185];
    assign layer4_out[5513] = ~layer3_out[740];
    assign layer4_out[5514] = layer3_out[828];
    assign layer4_out[5515] = ~layer3_out[4891];
    assign layer4_out[5516] = layer3_out[4786];
    assign layer4_out[5517] = ~layer3_out[4160] | layer3_out[4159];
    assign layer4_out[5518] = layer3_out[7012] & ~layer3_out[7013];
    assign layer4_out[5519] = layer3_out[6438];
    assign layer4_out[5520] = ~(layer3_out[3040] & layer3_out[3041]);
    assign layer4_out[5521] = layer3_out[4563] & ~layer3_out[4562];
    assign layer4_out[5522] = layer3_out[6237] & ~layer3_out[6238];
    assign layer4_out[5523] = ~layer3_out[195];
    assign layer4_out[5524] = layer3_out[390] | layer3_out[391];
    assign layer4_out[5525] = layer3_out[2391] & ~layer3_out[2390];
    assign layer4_out[5526] = ~(layer3_out[2672] ^ layer3_out[2673]);
    assign layer4_out[5527] = layer3_out[5217] ^ layer3_out[5218];
    assign layer4_out[5528] = layer3_out[3504];
    assign layer4_out[5529] = layer3_out[2082] & layer3_out[2083];
    assign layer4_out[5530] = ~(layer3_out[2844] & layer3_out[2845]);
    assign layer4_out[5531] = ~layer3_out[734];
    assign layer4_out[5532] = ~layer3_out[4941];
    assign layer4_out[5533] = ~(layer3_out[643] & layer3_out[644]);
    assign layer4_out[5534] = ~layer3_out[6532] | layer3_out[6531];
    assign layer4_out[5535] = ~layer3_out[4715] | layer3_out[4716];
    assign layer4_out[5536] = layer3_out[2235];
    assign layer4_out[5537] = layer3_out[4055] & ~layer3_out[4056];
    assign layer4_out[5538] = layer3_out[881];
    assign layer4_out[5539] = layer3_out[3400];
    assign layer4_out[5540] = ~layer3_out[3338];
    assign layer4_out[5541] = ~layer3_out[1206];
    assign layer4_out[5542] = layer3_out[1308] & layer3_out[1309];
    assign layer4_out[5543] = ~(layer3_out[597] & layer3_out[598]);
    assign layer4_out[5544] = ~(layer3_out[5309] & layer3_out[5310]);
    assign layer4_out[5545] = ~layer3_out[2227];
    assign layer4_out[5546] = ~layer3_out[6415];
    assign layer4_out[5547] = layer3_out[516];
    assign layer4_out[5548] = ~(layer3_out[5690] | layer3_out[5691]);
    assign layer4_out[5549] = layer3_out[1382] & ~layer3_out[1383];
    assign layer4_out[5550] = layer3_out[6971];
    assign layer4_out[5551] = layer3_out[3029];
    assign layer4_out[5552] = ~layer3_out[790];
    assign layer4_out[5553] = ~layer3_out[3214];
    assign layer4_out[5554] = ~(layer3_out[4107] ^ layer3_out[4108]);
    assign layer4_out[5555] = layer3_out[4189] & ~layer3_out[4190];
    assign layer4_out[5556] = layer3_out[4438];
    assign layer4_out[5557] = layer3_out[1649] & ~layer3_out[1650];
    assign layer4_out[5558] = layer3_out[1100] ^ layer3_out[1101];
    assign layer4_out[5559] = layer3_out[5895] & layer3_out[5896];
    assign layer4_out[5560] = layer3_out[5787];
    assign layer4_out[5561] = layer3_out[2380] & ~layer3_out[2379];
    assign layer4_out[5562] = ~layer3_out[2725];
    assign layer4_out[5563] = ~layer3_out[6384] | layer3_out[6383];
    assign layer4_out[5564] = ~layer3_out[1587] | layer3_out[1586];
    assign layer4_out[5565] = layer3_out[3631];
    assign layer4_out[5566] = layer3_out[5545] & ~layer3_out[5546];
    assign layer4_out[5567] = layer3_out[3748] & ~layer3_out[3747];
    assign layer4_out[5568] = ~layer3_out[7302];
    assign layer4_out[5569] = layer3_out[3817];
    assign layer4_out[5570] = ~(layer3_out[5717] ^ layer3_out[5718]);
    assign layer4_out[5571] = ~layer3_out[5570];
    assign layer4_out[5572] = layer3_out[1191] ^ layer3_out[1192];
    assign layer4_out[5573] = layer3_out[7559];
    assign layer4_out[5574] = layer3_out[1151];
    assign layer4_out[5575] = ~layer3_out[4733] | layer3_out[4734];
    assign layer4_out[5576] = ~(layer3_out[1740] ^ layer3_out[1741]);
    assign layer4_out[5577] = layer3_out[41];
    assign layer4_out[5578] = ~(layer3_out[2369] ^ layer3_out[2370]);
    assign layer4_out[5579] = ~layer3_out[1251] | layer3_out[1250];
    assign layer4_out[5580] = ~layer3_out[2443];
    assign layer4_out[5581] = layer3_out[6696] & layer3_out[6697];
    assign layer4_out[5582] = layer3_out[6022] & ~layer3_out[6021];
    assign layer4_out[5583] = layer3_out[4223] ^ layer3_out[4224];
    assign layer4_out[5584] = layer3_out[5257];
    assign layer4_out[5585] = layer3_out[7531];
    assign layer4_out[5586] = ~(layer3_out[7512] ^ layer3_out[7513]);
    assign layer4_out[5587] = layer3_out[4502] & layer3_out[4503];
    assign layer4_out[5588] = layer3_out[4762] ^ layer3_out[4763];
    assign layer4_out[5589] = layer3_out[2968];
    assign layer4_out[5590] = ~(layer3_out[2745] | layer3_out[2746]);
    assign layer4_out[5591] = ~layer3_out[6757];
    assign layer4_out[5592] = layer3_out[2613] & layer3_out[2614];
    assign layer4_out[5593] = ~(layer3_out[1718] | layer3_out[1719]);
    assign layer4_out[5594] = layer3_out[7655] | layer3_out[7656];
    assign layer4_out[5595] = layer3_out[5535] & ~layer3_out[5534];
    assign layer4_out[5596] = layer3_out[5678] & ~layer3_out[5679];
    assign layer4_out[5597] = layer3_out[692];
    assign layer4_out[5598] = ~layer3_out[3104];
    assign layer4_out[5599] = ~(layer3_out[3834] | layer3_out[3835]);
    assign layer4_out[5600] = ~layer3_out[6831];
    assign layer4_out[5601] = ~layer3_out[7473];
    assign layer4_out[5602] = layer3_out[3399] & ~layer3_out[3400];
    assign layer4_out[5603] = ~layer3_out[4183] | layer3_out[4182];
    assign layer4_out[5604] = ~(layer3_out[5907] ^ layer3_out[5908]);
    assign layer4_out[5605] = layer3_out[7654];
    assign layer4_out[5606] = ~layer3_out[7417];
    assign layer4_out[5607] = ~layer3_out[7678] | layer3_out[7677];
    assign layer4_out[5608] = ~(layer3_out[5348] ^ layer3_out[5349]);
    assign layer4_out[5609] = ~layer3_out[4271];
    assign layer4_out[5610] = ~(layer3_out[2957] ^ layer3_out[2958]);
    assign layer4_out[5611] = layer3_out[3351];
    assign layer4_out[5612] = layer3_out[2508] & ~layer3_out[2507];
    assign layer4_out[5613] = layer3_out[3300] ^ layer3_out[3301];
    assign layer4_out[5614] = ~layer3_out[1314];
    assign layer4_out[5615] = layer3_out[4479] & ~layer3_out[4478];
    assign layer4_out[5616] = ~(layer3_out[6613] ^ layer3_out[6614]);
    assign layer4_out[5617] = ~layer3_out[5354];
    assign layer4_out[5618] = ~(layer3_out[7465] ^ layer3_out[7466]);
    assign layer4_out[5619] = ~layer3_out[2063] | layer3_out[2062];
    assign layer4_out[5620] = layer3_out[3020];
    assign layer4_out[5621] = ~layer3_out[1550];
    assign layer4_out[5622] = layer3_out[7007] & ~layer3_out[7008];
    assign layer4_out[5623] = layer3_out[2118];
    assign layer4_out[5624] = ~layer3_out[5863] | layer3_out[5864];
    assign layer4_out[5625] = ~layer3_out[173] | layer3_out[172];
    assign layer4_out[5626] = ~layer3_out[3534];
    assign layer4_out[5627] = ~layer3_out[849] | layer3_out[848];
    assign layer4_out[5628] = ~(layer3_out[1767] | layer3_out[1768]);
    assign layer4_out[5629] = ~layer3_out[5035] | layer3_out[5034];
    assign layer4_out[5630] = ~(layer3_out[7814] & layer3_out[7815]);
    assign layer4_out[5631] = layer3_out[2887];
    assign layer4_out[5632] = ~(layer3_out[4499] & layer3_out[4500]);
    assign layer4_out[5633] = ~layer3_out[5439];
    assign layer4_out[5634] = layer3_out[3697] | layer3_out[3698];
    assign layer4_out[5635] = ~layer3_out[4518] | layer3_out[4517];
    assign layer4_out[5636] = layer3_out[4546];
    assign layer4_out[5637] = layer3_out[332];
    assign layer4_out[5638] = layer3_out[973] ^ layer3_out[974];
    assign layer4_out[5639] = layer3_out[4509];
    assign layer4_out[5640] = ~layer3_out[7818];
    assign layer4_out[5641] = layer3_out[2283] | layer3_out[2284];
    assign layer4_out[5642] = ~layer3_out[6863];
    assign layer4_out[5643] = layer3_out[2245] | layer3_out[2246];
    assign layer4_out[5644] = ~layer3_out[1195];
    assign layer4_out[5645] = ~layer3_out[7010];
    assign layer4_out[5646] = ~layer3_out[472];
    assign layer4_out[5647] = ~(layer3_out[4163] ^ layer3_out[4164]);
    assign layer4_out[5648] = ~(layer3_out[7482] ^ layer3_out[7483]);
    assign layer4_out[5649] = layer3_out[91] | layer3_out[92];
    assign layer4_out[5650] = ~layer3_out[159];
    assign layer4_out[5651] = ~layer3_out[2873];
    assign layer4_out[5652] = layer3_out[2748];
    assign layer4_out[5653] = ~layer3_out[7138];
    assign layer4_out[5654] = layer3_out[3334] & ~layer3_out[3333];
    assign layer4_out[5655] = layer3_out[6189];
    assign layer4_out[5656] = ~(layer3_out[6681] ^ layer3_out[6682]);
    assign layer4_out[5657] = layer3_out[4621];
    assign layer4_out[5658] = ~layer3_out[6088] | layer3_out[6089];
    assign layer4_out[5659] = 1'b1;
    assign layer4_out[5660] = ~layer3_out[6973] | layer3_out[6974];
    assign layer4_out[5661] = layer3_out[7935] ^ layer3_out[7936];
    assign layer4_out[5662] = ~layer3_out[6086];
    assign layer4_out[5663] = ~layer3_out[3025];
    assign layer4_out[5664] = ~layer3_out[5692];
    assign layer4_out[5665] = layer3_out[6381] & ~layer3_out[6380];
    assign layer4_out[5666] = ~layer3_out[7462] | layer3_out[7463];
    assign layer4_out[5667] = layer3_out[2485];
    assign layer4_out[5668] = ~(layer3_out[1052] ^ layer3_out[1053]);
    assign layer4_out[5669] = 1'b1;
    assign layer4_out[5670] = layer3_out[1611] ^ layer3_out[1612];
    assign layer4_out[5671] = layer3_out[1566];
    assign layer4_out[5672] = ~layer3_out[2006];
    assign layer4_out[5673] = ~layer3_out[894];
    assign layer4_out[5674] = ~(layer3_out[3846] & layer3_out[3847]);
    assign layer4_out[5675] = layer3_out[4657] & ~layer3_out[4656];
    assign layer4_out[5676] = layer3_out[6843] & ~layer3_out[6842];
    assign layer4_out[5677] = layer3_out[1174];
    assign layer4_out[5678] = ~(layer3_out[3700] | layer3_out[3701]);
    assign layer4_out[5679] = layer3_out[4807];
    assign layer4_out[5680] = ~(layer3_out[5519] | layer3_out[5520]);
    assign layer4_out[5681] = ~layer3_out[4042] | layer3_out[4043];
    assign layer4_out[5682] = ~(layer3_out[415] & layer3_out[416]);
    assign layer4_out[5683] = layer3_out[6623] & ~layer3_out[6622];
    assign layer4_out[5684] = layer3_out[2066];
    assign layer4_out[5685] = ~(layer3_out[7917] ^ layer3_out[7918]);
    assign layer4_out[5686] = layer3_out[3826] & ~layer3_out[3827];
    assign layer4_out[5687] = ~layer3_out[1457] | layer3_out[1456];
    assign layer4_out[5688] = layer3_out[7043];
    assign layer4_out[5689] = layer3_out[4410] & ~layer3_out[4411];
    assign layer4_out[5690] = ~layer3_out[1453];
    assign layer4_out[5691] = ~layer3_out[4329];
    assign layer4_out[5692] = layer3_out[3705];
    assign layer4_out[5693] = layer3_out[7296] ^ layer3_out[7297];
    assign layer4_out[5694] = layer3_out[2099];
    assign layer4_out[5695] = layer3_out[1726];
    assign layer4_out[5696] = ~layer3_out[2633] | layer3_out[2632];
    assign layer4_out[5697] = ~(layer3_out[2986] & layer3_out[2987]);
    assign layer4_out[5698] = ~layer3_out[4340] | layer3_out[4341];
    assign layer4_out[5699] = ~layer3_out[5677];
    assign layer4_out[5700] = layer3_out[3043];
    assign layer4_out[5701] = layer3_out[6665] & ~layer3_out[6664];
    assign layer4_out[5702] = ~(layer3_out[2760] | layer3_out[2761]);
    assign layer4_out[5703] = layer3_out[3509] ^ layer3_out[3510];
    assign layer4_out[5704] = layer3_out[3662];
    assign layer4_out[5705] = ~(layer3_out[3572] | layer3_out[3573]);
    assign layer4_out[5706] = layer3_out[7887] & ~layer3_out[7888];
    assign layer4_out[5707] = ~(layer3_out[6057] | layer3_out[6058]);
    assign layer4_out[5708] = ~(layer3_out[2192] ^ layer3_out[2193]);
    assign layer4_out[5709] = ~(layer3_out[6279] & layer3_out[6280]);
    assign layer4_out[5710] = ~layer3_out[2761];
    assign layer4_out[5711] = ~layer3_out[3430] | layer3_out[3429];
    assign layer4_out[5712] = layer3_out[2797] ^ layer3_out[2798];
    assign layer4_out[5713] = layer3_out[3183] & layer3_out[3184];
    assign layer4_out[5714] = layer3_out[946];
    assign layer4_out[5715] = layer3_out[4459] & ~layer3_out[4458];
    assign layer4_out[5716] = layer3_out[1221];
    assign layer4_out[5717] = layer3_out[1641] ^ layer3_out[1642];
    assign layer4_out[5718] = layer3_out[4452] & ~layer3_out[4451];
    assign layer4_out[5719] = layer3_out[1716];
    assign layer4_out[5720] = ~(layer3_out[5165] & layer3_out[5166]);
    assign layer4_out[5721] = ~layer3_out[4263];
    assign layer4_out[5722] = ~(layer3_out[826] & layer3_out[827]);
    assign layer4_out[5723] = layer3_out[929] & ~layer3_out[930];
    assign layer4_out[5724] = layer3_out[7456];
    assign layer4_out[5725] = layer3_out[5946] & layer3_out[5947];
    assign layer4_out[5726] = ~(layer3_out[1073] | layer3_out[1074]);
    assign layer4_out[5727] = ~layer3_out[7043];
    assign layer4_out[5728] = ~layer3_out[2180];
    assign layer4_out[5729] = layer3_out[3571] & ~layer3_out[3572];
    assign layer4_out[5730] = ~layer3_out[7097] | layer3_out[7098];
    assign layer4_out[5731] = ~(layer3_out[2352] & layer3_out[2353]);
    assign layer4_out[5732] = ~layer3_out[3923];
    assign layer4_out[5733] = ~(layer3_out[5507] | layer3_out[5508]);
    assign layer4_out[5734] = layer3_out[2514];
    assign layer4_out[5735] = layer3_out[2090] & layer3_out[2091];
    assign layer4_out[5736] = ~layer3_out[5983] | layer3_out[5984];
    assign layer4_out[5737] = layer3_out[6991] | layer3_out[6992];
    assign layer4_out[5738] = layer3_out[5966] ^ layer3_out[5967];
    assign layer4_out[5739] = layer3_out[962] ^ layer3_out[963];
    assign layer4_out[5740] = layer3_out[446];
    assign layer4_out[5741] = layer3_out[7787];
    assign layer4_out[5742] = ~layer3_out[475];
    assign layer4_out[5743] = layer3_out[2240] & ~layer3_out[2241];
    assign layer4_out[5744] = layer3_out[4274] | layer3_out[4275];
    assign layer4_out[5745] = ~layer3_out[5639];
    assign layer4_out[5746] = ~layer3_out[7360] | layer3_out[7359];
    assign layer4_out[5747] = ~layer3_out[5552];
    assign layer4_out[5748] = ~layer3_out[3797];
    assign layer4_out[5749] = layer3_out[6940] ^ layer3_out[6941];
    assign layer4_out[5750] = ~(layer3_out[4464] & layer3_out[4465]);
    assign layer4_out[5751] = layer3_out[6645];
    assign layer4_out[5752] = ~layer3_out[6262];
    assign layer4_out[5753] = ~(layer3_out[2336] ^ layer3_out[2337]);
    assign layer4_out[5754] = layer3_out[4827];
    assign layer4_out[5755] = layer3_out[1835] & ~layer3_out[1834];
    assign layer4_out[5756] = ~layer3_out[4552];
    assign layer4_out[5757] = ~layer3_out[3954];
    assign layer4_out[5758] = layer3_out[5173];
    assign layer4_out[5759] = ~(layer3_out[4874] | layer3_out[4875]);
    assign layer4_out[5760] = layer3_out[6890];
    assign layer4_out[5761] = layer3_out[6520] | layer3_out[6521];
    assign layer4_out[5762] = layer3_out[6386] & ~layer3_out[6387];
    assign layer4_out[5763] = layer3_out[5065];
    assign layer4_out[5764] = ~(layer3_out[6515] ^ layer3_out[6516]);
    assign layer4_out[5765] = ~(layer3_out[6381] ^ layer3_out[6382]);
    assign layer4_out[5766] = ~layer3_out[5426];
    assign layer4_out[5767] = ~layer3_out[7268];
    assign layer4_out[5768] = layer3_out[1048];
    assign layer4_out[5769] = layer3_out[5802] & ~layer3_out[5801];
    assign layer4_out[5770] = ~layer3_out[4378];
    assign layer4_out[5771] = 1'b1;
    assign layer4_out[5772] = ~(layer3_out[2161] ^ layer3_out[2162]);
    assign layer4_out[5773] = layer3_out[1639] ^ layer3_out[1640];
    assign layer4_out[5774] = ~(layer3_out[6451] & layer3_out[6452]);
    assign layer4_out[5775] = ~layer3_out[2635] | layer3_out[2636];
    assign layer4_out[5776] = layer3_out[1667];
    assign layer4_out[5777] = layer3_out[1547] ^ layer3_out[1548];
    assign layer4_out[5778] = layer3_out[2286];
    assign layer4_out[5779] = layer3_out[877];
    assign layer4_out[5780] = layer3_out[5125] | layer3_out[5126];
    assign layer4_out[5781] = layer3_out[5086] | layer3_out[5087];
    assign layer4_out[5782] = layer3_out[7333];
    assign layer4_out[5783] = layer3_out[3304] & layer3_out[3305];
    assign layer4_out[5784] = ~layer3_out[3508];
    assign layer4_out[5785] = layer3_out[5042] | layer3_out[5043];
    assign layer4_out[5786] = ~(layer3_out[6980] & layer3_out[6981]);
    assign layer4_out[5787] = ~layer3_out[681];
    assign layer4_out[5788] = layer3_out[7124] ^ layer3_out[7125];
    assign layer4_out[5789] = ~layer3_out[6405];
    assign layer4_out[5790] = layer3_out[5905];
    assign layer4_out[5791] = layer3_out[4038] | layer3_out[4039];
    assign layer4_out[5792] = ~(layer3_out[2894] | layer3_out[2895]);
    assign layer4_out[5793] = layer3_out[3075] & ~layer3_out[3076];
    assign layer4_out[5794] = ~layer3_out[805];
    assign layer4_out[5795] = layer3_out[6163] ^ layer3_out[6164];
    assign layer4_out[5796] = ~layer3_out[1106] | layer3_out[1107];
    assign layer4_out[5797] = ~layer3_out[5532];
    assign layer4_out[5798] = layer3_out[5272];
    assign layer4_out[5799] = layer3_out[3056] & ~layer3_out[3055];
    assign layer4_out[5800] = ~layer3_out[6526];
    assign layer4_out[5801] = layer3_out[5225];
    assign layer4_out[5802] = ~layer3_out[4899];
    assign layer4_out[5803] = ~(layer3_out[4957] ^ layer3_out[4958]);
    assign layer4_out[5804] = layer3_out[1758];
    assign layer4_out[5805] = ~layer3_out[7597];
    assign layer4_out[5806] = ~layer3_out[7763];
    assign layer4_out[5807] = ~(layer3_out[7472] | layer3_out[7473]);
    assign layer4_out[5808] = layer3_out[6833] ^ layer3_out[6834];
    assign layer4_out[5809] = layer3_out[4681] | layer3_out[4682];
    assign layer4_out[5810] = ~(layer3_out[320] | layer3_out[321]);
    assign layer4_out[5811] = layer3_out[7689] | layer3_out[7690];
    assign layer4_out[5812] = ~layer3_out[5367];
    assign layer4_out[5813] = ~layer3_out[2558];
    assign layer4_out[5814] = layer3_out[3248] & ~layer3_out[3249];
    assign layer4_out[5815] = ~(layer3_out[3137] & layer3_out[3138]);
    assign layer4_out[5816] = ~layer3_out[2496] | layer3_out[2497];
    assign layer4_out[5817] = layer3_out[4728];
    assign layer4_out[5818] = layer3_out[3184];
    assign layer4_out[5819] = layer3_out[1036] ^ layer3_out[1037];
    assign layer4_out[5820] = layer3_out[423] ^ layer3_out[424];
    assign layer4_out[5821] = ~layer3_out[7382] | layer3_out[7383];
    assign layer4_out[5822] = layer3_out[192];
    assign layer4_out[5823] = ~layer3_out[2395];
    assign layer4_out[5824] = ~(layer3_out[6040] ^ layer3_out[6041]);
    assign layer4_out[5825] = layer3_out[5044] & ~layer3_out[5043];
    assign layer4_out[5826] = ~layer3_out[3177] | layer3_out[3176];
    assign layer4_out[5827] = layer3_out[2410];
    assign layer4_out[5828] = ~layer3_out[2642];
    assign layer4_out[5829] = layer3_out[1992] & ~layer3_out[1993];
    assign layer4_out[5830] = layer3_out[849] & ~layer3_out[850];
    assign layer4_out[5831] = ~(layer3_out[7745] ^ layer3_out[7746]);
    assign layer4_out[5832] = layer3_out[6444] ^ layer3_out[6445];
    assign layer4_out[5833] = layer3_out[3309] | layer3_out[3310];
    assign layer4_out[5834] = layer3_out[2285] & ~layer3_out[2284];
    assign layer4_out[5835] = ~layer3_out[6082];
    assign layer4_out[5836] = layer3_out[4080] & layer3_out[4081];
    assign layer4_out[5837] = ~layer3_out[5254];
    assign layer4_out[5838] = layer3_out[1436];
    assign layer4_out[5839] = layer3_out[5007];
    assign layer4_out[5840] = layer3_out[7127] & layer3_out[7128];
    assign layer4_out[5841] = layer3_out[2905] & ~layer3_out[2906];
    assign layer4_out[5842] = 1'b0;
    assign layer4_out[5843] = layer3_out[5698];
    assign layer4_out[5844] = ~layer3_out[3212];
    assign layer4_out[5845] = layer3_out[4915] & ~layer3_out[4914];
    assign layer4_out[5846] = layer3_out[200];
    assign layer4_out[5847] = layer3_out[6028] & ~layer3_out[6027];
    assign layer4_out[5848] = layer3_out[2361] ^ layer3_out[2362];
    assign layer4_out[5849] = layer3_out[5400] ^ layer3_out[5401];
    assign layer4_out[5850] = ~(layer3_out[3037] ^ layer3_out[3038]);
    assign layer4_out[5851] = ~(layer3_out[2279] & layer3_out[2280]);
    assign layer4_out[5852] = ~(layer3_out[1994] & layer3_out[1995]);
    assign layer4_out[5853] = ~(layer3_out[720] ^ layer3_out[721]);
    assign layer4_out[5854] = layer3_out[724] & layer3_out[725];
    assign layer4_out[5855] = layer3_out[1350] ^ layer3_out[1351];
    assign layer4_out[5856] = ~layer3_out[7547] | layer3_out[7548];
    assign layer4_out[5857] = ~layer3_out[630];
    assign layer4_out[5858] = layer3_out[1413] & ~layer3_out[1414];
    assign layer4_out[5859] = layer3_out[2412] ^ layer3_out[2413];
    assign layer4_out[5860] = layer3_out[5924];
    assign layer4_out[5861] = ~layer3_out[3060];
    assign layer4_out[5862] = ~layer3_out[4398];
    assign layer4_out[5863] = ~(layer3_out[1460] ^ layer3_out[1461]);
    assign layer4_out[5864] = layer3_out[612] & ~layer3_out[611];
    assign layer4_out[5865] = layer3_out[3935];
    assign layer4_out[5866] = ~layer3_out[3003];
    assign layer4_out[5867] = layer3_out[5041] & ~layer3_out[5042];
    assign layer4_out[5868] = ~layer3_out[3169];
    assign layer4_out[5869] = layer3_out[4372] & layer3_out[4373];
    assign layer4_out[5870] = layer3_out[1873] & layer3_out[1874];
    assign layer4_out[5871] = layer3_out[1509];
    assign layer4_out[5872] = ~(layer3_out[6182] | layer3_out[6183]);
    assign layer4_out[5873] = ~(layer3_out[1163] & layer3_out[1164]);
    assign layer4_out[5874] = layer3_out[363];
    assign layer4_out[5875] = layer3_out[2535] & layer3_out[2536];
    assign layer4_out[5876] = layer3_out[6261] ^ layer3_out[6262];
    assign layer4_out[5877] = layer3_out[3960] & layer3_out[3961];
    assign layer4_out[5878] = layer3_out[5382] ^ layer3_out[5383];
    assign layer4_out[5879] = ~(layer3_out[5252] | layer3_out[5253]);
    assign layer4_out[5880] = layer3_out[179] | layer3_out[180];
    assign layer4_out[5881] = layer3_out[6697] & ~layer3_out[6698];
    assign layer4_out[5882] = layer3_out[4820];
    assign layer4_out[5883] = ~(layer3_out[757] & layer3_out[758]);
    assign layer4_out[5884] = ~(layer3_out[2151] | layer3_out[2152]);
    assign layer4_out[5885] = ~layer3_out[4233];
    assign layer4_out[5886] = ~layer3_out[4457];
    assign layer4_out[5887] = layer3_out[2357];
    assign layer4_out[5888] = layer3_out[2425] | layer3_out[2426];
    assign layer4_out[5889] = ~layer3_out[4992];
    assign layer4_out[5890] = layer3_out[5907] & ~layer3_out[5906];
    assign layer4_out[5891] = layer3_out[5664];
    assign layer4_out[5892] = layer3_out[2790] ^ layer3_out[2791];
    assign layer4_out[5893] = layer3_out[6092];
    assign layer4_out[5894] = layer3_out[4000];
    assign layer4_out[5895] = layer3_out[7320] ^ layer3_out[7321];
    assign layer4_out[5896] = ~(layer3_out[5465] & layer3_out[5466]);
    assign layer4_out[5897] = ~layer3_out[1150];
    assign layer4_out[5898] = layer3_out[4574];
    assign layer4_out[5899] = layer3_out[5112];
    assign layer4_out[5900] = ~(layer3_out[7437] ^ layer3_out[7438]);
    assign layer4_out[5901] = ~layer3_out[5007] | layer3_out[5006];
    assign layer4_out[5902] = ~layer3_out[185] | layer3_out[184];
    assign layer4_out[5903] = ~layer3_out[5487];
    assign layer4_out[5904] = ~layer3_out[7619];
    assign layer4_out[5905] = ~layer3_out[4048];
    assign layer4_out[5906] = ~layer3_out[5736];
    assign layer4_out[5907] = layer3_out[3200] | layer3_out[3201];
    assign layer4_out[5908] = ~(layer3_out[3257] | layer3_out[3258]);
    assign layer4_out[5909] = ~layer3_out[6485];
    assign layer4_out[5910] = ~layer3_out[7472];
    assign layer4_out[5911] = layer3_out[1744] & layer3_out[1745];
    assign layer4_out[5912] = layer3_out[1618];
    assign layer4_out[5913] = ~layer3_out[5314];
    assign layer4_out[5914] = ~(layer3_out[5846] ^ layer3_out[5847]);
    assign layer4_out[5915] = layer3_out[1959] | layer3_out[1960];
    assign layer4_out[5916] = ~(layer3_out[4119] | layer3_out[4120]);
    assign layer4_out[5917] = layer3_out[3132] & layer3_out[3133];
    assign layer4_out[5918] = ~(layer3_out[7261] ^ layer3_out[7262]);
    assign layer4_out[5919] = layer3_out[1591] & ~layer3_out[1590];
    assign layer4_out[5920] = layer3_out[5798] & ~layer3_out[5797];
    assign layer4_out[5921] = ~layer3_out[4814];
    assign layer4_out[5922] = layer3_out[1923] & ~layer3_out[1924];
    assign layer4_out[5923] = ~layer3_out[2674];
    assign layer4_out[5924] = ~layer3_out[900] | layer3_out[901];
    assign layer4_out[5925] = layer3_out[4473];
    assign layer4_out[5926] = ~(layer3_out[3162] & layer3_out[3163]);
    assign layer4_out[5927] = layer3_out[6095];
    assign layer4_out[5928] = layer3_out[6460] & ~layer3_out[6459];
    assign layer4_out[5929] = layer3_out[5258];
    assign layer4_out[5930] = ~layer3_out[2393];
    assign layer4_out[5931] = ~layer3_out[6432] | layer3_out[6433];
    assign layer4_out[5932] = ~(layer3_out[7102] ^ layer3_out[7103]);
    assign layer4_out[5933] = ~layer3_out[645] | layer3_out[646];
    assign layer4_out[5934] = ~layer3_out[4221];
    assign layer4_out[5935] = layer3_out[4581] & ~layer3_out[4582];
    assign layer4_out[5936] = ~(layer3_out[2628] | layer3_out[2629]);
    assign layer4_out[5937] = layer3_out[2671];
    assign layer4_out[5938] = layer3_out[7806] ^ layer3_out[7807];
    assign layer4_out[5939] = layer3_out[4038];
    assign layer4_out[5940] = layer3_out[7449] | layer3_out[7450];
    assign layer4_out[5941] = layer3_out[5239];
    assign layer4_out[5942] = ~(layer3_out[6578] | layer3_out[6579]);
    assign layer4_out[5943] = ~layer3_out[2918];
    assign layer4_out[5944] = ~layer3_out[7558];
    assign layer4_out[5945] = ~layer3_out[5720] | layer3_out[5721];
    assign layer4_out[5946] = 1'b0;
    assign layer4_out[5947] = layer3_out[6062] & ~layer3_out[6061];
    assign layer4_out[5948] = layer3_out[3010] | layer3_out[3011];
    assign layer4_out[5949] = ~layer3_out[4572];
    assign layer4_out[5950] = layer3_out[6465] | layer3_out[6466];
    assign layer4_out[5951] = ~layer3_out[1043];
    assign layer4_out[5952] = layer3_out[2030];
    assign layer4_out[5953] = ~layer3_out[1161] | layer3_out[1160];
    assign layer4_out[5954] = ~(layer3_out[7551] & layer3_out[7552]);
    assign layer4_out[5955] = ~(layer3_out[7571] | layer3_out[7572]);
    assign layer4_out[5956] = ~(layer3_out[1909] & layer3_out[1910]);
    assign layer4_out[5957] = ~layer3_out[1759] | layer3_out[1760];
    assign layer4_out[5958] = ~layer3_out[6480] | layer3_out[6481];
    assign layer4_out[5959] = layer3_out[3896];
    assign layer4_out[5960] = ~layer3_out[6087];
    assign layer4_out[5961] = ~(layer3_out[765] & layer3_out[766]);
    assign layer4_out[5962] = ~(layer3_out[6070] | layer3_out[6071]);
    assign layer4_out[5963] = layer3_out[16] & layer3_out[17];
    assign layer4_out[5964] = ~(layer3_out[2497] ^ layer3_out[2498]);
    assign layer4_out[5965] = ~(layer3_out[7354] & layer3_out[7355]);
    assign layer4_out[5966] = ~layer3_out[4179] | layer3_out[4178];
    assign layer4_out[5967] = ~layer3_out[7244] | layer3_out[7245];
    assign layer4_out[5968] = layer3_out[3352] | layer3_out[3353];
    assign layer4_out[5969] = ~layer3_out[7871];
    assign layer4_out[5970] = ~layer3_out[3878];
    assign layer4_out[5971] = ~layer3_out[4514];
    assign layer4_out[5972] = ~(layer3_out[5918] ^ layer3_out[5919]);
    assign layer4_out[5973] = layer3_out[1925];
    assign layer4_out[5974] = layer3_out[2676];
    assign layer4_out[5975] = ~layer3_out[6044];
    assign layer4_out[5976] = ~layer3_out[2446] | layer3_out[2445];
    assign layer4_out[5977] = layer3_out[1048] & ~layer3_out[1049];
    assign layer4_out[5978] = ~layer3_out[5380];
    assign layer4_out[5979] = layer3_out[1455] & ~layer3_out[1456];
    assign layer4_out[5980] = layer3_out[4222] & ~layer3_out[4221];
    assign layer4_out[5981] = ~(layer3_out[3655] & layer3_out[3656]);
    assign layer4_out[5982] = ~layer3_out[1332];
    assign layer4_out[5983] = ~(layer3_out[2217] & layer3_out[2218]);
    assign layer4_out[5984] = layer3_out[5442] | layer3_out[5443];
    assign layer4_out[5985] = layer3_out[3742] & layer3_out[3743];
    assign layer4_out[5986] = layer3_out[6926];
    assign layer4_out[5987] = ~layer3_out[6141] | layer3_out[6140];
    assign layer4_out[5988] = ~layer3_out[4971];
    assign layer4_out[5989] = layer3_out[5281] ^ layer3_out[5282];
    assign layer4_out[5990] = ~layer3_out[6440];
    assign layer4_out[5991] = ~layer3_out[2627];
    assign layer4_out[5992] = layer3_out[498];
    assign layer4_out[5993] = layer3_out[6734];
    assign layer4_out[5994] = ~layer3_out[7497];
    assign layer4_out[5995] = layer3_out[7201] | layer3_out[7202];
    assign layer4_out[5996] = layer3_out[3194] ^ layer3_out[3195];
    assign layer4_out[5997] = ~layer3_out[1545];
    assign layer4_out[5998] = ~layer3_out[5095];
    assign layer4_out[5999] = ~layer3_out[1730] | layer3_out[1729];
    assign layer4_out[6000] = ~layer3_out[6634];
    assign layer4_out[6001] = ~layer3_out[4999];
    assign layer4_out[6002] = layer3_out[7627];
    assign layer4_out[6003] = ~layer3_out[5147];
    assign layer4_out[6004] = layer3_out[4327];
    assign layer4_out[6005] = ~(layer3_out[5011] ^ layer3_out[5012]);
    assign layer4_out[6006] = ~layer3_out[4358];
    assign layer4_out[6007] = ~(layer3_out[5597] | layer3_out[5598]);
    assign layer4_out[6008] = ~layer3_out[5772];
    assign layer4_out[6009] = layer3_out[6433] & layer3_out[6434];
    assign layer4_out[6010] = ~layer3_out[2929];
    assign layer4_out[6011] = ~layer3_out[5384];
    assign layer4_out[6012] = ~(layer3_out[7617] ^ layer3_out[7618]);
    assign layer4_out[6013] = ~layer3_out[2677];
    assign layer4_out[6014] = layer3_out[5390];
    assign layer4_out[6015] = ~layer3_out[2913] | layer3_out[2914];
    assign layer4_out[6016] = ~(layer3_out[7277] & layer3_out[7278]);
    assign layer4_out[6017] = ~layer3_out[2717] | layer3_out[2716];
    assign layer4_out[6018] = ~layer3_out[2290];
    assign layer4_out[6019] = ~layer3_out[6988] | layer3_out[6989];
    assign layer4_out[6020] = layer3_out[3990] & ~layer3_out[3991];
    assign layer4_out[6021] = layer3_out[5763] & ~layer3_out[5764];
    assign layer4_out[6022] = ~(layer3_out[6199] & layer3_out[6200]);
    assign layer4_out[6023] = layer3_out[3115];
    assign layer4_out[6024] = layer3_out[971] | layer3_out[972];
    assign layer4_out[6025] = layer3_out[463] & ~layer3_out[462];
    assign layer4_out[6026] = ~(layer3_out[1804] ^ layer3_out[1805]);
    assign layer4_out[6027] = ~layer3_out[3818] | layer3_out[3817];
    assign layer4_out[6028] = layer3_out[6188] & layer3_out[6189];
    assign layer4_out[6029] = layer3_out[7511] ^ layer3_out[7512];
    assign layer4_out[6030] = layer3_out[4225];
    assign layer4_out[6031] = ~(layer3_out[3570] & layer3_out[3571]);
    assign layer4_out[6032] = layer3_out[3181];
    assign layer4_out[6033] = ~layer3_out[2267];
    assign layer4_out[6034] = ~(layer3_out[6033] | layer3_out[6034]);
    assign layer4_out[6035] = layer3_out[1434] ^ layer3_out[1435];
    assign layer4_out[6036] = ~(layer3_out[1886] | layer3_out[1887]);
    assign layer4_out[6037] = layer3_out[1599] ^ layer3_out[1600];
    assign layer4_out[6038] = ~layer3_out[7] | layer3_out[6];
    assign layer4_out[6039] = layer3_out[1426] ^ layer3_out[1427];
    assign layer4_out[6040] = ~layer3_out[1598];
    assign layer4_out[6041] = layer3_out[3327] & ~layer3_out[3326];
    assign layer4_out[6042] = ~(layer3_out[4049] ^ layer3_out[4050]);
    assign layer4_out[6043] = ~layer3_out[2265] | layer3_out[2266];
    assign layer4_out[6044] = ~layer3_out[5580];
    assign layer4_out[6045] = ~(layer3_out[3797] | layer3_out[3798]);
    assign layer4_out[6046] = ~layer3_out[2218] | layer3_out[2219];
    assign layer4_out[6047] = layer3_out[769];
    assign layer4_out[6048] = layer3_out[1626];
    assign layer4_out[6049] = ~layer3_out[6628];
    assign layer4_out[6050] = ~layer3_out[4784];
    assign layer4_out[6051] = ~layer3_out[4945];
    assign layer4_out[6052] = layer3_out[2708] & layer3_out[2709];
    assign layer4_out[6053] = ~layer3_out[2556] | layer3_out[2557];
    assign layer4_out[6054] = layer3_out[6835] ^ layer3_out[6836];
    assign layer4_out[6055] = layer3_out[127] | layer3_out[128];
    assign layer4_out[6056] = layer3_out[10] ^ layer3_out[11];
    assign layer4_out[6057] = layer3_out[211];
    assign layer4_out[6058] = ~(layer3_out[476] & layer3_out[477]);
    assign layer4_out[6059] = layer3_out[4779] ^ layer3_out[4780];
    assign layer4_out[6060] = ~(layer3_out[3387] | layer3_out[3388]);
    assign layer4_out[6061] = layer3_out[3893] ^ layer3_out[3894];
    assign layer4_out[6062] = ~layer3_out[4669];
    assign layer4_out[6063] = ~(layer3_out[472] & layer3_out[473]);
    assign layer4_out[6064] = layer3_out[2083] ^ layer3_out[2084];
    assign layer4_out[6065] = layer3_out[3784] ^ layer3_out[3785];
    assign layer4_out[6066] = layer3_out[809] ^ layer3_out[810];
    assign layer4_out[6067] = layer3_out[5929];
    assign layer4_out[6068] = layer3_out[6265];
    assign layer4_out[6069] = layer3_out[2751] | layer3_out[2752];
    assign layer4_out[6070] = layer3_out[4749] & layer3_out[4750];
    assign layer4_out[6071] = ~layer3_out[737] | layer3_out[738];
    assign layer4_out[6072] = ~layer3_out[5882];
    assign layer4_out[6073] = layer3_out[3712];
    assign layer4_out[6074] = ~layer3_out[888];
    assign layer4_out[6075] = ~layer3_out[6487] | layer3_out[6486];
    assign layer4_out[6076] = layer3_out[7997] & layer3_out[7998];
    assign layer4_out[6077] = layer3_out[4560];
    assign layer4_out[6078] = layer3_out[7636] & ~layer3_out[7635];
    assign layer4_out[6079] = ~layer3_out[5620];
    assign layer4_out[6080] = layer3_out[2143];
    assign layer4_out[6081] = layer3_out[2705];
    assign layer4_out[6082] = ~layer3_out[992];
    assign layer4_out[6083] = layer3_out[7037] & layer3_out[7038];
    assign layer4_out[6084] = ~layer3_out[6036];
    assign layer4_out[6085] = ~(layer3_out[6009] ^ layer3_out[6010]);
    assign layer4_out[6086] = ~(layer3_out[6826] ^ layer3_out[6827]);
    assign layer4_out[6087] = ~layer3_out[4580];
    assign layer4_out[6088] = ~layer3_out[7077];
    assign layer4_out[6089] = layer3_out[2771] & ~layer3_out[2770];
    assign layer4_out[6090] = ~(layer3_out[7336] & layer3_out[7337]);
    assign layer4_out[6091] = ~layer3_out[7871];
    assign layer4_out[6092] = layer3_out[6686] & ~layer3_out[6687];
    assign layer4_out[6093] = layer3_out[5816];
    assign layer4_out[6094] = ~(layer3_out[4677] ^ layer3_out[4678]);
    assign layer4_out[6095] = ~layer3_out[261] | layer3_out[260];
    assign layer4_out[6096] = layer3_out[6344];
    assign layer4_out[6097] = layer3_out[574] & ~layer3_out[575];
    assign layer4_out[6098] = ~layer3_out[605];
    assign layer4_out[6099] = ~layer3_out[5629];
    assign layer4_out[6100] = layer3_out[2075] & ~layer3_out[2076];
    assign layer4_out[6101] = layer3_out[7449] & ~layer3_out[7448];
    assign layer4_out[6102] = ~layer3_out[5353] | layer3_out[5352];
    assign layer4_out[6103] = layer3_out[7203] & ~layer3_out[7202];
    assign layer4_out[6104] = layer3_out[5141];
    assign layer4_out[6105] = layer3_out[2706] ^ layer3_out[2707];
    assign layer4_out[6106] = layer3_out[4792];
    assign layer4_out[6107] = ~(layer3_out[6193] ^ layer3_out[6194]);
    assign layer4_out[6108] = ~(layer3_out[1480] & layer3_out[1481]);
    assign layer4_out[6109] = ~(layer3_out[943] ^ layer3_out[944]);
    assign layer4_out[6110] = ~layer3_out[1351];
    assign layer4_out[6111] = layer3_out[3410] | layer3_out[3411];
    assign layer4_out[6112] = layer3_out[6563];
    assign layer4_out[6113] = ~layer3_out[7540];
    assign layer4_out[6114] = layer3_out[4215];
    assign layer4_out[6115] = ~layer3_out[2287] | layer3_out[2288];
    assign layer4_out[6116] = layer3_out[3403];
    assign layer4_out[6117] = ~layer3_out[7180];
    assign layer4_out[6118] = ~layer3_out[1421];
    assign layer4_out[6119] = layer3_out[2333];
    assign layer4_out[6120] = ~(layer3_out[3746] ^ layer3_out[3747]);
    assign layer4_out[6121] = layer3_out[5542] ^ layer3_out[5543];
    assign layer4_out[6122] = layer3_out[5384] | layer3_out[5385];
    assign layer4_out[6123] = layer3_out[342] & ~layer3_out[343];
    assign layer4_out[6124] = ~layer3_out[2088];
    assign layer4_out[6125] = layer3_out[3586] ^ layer3_out[3587];
    assign layer4_out[6126] = layer3_out[51];
    assign layer4_out[6127] = layer3_out[5511];
    assign layer4_out[6128] = ~layer3_out[4392] | layer3_out[4393];
    assign layer4_out[6129] = layer3_out[6315] & ~layer3_out[6314];
    assign layer4_out[6130] = layer3_out[163] & ~layer3_out[164];
    assign layer4_out[6131] = ~(layer3_out[7185] | layer3_out[7186]);
    assign layer4_out[6132] = layer3_out[7452] ^ layer3_out[7453];
    assign layer4_out[6133] = layer3_out[700] | layer3_out[701];
    assign layer4_out[6134] = layer3_out[2229] & ~layer3_out[2228];
    assign layer4_out[6135] = 1'b0;
    assign layer4_out[6136] = ~layer3_out[897] | layer3_out[898];
    assign layer4_out[6137] = layer3_out[94] ^ layer3_out[95];
    assign layer4_out[6138] = ~(layer3_out[1894] | layer3_out[1895]);
    assign layer4_out[6139] = ~layer3_out[2823];
    assign layer4_out[6140] = layer3_out[1986] ^ layer3_out[1987];
    assign layer4_out[6141] = layer3_out[5619] & ~layer3_out[5618];
    assign layer4_out[6142] = layer3_out[4185];
    assign layer4_out[6143] = layer3_out[253] & ~layer3_out[254];
    assign layer4_out[6144] = layer3_out[7397];
    assign layer4_out[6145] = layer3_out[1023];
    assign layer4_out[6146] = layer3_out[1899];
    assign layer4_out[6147] = layer3_out[4841] & ~layer3_out[4842];
    assign layer4_out[6148] = layer3_out[7839] & ~layer3_out[7840];
    assign layer4_out[6149] = layer3_out[2708] & ~layer3_out[2707];
    assign layer4_out[6150] = layer3_out[4752] | layer3_out[4753];
    assign layer4_out[6151] = layer3_out[6882] ^ layer3_out[6883];
    assign layer4_out[6152] = layer3_out[7686];
    assign layer4_out[6153] = ~(layer3_out[5413] ^ layer3_out[5414]);
    assign layer4_out[6154] = layer3_out[7458] & ~layer3_out[7457];
    assign layer4_out[6155] = layer3_out[7658] & layer3_out[7659];
    assign layer4_out[6156] = layer3_out[7835] & ~layer3_out[7836];
    assign layer4_out[6157] = layer3_out[3240] & ~layer3_out[3241];
    assign layer4_out[6158] = 1'b0;
    assign layer4_out[6159] = ~(layer3_out[6550] & layer3_out[6551]);
    assign layer4_out[6160] = layer3_out[6709] ^ layer3_out[6710];
    assign layer4_out[6161] = layer3_out[3600];
    assign layer4_out[6162] = ~(layer3_out[4234] ^ layer3_out[4235]);
    assign layer4_out[6163] = 1'b1;
    assign layer4_out[6164] = layer3_out[7188] ^ layer3_out[7189];
    assign layer4_out[6165] = layer3_out[6057];
    assign layer4_out[6166] = ~(layer3_out[5659] & layer3_out[5660]);
    assign layer4_out[6167] = ~layer3_out[317];
    assign layer4_out[6168] = layer3_out[5049];
    assign layer4_out[6169] = ~layer3_out[239] | layer3_out[238];
    assign layer4_out[6170] = ~layer3_out[5483] | layer3_out[5484];
    assign layer4_out[6171] = ~layer3_out[2231];
    assign layer4_out[6172] = layer3_out[5595];
    assign layer4_out[6173] = ~layer3_out[5267] | layer3_out[5268];
    assign layer4_out[6174] = layer3_out[3602] & layer3_out[3603];
    assign layer4_out[6175] = ~layer3_out[6295];
    assign layer4_out[6176] = ~layer3_out[7619];
    assign layer4_out[6177] = ~layer3_out[3981] | layer3_out[3980];
    assign layer4_out[6178] = ~(layer3_out[5110] ^ layer3_out[5111]);
    assign layer4_out[6179] = layer3_out[7659] | layer3_out[7660];
    assign layer4_out[6180] = layer3_out[3411];
    assign layer4_out[6181] = ~(layer3_out[6307] & layer3_out[6308]);
    assign layer4_out[6182] = ~layer3_out[771];
    assign layer4_out[6183] = layer3_out[2271] & ~layer3_out[2270];
    assign layer4_out[6184] = layer3_out[7026] ^ layer3_out[7027];
    assign layer4_out[6185] = layer3_out[1534] ^ layer3_out[1535];
    assign layer4_out[6186] = ~layer3_out[641] | layer3_out[640];
    assign layer4_out[6187] = ~(layer3_out[687] | layer3_out[688]);
    assign layer4_out[6188] = layer3_out[835];
    assign layer4_out[6189] = layer3_out[7222];
    assign layer4_out[6190] = ~layer3_out[6257];
    assign layer4_out[6191] = ~(layer3_out[3617] ^ layer3_out[3618]);
    assign layer4_out[6192] = ~(layer3_out[7793] ^ layer3_out[7794]);
    assign layer4_out[6193] = ~(layer3_out[2762] ^ layer3_out[2763]);
    assign layer4_out[6194] = layer3_out[2819] | layer3_out[2820];
    assign layer4_out[6195] = layer3_out[5444] & ~layer3_out[5445];
    assign layer4_out[6196] = ~(layer3_out[634] ^ layer3_out[635]);
    assign layer4_out[6197] = layer3_out[5533];
    assign layer4_out[6198] = ~layer3_out[7625];
    assign layer4_out[6199] = ~layer3_out[7422] | layer3_out[7423];
    assign layer4_out[6200] = ~layer3_out[1347] | layer3_out[1346];
    assign layer4_out[6201] = ~(layer3_out[7287] | layer3_out[7288]);
    assign layer4_out[6202] = layer3_out[3647];
    assign layer4_out[6203] = layer3_out[920];
    assign layer4_out[6204] = ~layer3_out[2158];
    assign layer4_out[6205] = layer3_out[1806] & ~layer3_out[1807];
    assign layer4_out[6206] = layer3_out[5661];
    assign layer4_out[6207] = layer3_out[3231] & ~layer3_out[3232];
    assign layer4_out[6208] = ~(layer3_out[5005] | layer3_out[5006]);
    assign layer4_out[6209] = ~layer3_out[4222];
    assign layer4_out[6210] = ~(layer3_out[711] ^ layer3_out[712]);
    assign layer4_out[6211] = ~layer3_out[886];
    assign layer4_out[6212] = ~(layer3_out[1807] | layer3_out[1808]);
    assign layer4_out[6213] = ~(layer3_out[5139] & layer3_out[5140]);
    assign layer4_out[6214] = ~layer3_out[6426] | layer3_out[6427];
    assign layer4_out[6215] = layer3_out[77] & ~layer3_out[76];
    assign layer4_out[6216] = ~layer3_out[5457];
    assign layer4_out[6217] = ~(layer3_out[5996] ^ layer3_out[5997]);
    assign layer4_out[6218] = ~layer3_out[7422] | layer3_out[7421];
    assign layer4_out[6219] = layer3_out[4679];
    assign layer4_out[6220] = layer3_out[5959] & ~layer3_out[5960];
    assign layer4_out[6221] = layer3_out[4259] ^ layer3_out[4260];
    assign layer4_out[6222] = layer3_out[1131] ^ layer3_out[1132];
    assign layer4_out[6223] = ~layer3_out[7697];
    assign layer4_out[6224] = layer3_out[2698];
    assign layer4_out[6225] = layer3_out[6756] & layer3_out[6757];
    assign layer4_out[6226] = ~layer3_out[5233];
    assign layer4_out[6227] = layer3_out[4174] | layer3_out[4175];
    assign layer4_out[6228] = layer3_out[7779] ^ layer3_out[7780];
    assign layer4_out[6229] = ~layer3_out[3557];
    assign layer4_out[6230] = ~(layer3_out[3866] ^ layer3_out[3867]);
    assign layer4_out[6231] = ~(layer3_out[2101] ^ layer3_out[2102]);
    assign layer4_out[6232] = layer3_out[5317] & layer3_out[5318];
    assign layer4_out[6233] = layer3_out[2340] & ~layer3_out[2339];
    assign layer4_out[6234] = layer3_out[5680];
    assign layer4_out[6235] = ~layer3_out[1431];
    assign layer4_out[6236] = layer3_out[4333];
    assign layer4_out[6237] = ~(layer3_out[3908] | layer3_out[3909]);
    assign layer4_out[6238] = layer3_out[2731];
    assign layer4_out[6239] = layer3_out[4399];
    assign layer4_out[6240] = ~layer3_out[1621] | layer3_out[1620];
    assign layer4_out[6241] = layer3_out[6750];
    assign layer4_out[6242] = layer3_out[346];
    assign layer4_out[6243] = layer3_out[3831] ^ layer3_out[3832];
    assign layer4_out[6244] = layer3_out[5530];
    assign layer4_out[6245] = layer3_out[1251];
    assign layer4_out[6246] = ~layer3_out[2835];
    assign layer4_out[6247] = ~(layer3_out[6123] & layer3_out[6124]);
    assign layer4_out[6248] = ~layer3_out[4562];
    assign layer4_out[6249] = layer3_out[1447] & ~layer3_out[1448];
    assign layer4_out[6250] = ~layer3_out[7653] | layer3_out[7654];
    assign layer4_out[6251] = ~layer3_out[6794] | layer3_out[6793];
    assign layer4_out[6252] = layer3_out[1316];
    assign layer4_out[6253] = ~(layer3_out[629] & layer3_out[630]);
    assign layer4_out[6254] = ~(layer3_out[3583] & layer3_out[3584]);
    assign layer4_out[6255] = layer3_out[2950];
    assign layer4_out[6256] = layer3_out[5073];
    assign layer4_out[6257] = ~(layer3_out[5675] ^ layer3_out[5676]);
    assign layer4_out[6258] = layer3_out[7695] & ~layer3_out[7696];
    assign layer4_out[6259] = layer3_out[642];
    assign layer4_out[6260] = layer3_out[1585];
    assign layer4_out[6261] = ~(layer3_out[7891] ^ layer3_out[7892]);
    assign layer4_out[6262] = layer3_out[6582] ^ layer3_out[6583];
    assign layer4_out[6263] = ~(layer3_out[5020] & layer3_out[5021]);
    assign layer4_out[6264] = ~layer3_out[2584];
    assign layer4_out[6265] = ~layer3_out[7103] | layer3_out[7104];
    assign layer4_out[6266] = layer3_out[5980] & ~layer3_out[5979];
    assign layer4_out[6267] = layer3_out[5574];
    assign layer4_out[6268] = layer3_out[6326] ^ layer3_out[6327];
    assign layer4_out[6269] = layer3_out[2718] & layer3_out[2719];
    assign layer4_out[6270] = ~layer3_out[5551] | layer3_out[5552];
    assign layer4_out[6271] = layer3_out[2235] & layer3_out[2236];
    assign layer4_out[6272] = layer3_out[2922];
    assign layer4_out[6273] = ~(layer3_out[3319] & layer3_out[3320]);
    assign layer4_out[6274] = layer3_out[2806] & ~layer3_out[2807];
    assign layer4_out[6275] = ~(layer3_out[4206] | layer3_out[4207]);
    assign layer4_out[6276] = layer3_out[825] | layer3_out[826];
    assign layer4_out[6277] = ~layer3_out[6862] | layer3_out[6861];
    assign layer4_out[6278] = layer3_out[3413];
    assign layer4_out[6279] = ~(layer3_out[1781] & layer3_out[1782]);
    assign layer4_out[6280] = layer3_out[1637] ^ layer3_out[1638];
    assign layer4_out[6281] = layer3_out[4870] | layer3_out[4871];
    assign layer4_out[6282] = layer3_out[5044];
    assign layer4_out[6283] = layer3_out[4926];
    assign layer4_out[6284] = ~(layer3_out[4597] ^ layer3_out[4598]);
    assign layer4_out[6285] = ~(layer3_out[4785] ^ layer3_out[4786]);
    assign layer4_out[6286] = layer3_out[5564] & layer3_out[5565];
    assign layer4_out[6287] = layer3_out[3690];
    assign layer4_out[6288] = layer3_out[7025] | layer3_out[7026];
    assign layer4_out[6289] = ~(layer3_out[7998] | layer3_out[7999]);
    assign layer4_out[6290] = ~layer3_out[1958];
    assign layer4_out[6291] = ~layer3_out[5758];
    assign layer4_out[6292] = layer3_out[3895] & ~layer3_out[3896];
    assign layer4_out[6293] = ~layer3_out[7349] | layer3_out[7348];
    assign layer4_out[6294] = ~layer3_out[4461] | layer3_out[4462];
    assign layer4_out[6295] = ~layer3_out[6135] | layer3_out[6134];
    assign layer4_out[6296] = layer3_out[7710] ^ layer3_out[7711];
    assign layer4_out[6297] = ~(layer3_out[745] | layer3_out[746]);
    assign layer4_out[6298] = ~layer3_out[5944];
    assign layer4_out[6299] = ~layer3_out[7824];
    assign layer4_out[6300] = ~(layer3_out[1696] | layer3_out[1697]);
    assign layer4_out[6301] = ~layer3_out[2981];
    assign layer4_out[6302] = layer3_out[4061];
    assign layer4_out[6303] = ~(layer3_out[1252] & layer3_out[1253]);
    assign layer4_out[6304] = ~(layer3_out[1418] & layer3_out[1419]);
    assign layer4_out[6305] = layer3_out[2061];
    assign layer4_out[6306] = layer3_out[4550];
    assign layer4_out[6307] = layer3_out[25];
    assign layer4_out[6308] = layer3_out[5554] ^ layer3_out[5555];
    assign layer4_out[6309] = layer3_out[6899] ^ layer3_out[6900];
    assign layer4_out[6310] = layer3_out[1248];
    assign layer4_out[6311] = layer3_out[3177] ^ layer3_out[3178];
    assign layer4_out[6312] = layer3_out[222] & layer3_out[223];
    assign layer4_out[6313] = layer3_out[3823] ^ layer3_out[3824];
    assign layer4_out[6314] = ~layer3_out[7885];
    assign layer4_out[6315] = ~layer3_out[2681];
    assign layer4_out[6316] = layer3_out[2956] | layer3_out[2957];
    assign layer4_out[6317] = ~layer3_out[4696];
    assign layer4_out[6318] = ~layer3_out[355] | layer3_out[356];
    assign layer4_out[6319] = layer3_out[6664];
    assign layer4_out[6320] = layer3_out[6282];
    assign layer4_out[6321] = layer3_out[6473] & layer3_out[6474];
    assign layer4_out[6322] = 1'b1;
    assign layer4_out[6323] = ~(layer3_out[1140] ^ layer3_out[1141]);
    assign layer4_out[6324] = layer3_out[7650];
    assign layer4_out[6325] = layer3_out[325] ^ layer3_out[326];
    assign layer4_out[6326] = ~layer3_out[7017];
    assign layer4_out[6327] = layer3_out[7882] & ~layer3_out[7883];
    assign layer4_out[6328] = layer3_out[1470];
    assign layer4_out[6329] = layer3_out[3159];
    assign layer4_out[6330] = ~(layer3_out[2631] & layer3_out[2632]);
    assign layer4_out[6331] = layer3_out[957];
    assign layer4_out[6332] = ~layer3_out[7504];
    assign layer4_out[6333] = ~(layer3_out[5544] & layer3_out[5545]);
    assign layer4_out[6334] = ~layer3_out[250];
    assign layer4_out[6335] = layer3_out[5696];
    assign layer4_out[6336] = layer3_out[4402];
    assign layer4_out[6337] = layer3_out[599] & ~layer3_out[600];
    assign layer4_out[6338] = layer3_out[6000] & ~layer3_out[6001];
    assign layer4_out[6339] = layer3_out[3324];
    assign layer4_out[6340] = layer3_out[7306];
    assign layer4_out[6341] = layer3_out[7168] & layer3_out[7169];
    assign layer4_out[6342] = ~(layer3_out[6577] ^ layer3_out[6578]);
    assign layer4_out[6343] = ~layer3_out[2253];
    assign layer4_out[6344] = ~(layer3_out[1099] & layer3_out[1100]);
    assign layer4_out[6345] = layer3_out[3988] & layer3_out[3989];
    assign layer4_out[6346] = ~(layer3_out[5248] ^ layer3_out[5249]);
    assign layer4_out[6347] = layer3_out[6866] ^ layer3_out[6867];
    assign layer4_out[6348] = layer3_out[5755] ^ layer3_out[5756];
    assign layer4_out[6349] = layer3_out[4430] | layer3_out[4431];
    assign layer4_out[6350] = ~layer3_out[5663];
    assign layer4_out[6351] = layer3_out[5304];
    assign layer4_out[6352] = layer3_out[6030] & ~layer3_out[6029];
    assign layer4_out[6353] = ~(layer3_out[6252] | layer3_out[6253]);
    assign layer4_out[6354] = layer3_out[4203] & ~layer3_out[4202];
    assign layer4_out[6355] = layer3_out[6073];
    assign layer4_out[6356] = layer3_out[6179] & ~layer3_out[6178];
    assign layer4_out[6357] = 1'b0;
    assign layer4_out[6358] = layer3_out[86] & ~layer3_out[85];
    assign layer4_out[6359] = ~layer3_out[3486];
    assign layer4_out[6360] = layer3_out[5877] ^ layer3_out[5878];
    assign layer4_out[6361] = 1'b0;
    assign layer4_out[6362] = layer3_out[4642] & ~layer3_out[4641];
    assign layer4_out[6363] = ~layer3_out[3208] | layer3_out[3209];
    assign layer4_out[6364] = ~(layer3_out[1616] | layer3_out[1617]);
    assign layer4_out[6365] = ~(layer3_out[6293] | layer3_out[6294]);
    assign layer4_out[6366] = layer3_out[4579] ^ layer3_out[4580];
    assign layer4_out[6367] = ~layer3_out[1488];
    assign layer4_out[6368] = layer3_out[3409] & ~layer3_out[3408];
    assign layer4_out[6369] = layer3_out[3276] ^ layer3_out[3277];
    assign layer4_out[6370] = ~(layer3_out[7764] & layer3_out[7765]);
    assign layer4_out[6371] = layer3_out[3167] & ~layer3_out[3168];
    assign layer4_out[6372] = layer3_out[3740] & layer3_out[3741];
    assign layer4_out[6373] = ~layer3_out[7941];
    assign layer4_out[6374] = ~layer3_out[413];
    assign layer4_out[6375] = layer3_out[556];
    assign layer4_out[6376] = layer3_out[4544] ^ layer3_out[4545];
    assign layer4_out[6377] = ~layer3_out[644] | layer3_out[645];
    assign layer4_out[6378] = layer3_out[855];
    assign layer4_out[6379] = layer3_out[7607];
    assign layer4_out[6380] = layer3_out[6767];
    assign layer4_out[6381] = ~(layer3_out[6094] ^ layer3_out[6095]);
    assign layer4_out[6382] = ~(layer3_out[2238] ^ layer3_out[2239]);
    assign layer4_out[6383] = 1'b0;
    assign layer4_out[6384] = ~(layer3_out[3670] ^ layer3_out[3671]);
    assign layer4_out[6385] = ~layer3_out[5726];
    assign layer4_out[6386] = layer3_out[2345] | layer3_out[2346];
    assign layer4_out[6387] = ~(layer3_out[7108] & layer3_out[7109]);
    assign layer4_out[6388] = ~layer3_out[6371];
    assign layer4_out[6389] = ~(layer3_out[2982] ^ layer3_out[2983]);
    assign layer4_out[6390] = ~(layer3_out[2646] & layer3_out[2647]);
    assign layer4_out[6391] = layer3_out[5976];
    assign layer4_out[6392] = layer3_out[171] ^ layer3_out[172];
    assign layer4_out[6393] = ~layer3_out[3451];
    assign layer4_out[6394] = layer3_out[3370];
    assign layer4_out[6395] = ~(layer3_out[5250] ^ layer3_out[5251]);
    assign layer4_out[6396] = ~layer3_out[6183] | layer3_out[6184];
    assign layer4_out[6397] = layer3_out[5474] | layer3_out[5475];
    assign layer4_out[6398] = ~layer3_out[982];
    assign layer4_out[6399] = layer3_out[7003];
    assign layer4_out[6400] = layer3_out[546] ^ layer3_out[547];
    assign layer4_out[6401] = layer3_out[1551] | layer3_out[1552];
    assign layer4_out[6402] = layer3_out[6395];
    assign layer4_out[6403] = ~layer3_out[3576];
    assign layer4_out[6404] = ~layer3_out[6898] | layer3_out[6897];
    assign layer4_out[6405] = ~(layer3_out[90] | layer3_out[91]);
    assign layer4_out[6406] = ~layer3_out[4799] | layer3_out[4800];
    assign layer4_out[6407] = layer3_out[443];
    assign layer4_out[6408] = ~layer3_out[7475];
    assign layer4_out[6409] = layer3_out[142];
    assign layer4_out[6410] = layer3_out[1946] & ~layer3_out[1945];
    assign layer4_out[6411] = layer3_out[1069] & layer3_out[1070];
    assign layer4_out[6412] = layer3_out[1706] ^ layer3_out[1707];
    assign layer4_out[6413] = 1'b1;
    assign layer4_out[6414] = layer3_out[4971] ^ layer3_out[4972];
    assign layer4_out[6415] = ~(layer3_out[4060] ^ layer3_out[4061]);
    assign layer4_out[6416] = layer3_out[521];
    assign layer4_out[6417] = ~layer3_out[7501];
    assign layer4_out[6418] = ~layer3_out[6987];
    assign layer4_out[6419] = ~layer3_out[2659];
    assign layer4_out[6420] = layer3_out[4154] | layer3_out[4155];
    assign layer4_out[6421] = ~layer3_out[4447];
    assign layer4_out[6422] = ~layer3_out[1896];
    assign layer4_out[6423] = layer3_out[7518];
    assign layer4_out[6424] = ~(layer3_out[1000] & layer3_out[1001]);
    assign layer4_out[6425] = layer3_out[7914];
    assign layer4_out[6426] = ~(layer3_out[557] & layer3_out[558]);
    assign layer4_out[6427] = layer3_out[7813];
    assign layer4_out[6428] = ~layer3_out[7130] | layer3_out[7129];
    assign layer4_out[6429] = ~(layer3_out[7808] ^ layer3_out[7809]);
    assign layer4_out[6430] = layer3_out[2856];
    assign layer4_out[6431] = layer3_out[500] ^ layer3_out[501];
    assign layer4_out[6432] = ~layer3_out[806];
    assign layer4_out[6433] = ~layer3_out[3011];
    assign layer4_out[6434] = ~layer3_out[4536];
    assign layer4_out[6435] = ~layer3_out[1056];
    assign layer4_out[6436] = layer3_out[3362] | layer3_out[3363];
    assign layer4_out[6437] = ~layer3_out[4939];
    assign layer4_out[6438] = ~layer3_out[5523];
    assign layer4_out[6439] = ~(layer3_out[6264] & layer3_out[6265]);
    assign layer4_out[6440] = ~layer3_out[2764];
    assign layer4_out[6441] = layer3_out[267] ^ layer3_out[268];
    assign layer4_out[6442] = layer3_out[4500] ^ layer3_out[4501];
    assign layer4_out[6443] = layer3_out[1255];
    assign layer4_out[6444] = layer3_out[1993] | layer3_out[1994];
    assign layer4_out[6445] = ~layer3_out[6428];
    assign layer4_out[6446] = layer3_out[6652];
    assign layer4_out[6447] = ~(layer3_out[1566] | layer3_out[1567]);
    assign layer4_out[6448] = layer3_out[1924] & ~layer3_out[1925];
    assign layer4_out[6449] = layer3_out[3867] & layer3_out[3868];
    assign layer4_out[6450] = ~(layer3_out[2459] | layer3_out[2460]);
    assign layer4_out[6451] = layer3_out[5968];
    assign layer4_out[6452] = layer3_out[7536];
    assign layer4_out[6453] = ~(layer3_out[2465] ^ layer3_out[2466]);
    assign layer4_out[6454] = layer3_out[6107];
    assign layer4_out[6455] = layer3_out[635] & ~layer3_out[636];
    assign layer4_out[6456] = layer3_out[2703] & ~layer3_out[2702];
    assign layer4_out[6457] = ~(layer3_out[1852] ^ layer3_out[1853]);
    assign layer4_out[6458] = layer3_out[5769] & ~layer3_out[5768];
    assign layer4_out[6459] = layer3_out[2446] & layer3_out[2447];
    assign layer4_out[6460] = ~(layer3_out[3165] & layer3_out[3166]);
    assign layer4_out[6461] = ~(layer3_out[2699] | layer3_out[2700]);
    assign layer4_out[6462] = 1'b1;
    assign layer4_out[6463] = layer3_out[7581] & ~layer3_out[7580];
    assign layer4_out[6464] = layer3_out[7530];
    assign layer4_out[6465] = ~(layer3_out[731] & layer3_out[732]);
    assign layer4_out[6466] = ~layer3_out[1417];
    assign layer4_out[6467] = layer3_out[7658];
    assign layer4_out[6468] = layer3_out[2526] & layer3_out[2527];
    assign layer4_out[6469] = layer3_out[5810] ^ layer3_out[5811];
    assign layer4_out[6470] = layer3_out[3691] ^ layer3_out[3692];
    assign layer4_out[6471] = ~layer3_out[6147];
    assign layer4_out[6472] = layer3_out[5392] & layer3_out[5393];
    assign layer4_out[6473] = layer3_out[11];
    assign layer4_out[6474] = ~(layer3_out[6274] & layer3_out[6275]);
    assign layer4_out[6475] = layer3_out[1404] & layer3_out[1405];
    assign layer4_out[6476] = ~layer3_out[3167];
    assign layer4_out[6477] = layer3_out[3643];
    assign layer4_out[6478] = layer3_out[906];
    assign layer4_out[6479] = ~(layer3_out[2450] | layer3_out[2451]);
    assign layer4_out[6480] = ~(layer3_out[4213] ^ layer3_out[4214]);
    assign layer4_out[6481] = layer3_out[1673];
    assign layer4_out[6482] = layer3_out[7366] | layer3_out[7367];
    assign layer4_out[6483] = layer3_out[5142];
    assign layer4_out[6484] = ~(layer3_out[3340] ^ layer3_out[3341]);
    assign layer4_out[6485] = ~layer3_out[2467] | layer3_out[2466];
    assign layer4_out[6486] = layer3_out[536];
    assign layer4_out[6487] = layer3_out[5591];
    assign layer4_out[6488] = layer3_out[6930];
    assign layer4_out[6489] = layer3_out[966] & ~layer3_out[965];
    assign layer4_out[6490] = ~layer3_out[387];
    assign layer4_out[6491] = ~layer3_out[7073];
    assign layer4_out[6492] = ~(layer3_out[6034] | layer3_out[6035]);
    assign layer4_out[6493] = layer3_out[7524];
    assign layer4_out[6494] = ~layer3_out[4370];
    assign layer4_out[6495] = layer3_out[5586] & ~layer3_out[5585];
    assign layer4_out[6496] = ~layer3_out[6093];
    assign layer4_out[6497] = ~layer3_out[7611];
    assign layer4_out[6498] = layer3_out[5270] | layer3_out[5271];
    assign layer4_out[6499] = ~layer3_out[1167];
    assign layer4_out[6500] = layer3_out[964] & ~layer3_out[965];
    assign layer4_out[6501] = ~(layer3_out[1305] ^ layer3_out[1306]);
    assign layer4_out[6502] = ~layer3_out[60];
    assign layer4_out[6503] = ~layer3_out[559];
    assign layer4_out[6504] = ~(layer3_out[3395] ^ layer3_out[3396]);
    assign layer4_out[6505] = layer3_out[7727] & ~layer3_out[7728];
    assign layer4_out[6506] = ~layer3_out[4375];
    assign layer4_out[6507] = ~(layer3_out[5008] & layer3_out[5009]);
    assign layer4_out[6508] = layer3_out[4766];
    assign layer4_out[6509] = ~layer3_out[2041] | layer3_out[2040];
    assign layer4_out[6510] = layer3_out[3115];
    assign layer4_out[6511] = layer3_out[5176] | layer3_out[5177];
    assign layer4_out[6512] = ~(layer3_out[7900] ^ layer3_out[7901]);
    assign layer4_out[6513] = ~layer3_out[7737];
    assign layer4_out[6514] = ~layer3_out[5583] | layer3_out[5584];
    assign layer4_out[6515] = layer3_out[6925] ^ layer3_out[6926];
    assign layer4_out[6516] = ~(layer3_out[4367] | layer3_out[4368]);
    assign layer4_out[6517] = layer3_out[3050];
    assign layer4_out[6518] = ~layer3_out[1329];
    assign layer4_out[6519] = ~layer3_out[6590];
    assign layer4_out[6520] = layer3_out[5029] | layer3_out[5030];
    assign layer4_out[6521] = layer3_out[4258] & ~layer3_out[4259];
    assign layer4_out[6522] = layer3_out[4400] | layer3_out[4401];
    assign layer4_out[6523] = ~layer3_out[1145] | layer3_out[1146];
    assign layer4_out[6524] = layer3_out[4895] ^ layer3_out[4896];
    assign layer4_out[6525] = ~layer3_out[7167];
    assign layer4_out[6526] = layer3_out[3432];
    assign layer4_out[6527] = layer3_out[7635];
    assign layer4_out[6528] = layer3_out[3263];
    assign layer4_out[6529] = layer3_out[3544] | layer3_out[3545];
    assign layer4_out[6530] = ~layer3_out[753] | layer3_out[754];
    assign layer4_out[6531] = ~layer3_out[6977];
    assign layer4_out[6532] = layer3_out[1118];
    assign layer4_out[6533] = ~(layer3_out[6305] & layer3_out[6306]);
    assign layer4_out[6534] = ~layer3_out[4981] | layer3_out[4982];
    assign layer4_out[6535] = ~layer3_out[6295];
    assign layer4_out[6536] = ~(layer3_out[2391] & layer3_out[2392]);
    assign layer4_out[6537] = ~layer3_out[2409] | layer3_out[2408];
    assign layer4_out[6538] = ~layer3_out[4168];
    assign layer4_out[6539] = ~(layer3_out[5458] & layer3_out[5459]);
    assign layer4_out[6540] = ~(layer3_out[6387] | layer3_out[6388]);
    assign layer4_out[6541] = ~layer3_out[284];
    assign layer4_out[6542] = layer3_out[7877] ^ layer3_out[7878];
    assign layer4_out[6543] = layer3_out[5245];
    assign layer4_out[6544] = layer3_out[7953];
    assign layer4_out[6545] = ~layer3_out[3657];
    assign layer4_out[6546] = layer3_out[45];
    assign layer4_out[6547] = ~layer3_out[3849];
    assign layer4_out[6548] = ~layer3_out[4289];
    assign layer4_out[6549] = layer3_out[1020];
    assign layer4_out[6550] = ~layer3_out[7198];
    assign layer4_out[6551] = ~layer3_out[6636];
    assign layer4_out[6552] = layer3_out[7400] & ~layer3_out[7399];
    assign layer4_out[6553] = layer3_out[577];
    assign layer4_out[6554] = layer3_out[4541];
    assign layer4_out[6555] = ~layer3_out[4460] | layer3_out[4459];
    assign layer4_out[6556] = ~layer3_out[1164] | layer3_out[1165];
    assign layer4_out[6557] = layer3_out[1237];
    assign layer4_out[6558] = ~layer3_out[2845];
    assign layer4_out[6559] = layer3_out[5878];
    assign layer4_out[6560] = layer3_out[1628] & ~layer3_out[1627];
    assign layer4_out[6561] = ~layer3_out[2602];
    assign layer4_out[6562] = ~layer3_out[1916];
    assign layer4_out[6563] = ~layer3_out[5656];
    assign layer4_out[6564] = layer3_out[255];
    assign layer4_out[6565] = ~(layer3_out[722] | layer3_out[723]);
    assign layer4_out[6566] = layer3_out[2637] ^ layer3_out[2638];
    assign layer4_out[6567] = layer3_out[4254] & ~layer3_out[4255];
    assign layer4_out[6568] = layer3_out[7964] & ~layer3_out[7963];
    assign layer4_out[6569] = ~layer3_out[7769] | layer3_out[7768];
    assign layer4_out[6570] = layer3_out[5711];
    assign layer4_out[6571] = ~layer3_out[7282];
    assign layer4_out[6572] = ~layer3_out[1149];
    assign layer4_out[6573] = ~layer3_out[4918];
    assign layer4_out[6574] = layer3_out[2106] ^ layer3_out[2107];
    assign layer4_out[6575] = layer3_out[3424] | layer3_out[3425];
    assign layer4_out[6576] = ~layer3_out[3515];
    assign layer4_out[6577] = ~(layer3_out[490] ^ layer3_out[491]);
    assign layer4_out[6578] = layer3_out[6992] ^ layer3_out[6993];
    assign layer4_out[6579] = layer3_out[1949] | layer3_out[1950];
    assign layer4_out[6580] = ~layer3_out[3676] | layer3_out[3675];
    assign layer4_out[6581] = layer3_out[1699];
    assign layer4_out[6582] = ~(layer3_out[6996] ^ layer3_out[6997]);
    assign layer4_out[6583] = layer3_out[7569] & layer3_out[7570];
    assign layer4_out[6584] = ~layer3_out[5965] | layer3_out[5964];
    assign layer4_out[6585] = ~(layer3_out[3928] & layer3_out[3929]);
    assign layer4_out[6586] = layer3_out[6491] ^ layer3_out[6492];
    assign layer4_out[6587] = ~layer3_out[4379];
    assign layer4_out[6588] = ~layer3_out[3378];
    assign layer4_out[6589] = ~(layer3_out[7361] & layer3_out[7362]);
    assign layer4_out[6590] = layer3_out[6859] | layer3_out[6860];
    assign layer4_out[6591] = layer3_out[3499];
    assign layer4_out[6592] = layer3_out[7554];
    assign layer4_out[6593] = ~(layer3_out[18] & layer3_out[19]);
    assign layer4_out[6594] = layer3_out[1908] | layer3_out[1909];
    assign layer4_out[6595] = layer3_out[6996] & ~layer3_out[6995];
    assign layer4_out[6596] = ~layer3_out[7303];
    assign layer4_out[6597] = ~layer3_out[2522];
    assign layer4_out[6598] = ~layer3_out[925] | layer3_out[926];
    assign layer4_out[6599] = ~layer3_out[5999];
    assign layer4_out[6600] = layer3_out[1966] & layer3_out[1967];
    assign layer4_out[6601] = layer3_out[72];
    assign layer4_out[6602] = layer3_out[7760] & ~layer3_out[7761];
    assign layer4_out[6603] = ~(layer3_out[4532] | layer3_out[4533]);
    assign layer4_out[6604] = layer3_out[3390];
    assign layer4_out[6605] = ~(layer3_out[5431] ^ layer3_out[5432]);
    assign layer4_out[6606] = layer3_out[495];
    assign layer4_out[6607] = layer3_out[6101];
    assign layer4_out[6608] = layer3_out[2650];
    assign layer4_out[6609] = ~layer3_out[4677];
    assign layer4_out[6610] = layer3_out[4743] & layer3_out[4744];
    assign layer4_out[6611] = layer3_out[6642] ^ layer3_out[6643];
    assign layer4_out[6612] = ~layer3_out[1536];
    assign layer4_out[6613] = layer3_out[6567];
    assign layer4_out[6614] = layer3_out[2940];
    assign layer4_out[6615] = ~layer3_out[3142];
    assign layer4_out[6616] = ~layer3_out[6047] | layer3_out[6046];
    assign layer4_out[6617] = layer3_out[5649];
    assign layer4_out[6618] = ~layer3_out[1066];
    assign layer4_out[6619] = layer3_out[5242];
    assign layer4_out[6620] = ~(layer3_out[2923] & layer3_out[2924]);
    assign layer4_out[6621] = layer3_out[4363];
    assign layer4_out[6622] = ~layer3_out[4150];
    assign layer4_out[6623] = layer3_out[603] | layer3_out[604];
    assign layer4_out[6624] = ~layer3_out[861];
    assign layer4_out[6625] = ~(layer3_out[2222] | layer3_out[2223]);
    assign layer4_out[6626] = ~layer3_out[1863];
    assign layer4_out[6627] = layer3_out[2823] & ~layer3_out[2824];
    assign layer4_out[6628] = ~layer3_out[2481] | layer3_out[2482];
    assign layer4_out[6629] = layer3_out[2402] ^ layer3_out[2403];
    assign layer4_out[6630] = layer3_out[703];
    assign layer4_out[6631] = layer3_out[6313] & ~layer3_out[6314];
    assign layer4_out[6632] = ~(layer3_out[6202] ^ layer3_out[6203]);
    assign layer4_out[6633] = layer3_out[2128] & layer3_out[2129];
    assign layer4_out[6634] = layer3_out[518];
    assign layer4_out[6635] = ~(layer3_out[3470] ^ layer3_out[3471]);
    assign layer4_out[6636] = layer3_out[6417] ^ layer3_out[6418];
    assign layer4_out[6637] = layer3_out[6542] & ~layer3_out[6543];
    assign layer4_out[6638] = layer3_out[1493] & layer3_out[1494];
    assign layer4_out[6639] = layer3_out[5771];
    assign layer4_out[6640] = layer3_out[7178] | layer3_out[7179];
    assign layer4_out[6641] = ~layer3_out[2458] | layer3_out[2457];
    assign layer4_out[6642] = layer3_out[2476] & layer3_out[2477];
    assign layer4_out[6643] = ~layer3_out[3731];
    assign layer4_out[6644] = layer3_out[6158] & ~layer3_out[6159];
    assign layer4_out[6645] = layer3_out[1067];
    assign layer4_out[6646] = ~layer3_out[5782];
    assign layer4_out[6647] = ~layer3_out[2026];
    assign layer4_out[6648] = layer3_out[2735] | layer3_out[2736];
    assign layer4_out[6649] = ~layer3_out[365];
    assign layer4_out[6650] = ~(layer3_out[1732] | layer3_out[1733]);
    assign layer4_out[6651] = layer3_out[2834] & layer3_out[2835];
    assign layer4_out[6652] = layer3_out[1154];
    assign layer4_out[6653] = ~(layer3_out[7295] & layer3_out[7296]);
    assign layer4_out[6654] = layer3_out[3219] & ~layer3_out[3218];
    assign layer4_out[6655] = ~layer3_out[1806];
    assign layer4_out[6656] = ~layer3_out[2671];
    assign layer4_out[6657] = layer3_out[114];
    assign layer4_out[6658] = layer3_out[3302] ^ layer3_out[3303];
    assign layer4_out[6659] = layer3_out[5082];
    assign layer4_out[6660] = layer3_out[6195] & ~layer3_out[6196];
    assign layer4_out[6661] = layer3_out[5353] ^ layer3_out[5354];
    assign layer4_out[6662] = 1'b0;
    assign layer4_out[6663] = layer3_out[4192];
    assign layer4_out[6664] = ~(layer3_out[7788] ^ layer3_out[7789]);
    assign layer4_out[6665] = ~layer3_out[1812];
    assign layer4_out[6666] = ~layer3_out[5550] | layer3_out[5549];
    assign layer4_out[6667] = ~layer3_out[6002] | layer3_out[6001];
    assign layer4_out[6668] = ~layer3_out[3480] | layer3_out[3479];
    assign layer4_out[6669] = layer3_out[4083] ^ layer3_out[4084];
    assign layer4_out[6670] = ~(layer3_out[3761] | layer3_out[3762]);
    assign layer4_out[6671] = layer3_out[2008];
    assign layer4_out[6672] = ~(layer3_out[7160] & layer3_out[7161]);
    assign layer4_out[6673] = layer3_out[7044] ^ layer3_out[7045];
    assign layer4_out[6674] = ~(layer3_out[7762] | layer3_out[7763]);
    assign layer4_out[6675] = ~(layer3_out[5347] ^ layer3_out[5348]);
    assign layer4_out[6676] = layer3_out[6662];
    assign layer4_out[6677] = ~layer3_out[2187] | layer3_out[2186];
    assign layer4_out[6678] = ~layer3_out[980];
    assign layer4_out[6679] = ~(layer3_out[4444] | layer3_out[4445]);
    assign layer4_out[6680] = ~layer3_out[2935];
    assign layer4_out[6681] = layer3_out[5742];
    assign layer4_out[6682] = ~layer3_out[7942];
    assign layer4_out[6683] = ~(layer3_out[5084] | layer3_out[5085]);
    assign layer4_out[6684] = ~(layer3_out[4304] ^ layer3_out[4305]);
    assign layer4_out[6685] = ~layer3_out[1402];
    assign layer4_out[6686] = layer3_out[5657] & layer3_out[5658];
    assign layer4_out[6687] = layer3_out[7137] & ~layer3_out[7136];
    assign layer4_out[6688] = ~(layer3_out[6165] | layer3_out[6166]);
    assign layer4_out[6689] = ~layer3_out[3015] | layer3_out[3014];
    assign layer4_out[6690] = layer3_out[6333] & ~layer3_out[6332];
    assign layer4_out[6691] = ~(layer3_out[5684] ^ layer3_out[5685]);
    assign layer4_out[6692] = layer3_out[5235];
    assign layer4_out[6693] = ~layer3_out[6680] | layer3_out[6679];
    assign layer4_out[6694] = layer3_out[2927] & layer3_out[2928];
    assign layer4_out[6695] = ~layer3_out[4977];
    assign layer4_out[6696] = layer3_out[2775] ^ layer3_out[2776];
    assign layer4_out[6697] = ~(layer3_out[3190] | layer3_out[3191]);
    assign layer4_out[6698] = layer3_out[2909] | layer3_out[2910];
    assign layer4_out[6699] = layer3_out[7270] ^ layer3_out[7271];
    assign layer4_out[6700] = layer3_out[6907];
    assign layer4_out[6701] = ~layer3_out[5448];
    assign layer4_out[6702] = layer3_out[4427];
    assign layer4_out[6703] = ~(layer3_out[5677] & layer3_out[5678]);
    assign layer4_out[6704] = layer3_out[2423];
    assign layer4_out[6705] = layer3_out[5933] ^ layer3_out[5934];
    assign layer4_out[6706] = layer3_out[7486];
    assign layer4_out[6707] = layer3_out[1171];
    assign layer4_out[6708] = ~(layer3_out[5296] ^ layer3_out[5297]);
    assign layer4_out[6709] = ~layer3_out[987];
    assign layer4_out[6710] = 1'b0;
    assign layer4_out[6711] = layer3_out[4328] ^ layer3_out[4329];
    assign layer4_out[6712] = ~(layer3_out[7856] | layer3_out[7857]);
    assign layer4_out[6713] = layer3_out[331];
    assign layer4_out[6714] = ~layer3_out[3794] | layer3_out[3795];
    assign layer4_out[6715] = ~layer3_out[1293] | layer3_out[1292];
    assign layer4_out[6716] = layer3_out[1498] | layer3_out[1499];
    assign layer4_out[6717] = ~layer3_out[61];
    assign layer4_out[6718] = layer3_out[6721] ^ layer3_out[6722];
    assign layer4_out[6719] = ~layer3_out[3685];
    assign layer4_out[6720] = layer3_out[1703] & layer3_out[1704];
    assign layer4_out[6721] = layer3_out[7983];
    assign layer4_out[6722] = layer3_out[7148] ^ layer3_out[7149];
    assign layer4_out[6723] = ~layer3_out[3009];
    assign layer4_out[6724] = ~(layer3_out[6905] & layer3_out[6906]);
    assign layer4_out[6725] = layer3_out[399] & layer3_out[400];
    assign layer4_out[6726] = ~(layer3_out[3878] ^ layer3_out[3879]);
    assign layer4_out[6727] = ~(layer3_out[3067] & layer3_out[3068]);
    assign layer4_out[6728] = layer3_out[1085] & ~layer3_out[1084];
    assign layer4_out[6729] = ~layer3_out[2653];
    assign layer4_out[6730] = ~(layer3_out[5249] | layer3_out[5250]);
    assign layer4_out[6731] = layer3_out[4664] | layer3_out[4665];
    assign layer4_out[6732] = ~layer3_out[66];
    assign layer4_out[6733] = layer3_out[5876] & ~layer3_out[5875];
    assign layer4_out[6734] = ~layer3_out[7471];
    assign layer4_out[6735] = ~layer3_out[7755];
    assign layer4_out[6736] = ~layer3_out[5027];
    assign layer4_out[6737] = layer3_out[4085] & ~layer3_out[4084];
    assign layer4_out[6738] = ~layer3_out[776] | layer3_out[775];
    assign layer4_out[6739] = ~layer3_out[3699] | layer3_out[3700];
    assign layer4_out[6740] = ~(layer3_out[7534] | layer3_out[7535]);
    assign layer4_out[6741] = ~layer3_out[416];
    assign layer4_out[6742] = layer3_out[732] & ~layer3_out[733];
    assign layer4_out[6743] = ~layer3_out[4849] | layer3_out[4850];
    assign layer4_out[6744] = layer3_out[7667];
    assign layer4_out[6745] = layer3_out[7379] & ~layer3_out[7380];
    assign layer4_out[6746] = layer3_out[6551] & ~layer3_out[6552];
    assign layer4_out[6747] = ~(layer3_out[5202] & layer3_out[5203]);
    assign layer4_out[6748] = ~layer3_out[803];
    assign layer4_out[6749] = ~layer3_out[4999] | layer3_out[5000];
    assign layer4_out[6750] = layer3_out[1241] & layer3_out[1242];
    assign layer4_out[6751] = layer3_out[3002] & layer3_out[3003];
    assign layer4_out[6752] = layer3_out[4204];
    assign layer4_out[6753] = layer3_out[297] & ~layer3_out[296];
    assign layer4_out[6754] = layer3_out[2281];
    assign layer4_out[6755] = layer3_out[4429];
    assign layer4_out[6756] = ~layer3_out[718] | layer3_out[717];
    assign layer4_out[6757] = ~layer3_out[2296] | layer3_out[2297];
    assign layer4_out[6758] = layer3_out[648];
    assign layer4_out[6759] = layer3_out[4419];
    assign layer4_out[6760] = layer3_out[2437];
    assign layer4_out[6761] = layer3_out[7085];
    assign layer4_out[6762] = layer3_out[5406] ^ layer3_out[5407];
    assign layer4_out[6763] = ~layer3_out[6342] | layer3_out[6343];
    assign layer4_out[6764] = layer3_out[7627];
    assign layer4_out[6765] = ~layer3_out[3616];
    assign layer4_out[6766] = ~layer3_out[5834];
    assign layer4_out[6767] = ~layer3_out[1263];
    assign layer4_out[6768] = layer3_out[4433] | layer3_out[4434];
    assign layer4_out[6769] = ~(layer3_out[1918] ^ layer3_out[1919]);
    assign layer4_out[6770] = ~layer3_out[6702] | layer3_out[6701];
    assign layer4_out[6771] = 1'b1;
    assign layer4_out[6772] = ~(layer3_out[1996] | layer3_out[1997]);
    assign layer4_out[6773] = ~layer3_out[3872] | layer3_out[3873];
    assign layer4_out[6774] = layer3_out[2397];
    assign layer4_out[6775] = layer3_out[6987] ^ layer3_out[6988];
    assign layer4_out[6776] = layer3_out[7059];
    assign layer4_out[6777] = ~layer3_out[148] | layer3_out[149];
    assign layer4_out[6778] = layer3_out[7075];
    assign layer4_out[6779] = 1'b1;
    assign layer4_out[6780] = layer3_out[5999] ^ layer3_out[6000];
    assign layer4_out[6781] = ~(layer3_out[7588] | layer3_out[7589]);
    assign layer4_out[6782] = layer3_out[3559];
    assign layer4_out[6783] = layer3_out[4629];
    assign layer4_out[6784] = ~layer3_out[1742];
    assign layer4_out[6785] = layer3_out[5275];
    assign layer4_out[6786] = layer3_out[1289] ^ layer3_out[1290];
    assign layer4_out[6787] = ~layer3_out[6541];
    assign layer4_out[6788] = layer3_out[3940] ^ layer3_out[3941];
    assign layer4_out[6789] = layer3_out[7041] & layer3_out[7042];
    assign layer4_out[6790] = layer3_out[3762] ^ layer3_out[3763];
    assign layer4_out[6791] = 1'b1;
    assign layer4_out[6792] = ~layer3_out[6243];
    assign layer4_out[6793] = layer3_out[1497];
    assign layer4_out[6794] = ~layer3_out[7914] | layer3_out[7915];
    assign layer4_out[6795] = ~layer3_out[7259] | layer3_out[7258];
    assign layer4_out[6796] = ~layer3_out[4330];
    assign layer4_out[6797] = layer3_out[1389];
    assign layer4_out[6798] = layer3_out[5361];
    assign layer4_out[6799] = layer3_out[4108] ^ layer3_out[4109];
    assign layer4_out[6800] = ~layer3_out[4133] | layer3_out[4134];
    assign layer4_out[6801] = ~(layer3_out[1176] ^ layer3_out[1177]);
    assign layer4_out[6802] = ~(layer3_out[6105] ^ layer3_out[6106]);
    assign layer4_out[6803] = layer3_out[3208];
    assign layer4_out[6804] = ~(layer3_out[4977] ^ layer3_out[4978]);
    assign layer4_out[6805] = layer3_out[6210] & ~layer3_out[6211];
    assign layer4_out[6806] = layer3_out[1780] | layer3_out[1781];
    assign layer4_out[6807] = ~layer3_out[3987];
    assign layer4_out[6808] = layer3_out[4913];
    assign layer4_out[6809] = layer3_out[7517] & layer3_out[7518];
    assign layer4_out[6810] = layer3_out[1956];
    assign layer4_out[6811] = ~layer3_out[2840];
    assign layer4_out[6812] = ~(layer3_out[7784] & layer3_out[7785]);
    assign layer4_out[6813] = ~(layer3_out[3391] ^ layer3_out[3392]);
    assign layer4_out[6814] = layer3_out[730];
    assign layer4_out[6815] = layer3_out[3967];
    assign layer4_out[6816] = layer3_out[3659] & ~layer3_out[3660];
    assign layer4_out[6817] = ~(layer3_out[6809] ^ layer3_out[6810]);
    assign layer4_out[6818] = ~(layer3_out[2448] ^ layer3_out[2449]);
    assign layer4_out[6819] = ~layer3_out[5748] | layer3_out[5747];
    assign layer4_out[6820] = ~layer3_out[7691] | layer3_out[7692];
    assign layer4_out[6821] = layer3_out[4377] | layer3_out[4378];
    assign layer4_out[6822] = layer3_out[4717] & ~layer3_out[4716];
    assign layer4_out[6823] = ~layer3_out[7333];
    assign layer4_out[6824] = ~layer3_out[7755];
    assign layer4_out[6825] = layer3_out[2758] & ~layer3_out[2759];
    assign layer4_out[6826] = ~layer3_out[1543] | layer3_out[1544];
    assign layer4_out[6827] = ~layer3_out[2745];
    assign layer4_out[6828] = layer3_out[5346] ^ layer3_out[5347];
    assign layer4_out[6829] = layer3_out[3861];
    assign layer4_out[6830] = ~layer3_out[4130];
    assign layer4_out[6831] = layer3_out[3309] & ~layer3_out[3308];
    assign layer4_out[6832] = layer3_out[5267];
    assign layer4_out[6833] = layer3_out[4797];
    assign layer4_out[6834] = ~(layer3_out[6637] ^ layer3_out[6638]);
    assign layer4_out[6835] = ~(layer3_out[6083] ^ layer3_out[6084]);
    assign layer4_out[6836] = layer3_out[5408];
    assign layer4_out[6837] = ~(layer3_out[5746] ^ layer3_out[5747]);
    assign layer4_out[6838] = ~layer3_out[2677];
    assign layer4_out[6839] = ~(layer3_out[4528] ^ layer3_out[4529]);
    assign layer4_out[6840] = ~(layer3_out[727] ^ layer3_out[728]);
    assign layer4_out[6841] = ~(layer3_out[5506] | layer3_out[5507]);
    assign layer4_out[6842] = ~layer3_out[7233];
    assign layer4_out[6843] = layer3_out[2951];
    assign layer4_out[6844] = layer3_out[4970];
    assign layer4_out[6845] = ~layer3_out[1609];
    assign layer4_out[6846] = layer3_out[7133];
    assign layer4_out[6847] = ~layer3_out[4334];
    assign layer4_out[6848] = layer3_out[569] | layer3_out[570];
    assign layer4_out[6849] = layer3_out[857] ^ layer3_out[858];
    assign layer4_out[6850] = ~layer3_out[1064] | layer3_out[1065];
    assign layer4_out[6851] = ~(layer3_out[2869] | layer3_out[2870]);
    assign layer4_out[6852] = layer3_out[591] ^ layer3_out[592];
    assign layer4_out[6853] = ~layer3_out[7370];
    assign layer4_out[6854] = layer3_out[4819];
    assign layer4_out[6855] = ~layer3_out[2931];
    assign layer4_out[6856] = layer3_out[1058] | layer3_out[1059];
    assign layer4_out[6857] = ~layer3_out[6301];
    assign layer4_out[6858] = ~layer3_out[3266] | layer3_out[3265];
    assign layer4_out[6859] = layer3_out[534] ^ layer3_out[535];
    assign layer4_out[6860] = ~layer3_out[3930];
    assign layer4_out[6861] = ~(layer3_out[5800] | layer3_out[5801]);
    assign layer4_out[6862] = layer3_out[1306] ^ layer3_out[1307];
    assign layer4_out[6863] = layer3_out[4469];
    assign layer4_out[6864] = ~(layer3_out[3856] & layer3_out[3857]);
    assign layer4_out[6865] = layer3_out[5103];
    assign layer4_out[6866] = ~layer3_out[5567];
    assign layer4_out[6867] = ~(layer3_out[2892] ^ layer3_out[2893]);
    assign layer4_out[6868] = layer3_out[4015];
    assign layer4_out[6869] = layer3_out[7827] & ~layer3_out[7826];
    assign layer4_out[6870] = layer3_out[7717] & layer3_out[7718];
    assign layer4_out[6871] = ~layer3_out[1459];
    assign layer4_out[6872] = ~layer3_out[3979];
    assign layer4_out[6873] = layer3_out[3355];
    assign layer4_out[6874] = ~layer3_out[1224];
    assign layer4_out[6875] = ~layer3_out[3105];
    assign layer4_out[6876] = ~layer3_out[7261] | layer3_out[7260];
    assign layer4_out[6877] = layer3_out[5161];
    assign layer4_out[6878] = layer3_out[1285];
    assign layer4_out[6879] = layer3_out[5078] ^ layer3_out[5079];
    assign layer4_out[6880] = ~layer3_out[1769];
    assign layer4_out[6881] = 1'b0;
    assign layer4_out[6882] = layer3_out[160] ^ layer3_out[161];
    assign layer4_out[6883] = layer3_out[3422];
    assign layer4_out[6884] = layer3_out[2959];
    assign layer4_out[6885] = layer3_out[7882];
    assign layer4_out[6886] = layer3_out[7662] ^ layer3_out[7663];
    assign layer4_out[6887] = layer3_out[3150] ^ layer3_out[3151];
    assign layer4_out[6888] = ~layer3_out[4385];
    assign layer4_out[6889] = layer3_out[2736];
    assign layer4_out[6890] = layer3_out[6240] & ~layer3_out[6241];
    assign layer4_out[6891] = layer3_out[977] & ~layer3_out[976];
    assign layer4_out[6892] = layer3_out[1093];
    assign layer4_out[6893] = ~layer3_out[1588] | layer3_out[1589];
    assign layer4_out[6894] = ~layer3_out[2844];
    assign layer4_out[6895] = layer3_out[4302] | layer3_out[4303];
    assign layer4_out[6896] = layer3_out[6561] & layer3_out[6562];
    assign layer4_out[6897] = ~(layer3_out[309] ^ layer3_out[310]);
    assign layer4_out[6898] = ~layer3_out[1803];
    assign layer4_out[6899] = layer3_out[4415] ^ layer3_out[4416];
    assign layer4_out[6900] = layer3_out[3492];
    assign layer4_out[6901] = layer3_out[6564] & layer3_out[6565];
    assign layer4_out[6902] = ~layer3_out[7940];
    assign layer4_out[6903] = layer3_out[1428];
    assign layer4_out[6904] = layer3_out[2574];
    assign layer4_out[6905] = ~layer3_out[3186];
    assign layer4_out[6906] = layer3_out[7463] ^ layer3_out[7464];
    assign layer4_out[6907] = ~(layer3_out[2765] & layer3_out[2766]);
    assign layer4_out[6908] = ~(layer3_out[3812] ^ layer3_out[3813]);
    assign layer4_out[6909] = ~(layer3_out[4576] ^ layer3_out[4577]);
    assign layer4_out[6910] = layer3_out[6268];
    assign layer4_out[6911] = layer3_out[2767] & layer3_out[2768];
    assign layer4_out[6912] = ~(layer3_out[1038] | layer3_out[1039]);
    assign layer4_out[6913] = ~(layer3_out[2295] | layer3_out[2296]);
    assign layer4_out[6914] = ~layer3_out[5594] | layer3_out[5593];
    assign layer4_out[6915] = 1'b1;
    assign layer4_out[6916] = ~layer3_out[3114];
    assign layer4_out[6917] = ~layer3_out[6793] | layer3_out[6792];
    assign layer4_out[6918] = layer3_out[1846];
    assign layer4_out[6919] = layer3_out[3734] & ~layer3_out[3733];
    assign layer4_out[6920] = ~(layer3_out[3434] | layer3_out[3435]);
    assign layer4_out[6921] = ~(layer3_out[6677] | layer3_out[6678]);
    assign layer4_out[6922] = layer3_out[6037];
    assign layer4_out[6923] = ~layer3_out[394];
    assign layer4_out[6924] = layer3_out[2618];
    assign layer4_out[6925] = layer3_out[6659];
    assign layer4_out[6926] = ~(layer3_out[4709] ^ layer3_out[4710]);
    assign layer4_out[6927] = ~layer3_out[7174] | layer3_out[7173];
    assign layer4_out[6928] = ~layer3_out[2402];
    assign layer4_out[6929] = layer3_out[1441];
    assign layer4_out[6930] = ~layer3_out[311];
    assign layer4_out[6931] = ~layer3_out[4794] | layer3_out[4793];
    assign layer4_out[6932] = layer3_out[3418] & ~layer3_out[3419];
    assign layer4_out[6933] = layer3_out[2292];
    assign layer4_out[6934] = ~layer3_out[6743];
    assign layer4_out[6935] = ~layer3_out[5647];
    assign layer4_out[6936] = ~layer3_out[4690];
    assign layer4_out[6937] = ~(layer3_out[1546] | layer3_out[1547]);
    assign layer4_out[6938] = layer3_out[191];
    assign layer4_out[6939] = ~(layer3_out[5879] ^ layer3_out[5880]);
    assign layer4_out[6940] = ~(layer3_out[5304] ^ layer3_out[5305]);
    assign layer4_out[6941] = ~layer3_out[3200];
    assign layer4_out[6942] = layer3_out[3006];
    assign layer4_out[6943] = ~(layer3_out[1068] ^ layer3_out[1069]);
    assign layer4_out[6944] = ~layer3_out[6770];
    assign layer4_out[6945] = ~(layer3_out[2191] & layer3_out[2192]);
    assign layer4_out[6946] = layer3_out[2576] ^ layer3_out[2577];
    assign layer4_out[6947] = ~layer3_out[55];
    assign layer4_out[6948] = ~layer3_out[93];
    assign layer4_out[6949] = layer3_out[4722];
    assign layer4_out[6950] = ~(layer3_out[4197] ^ layer3_out[4198]);
    assign layer4_out[6951] = layer3_out[5499] & layer3_out[5500];
    assign layer4_out[6952] = ~layer3_out[3688];
    assign layer4_out[6953] = ~layer3_out[814] | layer3_out[813];
    assign layer4_out[6954] = ~layer3_out[5542];
    assign layer4_out[6955] = ~layer3_out[1849];
    assign layer4_out[6956] = layer3_out[7792];
    assign layer4_out[6957] = ~(layer3_out[5992] | layer3_out[5993]);
    assign layer4_out[6958] = layer3_out[4396] ^ layer3_out[4397];
    assign layer4_out[6959] = layer3_out[3610] | layer3_out[3611];
    assign layer4_out[6960] = ~(layer3_out[3875] | layer3_out[3876]);
    assign layer4_out[6961] = ~layer3_out[1214];
    assign layer4_out[6962] = layer3_out[3512];
    assign layer4_out[6963] = ~(layer3_out[1851] ^ layer3_out[1852]);
    assign layer4_out[6964] = layer3_out[812];
    assign layer4_out[6965] = layer3_out[2116];
    assign layer4_out[6966] = layer3_out[2840] & ~layer3_out[2841];
    assign layer4_out[6967] = layer3_out[3977] & layer3_out[3978];
    assign layer4_out[6968] = layer3_out[4353];
    assign layer4_out[6969] = ~(layer3_out[5715] | layer3_out[5716]);
    assign layer4_out[6970] = layer3_out[158];
    assign layer4_out[6971] = layer3_out[927];
    assign layer4_out[6972] = ~(layer3_out[7802] ^ layer3_out[7803]);
    assign layer4_out[6973] = layer3_out[5959] & ~layer3_out[5958];
    assign layer4_out[6974] = ~layer3_out[683];
    assign layer4_out[6975] = layer3_out[210];
    assign layer4_out[6976] = layer3_out[4646];
    assign layer4_out[6977] = ~layer3_out[2743];
    assign layer4_out[6978] = ~layer3_out[1679] | layer3_out[1680];
    assign layer4_out[6979] = ~layer3_out[2167] | layer3_out[2168];
    assign layer4_out[6980] = layer3_out[207];
    assign layer4_out[6981] = ~layer3_out[3754] | layer3_out[3755];
    assign layer4_out[6982] = ~layer3_out[1253] | layer3_out[1254];
    assign layer4_out[6983] = ~layer3_out[4521];
    assign layer4_out[6984] = ~layer3_out[4193];
    assign layer4_out[6985] = layer3_out[3478] & ~layer3_out[3479];
    assign layer4_out[6986] = ~(layer3_out[2664] ^ layer3_out[2665]);
    assign layer4_out[6987] = ~layer3_out[6168];
    assign layer4_out[6988] = ~layer3_out[6857];
    assign layer4_out[6989] = ~layer3_out[4190];
    assign layer4_out[6990] = layer3_out[2324] ^ layer3_out[2325];
    assign layer4_out[6991] = layer3_out[2350] | layer3_out[2351];
    assign layer4_out[6992] = ~(layer3_out[3271] & layer3_out[3272]);
    assign layer4_out[6993] = layer3_out[5051] & layer3_out[5052];
    assign layer4_out[6994] = ~(layer3_out[2494] & layer3_out[2495]);
    assign layer4_out[6995] = ~layer3_out[2302];
    assign layer4_out[6996] = layer3_out[1072];
    assign layer4_out[6997] = layer3_out[507];
    assign layer4_out[6998] = ~layer3_out[2214];
    assign layer4_out[6999] = layer3_out[6097];
    assign layer4_out[7000] = ~(layer3_out[695] ^ layer3_out[696]);
    assign layer4_out[7001] = layer3_out[5633];
    assign layer4_out[7002] = layer3_out[1159];
    assign layer4_out[7003] = ~(layer3_out[318] ^ layer3_out[319]);
    assign layer4_out[7004] = layer3_out[2893] ^ layer3_out[2894];
    assign layer4_out[7005] = ~(layer3_out[3201] ^ layer3_out[3202]);
    assign layer4_out[7006] = layer3_out[309];
    assign layer4_out[7007] = ~(layer3_out[2907] | layer3_out[2908]);
    assign layer4_out[7008] = layer3_out[7088];
    assign layer4_out[7009] = layer3_out[591];
    assign layer4_out[7010] = ~layer3_out[6929];
    assign layer4_out[7011] = ~layer3_out[1652] | layer3_out[1651];
    assign layer4_out[7012] = ~layer3_out[1866];
    assign layer4_out[7013] = layer3_out[1844];
    assign layer4_out[7014] = layer3_out[6556] & ~layer3_out[6557];
    assign layer4_out[7015] = layer3_out[2767] & ~layer3_out[2766];
    assign layer4_out[7016] = layer3_out[2473];
    assign layer4_out[7017] = ~(layer3_out[2774] & layer3_out[2775]);
    assign layer4_out[7018] = layer3_out[4313] & layer3_out[4314];
    assign layer4_out[7019] = ~(layer3_out[2764] | layer3_out[2765]);
    assign layer4_out[7020] = layer3_out[6159];
    assign layer4_out[7021] = layer3_out[5356] ^ layer3_out[5357];
    assign layer4_out[7022] = ~layer3_out[3669] | layer3_out[3670];
    assign layer4_out[7023] = layer3_out[6590];
    assign layer4_out[7024] = ~layer3_out[1193];
    assign layer4_out[7025] = layer3_out[7418];
    assign layer4_out[7026] = ~(layer3_out[1593] & layer3_out[1594]);
    assign layer4_out[7027] = layer3_out[841] & ~layer3_out[840];
    assign layer4_out[7028] = ~(layer3_out[7460] | layer3_out[7461]);
    assign layer4_out[7029] = ~(layer3_out[1390] ^ layer3_out[1391]);
    assign layer4_out[7030] = ~layer3_out[6585];
    assign layer4_out[7031] = layer3_out[5728];
    assign layer4_out[7032] = ~layer3_out[6513];
    assign layer4_out[7033] = ~(layer3_out[3804] | layer3_out[3805]);
    assign layer4_out[7034] = layer3_out[7816] & ~layer3_out[7817];
    assign layer4_out[7035] = layer3_out[7495] & layer3_out[7496];
    assign layer4_out[7036] = layer3_out[3703] | layer3_out[3704];
    assign layer4_out[7037] = ~layer3_out[7113];
    assign layer4_out[7038] = layer3_out[106];
    assign layer4_out[7039] = layer3_out[1918];
    assign layer4_out[7040] = ~(layer3_out[6345] | layer3_out[6346]);
    assign layer4_out[7041] = layer3_out[5151] & layer3_out[5152];
    assign layer4_out[7042] = ~layer3_out[4169];
    assign layer4_out[7043] = layer3_out[6434] | layer3_out[6435];
    assign layer4_out[7044] = layer3_out[3039] | layer3_out[3040];
    assign layer4_out[7045] = layer3_out[1603] & ~layer3_out[1602];
    assign layer4_out[7046] = ~layer3_out[4777];
    assign layer4_out[7047] = layer3_out[4261];
    assign layer4_out[7048] = layer3_out[5440] & ~layer3_out[5441];
    assign layer4_out[7049] = ~layer3_out[6386];
    assign layer4_out[7050] = layer3_out[4651] | layer3_out[4652];
    assign layer4_out[7051] = ~(layer3_out[6640] & layer3_out[6641]);
    assign layer4_out[7052] = ~layer3_out[3778];
    assign layer4_out[7053] = ~layer3_out[6765];
    assign layer4_out[7054] = ~(layer3_out[4806] | layer3_out[4807]);
    assign layer4_out[7055] = ~(layer3_out[1422] & layer3_out[1423]);
    assign layer4_out[7056] = ~(layer3_out[5027] | layer3_out[5028]);
    assign layer4_out[7057] = ~(layer3_out[2597] ^ layer3_out[2598]);
    assign layer4_out[7058] = layer3_out[4962];
    assign layer4_out[7059] = ~(layer3_out[7972] & layer3_out[7973]);
    assign layer4_out[7060] = layer3_out[3039];
    assign layer4_out[7061] = ~layer3_out[3330] | layer3_out[3331];
    assign layer4_out[7062] = layer3_out[1926];
    assign layer4_out[7063] = ~(layer3_out[3372] | layer3_out[3373]);
    assign layer4_out[7064] = ~(layer3_out[2838] ^ layer3_out[2839]);
    assign layer4_out[7065] = layer3_out[3657] ^ layer3_out[3658];
    assign layer4_out[7066] = ~layer3_out[2136] | layer3_out[2137];
    assign layer4_out[7067] = ~(layer3_out[7811] & layer3_out[7812]);
    assign layer4_out[7068] = layer3_out[3933] & ~layer3_out[3932];
    assign layer4_out[7069] = ~layer3_out[2987];
    assign layer4_out[7070] = ~layer3_out[4443];
    assign layer4_out[7071] = ~(layer3_out[5822] ^ layer3_out[5823]);
    assign layer4_out[7072] = ~layer3_out[5363] | layer3_out[5362];
    assign layer4_out[7073] = layer3_out[1620] & ~layer3_out[1619];
    assign layer4_out[7074] = ~layer3_out[6800] | layer3_out[6801];
    assign layer4_out[7075] = ~(layer3_out[4027] ^ layer3_out[4028]);
    assign layer4_out[7076] = ~layer3_out[3097] | layer3_out[3098];
    assign layer4_out[7077] = layer3_out[1931] | layer3_out[1932];
    assign layer4_out[7078] = ~(layer3_out[5673] ^ layer3_out[5674]);
    assign layer4_out[7079] = 1'b1;
    assign layer4_out[7080] = ~(layer3_out[4116] ^ layer3_out[4117]);
    assign layer4_out[7081] = ~layer3_out[5775];
    assign layer4_out[7082] = ~layer3_out[1276];
    assign layer4_out[7083] = ~layer3_out[873] | layer3_out[872];
    assign layer4_out[7084] = layer3_out[4530];
    assign layer4_out[7085] = layer3_out[5631] | layer3_out[5632];
    assign layer4_out[7086] = layer3_out[3220] ^ layer3_out[3221];
    assign layer4_out[7087] = ~layer3_out[6068] | layer3_out[6069];
    assign layer4_out[7088] = layer3_out[2723] & ~layer3_out[2722];
    assign layer4_out[7089] = layer3_out[1151];
    assign layer4_out[7090] = ~(layer3_out[4087] & layer3_out[4088]);
    assign layer4_out[7091] = ~layer3_out[197];
    assign layer4_out[7092] = layer3_out[7910] ^ layer3_out[7911];
    assign layer4_out[7093] = ~layer3_out[2502];
    assign layer4_out[7094] = layer3_out[7840] ^ layer3_out[7841];
    assign layer4_out[7095] = ~layer3_out[1761];
    assign layer4_out[7096] = layer3_out[5307] & layer3_out[5308];
    assign layer4_out[7097] = layer3_out[2611];
    assign layer4_out[7098] = ~(layer3_out[5455] ^ layer3_out[5456]);
    assign layer4_out[7099] = layer3_out[7331] ^ layer3_out[7332];
    assign layer4_out[7100] = ~(layer3_out[1919] ^ layer3_out[1920]);
    assign layer4_out[7101] = ~layer3_out[3021];
    assign layer4_out[7102] = ~layer3_out[5901];
    assign layer4_out[7103] = layer3_out[7944];
    assign layer4_out[7104] = ~layer3_out[3233];
    assign layer4_out[7105] = ~(layer3_out[4694] & layer3_out[4695]);
    assign layer4_out[7106] = layer3_out[2867];
    assign layer4_out[7107] = layer3_out[7499] ^ layer3_out[7500];
    assign layer4_out[7108] = layer3_out[6813] ^ layer3_out[6814];
    assign layer4_out[7109] = layer3_out[6132];
    assign layer4_out[7110] = ~layer3_out[7688] | layer3_out[7689];
    assign layer4_out[7111] = ~(layer3_out[2715] ^ layer3_out[2716]);
    assign layer4_out[7112] = ~layer3_out[7920] | layer3_out[7919];
    assign layer4_out[7113] = layer3_out[4315] | layer3_out[4316];
    assign layer4_out[7114] = ~layer3_out[2559];
    assign layer4_out[7115] = layer3_out[7239] & layer3_out[7240];
    assign layer4_out[7116] = ~layer3_out[5723] | layer3_out[5722];
    assign layer4_out[7117] = layer3_out[7943];
    assign layer4_out[7118] = ~(layer3_out[545] & layer3_out[546]);
    assign layer4_out[7119] = ~layer3_out[804];
    assign layer4_out[7120] = ~(layer3_out[5355] | layer3_out[5356]);
    assign layer4_out[7121] = ~layer3_out[2032];
    assign layer4_out[7122] = layer3_out[7064];
    assign layer4_out[7123] = layer3_out[7978];
    assign layer4_out[7124] = layer3_out[520] ^ layer3_out[521];
    assign layer4_out[7125] = layer3_out[1776] ^ layer3_out[1777];
    assign layer4_out[7126] = ~(layer3_out[686] ^ layer3_out[687]);
    assign layer4_out[7127] = ~layer3_out[5920];
    assign layer4_out[7128] = ~(layer3_out[5955] & layer3_out[5956]);
    assign layer4_out[7129] = layer3_out[3337];
    assign layer4_out[7130] = ~(layer3_out[4285] | layer3_out[4286]);
    assign layer4_out[7131] = ~layer3_out[5904] | layer3_out[5903];
    assign layer4_out[7132] = layer3_out[3820] & ~layer3_out[3819];
    assign layer4_out[7133] = layer3_out[6785];
    assign layer4_out[7134] = ~(layer3_out[4112] & layer3_out[4113]);
    assign layer4_out[7135] = ~(layer3_out[2780] ^ layer3_out[2781]);
    assign layer4_out[7136] = ~layer3_out[7029];
    assign layer4_out[7137] = ~(layer3_out[4165] | layer3_out[4166]);
    assign layer4_out[7138] = layer3_out[289] & layer3_out[290];
    assign layer4_out[7139] = ~(layer3_out[484] ^ layer3_out[485]);
    assign layer4_out[7140] = layer3_out[3031];
    assign layer4_out[7141] = ~layer3_out[3349];
    assign layer4_out[7142] = layer3_out[2293] & ~layer3_out[2294];
    assign layer4_out[7143] = ~(layer3_out[3972] ^ layer3_out[3973]);
    assign layer4_out[7144] = ~(layer3_out[2792] ^ layer3_out[2793]);
    assign layer4_out[7145] = ~layer3_out[7174];
    assign layer4_out[7146] = layer3_out[5312] ^ layer3_out[5313];
    assign layer4_out[7147] = ~layer3_out[6639];
    assign layer4_out[7148] = ~layer3_out[5119];
    assign layer4_out[7149] = layer3_out[4813] & ~layer3_out[4814];
    assign layer4_out[7150] = layer3_out[3381] & ~layer3_out[3380];
    assign layer4_out[7151] = layer3_out[1655] & ~layer3_out[1654];
    assign layer4_out[7152] = ~layer3_out[3713];
    assign layer4_out[7153] = layer3_out[468];
    assign layer4_out[7154] = ~layer3_out[3442];
    assign layer4_out[7155] = ~layer3_out[5784];
    assign layer4_out[7156] = ~layer3_out[4791];
    assign layer4_out[7157] = layer3_out[2007] & ~layer3_out[2008];
    assign layer4_out[7158] = layer3_out[4362] | layer3_out[4363];
    assign layer4_out[7159] = layer3_out[5107] & ~layer3_out[5108];
    assign layer4_out[7160] = ~(layer3_out[4149] ^ layer3_out[4150]);
    assign layer4_out[7161] = ~layer3_out[245];
    assign layer4_out[7162] = layer3_out[5681] & ~layer3_out[5682];
    assign layer4_out[7163] = layer3_out[519] & ~layer3_out[518];
    assign layer4_out[7164] = layer3_out[2750];
    assign layer4_out[7165] = ~layer3_out[3857];
    assign layer4_out[7166] = layer3_out[5125] & ~layer3_out[5124];
    assign layer4_out[7167] = ~(layer3_out[7128] ^ layer3_out[7129]);
    assign layer4_out[7168] = layer3_out[2086];
    assign layer4_out[7169] = layer3_out[1395] & layer3_out[1396];
    assign layer4_out[7170] = ~(layer3_out[4699] & layer3_out[4700]);
    assign layer4_out[7171] = ~(layer3_out[3721] | layer3_out[3722]);
    assign layer4_out[7172] = ~(layer3_out[2241] ^ layer3_out[2242]);
    assign layer4_out[7173] = ~(layer3_out[3555] ^ layer3_out[3556]);
    assign layer4_out[7174] = ~layer3_out[2776] | layer3_out[2777];
    assign layer4_out[7175] = ~layer3_out[2954];
    assign layer4_out[7176] = ~(layer3_out[1974] | layer3_out[1975]);
    assign layer4_out[7177] = ~(layer3_out[2880] | layer3_out[2881]);
    assign layer4_out[7178] = layer3_out[1946] | layer3_out[1947];
    assign layer4_out[7179] = layer3_out[5229];
    assign layer4_out[7180] = layer3_out[4960];
    assign layer4_out[7181] = layer3_out[4583] ^ layer3_out[4584];
    assign layer4_out[7182] = ~layer3_out[6003];
    assign layer4_out[7183] = layer3_out[3318] & layer3_out[3319];
    assign layer4_out[7184] = layer3_out[6846] & ~layer3_out[6845];
    assign layer4_out[7185] = layer3_out[2606];
    assign layer4_out[7186] = ~(layer3_out[3480] & layer3_out[3481]);
    assign layer4_out[7187] = layer3_out[1915];
    assign layer4_out[7188] = layer3_out[3341] & ~layer3_out[3342];
    assign layer4_out[7189] = layer3_out[5306] & ~layer3_out[5305];
    assign layer4_out[7190] = layer3_out[3917] & ~layer3_out[3916];
    assign layer4_out[7191] = layer3_out[6573] & layer3_out[6574];
    assign layer4_out[7192] = layer3_out[6654] ^ layer3_out[6655];
    assign layer4_out[7193] = ~layer3_out[3071] | layer3_out[3070];
    assign layer4_out[7194] = ~(layer3_out[2299] | layer3_out[2300]);
    assign layer4_out[7195] = layer3_out[6177] | layer3_out[6178];
    assign layer4_out[7196] = ~layer3_out[3594];
    assign layer4_out[7197] = ~layer3_out[5481];
    assign layer4_out[7198] = ~layer3_out[6487] | layer3_out[6488];
    assign layer4_out[7199] = layer3_out[1333];
    assign layer4_out[7200] = layer3_out[6510];
    assign layer4_out[7201] = ~layer3_out[3075] | layer3_out[3074];
    assign layer4_out[7202] = ~layer3_out[6157];
    assign layer4_out[7203] = layer3_out[932];
    assign layer4_out[7204] = layer3_out[4535] | layer3_out[4536];
    assign layer4_out[7205] = ~(layer3_out[2179] | layer3_out[2180]);
    assign layer4_out[7206] = ~layer3_out[6705] | layer3_out[6704];
    assign layer4_out[7207] = layer3_out[7876] ^ layer3_out[7877];
    assign layer4_out[7208] = ~layer3_out[2965];
    assign layer4_out[7209] = ~(layer3_out[7930] | layer3_out[7931]);
    assign layer4_out[7210] = layer3_out[4527] ^ layer3_out[4528];
    assign layer4_out[7211] = layer3_out[7926] | layer3_out[7927];
    assign layer4_out[7212] = layer3_out[3329];
    assign layer4_out[7213] = layer3_out[7555] ^ layer3_out[7556];
    assign layer4_out[7214] = layer3_out[4136] ^ layer3_out[4137];
    assign layer4_out[7215] = layer3_out[4295] | layer3_out[4296];
    assign layer4_out[7216] = ~layer3_out[1195];
    assign layer4_out[7217] = layer3_out[5987] | layer3_out[5988];
    assign layer4_out[7218] = layer3_out[1321];
    assign layer4_out[7219] = ~layer3_out[1650];
    assign layer4_out[7220] = layer3_out[1002] ^ layer3_out[1003];
    assign layer4_out[7221] = layer3_out[4727] ^ layer3_out[4728];
    assign layer4_out[7222] = ~(layer3_out[2482] | layer3_out[2483]);
    assign layer4_out[7223] = ~(layer3_out[3585] ^ layer3_out[3586]);
    assign layer4_out[7224] = layer3_out[3864] & ~layer3_out[3863];
    assign layer4_out[7225] = layer3_out[5004];
    assign layer4_out[7226] = ~(layer3_out[7023] ^ layer3_out[7024]);
    assign layer4_out[7227] = layer3_out[6400];
    assign layer4_out[7228] = layer3_out[7348] & ~layer3_out[7347];
    assign layer4_out[7229] = layer3_out[519] & layer3_out[520];
    assign layer4_out[7230] = layer3_out[3580] & layer3_out[3581];
    assign layer4_out[7231] = ~layer3_out[2116] | layer3_out[2117];
    assign layer4_out[7232] = ~(layer3_out[5668] | layer3_out[5669]);
    assign layer4_out[7233] = layer3_out[2298] | layer3_out[2299];
    assign layer4_out[7234] = ~layer3_out[5873];
    assign layer4_out[7235] = layer3_out[4936];
    assign layer4_out[7236] = layer3_out[3773];
    assign layer4_out[7237] = ~layer3_out[2728] | layer3_out[2727];
    assign layer4_out[7238] = ~(layer3_out[7843] | layer3_out[7844]);
    assign layer4_out[7239] = layer3_out[7549] ^ layer3_out[7550];
    assign layer4_out[7240] = layer3_out[4853] | layer3_out[4854];
    assign layer4_out[7241] = ~(layer3_out[2542] ^ layer3_out[2543]);
    assign layer4_out[7242] = layer3_out[2367];
    assign layer4_out[7243] = layer3_out[4063];
    assign layer4_out[7244] = layer3_out[7526];
    assign layer4_out[7245] = layer3_out[1271];
    assign layer4_out[7246] = ~layer3_out[6539] | layer3_out[6540];
    assign layer4_out[7247] = layer3_out[5186];
    assign layer4_out[7248] = ~layer3_out[3055];
    assign layer4_out[7249] = ~layer3_out[918];
    assign layer4_out[7250] = ~(layer3_out[5967] & layer3_out[5968]);
    assign layer4_out[7251] = layer3_out[5710] | layer3_out[5711];
    assign layer4_out[7252] = ~(layer3_out[4324] ^ layer3_out[4325]);
    assign layer4_out[7253] = ~(layer3_out[715] ^ layer3_out[716]);
    assign layer4_out[7254] = layer3_out[3102] & ~layer3_out[3103];
    assign layer4_out[7255] = layer3_out[7702] ^ layer3_out[7703];
    assign layer4_out[7256] = layer3_out[3297];
    assign layer4_out[7257] = ~layer3_out[6714] | layer3_out[6715];
    assign layer4_out[7258] = layer3_out[3719] ^ layer3_out[3720];
    assign layer4_out[7259] = ~layer3_out[2719];
    assign layer4_out[7260] = ~layer3_out[26];
    assign layer4_out[7261] = layer3_out[6997] ^ layer3_out[6998];
    assign layer4_out[7262] = layer3_out[37];
    assign layer4_out[7263] = layer3_out[3204] & ~layer3_out[3203];
    assign layer4_out[7264] = layer3_out[1482];
    assign layer4_out[7265] = ~layer3_out[3982] | layer3_out[3981];
    assign layer4_out[7266] = layer3_out[5112] ^ layer3_out[5113];
    assign layer4_out[7267] = ~(layer3_out[5315] & layer3_out[5316]);
    assign layer4_out[7268] = ~(layer3_out[2963] ^ layer3_out[2964]);
    assign layer4_out[7269] = layer3_out[4495] ^ layer3_out[4496];
    assign layer4_out[7270] = ~layer3_out[6916] | layer3_out[6915];
    assign layer4_out[7271] = layer3_out[3070];
    assign layer4_out[7272] = ~layer3_out[1683] | layer3_out[1684];
    assign layer4_out[7273] = layer3_out[7492] ^ layer3_out[7493];
    assign layer4_out[7274] = layer3_out[6358];
    assign layer4_out[7275] = ~layer3_out[5687];
    assign layer4_out[7276] = layer3_out[4702];
    assign layer4_out[7277] = ~(layer3_out[1288] & layer3_out[1289]);
    assign layer4_out[7278] = ~(layer3_out[3233] & layer3_out[3234]);
    assign layer4_out[7279] = ~(layer3_out[2683] ^ layer3_out[2684]);
    assign layer4_out[7280] = layer3_out[7181] & layer3_out[7182];
    assign layer4_out[7281] = layer3_out[7150] & layer3_out[7151];
    assign layer4_out[7282] = ~layer3_out[3161];
    assign layer4_out[7283] = ~(layer3_out[2973] | layer3_out[2974]);
    assign layer4_out[7284] = layer3_out[5221] ^ layer3_out[5222];
    assign layer4_out[7285] = ~layer3_out[2222] | layer3_out[2221];
    assign layer4_out[7286] = ~layer3_out[698];
    assign layer4_out[7287] = ~layer3_out[2233];
    assign layer4_out[7288] = ~layer3_out[1601];
    assign layer4_out[7289] = ~layer3_out[2261];
    assign layer4_out[7290] = layer3_out[466] & layer3_out[467];
    assign layer4_out[7291] = layer3_out[3732];
    assign layer4_out[7292] = layer3_out[7861] | layer3_out[7862];
    assign layer4_out[7293] = layer3_out[7875];
    assign layer4_out[7294] = ~layer3_out[5461] | layer3_out[5462];
    assign layer4_out[7295] = ~(layer3_out[6341] ^ layer3_out[6342]);
    assign layer4_out[7296] = layer3_out[2554] | layer3_out[2555];
    assign layer4_out[7297] = layer3_out[6423] | layer3_out[6424];
    assign layer4_out[7298] = ~layer3_out[5652] | layer3_out[5653];
    assign layer4_out[7299] = ~layer3_out[2791] | layer3_out[2792];
    assign layer4_out[7300] = layer3_out[3625] & layer3_out[3626];
    assign layer4_out[7301] = ~layer3_out[3082];
    assign layer4_out[7302] = ~(layer3_out[6271] & layer3_out[6272]);
    assign layer4_out[7303] = layer3_out[3339] & layer3_out[3340];
    assign layer4_out[7304] = layer3_out[5162];
    assign layer4_out[7305] = ~(layer3_out[5646] ^ layer3_out[5647]);
    assign layer4_out[7306] = layer3_out[389];
    assign layer4_out[7307] = layer3_out[1654];
    assign layer4_out[7308] = ~(layer3_out[3180] | layer3_out[3181]);
    assign layer4_out[7309] = layer3_out[4264];
    assign layer4_out[7310] = layer3_out[145] ^ layer3_out[146];
    assign layer4_out[7311] = ~layer3_out[3235] | layer3_out[3234];
    assign layer4_out[7312] = layer3_out[4654] ^ layer3_out[4655];
    assign layer4_out[7313] = ~(layer3_out[5527] & layer3_out[5528]);
    assign layer4_out[7314] = layer3_out[3846];
    assign layer4_out[7315] = layer3_out[6822] & layer3_out[6823];
    assign layer4_out[7316] = layer3_out[953] & ~layer3_out[952];
    assign layer4_out[7317] = layer3_out[5340] | layer3_out[5341];
    assign layer4_out[7318] = layer3_out[97] & layer3_out[98];
    assign layer4_out[7319] = ~(layer3_out[975] ^ layer3_out[976]);
    assign layer4_out[7320] = layer3_out[3760] | layer3_out[3761];
    assign layer4_out[7321] = ~layer3_out[7720];
    assign layer4_out[7322] = layer3_out[4283] | layer3_out[4284];
    assign layer4_out[7323] = ~(layer3_out[1322] & layer3_out[1323]);
    assign layer4_out[7324] = layer3_out[6568] | layer3_out[6569];
    assign layer4_out[7325] = ~(layer3_out[1009] & layer3_out[1010]);
    assign layer4_out[7326] = ~(layer3_out[2215] ^ layer3_out[2216]);
    assign layer4_out[7327] = ~(layer3_out[1988] | layer3_out[1989]);
    assign layer4_out[7328] = ~(layer3_out[1118] ^ layer3_out[1119]);
    assign layer4_out[7329] = ~layer3_out[483];
    assign layer4_out[7330] = layer3_out[5303];
    assign layer4_out[7331] = layer3_out[5255];
    assign layer4_out[7332] = ~layer3_out[1021];
    assign layer4_out[7333] = ~(layer3_out[6012] ^ layer3_out[6013]);
    assign layer4_out[7334] = ~layer3_out[7574];
    assign layer4_out[7335] = ~(layer3_out[6606] & layer3_out[6607]);
    assign layer4_out[7336] = ~layer3_out[7904] | layer3_out[7903];
    assign layer4_out[7337] = layer3_out[6067];
    assign layer4_out[7338] = ~layer3_out[2364] | layer3_out[2365];
    assign layer4_out[7339] = layer3_out[6363];
    assign layer4_out[7340] = layer3_out[1942] | layer3_out[1943];
    assign layer4_out[7341] = layer3_out[7595];
    assign layer4_out[7342] = layer3_out[2552];
    assign layer4_out[7343] = ~(layer3_out[5614] & layer3_out[5615]);
    assign layer4_out[7344] = ~layer3_out[7190];
    assign layer4_out[7345] = ~layer3_out[4123] | layer3_out[4124];
    assign layer4_out[7346] = layer3_out[4952] | layer3_out[4953];
    assign layer4_out[7347] = layer3_out[5740] & ~layer3_out[5739];
    assign layer4_out[7348] = ~layer3_out[792];
    assign layer4_out[7349] = layer3_out[23];
    assign layer4_out[7350] = layer3_out[5796] | layer3_out[5797];
    assign layer4_out[7351] = ~layer3_out[1827];
    assign layer4_out[7352] = layer3_out[7250] | layer3_out[7251];
    assign layer4_out[7353] = ~layer3_out[4417];
    assign layer4_out[7354] = ~(layer3_out[414] ^ layer3_out[415]);
    assign layer4_out[7355] = ~(layer3_out[378] & layer3_out[379]);
    assign layer4_out[7356] = ~(layer3_out[4335] ^ layer3_out[4336]);
    assign layer4_out[7357] = ~(layer3_out[5367] & layer3_out[5368]);
    assign layer4_out[7358] = ~(layer3_out[1430] | layer3_out[1431]);
    assign layer4_out[7359] = ~layer3_out[7741] | layer3_out[7740];
    assign layer4_out[7360] = layer3_out[944] & layer3_out[945];
    assign layer4_out[7361] = ~layer3_out[1584];
    assign layer4_out[7362] = ~layer3_out[647];
    assign layer4_out[7363] = layer3_out[1299] ^ layer3_out[1300];
    assign layer4_out[7364] = ~(layer3_out[53] ^ layer3_out[54]);
    assign layer4_out[7365] = layer3_out[1486] & ~layer3_out[1485];
    assign layer4_out[7366] = layer3_out[304] ^ layer3_out[305];
    assign layer4_out[7367] = ~(layer3_out[1854] | layer3_out[1855]);
    assign layer4_out[7368] = ~layer3_out[6959];
    assign layer4_out[7369] = layer3_out[1004] & ~layer3_out[1005];
    assign layer4_out[7370] = layer3_out[2478] ^ layer3_out[2479];
    assign layer4_out[7371] = layer3_out[7263];
    assign layer4_out[7372] = ~layer3_out[3636] | layer3_out[3637];
    assign layer4_out[7373] = ~layer3_out[5977] | layer3_out[5976];
    assign layer4_out[7374] = ~(layer3_out[104] | layer3_out[105]);
    assign layer4_out[7375] = ~layer3_out[6979] | layer3_out[6980];
    assign layer4_out[7376] = ~layer3_out[2710];
    assign layer4_out[7377] = ~(layer3_out[4534] & layer3_out[4535]);
    assign layer4_out[7378] = ~(layer3_out[3071] ^ layer3_out[3072]);
    assign layer4_out[7379] = ~layer3_out[4783];
    assign layer4_out[7380] = layer3_out[3545] ^ layer3_out[3546];
    assign layer4_out[7381] = ~layer3_out[1611] | layer3_out[1610];
    assign layer4_out[7382] = layer3_out[2828];
    assign layer4_out[7383] = ~layer3_out[7985];
    assign layer4_out[7384] = layer3_out[7846];
    assign layer4_out[7385] = layer3_out[6616] & ~layer3_out[6615];
    assign layer4_out[7386] = layer3_out[7751];
    assign layer4_out[7387] = ~layer3_out[3000];
    assign layer4_out[7388] = layer3_out[4505] & layer3_out[4506];
    assign layer4_out[7389] = ~(layer3_out[7532] | layer3_out[7533]);
    assign layer4_out[7390] = ~(layer3_out[2713] ^ layer3_out[2714]);
    assign layer4_out[7391] = layer3_out[4513] | layer3_out[4514];
    assign layer4_out[7392] = layer3_out[6476] & layer3_out[6477];
    assign layer4_out[7393] = ~layer3_out[5442];
    assign layer4_out[7394] = ~(layer3_out[4763] ^ layer3_out[4764]);
    assign layer4_out[7395] = ~(layer3_out[23] ^ layer3_out[24]);
    assign layer4_out[7396] = layer3_out[6325] ^ layer3_out[6326];
    assign layer4_out[7397] = layer3_out[6080] ^ layer3_out[6081];
    assign layer4_out[7398] = ~layer3_out[5974];
    assign layer4_out[7399] = ~(layer3_out[7058] | layer3_out[7059]);
    assign layer4_out[7400] = layer3_out[2925];
    assign layer4_out[7401] = ~layer3_out[954];
    assign layer4_out[7402] = layer3_out[4414] & layer3_out[4415];
    assign layer4_out[7403] = layer3_out[7224] | layer3_out[7225];
    assign layer4_out[7404] = ~(layer3_out[1660] & layer3_out[1661]);
    assign layer4_out[7405] = layer3_out[2169];
    assign layer4_out[7406] = ~(layer3_out[2779] | layer3_out[2780]);
    assign layer4_out[7407] = ~(layer3_out[4356] ^ layer3_out[4357]);
    assign layer4_out[7408] = layer3_out[3861];
    assign layer4_out[7409] = ~layer3_out[2896] | layer3_out[2895];
    assign layer4_out[7410] = ~(layer3_out[2610] & layer3_out[2611]);
    assign layer4_out[7411] = ~layer3_out[3596] | layer3_out[3597];
    assign layer4_out[7412] = layer3_out[465] & layer3_out[466];
    assign layer4_out[7413] = layer3_out[2552];
    assign layer4_out[7414] = ~layer3_out[657];
    assign layer4_out[7415] = layer3_out[6745];
    assign layer4_out[7416] = layer3_out[5095] & ~layer3_out[5094];
    assign layer4_out[7417] = layer3_out[1265] & layer3_out[1266];
    assign layer4_out[7418] = ~layer3_out[5524];
    assign layer4_out[7419] = layer3_out[4117];
    assign layer4_out[7420] = ~layer3_out[4006] | layer3_out[4007];
    assign layer4_out[7421] = ~layer3_out[504] | layer3_out[503];
    assign layer4_out[7422] = layer3_out[766] & layer3_out[767];
    assign layer4_out[7423] = ~layer3_out[4127] | layer3_out[4126];
    assign layer4_out[7424] = ~(layer3_out[4475] & layer3_out[4476]);
    assign layer4_out[7425] = layer3_out[2937] & ~layer3_out[2938];
    assign layer4_out[7426] = ~layer3_out[3685];
    assign layer4_out[7427] = ~(layer3_out[865] ^ layer3_out[866]);
    assign layer4_out[7428] = layer3_out[5133] ^ layer3_out[5134];
    assign layer4_out[7429] = layer3_out[4280] | layer3_out[4281];
    assign layer4_out[7430] = ~(layer3_out[2224] ^ layer3_out[2225]);
    assign layer4_out[7431] = 1'b1;
    assign layer4_out[7432] = layer3_out[7603];
    assign layer4_out[7433] = layer3_out[5181];
    assign layer4_out[7434] = ~layer3_out[1618];
    assign layer4_out[7435] = ~layer3_out[6229];
    assign layer4_out[7436] = ~layer3_out[2749] | layer3_out[2750];
    assign layer4_out[7437] = layer3_out[1173];
    assign layer4_out[7438] = ~(layer3_out[2679] & layer3_out[2680]);
    assign layer4_out[7439] = ~layer3_out[7629];
    assign layer4_out[7440] = layer3_out[215] & layer3_out[216];
    assign layer4_out[7441] = layer3_out[6552] & layer3_out[6553];
    assign layer4_out[7442] = layer3_out[3890] | layer3_out[3891];
    assign layer4_out[7443] = ~(layer3_out[5921] ^ layer3_out[5922]);
    assign layer4_out[7444] = layer3_out[3174] ^ layer3_out[3175];
    assign layer4_out[7445] = layer3_out[7470];
    assign layer4_out[7446] = ~(layer3_out[116] ^ layer3_out[117]);
    assign layer4_out[7447] = ~layer3_out[7845] | layer3_out[7846];
    assign layer4_out[7448] = ~layer3_out[2171];
    assign layer4_out[7449] = ~(layer3_out[7069] | layer3_out[7070]);
    assign layer4_out[7450] = layer3_out[3105] ^ layer3_out[3106];
    assign layer4_out[7451] = ~layer3_out[1248];
    assign layer4_out[7452] = layer3_out[5644] & layer3_out[5645];
    assign layer4_out[7453] = ~layer3_out[5123];
    assign layer4_out[7454] = layer3_out[215];
    assign layer4_out[7455] = ~layer3_out[7691];
    assign layer4_out[7456] = layer3_out[2068] | layer3_out[2069];
    assign layer4_out[7457] = ~layer3_out[2198];
    assign layer4_out[7458] = layer3_out[6205] | layer3_out[6206];
    assign layer4_out[7459] = ~layer3_out[6482];
    assign layer4_out[7460] = layer3_out[4594] & ~layer3_out[4593];
    assign layer4_out[7461] = ~(layer3_out[5379] ^ layer3_out[5380]);
    assign layer4_out[7462] = ~(layer3_out[2426] | layer3_out[2427]);
    assign layer4_out[7463] = layer3_out[3622];
    assign layer4_out[7464] = layer3_out[4280];
    assign layer4_out[7465] = layer3_out[2518];
    assign layer4_out[7466] = ~layer3_out[5226];
    assign layer4_out[7467] = layer3_out[5195];
    assign layer4_out[7468] = ~layer3_out[3959];
    assign layer4_out[7469] = ~(layer3_out[3492] | layer3_out[3493]);
    assign layer4_out[7470] = layer3_out[2678] ^ layer3_out[2679];
    assign layer4_out[7471] = ~layer3_out[1983] | layer3_out[1984];
    assign layer4_out[7472] = layer3_out[5621] & ~layer3_out[5622];
    assign layer4_out[7473] = ~layer3_out[2210];
    assign layer4_out[7474] = ~layer3_out[3164];
    assign layer4_out[7475] = ~(layer3_out[2329] | layer3_out[2330]);
    assign layer4_out[7476] = ~(layer3_out[5947] ^ layer3_out[5948]);
    assign layer4_out[7477] = ~layer3_out[1443];
    assign layer4_out[7478] = ~(layer3_out[7161] | layer3_out[7162]);
    assign layer4_out[7479] = layer3_out[4932] | layer3_out[4933];
    assign layer4_out[7480] = layer3_out[3278] ^ layer3_out[3279];
    assign layer4_out[7481] = ~layer3_out[4422];
    assign layer4_out[7482] = layer3_out[6212] & ~layer3_out[6211];
    assign layer4_out[7483] = layer3_out[556] ^ layer3_out[557];
    assign layer4_out[7484] = layer3_out[1972] & ~layer3_out[1971];
    assign layer4_out[7485] = layer3_out[7292] | layer3_out[7293];
    assign layer4_out[7486] = ~(layer3_out[1273] | layer3_out[1274]);
    assign layer4_out[7487] = ~layer3_out[3330] | layer3_out[3329];
    assign layer4_out[7488] = layer3_out[6751];
    assign layer4_out[7489] = ~(layer3_out[6547] | layer3_out[6548]);
    assign layer4_out[7490] = layer3_out[1153] & ~layer3_out[1154];
    assign layer4_out[7491] = layer3_out[7240];
    assign layer4_out[7492] = layer3_out[2580] ^ layer3_out[2581];
    assign layer4_out[7493] = ~layer3_out[3246];
    assign layer4_out[7494] = ~(layer3_out[920] & layer3_out[921]);
    assign layer4_out[7495] = ~layer3_out[3057];
    assign layer4_out[7496] = ~layer3_out[6719] | layer3_out[6720];
    assign layer4_out[7497] = layer3_out[5823] & layer3_out[5824];
    assign layer4_out[7498] = ~layer3_out[1999] | layer3_out[1998];
    assign layer4_out[7499] = layer3_out[728];
    assign layer4_out[7500] = layer3_out[6538];
    assign layer4_out[7501] = ~(layer3_out[6787] ^ layer3_out[6788]);
    assign layer4_out[7502] = ~layer3_out[6962];
    assign layer4_out[7503] = layer3_out[3898] ^ layer3_out[3899];
    assign layer4_out[7504] = layer3_out[6017] | layer3_out[6018];
    assign layer4_out[7505] = ~(layer3_out[499] ^ layer3_out[500]);
    assign layer4_out[7506] = ~(layer3_out[3195] & layer3_out[3196]);
    assign layer4_out[7507] = layer3_out[1772];
    assign layer4_out[7508] = layer3_out[4658];
    assign layer4_out[7509] = layer3_out[7390];
    assign layer4_out[7510] = ~layer3_out[861] | layer3_out[862];
    assign layer4_out[7511] = layer3_out[3345];
    assign layer4_out[7512] = ~layer3_out[3905];
    assign layer4_out[7513] = layer3_out[6685];
    assign layer4_out[7514] = layer3_out[1520] & layer3_out[1521];
    assign layer4_out[7515] = layer3_out[6354] & ~layer3_out[6353];
    assign layer4_out[7516] = layer3_out[7866];
    assign layer4_out[7517] = layer3_out[1450] & layer3_out[1451];
    assign layer4_out[7518] = layer3_out[4000] & ~layer3_out[4001];
    assign layer4_out[7519] = ~(layer3_out[2946] | layer3_out[2947]);
    assign layer4_out[7520] = ~(layer3_out[6359] | layer3_out[6360]);
    assign layer4_out[7521] = layer3_out[4904] | layer3_out[4905];
    assign layer4_out[7522] = ~layer3_out[5416] | layer3_out[5415];
    assign layer4_out[7523] = ~layer3_out[4377];
    assign layer4_out[7524] = layer3_out[764];
    assign layer4_out[7525] = ~layer3_out[7241];
    assign layer4_out[7526] = layer3_out[3599] & ~layer3_out[3598];
    assign layer4_out[7527] = layer3_out[3229];
    assign layer4_out[7528] = layer3_out[410] | layer3_out[411];
    assign layer4_out[7529] = ~layer3_out[7220];
    assign layer4_out[7530] = layer3_out[4];
    assign layer4_out[7531] = ~layer3_out[2170];
    assign layer4_out[7532] = layer3_out[3364] ^ layer3_out[3365];
    assign layer4_out[7533] = ~layer3_out[4479] | layer3_out[4480];
    assign layer4_out[7534] = ~layer3_out[583] | layer3_out[582];
    assign layer4_out[7535] = ~layer3_out[1060];
    assign layer4_out[7536] = ~(layer3_out[4180] ^ layer3_out[4181]);
    assign layer4_out[7537] = layer3_out[3509];
    assign layer4_out[7538] = layer3_out[293];
    assign layer4_out[7539] = layer3_out[6983] & layer3_out[6984];
    assign layer4_out[7540] = ~(layer3_out[620] ^ layer3_out[621]);
    assign layer4_out[7541] = ~layer3_out[1816] | layer3_out[1815];
    assign layer4_out[7542] = ~layer3_out[2313];
    assign layer4_out[7543] = ~layer3_out[5014] | layer3_out[5015];
    assign layer4_out[7544] = layer3_out[5115] & ~layer3_out[5114];
    assign layer4_out[7545] = layer3_out[3131];
    assign layer4_out[7546] = ~(layer3_out[5338] & layer3_out[5339]);
    assign layer4_out[7547] = layer3_out[3107] & layer3_out[3108];
    assign layer4_out[7548] = layer3_out[3559] & ~layer3_out[3558];
    assign layer4_out[7549] = ~(layer3_out[4740] ^ layer3_out[4741]);
    assign layer4_out[7550] = ~(layer3_out[1963] | layer3_out[1964]);
    assign layer4_out[7551] = layer3_out[7601] & layer3_out[7602];
    assign layer4_out[7552] = ~layer3_out[4425];
    assign layer4_out[7553] = ~layer3_out[989];
    assign layer4_out[7554] = layer3_out[1746];
    assign layer4_out[7555] = ~layer3_out[6508] | layer3_out[6507];
    assign layer4_out[7556] = ~layer3_out[288];
    assign layer4_out[7557] = layer3_out[6546];
    assign layer4_out[7558] = ~layer3_out[1200];
    assign layer4_out[7559] = layer3_out[5872];
    assign layer4_out[7560] = layer3_out[6971] & ~layer3_out[6972];
    assign layer4_out[7561] = layer3_out[2754] & layer3_out[2755];
    assign layer4_out[7562] = ~layer3_out[4036];
    assign layer4_out[7563] = ~layer3_out[5451] | layer3_out[5450];
    assign layer4_out[7564] = layer3_out[1885];
    assign layer4_out[7565] = layer3_out[7109] & layer3_out[7110];
    assign layer4_out[7566] = ~(layer3_out[2455] ^ layer3_out[2456]);
    assign layer4_out[7567] = layer3_out[709] | layer3_out[710];
    assign layer4_out[7568] = layer3_out[688] ^ layer3_out[689];
    assign layer4_out[7569] = ~layer3_out[5144];
    assign layer4_out[7570] = layer3_out[7879] & layer3_out[7880];
    assign layer4_out[7571] = ~layer3_out[3157];
    assign layer4_out[7572] = layer3_out[5016] | layer3_out[5017];
    assign layer4_out[7573] = ~layer3_out[2139];
    assign layer4_out[7574] = ~layer3_out[3300];
    assign layer4_out[7575] = layer3_out[58];
    assign layer4_out[7576] = layer3_out[3686] & layer3_out[3687];
    assign layer4_out[7577] = layer3_out[2561] & ~layer3_out[2560];
    assign layer4_out[7578] = layer3_out[477] & ~layer3_out[478];
    assign layer4_out[7579] = layer3_out[2979];
    assign layer4_out[7580] = layer3_out[242];
    assign layer4_out[7581] = layer3_out[2848];
    assign layer4_out[7582] = ~layer3_out[959];
    assign layer4_out[7583] = ~layer3_out[4474] | layer3_out[4475];
    assign layer4_out[7584] = ~(layer3_out[237] & layer3_out[238]);
    assign layer4_out[7585] = layer3_out[6819] & ~layer3_out[6820];
    assign layer4_out[7586] = ~(layer3_out[4093] | layer3_out[4094]);
    assign layer4_out[7587] = ~layer3_out[3428];
    assign layer4_out[7588] = layer3_out[6929] & ~layer3_out[6930];
    assign layer4_out[7589] = ~layer3_out[3498];
    assign layer4_out[7590] = ~layer3_out[3590];
    assign layer4_out[7591] = ~layer3_out[5805] | layer3_out[5806];
    assign layer4_out[7592] = layer3_out[4824];
    assign layer4_out[7593] = ~layer3_out[2105];
    assign layer4_out[7594] = layer3_out[4184];
    assign layer4_out[7595] = ~layer3_out[1949];
    assign layer4_out[7596] = layer3_out[1880] ^ layer3_out[1881];
    assign layer4_out[7597] = ~layer3_out[4986] | layer3_out[4985];
    assign layer4_out[7598] = ~layer3_out[2983] | layer3_out[2984];
    assign layer4_out[7599] = layer3_out[2971] & layer3_out[2972];
    assign layer4_out[7600] = ~layer3_out[3869];
    assign layer4_out[7601] = ~layer3_out[6776];
    assign layer4_out[7602] = layer3_out[3094];
    assign layer4_out[7603] = layer3_out[3222] ^ layer3_out[3223];
    assign layer4_out[7604] = ~(layer3_out[2772] ^ layer3_out[2773]);
    assign layer4_out[7605] = layer3_out[4469];
    assign layer4_out[7606] = layer3_out[7553] ^ layer3_out[7554];
    assign layer4_out[7607] = ~layer3_out[3749];
    assign layer4_out[7608] = layer3_out[3019] & ~layer3_out[3018];
    assign layer4_out[7609] = ~layer3_out[6248];
    assign layer4_out[7610] = ~layer3_out[3089];
    assign layer4_out[7611] = layer3_out[5825];
    assign layer4_out[7612] = ~(layer3_out[275] | layer3_out[276]);
    assign layer4_out[7613] = layer3_out[4839];
    assign layer4_out[7614] = ~layer3_out[7212] | layer3_out[7213];
    assign layer4_out[7615] = layer3_out[3626];
    assign layer4_out[7616] = layer3_out[4840] & ~layer3_out[4839];
    assign layer4_out[7617] = layer3_out[6609] & layer3_out[6610];
    assign layer4_out[7618] = ~layer3_out[2741];
    assign layer4_out[7619] = ~(layer3_out[5454] ^ layer3_out[5455]);
    assign layer4_out[7620] = layer3_out[5211] ^ layer3_out[5212];
    assign layer4_out[7621] = layer3_out[7479];
    assign layer4_out[7622] = layer3_out[987] & ~layer3_out[986];
    assign layer4_out[7623] = ~layer3_out[1415];
    assign layer4_out[7624] = ~layer3_out[7747];
    assign layer4_out[7625] = layer3_out[7533] | layer3_out[7534];
    assign layer4_out[7626] = layer3_out[2439] ^ layer3_out[2440];
    assign layer4_out[7627] = ~layer3_out[183];
    assign layer4_out[7628] = ~layer3_out[201];
    assign layer4_out[7629] = layer3_out[1398];
    assign layer4_out[7630] = layer3_out[6942] & ~layer3_out[6943];
    assign layer4_out[7631] = ~layer3_out[1045];
    assign layer4_out[7632] = layer3_out[56] & ~layer3_out[57];
    assign layer4_out[7633] = layer3_out[4425];
    assign layer4_out[7634] = layer3_out[3314];
    assign layer4_out[7635] = layer3_out[7870];
    assign layer4_out[7636] = layer3_out[5109];
    assign layer4_out[7637] = ~layer3_out[4091];
    assign layer4_out[7638] = ~layer3_out[4008] | layer3_out[4009];
    assign layer4_out[7639] = ~(layer3_out[311] | layer3_out[312]);
    assign layer4_out[7640] = ~(layer3_out[7330] | layer3_out[7331]);
    assign layer4_out[7641] = ~(layer3_out[7434] | layer3_out[7435]);
    assign layer4_out[7642] = layer3_out[2988] ^ layer3_out[2989];
    assign layer4_out[7643] = layer3_out[2870];
    assign layer4_out[7644] = ~layer3_out[790] | layer3_out[789];
    assign layer4_out[7645] = layer3_out[1667] & ~layer3_out[1668];
    assign layer4_out[7646] = layer3_out[101];
    assign layer4_out[7647] = ~(layer3_out[6949] ^ layer3_out[6950]);
    assign layer4_out[7648] = ~layer3_out[1387];
    assign layer4_out[7649] = ~layer3_out[454];
    assign layer4_out[7650] = ~(layer3_out[908] | layer3_out[909]);
    assign layer4_out[7651] = ~layer3_out[3763];
    assign layer4_out[7652] = ~(layer3_out[699] ^ layer3_out[700]);
    assign layer4_out[7653] = ~(layer3_out[7995] ^ layer3_out[7996]);
    assign layer4_out[7654] = ~layer3_out[6759];
    assign layer4_out[7655] = ~layer3_out[1366];
    assign layer4_out[7656] = ~layer3_out[7708] | layer3_out[7707];
    assign layer4_out[7657] = layer3_out[544] | layer3_out[545];
    assign layer4_out[7658] = layer3_out[460];
    assign layer4_out[7659] = ~layer3_out[2962];
    assign layer4_out[7660] = layer3_out[3116] ^ layer3_out[3117];
    assign layer4_out[7661] = ~(layer3_out[5896] ^ layer3_out[5897]);
    assign layer4_out[7662] = layer3_out[7537] & ~layer3_out[7538];
    assign layer4_out[7663] = ~layer3_out[4708];
    assign layer4_out[7664] = ~layer3_out[6968];
    assign layer4_out[7665] = ~(layer3_out[598] & layer3_out[599]);
    assign layer4_out[7666] = layer3_out[6540] ^ layer3_out[6541];
    assign layer4_out[7667] = layer3_out[966];
    assign layer4_out[7668] = layer3_out[307] ^ layer3_out[308];
    assign layer4_out[7669] = layer3_out[1680] & layer3_out[1681];
    assign layer4_out[7670] = ~layer3_out[6078] | layer3_out[6079];
    assign layer4_out[7671] = ~layer3_out[393];
    assign layer4_out[7672] = ~layer3_out[5389];
    assign layer4_out[7673] = ~layer3_out[6250];
    assign layer4_out[7674] = layer3_out[1205];
    assign layer4_out[7675] = ~(layer3_out[6243] | layer3_out[6244]);
    assign layer4_out[7676] = layer3_out[1034];
    assign layer4_out[7677] = layer3_out[4704] & ~layer3_out[4705];
    assign layer4_out[7678] = ~layer3_out[7335] | layer3_out[7334];
    assign layer4_out[7679] = ~layer3_out[7874];
    assign layer4_out[7680] = ~(layer3_out[3768] & layer3_out[3769]);
    assign layer4_out[7681] = layer3_out[2383];
    assign layer4_out[7682] = ~layer3_out[3189];
    assign layer4_out[7683] = layer3_out[1592];
    assign layer4_out[7684] = ~layer3_out[3592];
    assign layer4_out[7685] = layer3_out[5638];
    assign layer4_out[7686] = layer3_out[5945] | layer3_out[5946];
    assign layer4_out[7687] = ~layer3_out[5849] | layer3_out[5850];
    assign layer4_out[7688] = layer3_out[1121] ^ layer3_out[1122];
    assign layer4_out[7689] = layer3_out[4039] & ~layer3_out[4040];
    assign layer4_out[7690] = ~layer3_out[4555];
    assign layer4_out[7691] = ~layer3_out[6824];
    assign layer4_out[7692] = layer3_out[7064] & layer3_out[7065];
    assign layer4_out[7693] = layer3_out[3066];
    assign layer4_out[7694] = layer3_out[5890];
    assign layer4_out[7695] = layer3_out[439];
    assign layer4_out[7696] = 1'b0;
    assign layer4_out[7697] = ~layer3_out[1395];
    assign layer4_out[7698] = ~layer3_out[3607];
    assign layer4_out[7699] = layer3_out[5247];
    assign layer4_out[7700] = layer3_out[5412] | layer3_out[5413];
    assign layer4_out[7701] = ~layer3_out[4756] | layer3_out[4757];
    assign layer4_out[7702] = ~(layer3_out[1855] | layer3_out[1856]);
    assign layer4_out[7703] = layer3_out[5182] ^ layer3_out[5183];
    assign layer4_out[7704] = layer3_out[7480] & ~layer3_out[7481];
    assign layer4_out[7705] = layer3_out[3983];
    assign layer4_out[7706] = layer3_out[4157] ^ layer3_out[4158];
    assign layer4_out[7707] = layer3_out[7660] ^ layer3_out[7661];
    assign layer4_out[7708] = layer3_out[7987];
    assign layer4_out[7709] = ~(layer3_out[6406] & layer3_out[6407]);
    assign layer4_out[7710] = layer3_out[328] ^ layer3_out[329];
    assign layer4_out[7711] = ~layer3_out[75];
    assign layer4_out[7712] = ~layer3_out[3947] | layer3_out[3948];
    assign layer4_out[7713] = ~(layer3_out[7683] ^ layer3_out[7684]);
    assign layer4_out[7714] = ~layer3_out[6691];
    assign layer4_out[7715] = layer3_out[7450] ^ layer3_out[7451];
    assign layer4_out[7716] = layer3_out[7475];
    assign layer4_out[7717] = ~layer3_out[1819] | layer3_out[1820];
    assign layer4_out[7718] = ~(layer3_out[885] ^ layer3_out[886]);
    assign layer4_out[7719] = ~layer3_out[1189];
    assign layer4_out[7720] = layer3_out[4101] & layer3_out[4102];
    assign layer4_out[7721] = ~(layer3_out[7019] | layer3_out[7020]);
    assign layer4_out[7722] = ~layer3_out[2220];
    assign layer4_out[7723] = ~(layer3_out[7637] ^ layer3_out[7638]);
    assign layer4_out[7724] = ~layer3_out[1489];
    assign layer4_out[7725] = layer3_out[5091] & layer3_out[5092];
    assign layer4_out[7726] = layer3_out[6848];
    assign layer4_out[7727] = layer3_out[4509] | layer3_out[4510];
    assign layer4_out[7728] = layer3_out[2451] | layer3_out[2452];
    assign layer4_out[7729] = ~layer3_out[3430];
    assign layer4_out[7730] = layer3_out[2970] & ~layer3_out[2971];
    assign layer4_out[7731] = ~layer3_out[5307] | layer3_out[5306];
    assign layer4_out[7732] = ~layer3_out[7102];
    assign layer4_out[7733] = layer3_out[1241];
    assign layer4_out[7734] = ~layer3_out[7766] | layer3_out[7765];
    assign layer4_out[7735] = layer3_out[3017] & ~layer3_out[3016];
    assign layer4_out[7736] = layer3_out[3332] & ~layer3_out[3331];
    assign layer4_out[7737] = ~(layer3_out[3727] ^ layer3_out[3728]);
    assign layer4_out[7738] = layer3_out[3377] & layer3_out[3378];
    assign layer4_out[7739] = ~layer3_out[7482];
    assign layer4_out[7740] = ~(layer3_out[1529] | layer3_out[1530]);
    assign layer4_out[7741] = layer3_out[2281] & ~layer3_out[2280];
    assign layer4_out[7742] = layer3_out[7276] & ~layer3_out[7275];
    assign layer4_out[7743] = ~layer3_out[7375] | layer3_out[7376];
    assign layer4_out[7744] = layer3_out[1295] | layer3_out[1296];
    assign layer4_out[7745] = layer3_out[5766];
    assign layer4_out[7746] = ~layer3_out[2306] | layer3_out[2305];
    assign layer4_out[7747] = layer3_out[2670];
    assign layer4_out[7748] = layer3_out[170] | layer3_out[171];
    assign layer4_out[7749] = ~layer3_out[2326] | layer3_out[2325];
    assign layer4_out[7750] = layer3_out[3519];
    assign layer4_out[7751] = layer3_out[2054] & layer3_out[2055];
    assign layer4_out[7752] = ~layer3_out[3197] | layer3_out[3198];
    assign layer4_out[7753] = ~layer3_out[6145];
    assign layer4_out[7754] = layer3_out[6823];
    assign layer4_out[7755] = layer3_out[3996] & ~layer3_out[3997];
    assign layer4_out[7756] = ~layer3_out[2522];
    assign layer4_out[7757] = layer3_out[4629] & ~layer3_out[4630];
    assign layer4_out[7758] = layer3_out[5601] & ~layer3_out[5600];
    assign layer4_out[7759] = layer3_out[4742] & ~layer3_out[4741];
    assign layer4_out[7760] = layer3_out[270] ^ layer3_out[271];
    assign layer4_out[7761] = layer3_out[3619];
    assign layer4_out[7762] = ~layer3_out[7000];
    assign layer4_out[7763] = ~layer3_out[4624] | layer3_out[4623];
    assign layer4_out[7764] = ~layer3_out[6691];
    assign layer4_out[7765] = layer3_out[1324] ^ layer3_out[1325];
    assign layer4_out[7766] = ~layer3_out[5529];
    assign layer4_out[7767] = ~layer3_out[751];
    assign layer4_out[7768] = ~layer3_out[7159] | layer3_out[7158];
    assign layer4_out[7769] = layer3_out[4620];
    assign layer4_out[7770] = ~layer3_out[4592];
    assign layer4_out[7771] = layer3_out[6321];
    assign layer4_out[7772] = layer3_out[6241] | layer3_out[6242];
    assign layer4_out[7773] = ~(layer3_out[2568] | layer3_out[2569]);
    assign layer4_out[7774] = ~layer3_out[5855];
    assign layer4_out[7775] = ~layer3_out[7309];
    assign layer4_out[7776] = ~layer3_out[3679];
    assign layer4_out[7777] = layer3_out[6276] & layer3_out[6277];
    assign layer4_out[7778] = ~layer3_out[788];
    assign layer4_out[7779] = ~(layer3_out[935] ^ layer3_out[936]);
    assign layer4_out[7780] = ~(layer3_out[2510] | layer3_out[2511]);
    assign layer4_out[7781] = layer3_out[2160];
    assign layer4_out[7782] = layer3_out[3284] & ~layer3_out[3285];
    assign layer4_out[7783] = ~(layer3_out[5287] | layer3_out[5288]);
    assign layer4_out[7784] = ~layer3_out[4714];
    assign layer4_out[7785] = layer3_out[690] ^ layer3_out[691];
    assign layer4_out[7786] = ~(layer3_out[2811] & layer3_out[2812]);
    assign layer4_out[7787] = ~layer3_out[1637];
    assign layer4_out[7788] = layer3_out[4668];
    assign layer4_out[7789] = ~layer3_out[882];
    assign layer4_out[7790] = layer3_out[2488] ^ layer3_out[2489];
    assign layer4_out[7791] = ~layer3_out[5737];
    assign layer4_out[7792] = ~layer3_out[1581];
    assign layer4_out[7793] = layer3_out[515];
    assign layer4_out[7794] = layer3_out[7795];
    assign layer4_out[7795] = layer3_out[6603];
    assign layer4_out[7796] = layer3_out[1381] & ~layer3_out[1382];
    assign layer4_out[7797] = 1'b1;
    assign layer4_out[7798] = layer3_out[7403];
    assign layer4_out[7799] = layer3_out[2943] ^ layer3_out[2944];
    assign layer4_out[7800] = ~(layer3_out[428] ^ layer3_out[429]);
    assign layer4_out[7801] = ~layer3_out[608] | layer3_out[609];
    assign layer4_out[7802] = ~(layer3_out[5582] & layer3_out[5583]);
    assign layer4_out[7803] = ~layer3_out[2188] | layer3_out[2187];
    assign layer4_out[7804] = layer3_out[2734] & layer3_out[2735];
    assign layer4_out[7805] = layer3_out[1824] & layer3_out[1825];
    assign layer4_out[7806] = layer3_out[6895];
    assign layer4_out[7807] = layer3_out[2188] & layer3_out[2189];
    assign layer4_out[7808] = ~(layer3_out[6239] ^ layer3_out[6240]);
    assign layer4_out[7809] = ~(layer3_out[747] ^ layer3_out[748]);
    assign layer4_out[7810] = ~layer3_out[1779] | layer3_out[1780];
    assign layer4_out[7811] = layer3_out[7079] | layer3_out[7080];
    assign layer4_out[7812] = ~(layer3_out[945] & layer3_out[946]);
    assign layer4_out[7813] = ~layer3_out[851];
    assign layer4_out[7814] = ~(layer3_out[6902] & layer3_out[6903]);
    assign layer4_out[7815] = layer3_out[7387];
    assign layer4_out[7816] = layer3_out[5253] & ~layer3_out[5254];
    assign layer4_out[7817] = ~layer3_out[5065];
    assign layer4_out[7818] = layer3_out[1747] | layer3_out[1748];
    assign layer4_out[7819] = layer3_out[7924] & ~layer3_out[7923];
    assign layer4_out[7820] = ~layer3_out[1774] | layer3_out[1773];
    assign layer4_out[7821] = layer3_out[2021] & ~layer3_out[2022];
    assign layer4_out[7822] = layer3_out[4671] ^ layer3_out[4672];
    assign layer4_out[7823] = layer3_out[4017] & layer3_out[4018];
    assign layer4_out[7824] = layer3_out[7700];
    assign layer4_out[7825] = layer3_out[5021] ^ layer3_out[5022];
    assign layer4_out[7826] = layer3_out[8];
    assign layer4_out[7827] = layer3_out[35] | layer3_out[36];
    assign layer4_out[7828] = ~(layer3_out[6463] ^ layer3_out[6464]);
    assign layer4_out[7829] = ~(layer3_out[4460] ^ layer3_out[4461]);
    assign layer4_out[7830] = layer3_out[3648];
    assign layer4_out[7831] = ~layer3_out[2159];
    assign layer4_out[7832] = layer3_out[1323] & layer3_out[1324];
    assign layer4_out[7833] = layer3_out[7290] & ~layer3_out[7289];
    assign layer4_out[7834] = layer3_out[6782] & layer3_out[6783];
    assign layer4_out[7835] = layer3_out[3840] | layer3_out[3841];
    assign layer4_out[7836] = ~layer3_out[2063];
    assign layer4_out[7837] = ~layer3_out[7708];
    assign layer4_out[7838] = layer3_out[845];
    assign layer4_out[7839] = ~(layer3_out[3022] & layer3_out[3023]);
    assign layer4_out[7840] = ~(layer3_out[1258] ^ layer3_out[1259]);
    assign layer4_out[7841] = ~layer3_out[5077];
    assign layer4_out[7842] = layer3_out[2132];
    assign layer4_out[7843] = layer3_out[2794];
    assign layer4_out[7844] = ~layer3_out[3069];
    assign layer4_out[7845] = layer3_out[1908];
    assign layer4_out[7846] = ~(layer3_out[1168] & layer3_out[1169]);
    assign layer4_out[7847] = ~layer3_out[7354];
    assign layer4_out[7848] = layer3_out[5956] & layer3_out[5957];
    assign layer4_out[7849] = ~layer3_out[1349];
    assign layer4_out[7850] = ~layer3_out[4493] | layer3_out[4492];
    assign layer4_out[7851] = layer3_out[2575] & ~layer3_out[2576];
    assign layer4_out[7852] = 1'b1;
    assign layer4_out[7853] = layer3_out[2977];
    assign layer4_out[7854] = ~layer3_out[7761] | layer3_out[7762];
    assign layer4_out[7855] = layer3_out[853] & layer3_out[854];
    assign layer4_out[7856] = layer3_out[70];
    assign layer4_out[7857] = layer3_out[6585];
    assign layer4_out[7858] = layer3_out[2178] | layer3_out[2179];
    assign layer4_out[7859] = layer3_out[5099] ^ layer3_out[5100];
    assign layer4_out[7860] = ~(layer3_out[2182] ^ layer3_out[2183]);
    assign layer4_out[7861] = ~layer3_out[6297] | layer3_out[6296];
    assign layer4_out[7862] = ~layer3_out[4251] | layer3_out[4252];
    assign layer4_out[7863] = layer3_out[6944] & ~layer3_out[6945];
    assign layer4_out[7864] = layer3_out[3142];
    assign layer4_out[7865] = ~(layer3_out[357] ^ layer3_out[358]);
    assign layer4_out[7866] = ~layer3_out[6118];
    assign layer4_out[7867] = ~layer3_out[3252];
    assign layer4_out[7868] = ~layer3_out[1045];
    assign layer4_out[7869] = ~layer3_out[3520];
    assign layer4_out[7870] = layer3_out[884];
    assign layer4_out[7871] = layer3_out[4761] ^ layer3_out[4762];
    assign layer4_out[7872] = layer3_out[64];
    assign layer4_out[7873] = ~(layer3_out[288] | layer3_out[289]);
    assign layer4_out[7874] = 1'b1;
    assign layer4_out[7875] = layer3_out[6685] & ~layer3_out[6684];
    assign layer4_out[7876] = ~(layer3_out[7429] | layer3_out[7430]);
    assign layer4_out[7877] = layer3_out[6408] & ~layer3_out[6409];
    assign layer4_out[7878] = ~layer3_out[2534];
    assign layer4_out[7879] = ~(layer3_out[4342] & layer3_out[4343]);
    assign layer4_out[7880] = layer3_out[1563] ^ layer3_out[1564];
    assign layer4_out[7881] = ~layer3_out[1839] | layer3_out[1840];
    assign layer4_out[7882] = layer3_out[3845];
    assign layer4_out[7883] = layer3_out[3630];
    assign layer4_out[7884] = layer3_out[655];
    assign layer4_out[7885] = ~(layer3_out[136] ^ layer3_out[137]);
    assign layer4_out[7886] = layer3_out[4896];
    assign layer4_out[7887] = ~layer3_out[7464];
    assign layer4_out[7888] = 1'b1;
    assign layer4_out[7889] = layer3_out[5471] & ~layer3_out[5470];
    assign layer4_out[7890] = ~layer3_out[5602] | layer3_out[5603];
    assign layer4_out[7891] = layer3_out[4525];
    assign layer4_out[7892] = ~(layer3_out[697] & layer3_out[698]);
    assign layer4_out[7893] = layer3_out[1312];
    assign layer4_out[7894] = ~layer3_out[6394];
    assign layer4_out[7895] = layer3_out[1408];
    assign layer4_out[7896] = layer3_out[3697] & ~layer3_out[3696];
    assign layer4_out[7897] = layer3_out[7316];
    assign layer4_out[7898] = layer3_out[4406] | layer3_out[4407];
    assign layer4_out[7899] = ~(layer3_out[7756] ^ layer3_out[7757]);
    assign layer4_out[7900] = layer3_out[1457] ^ layer3_out[1458];
    assign layer4_out[7901] = ~layer3_out[4314];
    assign layer4_out[7902] = ~layer3_out[4630];
    assign layer4_out[7903] = ~layer3_out[7804] | layer3_out[7805];
    assign layer4_out[7904] = layer3_out[4359] & ~layer3_out[4358];
    assign layer4_out[7905] = ~layer3_out[5643] | layer3_out[5642];
    assign layer4_out[7906] = layer3_out[3924];
    assign layer4_out[7907] = layer3_out[1722];
    assign layer4_out[7908] = ~layer3_out[2538];
    assign layer4_out[7909] = layer3_out[6166] ^ layer3_out[6167];
    assign layer4_out[7910] = layer3_out[3414];
    assign layer4_out[7911] = layer3_out[1166];
    assign layer4_out[7912] = ~layer3_out[5713] | layer3_out[5714];
    assign layer4_out[7913] = layer3_out[968];
    assign layer4_out[7914] = ~layer3_out[2545] | layer3_out[2546];
    assign layer4_out[7915] = ~(layer3_out[6413] | layer3_out[6414]);
    assign layer4_out[7916] = layer3_out[7679] & ~layer3_out[7680];
    assign layer4_out[7917] = layer3_out[1143];
    assign layer4_out[7918] = layer3_out[5501] & ~layer3_out[5500];
    assign layer4_out[7919] = ~layer3_out[5342];
    assign layer4_out[7920] = ~layer3_out[904];
    assign layer4_out[7921] = ~layer3_out[775];
    assign layer4_out[7922] = ~layer3_out[2802];
    assign layer4_out[7923] = ~layer3_out[1492] | layer3_out[1491];
    assign layer4_out[7924] = ~layer3_out[134];
    assign layer4_out[7925] = layer3_out[3288];
    assign layer4_out[7926] = layer3_out[4032] & layer3_out[4033];
    assign layer4_out[7927] = layer3_out[3382] ^ layer3_out[3383];
    assign layer4_out[7928] = layer3_out[6287] & layer3_out[6288];
    assign layer4_out[7929] = layer3_out[5200];
    assign layer4_out[7930] = layer3_out[1364];
    assign layer4_out[7931] = ~(layer3_out[4923] & layer3_out[4924]);
    assign layer4_out[7932] = ~layer3_out[1961];
    assign layer4_out[7933] = ~(layer3_out[1026] ^ layer3_out[1027]);
    assign layer4_out[7934] = layer3_out[6634];
    assign layer4_out[7935] = ~(layer3_out[7027] ^ layer3_out[7028]);
    assign layer4_out[7936] = ~layer3_out[897] | layer3_out[896];
    assign layer4_out[7937] = layer3_out[44] & ~layer3_out[43];
    assign layer4_out[7938] = ~layer3_out[7142] | layer3_out[7141];
    assign layer4_out[7939] = layer3_out[7675] | layer3_out[7676];
    assign layer4_out[7940] = layer3_out[4454];
    assign layer4_out[7941] = ~(layer3_out[2908] ^ layer3_out[2909]);
    assign layer4_out[7942] = ~layer3_out[3814];
    assign layer4_out[7943] = ~layer3_out[4923];
    assign layer4_out[7944] = layer3_out[4238];
    assign layer4_out[7945] = ~(layer3_out[496] & layer3_out[497]);
    assign layer4_out[7946] = ~layer3_out[5981];
    assign layer4_out[7947] = layer3_out[3695] & layer3_out[3696];
    assign layer4_out[7948] = ~layer3_out[7547];
    assign layer4_out[7949] = layer3_out[6145];
    assign layer4_out[7950] = ~(layer3_out[5888] ^ layer3_out[5889]);
    assign layer4_out[7951] = layer3_out[5094] & ~layer3_out[5093];
    assign layer4_out[7952] = layer3_out[2127] & ~layer3_out[2126];
    assign layer4_out[7953] = ~layer3_out[2815];
    assign layer4_out[7954] = ~layer3_out[7796];
    assign layer4_out[7955] = ~layer3_out[5624];
    assign layer4_out[7956] = layer3_out[779];
    assign layer4_out[7957] = ~layer3_out[2643];
    assign layer4_out[7958] = layer3_out[2769];
    assign layer4_out[7959] = ~layer3_out[1209];
    assign layer4_out[7960] = layer3_out[7603];
    assign layer4_out[7961] = layer3_out[5838] & layer3_out[5839];
    assign layer4_out[7962] = layer3_out[5109];
    assign layer4_out[7963] = ~(layer3_out[5974] & layer3_out[5975]);
    assign layer4_out[7964] = ~layer3_out[2877];
    assign layer4_out[7965] = ~(layer3_out[38] ^ layer3_out[39]);
    assign layer4_out[7966] = ~layer3_out[353];
    assign layer4_out[7967] = layer3_out[505] & layer3_out[506];
    assign layer4_out[7968] = ~layer3_out[5950] | layer3_out[5949];
    assign layer4_out[7969] = ~layer3_out[97];
    assign layer4_out[7970] = layer3_out[6451];
    assign layer4_out[7971] = ~(layer3_out[2433] | layer3_out[2434]);
    assign layer4_out[7972] = ~layer3_out[4];
    assign layer4_out[7973] = ~(layer3_out[7577] ^ layer3_out[7578]);
    assign layer4_out[7974] = layer3_out[2035];
    assign layer4_out[7975] = layer3_out[2428] & layer3_out[2429];
    assign layer4_out[7976] = layer3_out[6891] ^ layer3_out[6892];
    assign layer4_out[7977] = ~layer3_out[2645];
    assign layer4_out[7978] = layer3_out[2484];
    assign layer4_out[7979] = layer3_out[3458];
    assign layer4_out[7980] = layer3_out[3189] | layer3_out[3190];
    assign layer4_out[7981] = ~layer3_out[4531];
    assign layer4_out[7982] = layer3_out[6904];
    assign layer4_out[7983] = ~layer3_out[7625];
    assign layer4_out[7984] = ~layer3_out[5571];
    assign layer4_out[7985] = layer3_out[3884];
    assign layer4_out[7986] = layer3_out[2077];
    assign layer4_out[7987] = layer3_out[1612];
    assign layer4_out[7988] = ~layer3_out[4006] | layer3_out[4005];
    assign layer4_out[7989] = layer3_out[2942] | layer3_out[2943];
    assign layer4_out[7990] = ~layer3_out[7807];
    assign layer4_out[7991] = ~(layer3_out[3123] & layer3_out[3124]);
    assign layer4_out[7992] = layer3_out[1519] ^ layer3_out[1520];
    assign layer4_out[7993] = ~layer3_out[2329];
    assign layer4_out[7994] = layer3_out[7875] | layer3_out[7876];
    assign layer4_out[7995] = layer3_out[190];
    assign layer4_out[7996] = layer3_out[7172] ^ layer3_out[7173];
    assign layer4_out[7997] = layer3_out[1589] | layer3_out[1590];
    assign layer4_out[7998] = ~layer3_out[3610];
    assign layer4_out[7999] = ~layer3_out[1802];
    assign layer5_out[0] = layer4_out[3971];
    assign layer5_out[1] = ~layer4_out[3119];
    assign layer5_out[2] = layer4_out[6604] & ~layer4_out[6605];
    assign layer5_out[3] = layer4_out[340] & ~layer4_out[339];
    assign layer5_out[4] = layer4_out[1405] & layer4_out[1406];
    assign layer5_out[5] = layer4_out[6655];
    assign layer5_out[6] = layer4_out[4883] ^ layer4_out[4884];
    assign layer5_out[7] = ~(layer4_out[827] ^ layer4_out[828]);
    assign layer5_out[8] = ~(layer4_out[1878] & layer4_out[1879]);
    assign layer5_out[9] = ~(layer4_out[1174] | layer4_out[1175]);
    assign layer5_out[10] = layer4_out[5528] | layer4_out[5529];
    assign layer5_out[11] = layer4_out[4400];
    assign layer5_out[12] = layer4_out[1925] ^ layer4_out[1926];
    assign layer5_out[13] = layer4_out[2215] & ~layer4_out[2216];
    assign layer5_out[14] = layer4_out[1672] & layer4_out[1673];
    assign layer5_out[15] = ~layer4_out[4557];
    assign layer5_out[16] = ~(layer4_out[5255] | layer4_out[5256]);
    assign layer5_out[17] = layer4_out[4646];
    assign layer5_out[18] = ~(layer4_out[5142] ^ layer4_out[5143]);
    assign layer5_out[19] = ~layer4_out[6880];
    assign layer5_out[20] = ~layer4_out[3895];
    assign layer5_out[21] = layer4_out[7791];
    assign layer5_out[22] = ~layer4_out[5005];
    assign layer5_out[23] = layer4_out[2397] ^ layer4_out[2398];
    assign layer5_out[24] = layer4_out[484] & ~layer4_out[483];
    assign layer5_out[25] = layer4_out[4113] & layer4_out[4114];
    assign layer5_out[26] = ~layer4_out[2311] | layer4_out[2312];
    assign layer5_out[27] = layer4_out[4035] ^ layer4_out[4036];
    assign layer5_out[28] = ~layer4_out[5486];
    assign layer5_out[29] = ~(layer4_out[1686] ^ layer4_out[1687]);
    assign layer5_out[30] = ~layer4_out[4279];
    assign layer5_out[31] = ~(layer4_out[5789] ^ layer4_out[5790]);
    assign layer5_out[32] = ~(layer4_out[2115] | layer4_out[2116]);
    assign layer5_out[33] = layer4_out[6208] ^ layer4_out[6209];
    assign layer5_out[34] = layer4_out[3465] & ~layer4_out[3464];
    assign layer5_out[35] = ~(layer4_out[7084] & layer4_out[7085]);
    assign layer5_out[36] = ~layer4_out[329];
    assign layer5_out[37] = layer4_out[597];
    assign layer5_out[38] = layer4_out[4680] & layer4_out[4681];
    assign layer5_out[39] = ~layer4_out[4];
    assign layer5_out[40] = layer4_out[1104] ^ layer4_out[1105];
    assign layer5_out[41] = layer4_out[7056];
    assign layer5_out[42] = layer4_out[2416];
    assign layer5_out[43] = layer4_out[7667];
    assign layer5_out[44] = ~layer4_out[3355];
    assign layer5_out[45] = ~(layer4_out[5534] ^ layer4_out[5535]);
    assign layer5_out[46] = layer4_out[3362] & ~layer4_out[3363];
    assign layer5_out[47] = layer4_out[2805];
    assign layer5_out[48] = ~(layer4_out[7308] | layer4_out[7309]);
    assign layer5_out[49] = ~layer4_out[7971];
    assign layer5_out[50] = layer4_out[3748] & layer4_out[3749];
    assign layer5_out[51] = layer4_out[6782] & ~layer4_out[6783];
    assign layer5_out[52] = ~layer4_out[3210];
    assign layer5_out[53] = ~layer4_out[1244];
    assign layer5_out[54] = ~layer4_out[1542] | layer4_out[1541];
    assign layer5_out[55] = layer4_out[2362] | layer4_out[2363];
    assign layer5_out[56] = layer4_out[4104] & ~layer4_out[4103];
    assign layer5_out[57] = layer4_out[6467];
    assign layer5_out[58] = layer4_out[27] ^ layer4_out[28];
    assign layer5_out[59] = ~layer4_out[4152];
    assign layer5_out[60] = layer4_out[1247];
    assign layer5_out[61] = ~layer4_out[5082];
    assign layer5_out[62] = layer4_out[7833];
    assign layer5_out[63] = layer4_out[5710] & layer4_out[5711];
    assign layer5_out[64] = ~layer4_out[6742];
    assign layer5_out[65] = layer4_out[6640];
    assign layer5_out[66] = ~layer4_out[403];
    assign layer5_out[67] = ~(layer4_out[5623] ^ layer4_out[5624]);
    assign layer5_out[68] = ~(layer4_out[241] ^ layer4_out[242]);
    assign layer5_out[69] = layer4_out[3991];
    assign layer5_out[70] = layer4_out[1435];
    assign layer5_out[71] = layer4_out[7127] ^ layer4_out[7128];
    assign layer5_out[72] = ~layer4_out[5257];
    assign layer5_out[73] = layer4_out[6807] & layer4_out[6808];
    assign layer5_out[74] = ~(layer4_out[410] & layer4_out[411]);
    assign layer5_out[75] = layer4_out[956] ^ layer4_out[957];
    assign layer5_out[76] = layer4_out[4975] ^ layer4_out[4976];
    assign layer5_out[77] = layer4_out[4967] & ~layer4_out[4966];
    assign layer5_out[78] = ~(layer4_out[7800] ^ layer4_out[7801]);
    assign layer5_out[79] = ~layer4_out[7335] | layer4_out[7336];
    assign layer5_out[80] = ~layer4_out[5906];
    assign layer5_out[81] = layer4_out[1330];
    assign layer5_out[82] = layer4_out[3001] ^ layer4_out[3002];
    assign layer5_out[83] = layer4_out[5992] ^ layer4_out[5993];
    assign layer5_out[84] = ~(layer4_out[5546] | layer4_out[5547]);
    assign layer5_out[85] = ~layer4_out[1827];
    assign layer5_out[86] = ~(layer4_out[4494] ^ layer4_out[4495]);
    assign layer5_out[87] = layer4_out[3121] & ~layer4_out[3122];
    assign layer5_out[88] = layer4_out[2732] ^ layer4_out[2733];
    assign layer5_out[89] = layer4_out[5204];
    assign layer5_out[90] = ~layer4_out[4480];
    assign layer5_out[91] = ~(layer4_out[6029] | layer4_out[6030]);
    assign layer5_out[92] = layer4_out[1917] & ~layer4_out[1916];
    assign layer5_out[93] = layer4_out[2734] & ~layer4_out[2735];
    assign layer5_out[94] = ~(layer4_out[2989] & layer4_out[2990]);
    assign layer5_out[95] = ~layer4_out[3954];
    assign layer5_out[96] = layer4_out[651];
    assign layer5_out[97] = ~layer4_out[2915];
    assign layer5_out[98] = ~layer4_out[6295];
    assign layer5_out[99] = ~(layer4_out[1594] ^ layer4_out[1595]);
    assign layer5_out[100] = ~(layer4_out[4723] | layer4_out[4724]);
    assign layer5_out[101] = layer4_out[3416] & layer4_out[3417];
    assign layer5_out[102] = ~layer4_out[3407];
    assign layer5_out[103] = layer4_out[7790] & ~layer4_out[7789];
    assign layer5_out[104] = layer4_out[5242] ^ layer4_out[5243];
    assign layer5_out[105] = layer4_out[4216];
    assign layer5_out[106] = ~(layer4_out[5952] & layer4_out[5953]);
    assign layer5_out[107] = layer4_out[5165] & ~layer4_out[5166];
    assign layer5_out[108] = layer4_out[2503] ^ layer4_out[2504];
    assign layer5_out[109] = layer4_out[6195] | layer4_out[6196];
    assign layer5_out[110] = ~layer4_out[313];
    assign layer5_out[111] = ~layer4_out[318];
    assign layer5_out[112] = ~layer4_out[4239] | layer4_out[4240];
    assign layer5_out[113] = layer4_out[1521];
    assign layer5_out[114] = ~layer4_out[2321];
    assign layer5_out[115] = layer4_out[2926] & ~layer4_out[2927];
    assign layer5_out[116] = layer4_out[3475] & ~layer4_out[3474];
    assign layer5_out[117] = layer4_out[6312];
    assign layer5_out[118] = layer4_out[554] ^ layer4_out[555];
    assign layer5_out[119] = layer4_out[6652];
    assign layer5_out[120] = layer4_out[6935] & ~layer4_out[6936];
    assign layer5_out[121] = layer4_out[6280] & ~layer4_out[6281];
    assign layer5_out[122] = layer4_out[5129];
    assign layer5_out[123] = layer4_out[499];
    assign layer5_out[124] = layer4_out[5675] & ~layer4_out[5674];
    assign layer5_out[125] = layer4_out[3221] & layer4_out[3222];
    assign layer5_out[126] = ~layer4_out[6355] | layer4_out[6356];
    assign layer5_out[127] = layer4_out[3815] & ~layer4_out[3816];
    assign layer5_out[128] = layer4_out[6418];
    assign layer5_out[129] = layer4_out[6021] ^ layer4_out[6022];
    assign layer5_out[130] = layer4_out[848];
    assign layer5_out[131] = ~layer4_out[1477] | layer4_out[1478];
    assign layer5_out[132] = layer4_out[3642];
    assign layer5_out[133] = ~layer4_out[7050];
    assign layer5_out[134] = layer4_out[7427] & ~layer4_out[7428];
    assign layer5_out[135] = layer4_out[7929] & layer4_out[7930];
    assign layer5_out[136] = ~(layer4_out[3880] | layer4_out[3881]);
    assign layer5_out[137] = ~(layer4_out[1862] | layer4_out[1863]);
    assign layer5_out[138] = layer4_out[2433] & layer4_out[2434];
    assign layer5_out[139] = ~(layer4_out[1633] ^ layer4_out[1634]);
    assign layer5_out[140] = layer4_out[963] ^ layer4_out[964];
    assign layer5_out[141] = ~layer4_out[5210];
    assign layer5_out[142] = layer4_out[2845];
    assign layer5_out[143] = layer4_out[1228] ^ layer4_out[1229];
    assign layer5_out[144] = layer4_out[7826] & ~layer4_out[7825];
    assign layer5_out[145] = ~layer4_out[4000];
    assign layer5_out[146] = layer4_out[3194] & ~layer4_out[3193];
    assign layer5_out[147] = ~layer4_out[882];
    assign layer5_out[148] = layer4_out[5462] ^ layer4_out[5463];
    assign layer5_out[149] = ~(layer4_out[7510] ^ layer4_out[7511]);
    assign layer5_out[150] = layer4_out[4508] & ~layer4_out[4509];
    assign layer5_out[151] = ~(layer4_out[7139] ^ layer4_out[7140]);
    assign layer5_out[152] = layer4_out[4774] & ~layer4_out[4775];
    assign layer5_out[153] = ~(layer4_out[3131] | layer4_out[3132]);
    assign layer5_out[154] = layer4_out[4024];
    assign layer5_out[155] = ~layer4_out[6657];
    assign layer5_out[156] = layer4_out[7350];
    assign layer5_out[157] = layer4_out[701];
    assign layer5_out[158] = layer4_out[4973] & ~layer4_out[4974];
    assign layer5_out[159] = layer4_out[1036] ^ layer4_out[1037];
    assign layer5_out[160] = layer4_out[6677] ^ layer4_out[6678];
    assign layer5_out[161] = layer4_out[7390];
    assign layer5_out[162] = ~(layer4_out[157] ^ layer4_out[158]);
    assign layer5_out[163] = ~layer4_out[5261];
    assign layer5_out[164] = ~layer4_out[2426];
    assign layer5_out[165] = ~(layer4_out[3827] ^ layer4_out[3828]);
    assign layer5_out[166] = ~(layer4_out[2387] ^ layer4_out[2388]);
    assign layer5_out[167] = layer4_out[925] & ~layer4_out[924];
    assign layer5_out[168] = ~layer4_out[7411];
    assign layer5_out[169] = ~(layer4_out[6861] | layer4_out[6862]);
    assign layer5_out[170] = ~(layer4_out[181] & layer4_out[182]);
    assign layer5_out[171] = ~(layer4_out[4388] ^ layer4_out[4389]);
    assign layer5_out[172] = layer4_out[5236] & ~layer4_out[5235];
    assign layer5_out[173] = ~(layer4_out[7099] | layer4_out[7100]);
    assign layer5_out[174] = ~layer4_out[5771] | layer4_out[5770];
    assign layer5_out[175] = layer4_out[5873] & layer4_out[5874];
    assign layer5_out[176] = layer4_out[4470] ^ layer4_out[4471];
    assign layer5_out[177] = ~(layer4_out[5146] | layer4_out[5147]);
    assign layer5_out[178] = layer4_out[3598] ^ layer4_out[3599];
    assign layer5_out[179] = ~layer4_out[1015];
    assign layer5_out[180] = ~layer4_out[4777];
    assign layer5_out[181] = layer4_out[291] & ~layer4_out[292];
    assign layer5_out[182] = ~layer4_out[108];
    assign layer5_out[183] = ~(layer4_out[3391] ^ layer4_out[3392]);
    assign layer5_out[184] = ~layer4_out[5138];
    assign layer5_out[185] = ~(layer4_out[2642] & layer4_out[2643]);
    assign layer5_out[186] = layer4_out[3409] & ~layer4_out[3410];
    assign layer5_out[187] = ~layer4_out[350];
    assign layer5_out[188] = ~layer4_out[7538] | layer4_out[7539];
    assign layer5_out[189] = ~(layer4_out[7348] ^ layer4_out[7349]);
    assign layer5_out[190] = layer4_out[4141];
    assign layer5_out[191] = layer4_out[4207] ^ layer4_out[4208];
    assign layer5_out[192] = ~(layer4_out[3042] ^ layer4_out[3043]);
    assign layer5_out[193] = layer4_out[7191] & ~layer4_out[7190];
    assign layer5_out[194] = layer4_out[4578] ^ layer4_out[4579];
    assign layer5_out[195] = ~(layer4_out[267] ^ layer4_out[268]);
    assign layer5_out[196] = ~layer4_out[3351] | layer4_out[3352];
    assign layer5_out[197] = layer4_out[7413];
    assign layer5_out[198] = ~layer4_out[1146];
    assign layer5_out[199] = layer4_out[5756] & ~layer4_out[5757];
    assign layer5_out[200] = layer4_out[1465];
    assign layer5_out[201] = ~(layer4_out[4270] ^ layer4_out[4271]);
    assign layer5_out[202] = layer4_out[484] & ~layer4_out[485];
    assign layer5_out[203] = ~layer4_out[6815];
    assign layer5_out[204] = ~(layer4_out[6644] ^ layer4_out[6645]);
    assign layer5_out[205] = ~layer4_out[6943];
    assign layer5_out[206] = ~layer4_out[5250];
    assign layer5_out[207] = layer4_out[3710];
    assign layer5_out[208] = ~(layer4_out[2921] | layer4_out[2922]);
    assign layer5_out[209] = ~layer4_out[4831];
    assign layer5_out[210] = layer4_out[3161];
    assign layer5_out[211] = ~(layer4_out[6613] | layer4_out[6614]);
    assign layer5_out[212] = layer4_out[6121] & layer4_out[6122];
    assign layer5_out[213] = layer4_out[4551] ^ layer4_out[4552];
    assign layer5_out[214] = ~(layer4_out[6507] | layer4_out[6508]);
    assign layer5_out[215] = ~(layer4_out[5929] ^ layer4_out[5930]);
    assign layer5_out[216] = layer4_out[1138];
    assign layer5_out[217] = layer4_out[3665];
    assign layer5_out[218] = ~layer4_out[4999];
    assign layer5_out[219] = ~layer4_out[2682];
    assign layer5_out[220] = ~layer4_out[3622];
    assign layer5_out[221] = layer4_out[1013] & ~layer4_out[1012];
    assign layer5_out[222] = layer4_out[1664] ^ layer4_out[1665];
    assign layer5_out[223] = ~(layer4_out[7140] ^ layer4_out[7141]);
    assign layer5_out[224] = layer4_out[491] ^ layer4_out[492];
    assign layer5_out[225] = ~(layer4_out[7853] | layer4_out[7854]);
    assign layer5_out[226] = ~layer4_out[2459];
    assign layer5_out[227] = layer4_out[226];
    assign layer5_out[228] = layer4_out[1233] ^ layer4_out[1234];
    assign layer5_out[229] = layer4_out[852] & layer4_out[853];
    assign layer5_out[230] = layer4_out[7008] | layer4_out[7009];
    assign layer5_out[231] = ~layer4_out[7837];
    assign layer5_out[232] = ~layer4_out[6835];
    assign layer5_out[233] = ~(layer4_out[682] ^ layer4_out[683]);
    assign layer5_out[234] = layer4_out[6820];
    assign layer5_out[235] = layer4_out[1148] ^ layer4_out[1149];
    assign layer5_out[236] = layer4_out[5645] & ~layer4_out[5646];
    assign layer5_out[237] = layer4_out[2772];
    assign layer5_out[238] = layer4_out[5854] & layer4_out[5855];
    assign layer5_out[239] = ~layer4_out[6042];
    assign layer5_out[240] = ~layer4_out[3523];
    assign layer5_out[241] = ~layer4_out[7812];
    assign layer5_out[242] = layer4_out[5178];
    assign layer5_out[243] = ~(layer4_out[2468] & layer4_out[2469]);
    assign layer5_out[244] = layer4_out[5139] & ~layer4_out[5140];
    assign layer5_out[245] = ~(layer4_out[7420] ^ layer4_out[7421]);
    assign layer5_out[246] = layer4_out[2746];
    assign layer5_out[247] = ~layer4_out[788];
    assign layer5_out[248] = ~layer4_out[338];
    assign layer5_out[249] = layer4_out[7928];
    assign layer5_out[250] = ~(layer4_out[4426] ^ layer4_out[4427]);
    assign layer5_out[251] = ~(layer4_out[7488] ^ layer4_out[7489]);
    assign layer5_out[252] = ~layer4_out[2528];
    assign layer5_out[253] = layer4_out[2834] & ~layer4_out[2835];
    assign layer5_out[254] = ~layer4_out[6572];
    assign layer5_out[255] = ~layer4_out[6018];
    assign layer5_out[256] = ~layer4_out[1164];
    assign layer5_out[257] = ~layer4_out[7062];
    assign layer5_out[258] = layer4_out[6770] & ~layer4_out[6769];
    assign layer5_out[259] = ~layer4_out[7375] | layer4_out[7376];
    assign layer5_out[260] = layer4_out[7429] & ~layer4_out[7428];
    assign layer5_out[261] = layer4_out[5087];
    assign layer5_out[262] = ~(layer4_out[5058] ^ layer4_out[5059]);
    assign layer5_out[263] = layer4_out[624];
    assign layer5_out[264] = ~(layer4_out[6783] & layer4_out[6784]);
    assign layer5_out[265] = ~(layer4_out[4625] ^ layer4_out[4626]);
    assign layer5_out[266] = layer4_out[7472];
    assign layer5_out[267] = layer4_out[7060];
    assign layer5_out[268] = ~layer4_out[7661];
    assign layer5_out[269] = layer4_out[881];
    assign layer5_out[270] = ~layer4_out[641] | layer4_out[642];
    assign layer5_out[271] = layer4_out[222] ^ layer4_out[223];
    assign layer5_out[272] = layer4_out[1083] & ~layer4_out[1082];
    assign layer5_out[273] = ~layer4_out[4792];
    assign layer5_out[274] = layer4_out[7905] ^ layer4_out[7906];
    assign layer5_out[275] = ~(layer4_out[4820] ^ layer4_out[4821]);
    assign layer5_out[276] = ~(layer4_out[5510] ^ layer4_out[5511]);
    assign layer5_out[277] = layer4_out[2802] ^ layer4_out[2803];
    assign layer5_out[278] = ~layer4_out[3759];
    assign layer5_out[279] = ~(layer4_out[6367] ^ layer4_out[6368]);
    assign layer5_out[280] = layer4_out[6490] ^ layer4_out[6491];
    assign layer5_out[281] = ~(layer4_out[5220] & layer4_out[5221]);
    assign layer5_out[282] = layer4_out[5864] & layer4_out[5865];
    assign layer5_out[283] = ~(layer4_out[5887] ^ layer4_out[5888]);
    assign layer5_out[284] = layer4_out[2363] & ~layer4_out[2364];
    assign layer5_out[285] = layer4_out[3957];
    assign layer5_out[286] = layer4_out[3032];
    assign layer5_out[287] = ~(layer4_out[3508] | layer4_out[3509]);
    assign layer5_out[288] = layer4_out[3611];
    assign layer5_out[289] = ~(layer4_out[7690] ^ layer4_out[7691]);
    assign layer5_out[290] = ~layer4_out[352] | layer4_out[353];
    assign layer5_out[291] = ~layer4_out[6026];
    assign layer5_out[292] = ~(layer4_out[3736] | layer4_out[3737]);
    assign layer5_out[293] = ~layer4_out[5684] | layer4_out[5683];
    assign layer5_out[294] = layer4_out[4162];
    assign layer5_out[295] = layer4_out[3709];
    assign layer5_out[296] = ~(layer4_out[7120] ^ layer4_out[7121]);
    assign layer5_out[297] = ~layer4_out[6660];
    assign layer5_out[298] = ~layer4_out[5531];
    assign layer5_out[299] = ~layer4_out[7829];
    assign layer5_out[300] = layer4_out[3710] & ~layer4_out[3711];
    assign layer5_out[301] = layer4_out[5639] ^ layer4_out[5640];
    assign layer5_out[302] = ~(layer4_out[7403] ^ layer4_out[7404]);
    assign layer5_out[303] = ~layer4_out[6950] | layer4_out[6949];
    assign layer5_out[304] = ~layer4_out[3418];
    assign layer5_out[305] = ~layer4_out[1294];
    assign layer5_out[306] = ~layer4_out[5678];
    assign layer5_out[307] = layer4_out[7643];
    assign layer5_out[308] = ~layer4_out[7239];
    assign layer5_out[309] = layer4_out[1780] & ~layer4_out[1779];
    assign layer5_out[310] = ~layer4_out[1014] | layer4_out[1013];
    assign layer5_out[311] = ~layer4_out[2159] | layer4_out[2160];
    assign layer5_out[312] = layer4_out[5200] ^ layer4_out[5201];
    assign layer5_out[313] = layer4_out[3613];
    assign layer5_out[314] = ~layer4_out[2684];
    assign layer5_out[315] = ~layer4_out[4107];
    assign layer5_out[316] = ~layer4_out[333];
    assign layer5_out[317] = layer4_out[2004];
    assign layer5_out[318] = layer4_out[3057] | layer4_out[3058];
    assign layer5_out[319] = layer4_out[753];
    assign layer5_out[320] = layer4_out[1863] ^ layer4_out[1864];
    assign layer5_out[321] = ~(layer4_out[4666] & layer4_out[4667]);
    assign layer5_out[322] = layer4_out[5354] & layer4_out[5355];
    assign layer5_out[323] = ~(layer4_out[7302] ^ layer4_out[7303]);
    assign layer5_out[324] = layer4_out[536];
    assign layer5_out[325] = ~layer4_out[6766];
    assign layer5_out[326] = layer4_out[3225] & ~layer4_out[3226];
    assign layer5_out[327] = layer4_out[3804] & layer4_out[3805];
    assign layer5_out[328] = ~layer4_out[5197];
    assign layer5_out[329] = layer4_out[668];
    assign layer5_out[330] = ~layer4_out[2569];
    assign layer5_out[331] = ~(layer4_out[7434] ^ layer4_out[7435]);
    assign layer5_out[332] = layer4_out[4565];
    assign layer5_out[333] = ~layer4_out[1749] | layer4_out[1748];
    assign layer5_out[334] = ~(layer4_out[1998] ^ layer4_out[1999]);
    assign layer5_out[335] = layer4_out[1198];
    assign layer5_out[336] = ~layer4_out[2694];
    assign layer5_out[337] = layer4_out[7324] & layer4_out[7325];
    assign layer5_out[338] = ~layer4_out[7655];
    assign layer5_out[339] = ~(layer4_out[4419] ^ layer4_out[4420]);
    assign layer5_out[340] = ~layer4_out[4499];
    assign layer5_out[341] = layer4_out[3588];
    assign layer5_out[342] = ~layer4_out[2720] | layer4_out[2721];
    assign layer5_out[343] = layer4_out[4222] ^ layer4_out[4223];
    assign layer5_out[344] = layer4_out[1795];
    assign layer5_out[345] = ~(layer4_out[7951] ^ layer4_out[7952]);
    assign layer5_out[346] = layer4_out[701];
    assign layer5_out[347] = layer4_out[3164] ^ layer4_out[3165];
    assign layer5_out[348] = layer4_out[3136];
    assign layer5_out[349] = layer4_out[5797] ^ layer4_out[5798];
    assign layer5_out[350] = layer4_out[385];
    assign layer5_out[351] = ~layer4_out[5246];
    assign layer5_out[352] = ~layer4_out[950];
    assign layer5_out[353] = ~layer4_out[2438];
    assign layer5_out[354] = ~layer4_out[4124];
    assign layer5_out[355] = layer4_out[1596] | layer4_out[1597];
    assign layer5_out[356] = ~layer4_out[7366] | layer4_out[7365];
    assign layer5_out[357] = layer4_out[4324] ^ layer4_out[4325];
    assign layer5_out[358] = ~layer4_out[3637] | layer4_out[3638];
    assign layer5_out[359] = layer4_out[2606];
    assign layer5_out[360] = ~(layer4_out[806] ^ layer4_out[807]);
    assign layer5_out[361] = ~layer4_out[819];
    assign layer5_out[362] = layer4_out[4265];
    assign layer5_out[363] = ~(layer4_out[6227] ^ layer4_out[6228]);
    assign layer5_out[364] = ~(layer4_out[6173] ^ layer4_out[6174]);
    assign layer5_out[365] = layer4_out[2703] & layer4_out[2704];
    assign layer5_out[366] = ~layer4_out[2094];
    assign layer5_out[367] = layer4_out[2779] & ~layer4_out[2780];
    assign layer5_out[368] = layer4_out[1974];
    assign layer5_out[369] = layer4_out[2237];
    assign layer5_out[370] = layer4_out[3506] & layer4_out[3507];
    assign layer5_out[371] = layer4_out[5711] & layer4_out[5712];
    assign layer5_out[372] = layer4_out[2633] ^ layer4_out[2634];
    assign layer5_out[373] = ~layer4_out[5594] | layer4_out[5595];
    assign layer5_out[374] = ~(layer4_out[5368] ^ layer4_out[5369]);
    assign layer5_out[375] = ~(layer4_out[5028] ^ layer4_out[5029]);
    assign layer5_out[376] = layer4_out[7530] & ~layer4_out[7531];
    assign layer5_out[377] = ~(layer4_out[7101] | layer4_out[7102]);
    assign layer5_out[378] = layer4_out[7798] ^ layer4_out[7799];
    assign layer5_out[379] = layer4_out[3276];
    assign layer5_out[380] = ~layer4_out[4180] | layer4_out[4181];
    assign layer5_out[381] = layer4_out[903];
    assign layer5_out[382] = layer4_out[2746];
    assign layer5_out[383] = layer4_out[2551] & ~layer4_out[2550];
    assign layer5_out[384] = ~(layer4_out[706] ^ layer4_out[707]);
    assign layer5_out[385] = ~layer4_out[3904];
    assign layer5_out[386] = layer4_out[884] & layer4_out[885];
    assign layer5_out[387] = layer4_out[1002];
    assign layer5_out[388] = layer4_out[4800] ^ layer4_out[4801];
    assign layer5_out[389] = layer4_out[2634] & ~layer4_out[2635];
    assign layer5_out[390] = layer4_out[5431] & ~layer4_out[5432];
    assign layer5_out[391] = ~layer4_out[6869];
    assign layer5_out[392] = ~layer4_out[7268] | layer4_out[7269];
    assign layer5_out[393] = layer4_out[1338];
    assign layer5_out[394] = ~(layer4_out[6040] ^ layer4_out[6041]);
    assign layer5_out[395] = ~layer4_out[777];
    assign layer5_out[396] = layer4_out[4642];
    assign layer5_out[397] = layer4_out[5740] ^ layer4_out[5741];
    assign layer5_out[398] = ~layer4_out[5568];
    assign layer5_out[399] = ~layer4_out[6895];
    assign layer5_out[400] = ~(layer4_out[6921] ^ layer4_out[6922]);
    assign layer5_out[401] = ~(layer4_out[1003] | layer4_out[1004]);
    assign layer5_out[402] = layer4_out[3988] & ~layer4_out[3987];
    assign layer5_out[403] = layer4_out[5393];
    assign layer5_out[404] = layer4_out[6533];
    assign layer5_out[405] = layer4_out[4637] & layer4_out[4638];
    assign layer5_out[406] = ~(layer4_out[2010] ^ layer4_out[2011]);
    assign layer5_out[407] = ~(layer4_out[5034] ^ layer4_out[5035]);
    assign layer5_out[408] = ~layer4_out[6022] | layer4_out[6023];
    assign layer5_out[409] = layer4_out[868];
    assign layer5_out[410] = layer4_out[6717] | layer4_out[6718];
    assign layer5_out[411] = ~layer4_out[830];
    assign layer5_out[412] = ~(layer4_out[2586] & layer4_out[2587]);
    assign layer5_out[413] = layer4_out[764];
    assign layer5_out[414] = layer4_out[6356];
    assign layer5_out[415] = ~layer4_out[2737];
    assign layer5_out[416] = layer4_out[2125] & ~layer4_out[2126];
    assign layer5_out[417] = ~(layer4_out[2341] ^ layer4_out[2342]);
    assign layer5_out[418] = layer4_out[3481] & ~layer4_out[3480];
    assign layer5_out[419] = ~layer4_out[3119];
    assign layer5_out[420] = ~(layer4_out[6944] ^ layer4_out[6945]);
    assign layer5_out[421] = ~(layer4_out[4329] & layer4_out[4330]);
    assign layer5_out[422] = ~(layer4_out[1090] ^ layer4_out[1091]);
    assign layer5_out[423] = layer4_out[7466] ^ layer4_out[7467];
    assign layer5_out[424] = layer4_out[4659];
    assign layer5_out[425] = ~layer4_out[5560];
    assign layer5_out[426] = layer4_out[3999] & ~layer4_out[3998];
    assign layer5_out[427] = layer4_out[2132] & ~layer4_out[2133];
    assign layer5_out[428] = ~layer4_out[7444];
    assign layer5_out[429] = ~layer4_out[3093];
    assign layer5_out[430] = ~layer4_out[3497] | layer4_out[3496];
    assign layer5_out[431] = layer4_out[7383];
    assign layer5_out[432] = layer4_out[4394];
    assign layer5_out[433] = layer4_out[2597];
    assign layer5_out[434] = ~(layer4_out[3156] | layer4_out[3157]);
    assign layer5_out[435] = layer4_out[6252] & layer4_out[6253];
    assign layer5_out[436] = ~layer4_out[3359];
    assign layer5_out[437] = layer4_out[7919] & ~layer4_out[7918];
    assign layer5_out[438] = ~(layer4_out[1425] & layer4_out[1426]);
    assign layer5_out[439] = ~(layer4_out[479] ^ layer4_out[480]);
    assign layer5_out[440] = layer4_out[7076];
    assign layer5_out[441] = layer4_out[2099];
    assign layer5_out[442] = ~(layer4_out[703] ^ layer4_out[704]);
    assign layer5_out[443] = layer4_out[290];
    assign layer5_out[444] = layer4_out[4340];
    assign layer5_out[445] = ~layer4_out[2723] | layer4_out[2722];
    assign layer5_out[446] = layer4_out[1618];
    assign layer5_out[447] = ~(layer4_out[3533] ^ layer4_out[3534]);
    assign layer5_out[448] = ~layer4_out[1875];
    assign layer5_out[449] = layer4_out[3371];
    assign layer5_out[450] = layer4_out[3276];
    assign layer5_out[451] = ~layer4_out[1287];
    assign layer5_out[452] = layer4_out[2196] ^ layer4_out[2197];
    assign layer5_out[453] = layer4_out[2980];
    assign layer5_out[454] = layer4_out[7264];
    assign layer5_out[455] = ~(layer4_out[249] ^ layer4_out[250]);
    assign layer5_out[456] = layer4_out[1120] & ~layer4_out[1119];
    assign layer5_out[457] = ~(layer4_out[3380] ^ layer4_out[3381]);
    assign layer5_out[458] = layer4_out[1566] & layer4_out[1567];
    assign layer5_out[459] = ~layer4_out[6130];
    assign layer5_out[460] = layer4_out[160] & ~layer4_out[159];
    assign layer5_out[461] = layer4_out[3018] ^ layer4_out[3019];
    assign layer5_out[462] = layer4_out[7481] ^ layer4_out[7482];
    assign layer5_out[463] = ~layer4_out[1052];
    assign layer5_out[464] = layer4_out[6516];
    assign layer5_out[465] = layer4_out[2938];
    assign layer5_out[466] = layer4_out[5025] ^ layer4_out[5026];
    assign layer5_out[467] = layer4_out[216] & ~layer4_out[217];
    assign layer5_out[468] = layer4_out[2583];
    assign layer5_out[469] = layer4_out[3183] ^ layer4_out[3184];
    assign layer5_out[470] = ~(layer4_out[732] ^ layer4_out[733]);
    assign layer5_out[471] = layer4_out[4715] & ~layer4_out[4714];
    assign layer5_out[472] = ~layer4_out[2092];
    assign layer5_out[473] = layer4_out[2977] ^ layer4_out[2978];
    assign layer5_out[474] = ~layer4_out[7335] | layer4_out[7334];
    assign layer5_out[475] = ~layer4_out[1058] | layer4_out[1057];
    assign layer5_out[476] = ~(layer4_out[4254] & layer4_out[4255]);
    assign layer5_out[477] = layer4_out[6230];
    assign layer5_out[478] = layer4_out[5293] ^ layer4_out[5294];
    assign layer5_out[479] = layer4_out[814] & layer4_out[815];
    assign layer5_out[480] = layer4_out[4421];
    assign layer5_out[481] = layer4_out[7585];
    assign layer5_out[482] = layer4_out[4181] ^ layer4_out[4182];
    assign layer5_out[483] = ~layer4_out[4430] | layer4_out[4431];
    assign layer5_out[484] = layer4_out[5334] | layer4_out[5335];
    assign layer5_out[485] = ~layer4_out[1622];
    assign layer5_out[486] = layer4_out[2774];
    assign layer5_out[487] = ~(layer4_out[907] | layer4_out[908]);
    assign layer5_out[488] = ~(layer4_out[2511] ^ layer4_out[2512]);
    assign layer5_out[489] = layer4_out[28] & ~layer4_out[29];
    assign layer5_out[490] = ~(layer4_out[7721] ^ layer4_out[7722]);
    assign layer5_out[491] = layer4_out[3099];
    assign layer5_out[492] = layer4_out[3829];
    assign layer5_out[493] = layer4_out[5591] & ~layer4_out[5590];
    assign layer5_out[494] = layer4_out[6074];
    assign layer5_out[495] = layer4_out[6232] & ~layer4_out[6233];
    assign layer5_out[496] = layer4_out[3877] | layer4_out[3878];
    assign layer5_out[497] = layer4_out[3829];
    assign layer5_out[498] = ~layer4_out[955] | layer4_out[954];
    assign layer5_out[499] = ~(layer4_out[4201] ^ layer4_out[4202]);
    assign layer5_out[500] = ~(layer4_out[101] ^ layer4_out[102]);
    assign layer5_out[501] = layer4_out[716] ^ layer4_out[717];
    assign layer5_out[502] = layer4_out[4768];
    assign layer5_out[503] = ~layer4_out[3156];
    assign layer5_out[504] = ~layer4_out[1115];
    assign layer5_out[505] = ~(layer4_out[857] ^ layer4_out[858]);
    assign layer5_out[506] = layer4_out[6009];
    assign layer5_out[507] = layer4_out[1921];
    assign layer5_out[508] = ~(layer4_out[5920] & layer4_out[5921]);
    assign layer5_out[509] = layer4_out[3516];
    assign layer5_out[510] = ~layer4_out[7102];
    assign layer5_out[511] = layer4_out[7517] & ~layer4_out[7518];
    assign layer5_out[512] = ~layer4_out[3926];
    assign layer5_out[513] = layer4_out[2302] & ~layer4_out[2301];
    assign layer5_out[514] = ~layer4_out[3577];
    assign layer5_out[515] = ~(layer4_out[3444] ^ layer4_out[3445]);
    assign layer5_out[516] = ~layer4_out[6841];
    assign layer5_out[517] = layer4_out[5341] ^ layer4_out[5342];
    assign layer5_out[518] = layer4_out[4511];
    assign layer5_out[519] = layer4_out[1526];
    assign layer5_out[520] = ~layer4_out[6406];
    assign layer5_out[521] = ~layer4_out[5839];
    assign layer5_out[522] = ~layer4_out[6148] | layer4_out[6147];
    assign layer5_out[523] = layer4_out[7935];
    assign layer5_out[524] = ~layer4_out[771] | layer4_out[772];
    assign layer5_out[525] = layer4_out[2800] & layer4_out[2801];
    assign layer5_out[526] = ~(layer4_out[1997] | layer4_out[1998]);
    assign layer5_out[527] = layer4_out[7307] & ~layer4_out[7308];
    assign layer5_out[528] = layer4_out[3741] & layer4_out[3742];
    assign layer5_out[529] = layer4_out[6798] & ~layer4_out[6797];
    assign layer5_out[530] = layer4_out[2526] | layer4_out[2527];
    assign layer5_out[531] = ~layer4_out[231];
    assign layer5_out[532] = ~layer4_out[3125];
    assign layer5_out[533] = layer4_out[4609];
    assign layer5_out[534] = layer4_out[1665] | layer4_out[1666];
    assign layer5_out[535] = ~(layer4_out[2914] | layer4_out[2915]);
    assign layer5_out[536] = layer4_out[4414];
    assign layer5_out[537] = ~(layer4_out[1046] | layer4_out[1047]);
    assign layer5_out[538] = layer4_out[1632] ^ layer4_out[1633];
    assign layer5_out[539] = layer4_out[570];
    assign layer5_out[540] = ~layer4_out[1899] | layer4_out[1898];
    assign layer5_out[541] = ~layer4_out[7036] | layer4_out[7035];
    assign layer5_out[542] = layer4_out[2862] & ~layer4_out[2863];
    assign layer5_out[543] = ~(layer4_out[5124] & layer4_out[5125]);
    assign layer5_out[544] = layer4_out[1903];
    assign layer5_out[545] = ~(layer4_out[7109] ^ layer4_out[7110]);
    assign layer5_out[546] = ~layer4_out[2438];
    assign layer5_out[547] = ~(layer4_out[4834] ^ layer4_out[4835]);
    assign layer5_out[548] = ~layer4_out[3093];
    assign layer5_out[549] = ~layer4_out[6675];
    assign layer5_out[550] = ~(layer4_out[177] ^ layer4_out[178]);
    assign layer5_out[551] = ~layer4_out[6596];
    assign layer5_out[552] = layer4_out[7680];
    assign layer5_out[553] = ~layer4_out[4516];
    assign layer5_out[554] = layer4_out[980];
    assign layer5_out[555] = layer4_out[5076];
    assign layer5_out[556] = ~layer4_out[4840];
    assign layer5_out[557] = layer4_out[2305] ^ layer4_out[2306];
    assign layer5_out[558] = ~layer4_out[2497];
    assign layer5_out[559] = ~layer4_out[5218];
    assign layer5_out[560] = layer4_out[40];
    assign layer5_out[561] = ~(layer4_out[7958] & layer4_out[7959]);
    assign layer5_out[562] = layer4_out[7327];
    assign layer5_out[563] = ~layer4_out[2089];
    assign layer5_out[564] = ~(layer4_out[7309] ^ layer4_out[7310]);
    assign layer5_out[565] = layer4_out[3466];
    assign layer5_out[566] = ~layer4_out[4772];
    assign layer5_out[567] = ~(layer4_out[5409] ^ layer4_out[5410]);
    assign layer5_out[568] = ~layer4_out[6295];
    assign layer5_out[569] = layer4_out[7928];
    assign layer5_out[570] = layer4_out[7156];
    assign layer5_out[571] = layer4_out[3267] & ~layer4_out[3268];
    assign layer5_out[572] = layer4_out[3796] | layer4_out[3797];
    assign layer5_out[573] = ~(layer4_out[7577] | layer4_out[7578]);
    assign layer5_out[574] = ~layer4_out[553];
    assign layer5_out[575] = ~(layer4_out[4228] & layer4_out[4229]);
    assign layer5_out[576] = layer4_out[5969] & layer4_out[5970];
    assign layer5_out[577] = layer4_out[7859] ^ layer4_out[7860];
    assign layer5_out[578] = layer4_out[4373] & ~layer4_out[4374];
    assign layer5_out[579] = layer4_out[2418] & ~layer4_out[2417];
    assign layer5_out[580] = ~(layer4_out[4717] ^ layer4_out[4718]);
    assign layer5_out[581] = layer4_out[5880] ^ layer4_out[5881];
    assign layer5_out[582] = layer4_out[3591];
    assign layer5_out[583] = layer4_out[4940] ^ layer4_out[4941];
    assign layer5_out[584] = layer4_out[820] & ~layer4_out[819];
    assign layer5_out[585] = layer4_out[2142] ^ layer4_out[2143];
    assign layer5_out[586] = layer4_out[2902] & ~layer4_out[2901];
    assign layer5_out[587] = ~(layer4_out[1419] | layer4_out[1420]);
    assign layer5_out[588] = ~layer4_out[6184] | layer4_out[6183];
    assign layer5_out[589] = ~(layer4_out[6413] ^ layer4_out[6414]);
    assign layer5_out[590] = layer4_out[4954];
    assign layer5_out[591] = ~layer4_out[6428] | layer4_out[6427];
    assign layer5_out[592] = ~layer4_out[610];
    assign layer5_out[593] = ~(layer4_out[3096] | layer4_out[3097]);
    assign layer5_out[594] = ~layer4_out[25];
    assign layer5_out[595] = ~layer4_out[4133];
    assign layer5_out[596] = layer4_out[7823];
    assign layer5_out[597] = ~layer4_out[1244];
    assign layer5_out[598] = layer4_out[5344] & ~layer4_out[5343];
    assign layer5_out[599] = ~(layer4_out[5305] & layer4_out[5306]);
    assign layer5_out[600] = ~(layer4_out[4777] | layer4_out[4778]);
    assign layer5_out[601] = layer4_out[4986] & ~layer4_out[4987];
    assign layer5_out[602] = layer4_out[2124] & ~layer4_out[2123];
    assign layer5_out[603] = ~layer4_out[5132] | layer4_out[5133];
    assign layer5_out[604] = layer4_out[87];
    assign layer5_out[605] = ~(layer4_out[6781] ^ layer4_out[6782]);
    assign layer5_out[606] = layer4_out[160] & layer4_out[161];
    assign layer5_out[607] = layer4_out[5714] & ~layer4_out[5713];
    assign layer5_out[608] = ~layer4_out[3407];
    assign layer5_out[609] = ~(layer4_out[2975] & layer4_out[2976]);
    assign layer5_out[610] = ~layer4_out[6907] | layer4_out[6908];
    assign layer5_out[611] = layer4_out[5940];
    assign layer5_out[612] = layer4_out[6568];
    assign layer5_out[613] = layer4_out[1412] ^ layer4_out[1413];
    assign layer5_out[614] = ~layer4_out[7812];
    assign layer5_out[615] = layer4_out[2293] ^ layer4_out[2294];
    assign layer5_out[616] = layer4_out[5503];
    assign layer5_out[617] = ~layer4_out[2110] | layer4_out[2109];
    assign layer5_out[618] = layer4_out[5822] & ~layer4_out[5823];
    assign layer5_out[619] = ~layer4_out[5008];
    assign layer5_out[620] = ~(layer4_out[7754] ^ layer4_out[7755]);
    assign layer5_out[621] = ~layer4_out[6713] | layer4_out[6712];
    assign layer5_out[622] = ~layer4_out[4770];
    assign layer5_out[623] = layer4_out[1691];
    assign layer5_out[624] = ~(layer4_out[2288] ^ layer4_out[2289]);
    assign layer5_out[625] = layer4_out[6842] ^ layer4_out[6843];
    assign layer5_out[626] = ~layer4_out[2106] | layer4_out[2105];
    assign layer5_out[627] = layer4_out[3507] & ~layer4_out[3508];
    assign layer5_out[628] = layer4_out[4200] & ~layer4_out[4199];
    assign layer5_out[629] = ~(layer4_out[4090] | layer4_out[4091]);
    assign layer5_out[630] = ~layer4_out[6620] | layer4_out[6619];
    assign layer5_out[631] = ~layer4_out[1787];
    assign layer5_out[632] = layer4_out[2558];
    assign layer5_out[633] = ~layer4_out[1219];
    assign layer5_out[634] = ~(layer4_out[5816] & layer4_out[5817]);
    assign layer5_out[635] = ~(layer4_out[7001] ^ layer4_out[7002]);
    assign layer5_out[636] = layer4_out[838] ^ layer4_out[839];
    assign layer5_out[637] = layer4_out[1655];
    assign layer5_out[638] = ~(layer4_out[4982] ^ layer4_out[4983]);
    assign layer5_out[639] = layer4_out[3378];
    assign layer5_out[640] = ~(layer4_out[4535] ^ layer4_out[4536]);
    assign layer5_out[641] = layer4_out[1208];
    assign layer5_out[642] = layer4_out[976];
    assign layer5_out[643] = layer4_out[5558] & ~layer4_out[5557];
    assign layer5_out[644] = layer4_out[3434];
    assign layer5_out[645] = ~layer4_out[4873];
    assign layer5_out[646] = layer4_out[1307] & ~layer4_out[1308];
    assign layer5_out[647] = ~(layer4_out[6338] ^ layer4_out[6339]);
    assign layer5_out[648] = layer4_out[2942] & layer4_out[2943];
    assign layer5_out[649] = ~layer4_out[7627];
    assign layer5_out[650] = layer4_out[6318] & layer4_out[6319];
    assign layer5_out[651] = layer4_out[6381] & ~layer4_out[6380];
    assign layer5_out[652] = layer4_out[7216];
    assign layer5_out[653] = layer4_out[5846];
    assign layer5_out[654] = ~(layer4_out[3803] ^ layer4_out[3804]);
    assign layer5_out[655] = layer4_out[29] ^ layer4_out[30];
    assign layer5_out[656] = ~(layer4_out[6204] ^ layer4_out[6205]);
    assign layer5_out[657] = layer4_out[2491] | layer4_out[2492];
    assign layer5_out[658] = layer4_out[7740] | layer4_out[7741];
    assign layer5_out[659] = ~(layer4_out[5904] & layer4_out[5905]);
    assign layer5_out[660] = ~(layer4_out[5799] ^ layer4_out[5800]);
    assign layer5_out[661] = ~(layer4_out[76] | layer4_out[77]);
    assign layer5_out[662] = layer4_out[4911];
    assign layer5_out[663] = ~layer4_out[7808];
    assign layer5_out[664] = layer4_out[7423];
    assign layer5_out[665] = layer4_out[2537] & ~layer4_out[2536];
    assign layer5_out[666] = ~layer4_out[1377];
    assign layer5_out[667] = layer4_out[5408];
    assign layer5_out[668] = ~layer4_out[4729] | layer4_out[4728];
    assign layer5_out[669] = layer4_out[1969] & ~layer4_out[1968];
    assign layer5_out[670] = ~(layer4_out[5652] ^ layer4_out[5653]);
    assign layer5_out[671] = layer4_out[6391] & ~layer4_out[6392];
    assign layer5_out[672] = ~layer4_out[4677];
    assign layer5_out[673] = layer4_out[1651];
    assign layer5_out[674] = layer4_out[6028] ^ layer4_out[6029];
    assign layer5_out[675] = layer4_out[6296] & ~layer4_out[6297];
    assign layer5_out[676] = ~layer4_out[2343] | layer4_out[2344];
    assign layer5_out[677] = layer4_out[3482];
    assign layer5_out[678] = ~layer4_out[5246];
    assign layer5_out[679] = layer4_out[6499];
    assign layer5_out[680] = layer4_out[3572] | layer4_out[3573];
    assign layer5_out[681] = ~layer4_out[6648] | layer4_out[6649];
    assign layer5_out[682] = layer4_out[2349];
    assign layer5_out[683] = layer4_out[6196];
    assign layer5_out[684] = ~layer4_out[185];
    assign layer5_out[685] = ~layer4_out[2195];
    assign layer5_out[686] = ~layer4_out[1167];
    assign layer5_out[687] = layer4_out[4327] ^ layer4_out[4328];
    assign layer5_out[688] = ~layer4_out[322];
    assign layer5_out[689] = ~layer4_out[3684];
    assign layer5_out[690] = layer4_out[798] & ~layer4_out[799];
    assign layer5_out[691] = layer4_out[6831];
    assign layer5_out[692] = ~layer4_out[7658];
    assign layer5_out[693] = ~layer4_out[106] | layer4_out[107];
    assign layer5_out[694] = layer4_out[2629] & layer4_out[2630];
    assign layer5_out[695] = ~(layer4_out[2538] ^ layer4_out[2539]);
    assign layer5_out[696] = ~layer4_out[6445];
    assign layer5_out[697] = layer4_out[2020] ^ layer4_out[2021];
    assign layer5_out[698] = ~layer4_out[3411] | layer4_out[3412];
    assign layer5_out[699] = ~(layer4_out[4784] & layer4_out[4785]);
    assign layer5_out[700] = ~layer4_out[2828];
    assign layer5_out[701] = ~(layer4_out[3054] ^ layer4_out[3055]);
    assign layer5_out[702] = layer4_out[7186];
    assign layer5_out[703] = ~layer4_out[7730];
    assign layer5_out[704] = layer4_out[7641] & ~layer4_out[7640];
    assign layer5_out[705] = layer4_out[4538];
    assign layer5_out[706] = layer4_out[3933];
    assign layer5_out[707] = layer4_out[3993];
    assign layer5_out[708] = layer4_out[6717];
    assign layer5_out[709] = layer4_out[2119] & layer4_out[2120];
    assign layer5_out[710] = layer4_out[3003] ^ layer4_out[3004];
    assign layer5_out[711] = layer4_out[6649] & ~layer4_out[6650];
    assign layer5_out[712] = ~layer4_out[322];
    assign layer5_out[713] = layer4_out[5067] & ~layer4_out[5066];
    assign layer5_out[714] = layer4_out[5872] & layer4_out[5873];
    assign layer5_out[715] = ~layer4_out[4988];
    assign layer5_out[716] = ~layer4_out[4822] | layer4_out[4823];
    assign layer5_out[717] = ~(layer4_out[4011] ^ layer4_out[4012]);
    assign layer5_out[718] = layer4_out[6637] | layer4_out[6638];
    assign layer5_out[719] = layer4_out[4221] ^ layer4_out[4222];
    assign layer5_out[720] = layer4_out[7014];
    assign layer5_out[721] = layer4_out[7867] & layer4_out[7868];
    assign layer5_out[722] = ~layer4_out[7759] | layer4_out[7758];
    assign layer5_out[723] = layer4_out[7025] & ~layer4_out[7024];
    assign layer5_out[724] = ~layer4_out[231];
    assign layer5_out[725] = ~layer4_out[6720];
    assign layer5_out[726] = ~layer4_out[3904];
    assign layer5_out[727] = layer4_out[355] | layer4_out[356];
    assign layer5_out[728] = ~(layer4_out[7945] & layer4_out[7946]);
    assign layer5_out[729] = layer4_out[681] ^ layer4_out[682];
    assign layer5_out[730] = ~layer4_out[973];
    assign layer5_out[731] = ~(layer4_out[3229] | layer4_out[3230]);
    assign layer5_out[732] = layer4_out[335] & layer4_out[336];
    assign layer5_out[733] = ~layer4_out[3536];
    assign layer5_out[734] = ~layer4_out[5795];
    assign layer5_out[735] = ~layer4_out[4798];
    assign layer5_out[736] = layer4_out[218] & ~layer4_out[217];
    assign layer5_out[737] = layer4_out[5810];
    assign layer5_out[738] = ~layer4_out[582];
    assign layer5_out[739] = layer4_out[3446] & ~layer4_out[3447];
    assign layer5_out[740] = layer4_out[628] & layer4_out[629];
    assign layer5_out[741] = layer4_out[3222] & layer4_out[3223];
    assign layer5_out[742] = layer4_out[7604];
    assign layer5_out[743] = layer4_out[3876] & layer4_out[3877];
    assign layer5_out[744] = ~layer4_out[2402] | layer4_out[2403];
    assign layer5_out[745] = ~layer4_out[2748];
    assign layer5_out[746] = layer4_out[6412];
    assign layer5_out[747] = layer4_out[2042];
    assign layer5_out[748] = layer4_out[3329] ^ layer4_out[3330];
    assign layer5_out[749] = ~layer4_out[7270] | layer4_out[7271];
    assign layer5_out[750] = ~layer4_out[1469];
    assign layer5_out[751] = ~layer4_out[3657] | layer4_out[3656];
    assign layer5_out[752] = ~layer4_out[1064] | layer4_out[1065];
    assign layer5_out[753] = layer4_out[519] ^ layer4_out[520];
    assign layer5_out[754] = layer4_out[5865] & layer4_out[5866];
    assign layer5_out[755] = layer4_out[6346];
    assign layer5_out[756] = ~(layer4_out[1297] ^ layer4_out[1298]);
    assign layer5_out[757] = layer4_out[6506] ^ layer4_out[6507];
    assign layer5_out[758] = ~(layer4_out[1225] & layer4_out[1226]);
    assign layer5_out[759] = layer4_out[4986];
    assign layer5_out[760] = ~(layer4_out[1707] & layer4_out[1708]);
    assign layer5_out[761] = ~(layer4_out[2100] ^ layer4_out[2101]);
    assign layer5_out[762] = layer4_out[1105] | layer4_out[1106];
    assign layer5_out[763] = ~layer4_out[6329];
    assign layer5_out[764] = ~layer4_out[3563];
    assign layer5_out[765] = ~(layer4_out[7028] ^ layer4_out[7029]);
    assign layer5_out[766] = ~(layer4_out[5109] ^ layer4_out[5110]);
    assign layer5_out[767] = layer4_out[7343] ^ layer4_out[7344];
    assign layer5_out[768] = ~layer4_out[7656];
    assign layer5_out[769] = ~(layer4_out[506] | layer4_out[507]);
    assign layer5_out[770] = layer4_out[7822] ^ layer4_out[7823];
    assign layer5_out[771] = layer4_out[6938] & layer4_out[6939];
    assign layer5_out[772] = ~(layer4_out[7245] ^ layer4_out[7246]);
    assign layer5_out[773] = layer4_out[6525];
    assign layer5_out[774] = ~(layer4_out[672] ^ layer4_out[673]);
    assign layer5_out[775] = layer4_out[6213];
    assign layer5_out[776] = layer4_out[704] ^ layer4_out[705];
    assign layer5_out[777] = layer4_out[5896] & ~layer4_out[5895];
    assign layer5_out[778] = layer4_out[42] ^ layer4_out[43];
    assign layer5_out[779] = layer4_out[6824];
    assign layer5_out[780] = ~(layer4_out[7086] ^ layer4_out[7087]);
    assign layer5_out[781] = ~layer4_out[4749];
    assign layer5_out[782] = layer4_out[4632] & layer4_out[4633];
    assign layer5_out[783] = ~(layer4_out[2863] | layer4_out[2864]);
    assign layer5_out[784] = layer4_out[1065];
    assign layer5_out[785] = layer4_out[3032];
    assign layer5_out[786] = layer4_out[2004];
    assign layer5_out[787] = layer4_out[3616];
    assign layer5_out[788] = layer4_out[5076];
    assign layer5_out[789] = ~(layer4_out[2974] ^ layer4_out[2975]);
    assign layer5_out[790] = layer4_out[2250];
    assign layer5_out[791] = layer4_out[6824];
    assign layer5_out[792] = ~layer4_out[7408];
    assign layer5_out[793] = ~layer4_out[2423];
    assign layer5_out[794] = layer4_out[4546];
    assign layer5_out[795] = ~(layer4_out[2786] | layer4_out[2787]);
    assign layer5_out[796] = layer4_out[4613];
    assign layer5_out[797] = ~(layer4_out[5513] ^ layer4_out[5514]);
    assign layer5_out[798] = ~layer4_out[1802];
    assign layer5_out[799] = layer4_out[47];
    assign layer5_out[800] = layer4_out[5195] | layer4_out[5196];
    assign layer5_out[801] = layer4_out[6832] & ~layer4_out[6831];
    assign layer5_out[802] = layer4_out[446] ^ layer4_out[447];
    assign layer5_out[803] = ~layer4_out[7606];
    assign layer5_out[804] = ~(layer4_out[747] | layer4_out[748]);
    assign layer5_out[805] = layer4_out[127] & layer4_out[128];
    assign layer5_out[806] = layer4_out[982] & ~layer4_out[981];
    assign layer5_out[807] = layer4_out[6268] & ~layer4_out[6267];
    assign layer5_out[808] = layer4_out[3071];
    assign layer5_out[809] = ~(layer4_out[52] ^ layer4_out[53]);
    assign layer5_out[810] = ~layer4_out[4966];
    assign layer5_out[811] = ~layer4_out[7336];
    assign layer5_out[812] = ~(layer4_out[7562] ^ layer4_out[7563]);
    assign layer5_out[813] = layer4_out[517] & ~layer4_out[516];
    assign layer5_out[814] = ~(layer4_out[6669] | layer4_out[6670]);
    assign layer5_out[815] = layer4_out[3047] & layer4_out[3048];
    assign layer5_out[816] = layer4_out[5908] ^ layer4_out[5909];
    assign layer5_out[817] = ~(layer4_out[3521] ^ layer4_out[3522]);
    assign layer5_out[818] = layer4_out[4119] ^ layer4_out[4120];
    assign layer5_out[819] = ~layer4_out[1941];
    assign layer5_out[820] = layer4_out[5115] ^ layer4_out[5116];
    assign layer5_out[821] = layer4_out[5808] ^ layer4_out[5809];
    assign layer5_out[822] = ~(layer4_out[1650] ^ layer4_out[1651]);
    assign layer5_out[823] = ~layer4_out[1743];
    assign layer5_out[824] = ~(layer4_out[6784] ^ layer4_out[6785]);
    assign layer5_out[825] = layer4_out[6381];
    assign layer5_out[826] = ~layer4_out[4598];
    assign layer5_out[827] = ~layer4_out[5361];
    assign layer5_out[828] = layer4_out[2378];
    assign layer5_out[829] = layer4_out[6100] ^ layer4_out[6101];
    assign layer5_out[830] = layer4_out[6680];
    assign layer5_out[831] = layer4_out[1131] & ~layer4_out[1130];
    assign layer5_out[832] = ~(layer4_out[6448] ^ layer4_out[6449]);
    assign layer5_out[833] = layer4_out[4556];
    assign layer5_out[834] = ~(layer4_out[5630] ^ layer4_out[5631]);
    assign layer5_out[835] = layer4_out[25] & ~layer4_out[26];
    assign layer5_out[836] = ~layer4_out[198];
    assign layer5_out[837] = layer4_out[6463] ^ layer4_out[6464];
    assign layer5_out[838] = layer4_out[2518];
    assign layer5_out[839] = ~layer4_out[1312] | layer4_out[1311];
    assign layer5_out[840] = layer4_out[762];
    assign layer5_out[841] = layer4_out[4905];
    assign layer5_out[842] = layer4_out[4203];
    assign layer5_out[843] = ~layer4_out[428];
    assign layer5_out[844] = layer4_out[4746] ^ layer4_out[4747];
    assign layer5_out[845] = ~layer4_out[5387];
    assign layer5_out[846] = ~layer4_out[2299];
    assign layer5_out[847] = ~(layer4_out[4976] ^ layer4_out[4977]);
    assign layer5_out[848] = ~layer4_out[7485] | layer4_out[7484];
    assign layer5_out[849] = ~layer4_out[2379];
    assign layer5_out[850] = ~(layer4_out[5260] ^ layer4_out[5261]);
    assign layer5_out[851] = layer4_out[5754] | layer4_out[5755];
    assign layer5_out[852] = ~layer4_out[1446];
    assign layer5_out[853] = ~layer4_out[6429] | layer4_out[6430];
    assign layer5_out[854] = ~layer4_out[6621];
    assign layer5_out[855] = ~layer4_out[2056];
    assign layer5_out[856] = layer4_out[4750];
    assign layer5_out[857] = ~(layer4_out[51] & layer4_out[52]);
    assign layer5_out[858] = ~layer4_out[6288];
    assign layer5_out[859] = ~layer4_out[3795] | layer4_out[3794];
    assign layer5_out[860] = layer4_out[4322] & ~layer4_out[4323];
    assign layer5_out[861] = layer4_out[4751] & ~layer4_out[4752];
    assign layer5_out[862] = layer4_out[93] ^ layer4_out[94];
    assign layer5_out[863] = layer4_out[496] & ~layer4_out[495];
    assign layer5_out[864] = layer4_out[539] & layer4_out[540];
    assign layer5_out[865] = ~layer4_out[2516];
    assign layer5_out[866] = layer4_out[3969] & layer4_out[3970];
    assign layer5_out[867] = layer4_out[6885] ^ layer4_out[6886];
    assign layer5_out[868] = ~(layer4_out[7514] ^ layer4_out[7515]);
    assign layer5_out[869] = layer4_out[1958] ^ layer4_out[1959];
    assign layer5_out[870] = layer4_out[4445] & ~layer4_out[4446];
    assign layer5_out[871] = ~(layer4_out[1076] ^ layer4_out[1077]);
    assign layer5_out[872] = layer4_out[892] & ~layer4_out[893];
    assign layer5_out[873] = layer4_out[6198];
    assign layer5_out[874] = ~layer4_out[6443];
    assign layer5_out[875] = layer4_out[180] ^ layer4_out[181];
    assign layer5_out[876] = layer4_out[1536];
    assign layer5_out[877] = layer4_out[332] & ~layer4_out[331];
    assign layer5_out[878] = layer4_out[1468];
    assign layer5_out[879] = ~layer4_out[1917];
    assign layer5_out[880] = ~layer4_out[1256] | layer4_out[1257];
    assign layer5_out[881] = layer4_out[4471] & layer4_out[4472];
    assign layer5_out[882] = layer4_out[3159];
    assign layer5_out[883] = ~(layer4_out[4286] ^ layer4_out[4287]);
    assign layer5_out[884] = layer4_out[7401] ^ layer4_out[7402];
    assign layer5_out[885] = layer4_out[5628] & layer4_out[5629];
    assign layer5_out[886] = layer4_out[4274] & ~layer4_out[4273];
    assign layer5_out[887] = ~(layer4_out[2031] & layer4_out[2032]);
    assign layer5_out[888] = ~(layer4_out[1447] ^ layer4_out[1448]);
    assign layer5_out[889] = layer4_out[4154] & ~layer4_out[4155];
    assign layer5_out[890] = ~(layer4_out[6694] & layer4_out[6695]);
    assign layer5_out[891] = layer4_out[1203] ^ layer4_out[1204];
    assign layer5_out[892] = ~(layer4_out[6785] | layer4_out[6786]);
    assign layer5_out[893] = layer4_out[5317] ^ layer4_out[5318];
    assign layer5_out[894] = layer4_out[6088];
    assign layer5_out[895] = ~(layer4_out[4348] & layer4_out[4349]);
    assign layer5_out[896] = ~(layer4_out[2313] | layer4_out[2314]);
    assign layer5_out[897] = layer4_out[406] | layer4_out[407];
    assign layer5_out[898] = ~(layer4_out[6809] ^ layer4_out[6810]);
    assign layer5_out[899] = layer4_out[4789];
    assign layer5_out[900] = layer4_out[1252] & layer4_out[1253];
    assign layer5_out[901] = ~layer4_out[2430] | layer4_out[2429];
    assign layer5_out[902] = layer4_out[7036] & layer4_out[7037];
    assign layer5_out[903] = ~layer4_out[4675] | layer4_out[4674];
    assign layer5_out[904] = layer4_out[5447] & ~layer4_out[5448];
    assign layer5_out[905] = layer4_out[1098];
    assign layer5_out[906] = layer4_out[5728];
    assign layer5_out[907] = layer4_out[7815] & ~layer4_out[7816];
    assign layer5_out[908] = layer4_out[7751] & layer4_out[7752];
    assign layer5_out[909] = ~layer4_out[2329] | layer4_out[2328];
    assign layer5_out[910] = layer4_out[6499] ^ layer4_out[6500];
    assign layer5_out[911] = layer4_out[5382];
    assign layer5_out[912] = ~layer4_out[7237] | layer4_out[7238];
    assign layer5_out[913] = layer4_out[6767] ^ layer4_out[6768];
    assign layer5_out[914] = layer4_out[5927] ^ layer4_out[5928];
    assign layer5_out[915] = layer4_out[1644];
    assign layer5_out[916] = ~(layer4_out[6417] ^ layer4_out[6418]);
    assign layer5_out[917] = layer4_out[6882] & ~layer4_out[6883];
    assign layer5_out[918] = ~(layer4_out[3730] ^ layer4_out[3731]);
    assign layer5_out[919] = layer4_out[759] ^ layer4_out[760];
    assign layer5_out[920] = layer4_out[7187] & ~layer4_out[7186];
    assign layer5_out[921] = layer4_out[7691] ^ layer4_out[7692];
    assign layer5_out[922] = layer4_out[4611] ^ layer4_out[4612];
    assign layer5_out[923] = layer4_out[5783];
    assign layer5_out[924] = layer4_out[5162];
    assign layer5_out[925] = layer4_out[5319] ^ layer4_out[5320];
    assign layer5_out[926] = layer4_out[4841];
    assign layer5_out[927] = ~(layer4_out[4917] ^ layer4_out[4918]);
    assign layer5_out[928] = ~layer4_out[6977] | layer4_out[6976];
    assign layer5_out[929] = layer4_out[7885] & ~layer4_out[7884];
    assign layer5_out[930] = ~(layer4_out[7356] ^ layer4_out[7357]);
    assign layer5_out[931] = ~(layer4_out[6538] ^ layer4_out[6539]);
    assign layer5_out[932] = ~layer4_out[2122] | layer4_out[2121];
    assign layer5_out[933] = layer4_out[896] & layer4_out[897];
    assign layer5_out[934] = ~(layer4_out[343] ^ layer4_out[344]);
    assign layer5_out[935] = layer4_out[1396];
    assign layer5_out[936] = ~layer4_out[7980];
    assign layer5_out[937] = layer4_out[20];
    assign layer5_out[938] = layer4_out[7880] ^ layer4_out[7881];
    assign layer5_out[939] = layer4_out[7743];
    assign layer5_out[940] = layer4_out[1719];
    assign layer5_out[941] = ~(layer4_out[2542] | layer4_out[2543]);
    assign layer5_out[942] = layer4_out[7802] ^ layer4_out[7803];
    assign layer5_out[943] = layer4_out[2167];
    assign layer5_out[944] = ~layer4_out[1224];
    assign layer5_out[945] = layer4_out[6202];
    assign layer5_out[946] = ~layer4_out[4074];
    assign layer5_out[947] = layer4_out[3367] ^ layer4_out[3368];
    assign layer5_out[948] = layer4_out[2068];
    assign layer5_out[949] = layer4_out[1159];
    assign layer5_out[950] = layer4_out[5660] ^ layer4_out[5661];
    assign layer5_out[951] = layer4_out[5262] & ~layer4_out[5263];
    assign layer5_out[952] = layer4_out[2749] | layer4_out[2750];
    assign layer5_out[953] = ~layer4_out[6653] | layer4_out[6654];
    assign layer5_out[954] = layer4_out[6951];
    assign layer5_out[955] = layer4_out[7395];
    assign layer5_out[956] = layer4_out[7710] & ~layer4_out[7711];
    assign layer5_out[957] = ~(layer4_out[6264] | layer4_out[6265]);
    assign layer5_out[958] = ~(layer4_out[727] ^ layer4_out[728]);
    assign layer5_out[959] = ~layer4_out[4654] | layer4_out[4655];
    assign layer5_out[960] = ~layer4_out[3201];
    assign layer5_out[961] = layer4_out[6699] & ~layer4_out[6700];
    assign layer5_out[962] = layer4_out[5077] ^ layer4_out[5078];
    assign layer5_out[963] = layer4_out[1536];
    assign layer5_out[964] = layer4_out[7866];
    assign layer5_out[965] = ~(layer4_out[1605] | layer4_out[1606]);
    assign layer5_out[966] = layer4_out[3518];
    assign layer5_out[967] = layer4_out[3985];
    assign layer5_out[968] = ~layer4_out[5349] | layer4_out[5348];
    assign layer5_out[969] = ~(layer4_out[7578] ^ layer4_out[7579]);
    assign layer5_out[970] = layer4_out[4670] ^ layer4_out[4671];
    assign layer5_out[971] = ~layer4_out[6681];
    assign layer5_out[972] = ~layer4_out[4243];
    assign layer5_out[973] = layer4_out[3214] & ~layer4_out[3213];
    assign layer5_out[974] = layer4_out[4235];
    assign layer5_out[975] = ~layer4_out[1506];
    assign layer5_out[976] = ~layer4_out[5228];
    assign layer5_out[977] = layer4_out[5078] | layer4_out[5079];
    assign layer5_out[978] = ~(layer4_out[1575] & layer4_out[1576]);
    assign layer5_out[979] = layer4_out[2326];
    assign layer5_out[980] = layer4_out[3086] ^ layer4_out[3087];
    assign layer5_out[981] = ~(layer4_out[5470] | layer4_out[5471]);
    assign layer5_out[982] = layer4_out[1258] ^ layer4_out[1259];
    assign layer5_out[983] = layer4_out[2923];
    assign layer5_out[984] = layer4_out[4861] ^ layer4_out[4862];
    assign layer5_out[985] = layer4_out[3071] & ~layer4_out[3070];
    assign layer5_out[986] = ~layer4_out[6536];
    assign layer5_out[987] = ~layer4_out[800];
    assign layer5_out[988] = layer4_out[1683] ^ layer4_out[1684];
    assign layer5_out[989] = layer4_out[4012] & layer4_out[4013];
    assign layer5_out[990] = ~(layer4_out[125] | layer4_out[126]);
    assign layer5_out[991] = ~layer4_out[804];
    assign layer5_out[992] = ~(layer4_out[1710] | layer4_out[1711]);
    assign layer5_out[993] = ~layer4_out[4484] | layer4_out[4483];
    assign layer5_out[994] = layer4_out[4553];
    assign layer5_out[995] = layer4_out[2931] & ~layer4_out[2932];
    assign layer5_out[996] = ~(layer4_out[2625] | layer4_out[2626]);
    assign layer5_out[997] = layer4_out[4361] ^ layer4_out[4362];
    assign layer5_out[998] = layer4_out[233] ^ layer4_out[234];
    assign layer5_out[999] = layer4_out[5643] ^ layer4_out[5644];
    assign layer5_out[1000] = ~layer4_out[6436];
    assign layer5_out[1001] = layer4_out[4010] & ~layer4_out[4011];
    assign layer5_out[1002] = ~(layer4_out[4122] ^ layer4_out[4123]);
    assign layer5_out[1003] = layer4_out[6984];
    assign layer5_out[1004] = layer4_out[3528];
    assign layer5_out[1005] = layer4_out[826] ^ layer4_out[827];
    assign layer5_out[1006] = layer4_out[7698] & layer4_out[7699];
    assign layer5_out[1007] = layer4_out[1931];
    assign layer5_out[1008] = layer4_out[3973] & ~layer4_out[3972];
    assign layer5_out[1009] = ~(layer4_out[1770] ^ layer4_out[1771]);
    assign layer5_out[1010] = ~layer4_out[4263] | layer4_out[4262];
    assign layer5_out[1011] = layer4_out[4719];
    assign layer5_out[1012] = layer4_out[6070];
    assign layer5_out[1013] = layer4_out[4378] ^ layer4_out[4379];
    assign layer5_out[1014] = layer4_out[3176];
    assign layer5_out[1015] = layer4_out[3594] & ~layer4_out[3593];
    assign layer5_out[1016] = ~(layer4_out[2441] ^ layer4_out[2442]);
    assign layer5_out[1017] = layer4_out[5543] ^ layer4_out[5544];
    assign layer5_out[1018] = ~(layer4_out[3671] ^ layer4_out[3672]);
    assign layer5_out[1019] = layer4_out[7027];
    assign layer5_out[1020] = layer4_out[409] & layer4_out[410];
    assign layer5_out[1021] = layer4_out[4607] & ~layer4_out[4606];
    assign layer5_out[1022] = layer4_out[3075] ^ layer4_out[3076];
    assign layer5_out[1023] = ~(layer4_out[7683] | layer4_out[7684]);
    assign layer5_out[1024] = ~(layer4_out[7718] ^ layer4_out[7719]);
    assign layer5_out[1025] = ~layer4_out[2715] | layer4_out[2714];
    assign layer5_out[1026] = layer4_out[4872];
    assign layer5_out[1027] = layer4_out[749] & ~layer4_out[750];
    assign layer5_out[1028] = layer4_out[6179] ^ layer4_out[6180];
    assign layer5_out[1029] = layer4_out[6973] | layer4_out[6974];
    assign layer5_out[1030] = layer4_out[2553];
    assign layer5_out[1031] = layer4_out[1196] ^ layer4_out[1197];
    assign layer5_out[1032] = layer4_out[3566] ^ layer4_out[3567];
    assign layer5_out[1033] = layer4_out[4627] ^ layer4_out[4628];
    assign layer5_out[1034] = ~(layer4_out[1328] & layer4_out[1329]);
    assign layer5_out[1035] = layer4_out[5957];
    assign layer5_out[1036] = layer4_out[3341];
    assign layer5_out[1037] = layer4_out[1810] & ~layer4_out[1809];
    assign layer5_out[1038] = layer4_out[351];
    assign layer5_out[1039] = layer4_out[4384];
    assign layer5_out[1040] = layer4_out[969] & layer4_out[970];
    assign layer5_out[1041] = ~(layer4_out[416] ^ layer4_out[417]);
    assign layer5_out[1042] = ~(layer4_out[2254] | layer4_out[2255]);
    assign layer5_out[1043] = ~layer4_out[3849];
    assign layer5_out[1044] = layer4_out[3921];
    assign layer5_out[1045] = layer4_out[6905] & ~layer4_out[6906];
    assign layer5_out[1046] = layer4_out[3530] ^ layer4_out[3531];
    assign layer5_out[1047] = layer4_out[124] & ~layer4_out[125];
    assign layer5_out[1048] = layer4_out[2455];
    assign layer5_out[1049] = layer4_out[1904];
    assign layer5_out[1050] = ~(layer4_out[3625] ^ layer4_out[3626]);
    assign layer5_out[1051] = layer4_out[4338];
    assign layer5_out[1052] = layer4_out[5159];
    assign layer5_out[1053] = layer4_out[7001] & ~layer4_out[7000];
    assign layer5_out[1054] = ~(layer4_out[4137] | layer4_out[4138]);
    assign layer5_out[1055] = ~(layer4_out[1240] ^ layer4_out[1241]);
    assign layer5_out[1056] = ~layer4_out[5352];
    assign layer5_out[1057] = ~layer4_out[4700];
    assign layer5_out[1058] = layer4_out[1031] & layer4_out[1032];
    assign layer5_out[1059] = ~(layer4_out[6739] ^ layer4_out[6740]);
    assign layer5_out[1060] = ~layer4_out[1962];
    assign layer5_out[1061] = layer4_out[6190] & ~layer4_out[6189];
    assign layer5_out[1062] = ~layer4_out[4963];
    assign layer5_out[1063] = layer4_out[5332];
    assign layer5_out[1064] = layer4_out[2565] ^ layer4_out[2566];
    assign layer5_out[1065] = layer4_out[829];
    assign layer5_out[1066] = layer4_out[2072];
    assign layer5_out[1067] = layer4_out[7664] & layer4_out[7665];
    assign layer5_out[1068] = layer4_out[6790];
    assign layer5_out[1069] = layer4_out[282] ^ layer4_out[283];
    assign layer5_out[1070] = layer4_out[7060];
    assign layer5_out[1071] = ~(layer4_out[1125] ^ layer4_out[1126]);
    assign layer5_out[1072] = layer4_out[2834] & ~layer4_out[2833];
    assign layer5_out[1073] = ~(layer4_out[6142] ^ layer4_out[6143]);
    assign layer5_out[1074] = layer4_out[1688] ^ layer4_out[1689];
    assign layer5_out[1075] = layer4_out[2017] & ~layer4_out[2018];
    assign layer5_out[1076] = layer4_out[6335] ^ layer4_out[6336];
    assign layer5_out[1077] = ~(layer4_out[5031] ^ layer4_out[5032]);
    assign layer5_out[1078] = layer4_out[4539] & layer4_out[4540];
    assign layer5_out[1079] = ~(layer4_out[58] ^ layer4_out[59]);
    assign layer5_out[1080] = ~layer4_out[3368];
    assign layer5_out[1081] = ~layer4_out[6599];
    assign layer5_out[1082] = ~(layer4_out[3090] ^ layer4_out[3091]);
    assign layer5_out[1083] = layer4_out[5247];
    assign layer5_out[1084] = ~(layer4_out[4028] ^ layer4_out[4029]);
    assign layer5_out[1085] = layer4_out[6732] & ~layer4_out[6733];
    assign layer5_out[1086] = ~layer4_out[722];
    assign layer5_out[1087] = ~(layer4_out[1183] ^ layer4_out[1184]);
    assign layer5_out[1088] = ~layer4_out[2310];
    assign layer5_out[1089] = ~layer4_out[7973];
    assign layer5_out[1090] = layer4_out[5742];
    assign layer5_out[1091] = ~(layer4_out[1948] ^ layer4_out[1949]);
    assign layer5_out[1092] = ~layer4_out[1370];
    assign layer5_out[1093] = layer4_out[2005] ^ layer4_out[2006];
    assign layer5_out[1094] = layer4_out[5525];
    assign layer5_out[1095] = ~layer4_out[310] | layer4_out[309];
    assign layer5_out[1096] = ~(layer4_out[1249] ^ layer4_out[1250]);
    assign layer5_out[1097] = ~(layer4_out[5184] ^ layer4_out[5185]);
    assign layer5_out[1098] = ~layer4_out[4909];
    assign layer5_out[1099] = ~(layer4_out[3747] ^ layer4_out[3748]);
    assign layer5_out[1100] = ~layer4_out[1971] | layer4_out[1970];
    assign layer5_out[1101] = layer4_out[38] ^ layer4_out[39];
    assign layer5_out[1102] = ~(layer4_out[1369] & layer4_out[1370]);
    assign layer5_out[1103] = layer4_out[3969];
    assign layer5_out[1104] = ~layer4_out[1661];
    assign layer5_out[1105] = ~layer4_out[7497];
    assign layer5_out[1106] = ~(layer4_out[4682] ^ layer4_out[4683]);
    assign layer5_out[1107] = layer4_out[3123] & ~layer4_out[3122];
    assign layer5_out[1108] = ~layer4_out[6879];
    assign layer5_out[1109] = ~layer4_out[4863];
    assign layer5_out[1110] = layer4_out[43];
    assign layer5_out[1111] = layer4_out[6207] ^ layer4_out[6208];
    assign layer5_out[1112] = layer4_out[5918];
    assign layer5_out[1113] = ~(layer4_out[1334] ^ layer4_out[1335]);
    assign layer5_out[1114] = layer4_out[7174] ^ layer4_out[7175];
    assign layer5_out[1115] = ~layer4_out[2506];
    assign layer5_out[1116] = ~(layer4_out[5675] | layer4_out[5676]);
    assign layer5_out[1117] = layer4_out[108] & ~layer4_out[109];
    assign layer5_out[1118] = ~layer4_out[6294];
    assign layer5_out[1119] = ~layer4_out[4677] | layer4_out[4676];
    assign layer5_out[1120] = layer4_out[1462] & ~layer4_out[1463];
    assign layer5_out[1121] = layer4_out[5664] & ~layer4_out[5665];
    assign layer5_out[1122] = ~(layer4_out[6316] ^ layer4_out[6317]);
    assign layer5_out[1123] = layer4_out[3681] & ~layer4_out[3680];
    assign layer5_out[1124] = layer4_out[3281];
    assign layer5_out[1125] = ~(layer4_out[1564] ^ layer4_out[1565]);
    assign layer5_out[1126] = layer4_out[2986] ^ layer4_out[2987];
    assign layer5_out[1127] = layer4_out[1331] | layer4_out[1332];
    assign layer5_out[1128] = layer4_out[7354];
    assign layer5_out[1129] = ~layer4_out[5724];
    assign layer5_out[1130] = layer4_out[1116] & layer4_out[1117];
    assign layer5_out[1131] = ~layer4_out[5815] | layer4_out[5814];
    assign layer5_out[1132] = layer4_out[960] ^ layer4_out[961];
    assign layer5_out[1133] = ~(layer4_out[2617] ^ layer4_out[2618]);
    assign layer5_out[1134] = ~(layer4_out[5995] & layer4_out[5996]);
    assign layer5_out[1135] = ~(layer4_out[4935] | layer4_out[4936]);
    assign layer5_out[1136] = layer4_out[1726] ^ layer4_out[1727];
    assign layer5_out[1137] = layer4_out[6359] & ~layer4_out[6360];
    assign layer5_out[1138] = layer4_out[2945] & layer4_out[2946];
    assign layer5_out[1139] = ~layer4_out[1333];
    assign layer5_out[1140] = layer4_out[2221] ^ layer4_out[2222];
    assign layer5_out[1141] = layer4_out[3973] | layer4_out[3974];
    assign layer5_out[1142] = layer4_out[5392];
    assign layer5_out[1143] = layer4_out[7723] ^ layer4_out[7724];
    assign layer5_out[1144] = ~layer4_out[2375];
    assign layer5_out[1145] = layer4_out[4047];
    assign layer5_out[1146] = layer4_out[3163] ^ layer4_out[3164];
    assign layer5_out[1147] = ~(layer4_out[4223] ^ layer4_out[4224]);
    assign layer5_out[1148] = layer4_out[590] & layer4_out[591];
    assign layer5_out[1149] = layer4_out[4816];
    assign layer5_out[1150] = ~layer4_out[3689];
    assign layer5_out[1151] = ~(layer4_out[3357] ^ layer4_out[3358]);
    assign layer5_out[1152] = layer4_out[143];
    assign layer5_out[1153] = ~(layer4_out[4531] | layer4_out[4532]);
    assign layer5_out[1154] = layer4_out[2453];
    assign layer5_out[1155] = ~layer4_out[1680];
    assign layer5_out[1156] = ~layer4_out[3666];
    assign layer5_out[1157] = layer4_out[3273] & layer4_out[3274];
    assign layer5_out[1158] = layer4_out[964] & layer4_out[965];
    assign layer5_out[1159] = layer4_out[799] & ~layer4_out[800];
    assign layer5_out[1160] = layer4_out[4853] ^ layer4_out[4854];
    assign layer5_out[1161] = layer4_out[3265];
    assign layer5_out[1162] = ~layer4_out[5089];
    assign layer5_out[1163] = layer4_out[6250] ^ layer4_out[6251];
    assign layer5_out[1164] = ~(layer4_out[976] ^ layer4_out[977]);
    assign layer5_out[1165] = ~(layer4_out[3955] ^ layer4_out[3956]);
    assign layer5_out[1166] = ~layer4_out[2497] | layer4_out[2496];
    assign layer5_out[1167] = layer4_out[1339] ^ layer4_out[1340];
    assign layer5_out[1168] = ~layer4_out[4468];
    assign layer5_out[1169] = ~(layer4_out[1430] ^ layer4_out[1431]);
    assign layer5_out[1170] = ~layer4_out[7178];
    assign layer5_out[1171] = layer4_out[5210];
    assign layer5_out[1172] = ~(layer4_out[821] | layer4_out[822]);
    assign layer5_out[1173] = layer4_out[6546] ^ layer4_out[6547];
    assign layer5_out[1174] = layer4_out[1764] ^ layer4_out[1765];
    assign layer5_out[1175] = ~(layer4_out[2490] ^ layer4_out[2491]);
    assign layer5_out[1176] = ~(layer4_out[2217] | layer4_out[2218]);
    assign layer5_out[1177] = layer4_out[2029] & layer4_out[2030];
    assign layer5_out[1178] = ~layer4_out[5591] | layer4_out[5592];
    assign layer5_out[1179] = ~layer4_out[6522];
    assign layer5_out[1180] = layer4_out[144];
    assign layer5_out[1181] = layer4_out[6985] & ~layer4_out[6986];
    assign layer5_out[1182] = ~(layer4_out[541] | layer4_out[542]);
    assign layer5_out[1183] = layer4_out[6470];
    assign layer5_out[1184] = layer4_out[6276] & ~layer4_out[6275];
    assign layer5_out[1185] = layer4_out[6537] ^ layer4_out[6538];
    assign layer5_out[1186] = layer4_out[2381] & ~layer4_out[2380];
    assign layer5_out[1187] = layer4_out[176];
    assign layer5_out[1188] = ~(layer4_out[5859] ^ layer4_out[5860]);
    assign layer5_out[1189] = layer4_out[4435] ^ layer4_out[4436];
    assign layer5_out[1190] = layer4_out[2443];
    assign layer5_out[1191] = ~layer4_out[3902];
    assign layer5_out[1192] = layer4_out[4578];
    assign layer5_out[1193] = layer4_out[3570] & ~layer4_out[3569];
    assign layer5_out[1194] = layer4_out[3030] ^ layer4_out[3031];
    assign layer5_out[1195] = ~layer4_out[6145];
    assign layer5_out[1196] = ~(layer4_out[6886] ^ layer4_out[6887]);
    assign layer5_out[1197] = ~(layer4_out[3561] ^ layer4_out[3562]);
    assign layer5_out[1198] = ~layer4_out[1819];
    assign layer5_out[1199] = layer4_out[6581];
    assign layer5_out[1200] = ~(layer4_out[2976] | layer4_out[2977]);
    assign layer5_out[1201] = layer4_out[7073];
    assign layer5_out[1202] = ~(layer4_out[5796] | layer4_out[5797]);
    assign layer5_out[1203] = layer4_out[5837] & ~layer4_out[5838];
    assign layer5_out[1204] = layer4_out[7143];
    assign layer5_out[1205] = layer4_out[431] ^ layer4_out[432];
    assign layer5_out[1206] = layer4_out[2222] ^ layer4_out[2223];
    assign layer5_out[1207] = layer4_out[7646] ^ layer4_out[7647];
    assign layer5_out[1208] = layer4_out[7393] & ~layer4_out[7392];
    assign layer5_out[1209] = layer4_out[2249];
    assign layer5_out[1210] = ~(layer4_out[4763] | layer4_out[4764]);
    assign layer5_out[1211] = ~(layer4_out[2624] ^ layer4_out[2625]);
    assign layer5_out[1212] = ~(layer4_out[4860] & layer4_out[4861]);
    assign layer5_out[1213] = ~(layer4_out[2668] ^ layer4_out[2669]);
    assign layer5_out[1214] = layer4_out[3307] ^ layer4_out[3308];
    assign layer5_out[1215] = layer4_out[3230];
    assign layer5_out[1216] = layer4_out[4156] & ~layer4_out[4157];
    assign layer5_out[1217] = ~(layer4_out[5472] | layer4_out[5473]);
    assign layer5_out[1218] = ~(layer4_out[7689] ^ layer4_out[7690]);
    assign layer5_out[1219] = layer4_out[2700] | layer4_out[2701];
    assign layer5_out[1220] = ~layer4_out[944];
    assign layer5_out[1221] = layer4_out[658] & ~layer4_out[657];
    assign layer5_out[1222] = layer4_out[4643] & ~layer4_out[4642];
    assign layer5_out[1223] = layer4_out[5063];
    assign layer5_out[1224] = ~layer4_out[60];
    assign layer5_out[1225] = layer4_out[5892] ^ layer4_out[5893];
    assign layer5_out[1226] = layer4_out[1923] & ~layer4_out[1924];
    assign layer5_out[1227] = ~layer4_out[529];
    assign layer5_out[1228] = layer4_out[4205] & layer4_out[4206];
    assign layer5_out[1229] = layer4_out[5155] & layer4_out[5156];
    assign layer5_out[1230] = ~(layer4_out[5977] | layer4_out[5978]);
    assign layer5_out[1231] = ~(layer4_out[5147] ^ layer4_out[5148]);
    assign layer5_out[1232] = ~layer4_out[7960];
    assign layer5_out[1233] = layer4_out[7634] & ~layer4_out[7635];
    assign layer5_out[1234] = layer4_out[1017] & ~layer4_out[1016];
    assign layer5_out[1235] = layer4_out[1101];
    assign layer5_out[1236] = layer4_out[4464] & ~layer4_out[4465];
    assign layer5_out[1237] = ~layer4_out[4360];
    assign layer5_out[1238] = ~layer4_out[3621];
    assign layer5_out[1239] = layer4_out[2295];
    assign layer5_out[1240] = ~(layer4_out[5540] | layer4_out[5541]);
    assign layer5_out[1241] = ~(layer4_out[6257] | layer4_out[6258]);
    assign layer5_out[1242] = ~(layer4_out[3575] ^ layer4_out[3576]);
    assign layer5_out[1243] = ~(layer4_out[1635] ^ layer4_out[1636]);
    assign layer5_out[1244] = ~layer4_out[1674];
    assign layer5_out[1245] = ~(layer4_out[7508] ^ layer4_out[7509]);
    assign layer5_out[1246] = layer4_out[1219];
    assign layer5_out[1247] = ~(layer4_out[3913] ^ layer4_out[3914]);
    assign layer5_out[1248] = ~(layer4_out[7944] ^ layer4_out[7945]);
    assign layer5_out[1249] = ~(layer4_out[7075] ^ layer4_out[7076]);
    assign layer5_out[1250] = layer4_out[5855] & ~layer4_out[5856];
    assign layer5_out[1251] = layer4_out[4516];
    assign layer5_out[1252] = ~layer4_out[3346] | layer4_out[3345];
    assign layer5_out[1253] = layer4_out[3930] & ~layer4_out[3929];
    assign layer5_out[1254] = ~(layer4_out[7735] | layer4_out[7736]);
    assign layer5_out[1255] = ~(layer4_out[5937] ^ layer4_out[5938]);
    assign layer5_out[1256] = layer4_out[472] & ~layer4_out[473];
    assign layer5_out[1257] = layer4_out[5617];
    assign layer5_out[1258] = layer4_out[7280];
    assign layer5_out[1259] = layer4_out[1704] & ~layer4_out[1705];
    assign layer5_out[1260] = layer4_out[2940] & layer4_out[2941];
    assign layer5_out[1261] = ~(layer4_out[303] ^ layer4_out[304]);
    assign layer5_out[1262] = ~layer4_out[4596];
    assign layer5_out[1263] = ~(layer4_out[696] ^ layer4_out[697]);
    assign layer5_out[1264] = layer4_out[7021] & ~layer4_out[7022];
    assign layer5_out[1265] = layer4_out[1342];
    assign layer5_out[1266] = ~layer4_out[558];
    assign layer5_out[1267] = ~layer4_out[6630];
    assign layer5_out[1268] = layer4_out[2150] ^ layer4_out[2151];
    assign layer5_out[1269] = layer4_out[5638];
    assign layer5_out[1270] = layer4_out[2365];
    assign layer5_out[1271] = layer4_out[6889] & ~layer4_out[6890];
    assign layer5_out[1272] = ~(layer4_out[7301] ^ layer4_out[7302]);
    assign layer5_out[1273] = layer4_out[1545];
    assign layer5_out[1274] = layer4_out[4865] & ~layer4_out[4864];
    assign layer5_out[1275] = layer4_out[6428] & ~layer4_out[6429];
    assign layer5_out[1276] = layer4_out[4066];
    assign layer5_out[1277] = ~(layer4_out[7318] ^ layer4_out[7319]);
    assign layer5_out[1278] = layer4_out[1491] | layer4_out[1492];
    assign layer5_out[1279] = ~(layer4_out[1028] ^ layer4_out[1029]);
    assign layer5_out[1280] = layer4_out[7418];
    assign layer5_out[1281] = ~(layer4_out[3493] & layer4_out[3494]);
    assign layer5_out[1282] = layer4_out[965] ^ layer4_out[966];
    assign layer5_out[1283] = ~(layer4_out[3256] | layer4_out[3257]);
    assign layer5_out[1284] = layer4_out[2290];
    assign layer5_out[1285] = ~(layer4_out[4875] ^ layer4_out[4876]);
    assign layer5_out[1286] = ~(layer4_out[5405] | layer4_out[5406]);
    assign layer5_out[1287] = ~layer4_out[1861] | layer4_out[1862];
    assign layer5_out[1288] = ~(layer4_out[5573] ^ layer4_out[5574]);
    assign layer5_out[1289] = layer4_out[7145] ^ layer4_out[7146];
    assign layer5_out[1290] = ~(layer4_out[807] | layer4_out[808]);
    assign layer5_out[1291] = ~layer4_out[6375];
    assign layer5_out[1292] = layer4_out[6454] & ~layer4_out[6455];
    assign layer5_out[1293] = layer4_out[3147];
    assign layer5_out[1294] = ~layer4_out[2907] | layer4_out[2908];
    assign layer5_out[1295] = ~layer4_out[7160] | layer4_out[7159];
    assign layer5_out[1296] = layer4_out[6465] ^ layer4_out[6466];
    assign layer5_out[1297] = layer4_out[5506];
    assign layer5_out[1298] = ~layer4_out[3475] | layer4_out[3476];
    assign layer5_out[1299] = ~layer4_out[1786] | layer4_out[1785];
    assign layer5_out[1300] = layer4_out[5867] & ~layer4_out[5868];
    assign layer5_out[1301] = layer4_out[4855] ^ layer4_out[4856];
    assign layer5_out[1302] = ~(layer4_out[6031] | layer4_out[6032]);
    assign layer5_out[1303] = ~layer4_out[1383];
    assign layer5_out[1304] = layer4_out[2453];
    assign layer5_out[1305] = ~(layer4_out[2025] ^ layer4_out[2026]);
    assign layer5_out[1306] = ~(layer4_out[7705] ^ layer4_out[7706]);
    assign layer5_out[1307] = ~(layer4_out[6185] ^ layer4_out[6186]);
    assign layer5_out[1308] = layer4_out[6314];
    assign layer5_out[1309] = layer4_out[6741] ^ layer4_out[6742];
    assign layer5_out[1310] = layer4_out[7363];
    assign layer5_out[1311] = layer4_out[5730] ^ layer4_out[5731];
    assign layer5_out[1312] = layer4_out[4417] & layer4_out[4418];
    assign layer5_out[1313] = ~layer4_out[7403] | layer4_out[7402];
    assign layer5_out[1314] = layer4_out[265] & ~layer4_out[264];
    assign layer5_out[1315] = layer4_out[4229] & layer4_out[4230];
    assign layer5_out[1316] = ~(layer4_out[2317] | layer4_out[2318]);
    assign layer5_out[1317] = ~layer4_out[4192];
    assign layer5_out[1318] = layer4_out[1512] & ~layer4_out[1513];
    assign layer5_out[1319] = ~(layer4_out[3427] | layer4_out[3428]);
    assign layer5_out[1320] = ~(layer4_out[468] ^ layer4_out[469]);
    assign layer5_out[1321] = layer4_out[4786] & ~layer4_out[4785];
    assign layer5_out[1322] = ~layer4_out[5533];
    assign layer5_out[1323] = layer4_out[725] & layer4_out[726];
    assign layer5_out[1324] = layer4_out[3808];
    assign layer5_out[1325] = layer4_out[7249] ^ layer4_out[7250];
    assign layer5_out[1326] = layer4_out[3443];
    assign layer5_out[1327] = ~layer4_out[2696];
    assign layer5_out[1328] = layer4_out[1314] ^ layer4_out[1315];
    assign layer5_out[1329] = layer4_out[2515] & ~layer4_out[2516];
    assign layer5_out[1330] = ~(layer4_out[6002] ^ layer4_out[6003]);
    assign layer5_out[1331] = ~(layer4_out[147] ^ layer4_out[148]);
    assign layer5_out[1332] = ~layer4_out[1699];
    assign layer5_out[1333] = layer4_out[5829];
    assign layer5_out[1334] = layer4_out[5841];
    assign layer5_out[1335] = ~layer4_out[4058];
    assign layer5_out[1336] = ~layer4_out[4148];
    assign layer5_out[1337] = ~layer4_out[1705];
    assign layer5_out[1338] = layer4_out[7015] ^ layer4_out[7016];
    assign layer5_out[1339] = ~layer4_out[5017];
    assign layer5_out[1340] = layer4_out[6170];
    assign layer5_out[1341] = layer4_out[7448];
    assign layer5_out[1342] = ~layer4_out[6754];
    assign layer5_out[1343] = ~(layer4_out[6366] | layer4_out[6367]);
    assign layer5_out[1344] = layer4_out[5991];
    assign layer5_out[1345] = layer4_out[7290] & ~layer4_out[7289];
    assign layer5_out[1346] = layer4_out[1102];
    assign layer5_out[1347] = layer4_out[3082];
    assign layer5_out[1348] = ~layer4_out[2379];
    assign layer5_out[1349] = layer4_out[7482] & layer4_out[7483];
    assign layer5_out[1350] = ~(layer4_out[1503] | layer4_out[1504]);
    assign layer5_out[1351] = layer4_out[2149] ^ layer4_out[2150];
    assign layer5_out[1352] = ~layer4_out[1128];
    assign layer5_out[1353] = ~layer4_out[1280];
    assign layer5_out[1354] = layer4_out[2107];
    assign layer5_out[1355] = layer4_out[2507] & layer4_out[2508];
    assign layer5_out[1356] = layer4_out[3875] ^ layer4_out[3876];
    assign layer5_out[1357] = ~layer4_out[1610];
    assign layer5_out[1358] = layer4_out[7535] ^ layer4_out[7536];
    assign layer5_out[1359] = layer4_out[3595];
    assign layer5_out[1360] = ~layer4_out[805];
    assign layer5_out[1361] = layer4_out[5300];
    assign layer5_out[1362] = layer4_out[2821] ^ layer4_out[2822];
    assign layer5_out[1363] = layer4_out[7788] ^ layer4_out[7789];
    assign layer5_out[1364] = ~layer4_out[3113];
    assign layer5_out[1365] = layer4_out[1451] ^ layer4_out[1452];
    assign layer5_out[1366] = layer4_out[2873] ^ layer4_out[2874];
    assign layer5_out[1367] = layer4_out[7803] ^ layer4_out[7804];
    assign layer5_out[1368] = ~layer4_out[576];
    assign layer5_out[1369] = ~(layer4_out[5535] ^ layer4_out[5536]);
    assign layer5_out[1370] = layer4_out[6627];
    assign layer5_out[1371] = layer4_out[6864] & layer4_out[6865];
    assign layer5_out[1372] = layer4_out[584] ^ layer4_out[585];
    assign layer5_out[1373] = layer4_out[636];
    assign layer5_out[1374] = layer4_out[5989];
    assign layer5_out[1375] = layer4_out[4131] ^ layer4_out[4132];
    assign layer5_out[1376] = ~(layer4_out[7601] ^ layer4_out[7602]);
    assign layer5_out[1377] = layer4_out[4811] ^ layer4_out[4812];
    assign layer5_out[1378] = layer4_out[4816] & ~layer4_out[4817];
    assign layer5_out[1379] = layer4_out[7411] & ~layer4_out[7410];
    assign layer5_out[1380] = layer4_out[749] & ~layer4_out[748];
    assign layer5_out[1381] = layer4_out[137] & ~layer4_out[136];
    assign layer5_out[1382] = ~(layer4_out[6629] ^ layer4_out[6630]);
    assign layer5_out[1383] = layer4_out[3142];
    assign layer5_out[1384] = layer4_out[4540] & ~layer4_out[4541];
    assign layer5_out[1385] = ~layer4_out[1136];
    assign layer5_out[1386] = ~(layer4_out[4731] | layer4_out[4732]);
    assign layer5_out[1387] = layer4_out[4478];
    assign layer5_out[1388] = ~(layer4_out[7776] ^ layer4_out[7777]);
    assign layer5_out[1389] = layer4_out[2485] ^ layer4_out[2486];
    assign layer5_out[1390] = ~(layer4_out[4308] ^ layer4_out[4309]);
    assign layer5_out[1391] = ~layer4_out[1815] | layer4_out[1814];
    assign layer5_out[1392] = layer4_out[6761] & layer4_out[6762];
    assign layer5_out[1393] = layer4_out[4803] ^ layer4_out[4804];
    assign layer5_out[1394] = ~(layer4_out[1619] ^ layer4_out[1620]);
    assign layer5_out[1395] = ~layer4_out[6870];
    assign layer5_out[1396] = ~(layer4_out[569] ^ layer4_out[570]);
    assign layer5_out[1397] = layer4_out[2754] ^ layer4_out[2755];
    assign layer5_out[1398] = layer4_out[5332] & ~layer4_out[5333];
    assign layer5_out[1399] = layer4_out[372] & ~layer4_out[371];
    assign layer5_out[1400] = layer4_out[4421];
    assign layer5_out[1401] = ~(layer4_out[7628] ^ layer4_out[7629]);
    assign layer5_out[1402] = layer4_out[301] & ~layer4_out[302];
    assign layer5_out[1403] = layer4_out[5488] ^ layer4_out[5489];
    assign layer5_out[1404] = ~(layer4_out[1641] | layer4_out[1642]);
    assign layer5_out[1405] = layer4_out[6192];
    assign layer5_out[1406] = ~(layer4_out[5231] ^ layer4_out[5232]);
    assign layer5_out[1407] = ~(layer4_out[2083] | layer4_out[2084]);
    assign layer5_out[1408] = ~(layer4_out[3916] ^ layer4_out[3917]);
    assign layer5_out[1409] = layer4_out[6704];
    assign layer5_out[1410] = layer4_out[2256] & ~layer4_out[2255];
    assign layer5_out[1411] = ~layer4_out[6211];
    assign layer5_out[1412] = ~layer4_out[7701];
    assign layer5_out[1413] = layer4_out[2995] ^ layer4_out[2996];
    assign layer5_out[1414] = ~layer4_out[6529] | layer4_out[6528];
    assign layer5_out[1415] = layer4_out[7054];
    assign layer5_out[1416] = ~(layer4_out[3899] ^ layer4_out[3900]);
    assign layer5_out[1417] = ~(layer4_out[6213] ^ layer4_out[6214]);
    assign layer5_out[1418] = layer4_out[4417];
    assign layer5_out[1419] = ~(layer4_out[5417] | layer4_out[5418]);
    assign layer5_out[1420] = layer4_out[3058] ^ layer4_out[3059];
    assign layer5_out[1421] = layer4_out[6056];
    assign layer5_out[1422] = ~layer4_out[628] | layer4_out[627];
    assign layer5_out[1423] = layer4_out[6540] & layer4_out[6541];
    assign layer5_out[1424] = ~layer4_out[7989] | layer4_out[7988];
    assign layer5_out[1425] = layer4_out[505];
    assign layer5_out[1426] = ~(layer4_out[6117] ^ layer4_out[6118]);
    assign layer5_out[1427] = layer4_out[2419] & layer4_out[2420];
    assign layer5_out[1428] = ~(layer4_out[1152] | layer4_out[1153]);
    assign layer5_out[1429] = layer4_out[5500] ^ layer4_out[5501];
    assign layer5_out[1430] = ~(layer4_out[831] ^ layer4_out[832]);
    assign layer5_out[1431] = layer4_out[2780];
    assign layer5_out[1432] = ~(layer4_out[5701] ^ layer4_out[5702]);
    assign layer5_out[1433] = layer4_out[1352] ^ layer4_out[1353];
    assign layer5_out[1434] = ~layer4_out[2626];
    assign layer5_out[1435] = ~(layer4_out[789] ^ layer4_out[790]);
    assign layer5_out[1436] = ~layer4_out[3859] | layer4_out[3858];
    assign layer5_out[1437] = ~layer4_out[7642] | layer4_out[7641];
    assign layer5_out[1438] = layer4_out[201] ^ layer4_out[202];
    assign layer5_out[1439] = layer4_out[4151];
    assign layer5_out[1440] = layer4_out[3365] ^ layer4_out[3366];
    assign layer5_out[1441] = layer4_out[3210] ^ layer4_out[3211];
    assign layer5_out[1442] = ~layer4_out[326];
    assign layer5_out[1443] = layer4_out[2729] & layer4_out[2730];
    assign layer5_out[1444] = ~layer4_out[5428];
    assign layer5_out[1445] = ~(layer4_out[6936] | layer4_out[6937]);
    assign layer5_out[1446] = layer4_out[6081];
    assign layer5_out[1447] = layer4_out[7143];
    assign layer5_out[1448] = layer4_out[968] ^ layer4_out[969];
    assign layer5_out[1449] = ~layer4_out[3252];
    assign layer5_out[1450] = ~(layer4_out[457] ^ layer4_out[458]);
    assign layer5_out[1451] = ~layer4_out[4742] | layer4_out[4741];
    assign layer5_out[1452] = ~(layer4_out[4490] & layer4_out[4491]);
    assign layer5_out[1453] = layer4_out[665] ^ layer4_out[666];
    assign layer5_out[1454] = layer4_out[1035] & layer4_out[1036];
    assign layer5_out[1455] = ~(layer4_out[4120] ^ layer4_out[4121]);
    assign layer5_out[1456] = layer4_out[5777] & layer4_out[5778];
    assign layer5_out[1457] = ~layer4_out[7253] | layer4_out[7254];
    assign layer5_out[1458] = ~layer4_out[1350];
    assign layer5_out[1459] = ~layer4_out[7761];
    assign layer5_out[1460] = ~layer4_out[2685];
    assign layer5_out[1461] = ~(layer4_out[5498] ^ layer4_out[5499]);
    assign layer5_out[1462] = layer4_out[1617];
    assign layer5_out[1463] = layer4_out[6225] ^ layer4_out[6226];
    assign layer5_out[1464] = ~(layer4_out[4650] | layer4_out[4651]);
    assign layer5_out[1465] = layer4_out[4469];
    assign layer5_out[1466] = ~layer4_out[7211];
    assign layer5_out[1467] = layer4_out[2759] & layer4_out[2760];
    assign layer5_out[1468] = ~(layer4_out[3810] & layer4_out[3811]);
    assign layer5_out[1469] = ~(layer4_out[5241] ^ layer4_out[5242]);
    assign layer5_out[1470] = layer4_out[7092];
    assign layer5_out[1471] = layer4_out[1226] ^ layer4_out[1227];
    assign layer5_out[1472] = ~(layer4_out[5496] | layer4_out[5497]);
    assign layer5_out[1473] = layer4_out[3800] & ~layer4_out[3801];
    assign layer5_out[1474] = layer4_out[3724];
    assign layer5_out[1475] = ~(layer4_out[349] ^ layer4_out[350]);
    assign layer5_out[1476] = layer4_out[466] ^ layer4_out[467];
    assign layer5_out[1477] = ~(layer4_out[7049] ^ layer4_out[7050]);
    assign layer5_out[1478] = ~layer4_out[7556];
    assign layer5_out[1479] = layer4_out[4998];
    assign layer5_out[1480] = layer4_out[5179] & layer4_out[5180];
    assign layer5_out[1481] = ~(layer4_out[654] ^ layer4_out[655]);
    assign layer5_out[1482] = layer4_out[990];
    assign layer5_out[1483] = ~(layer4_out[7780] ^ layer4_out[7781]);
    assign layer5_out[1484] = ~(layer4_out[5186] ^ layer4_out[5187]);
    assign layer5_out[1485] = ~(layer4_out[2790] ^ layer4_out[2791]);
    assign layer5_out[1486] = ~(layer4_out[6676] ^ layer4_out[6677]);
    assign layer5_out[1487] = layer4_out[299];
    assign layer5_out[1488] = ~(layer4_out[5830] | layer4_out[5831]);
    assign layer5_out[1489] = layer4_out[929] & ~layer4_out[928];
    assign layer5_out[1490] = ~(layer4_out[1373] & layer4_out[1374]);
    assign layer5_out[1491] = layer4_out[6488] & ~layer4_out[6489];
    assign layer5_out[1492] = ~layer4_out[2680];
    assign layer5_out[1493] = layer4_out[2154];
    assign layer5_out[1494] = layer4_out[3675] ^ layer4_out[3676];
    assign layer5_out[1495] = ~layer4_out[7933];
    assign layer5_out[1496] = layer4_out[1074] & layer4_out[1075];
    assign layer5_out[1497] = layer4_out[3048] ^ layer4_out[3049];
    assign layer5_out[1498] = ~(layer4_out[1305] ^ layer4_out[1306]);
    assign layer5_out[1499] = layer4_out[4476] ^ layer4_out[4477];
    assign layer5_out[1500] = layer4_out[5339];
    assign layer5_out[1501] = layer4_out[2553];
    assign layer5_out[1502] = ~(layer4_out[3000] ^ layer4_out[3001]);
    assign layer5_out[1503] = ~layer4_out[1944];
    assign layer5_out[1504] = ~(layer4_out[354] ^ layer4_out[355]);
    assign layer5_out[1505] = ~layer4_out[5655];
    assign layer5_out[1506] = layer4_out[6578] & ~layer4_out[6579];
    assign layer5_out[1507] = ~layer4_out[3257];
    assign layer5_out[1508] = layer4_out[1283];
    assign layer5_out[1509] = layer4_out[7256] & layer4_out[7257];
    assign layer5_out[1510] = layer4_out[7595] & layer4_out[7596];
    assign layer5_out[1511] = layer4_out[2835] ^ layer4_out[2836];
    assign layer5_out[1512] = layer4_out[3044] & ~layer4_out[3043];
    assign layer5_out[1513] = ~(layer4_out[1180] ^ layer4_out[1181]);
    assign layer5_out[1514] = layer4_out[3132];
    assign layer5_out[1515] = layer4_out[876] & layer4_out[877];
    assign layer5_out[1516] = layer4_out[1831] & ~layer4_out[1830];
    assign layer5_out[1517] = layer4_out[4195];
    assign layer5_out[1518] = layer4_out[2407] & layer4_out[2408];
    assign layer5_out[1519] = layer4_out[3644] | layer4_out[3645];
    assign layer5_out[1520] = layer4_out[5490];
    assign layer5_out[1521] = ~layer4_out[1538];
    assign layer5_out[1522] = ~(layer4_out[4576] ^ layer4_out[4577]);
    assign layer5_out[1523] = ~layer4_out[3554];
    assign layer5_out[1524] = ~layer4_out[3547] | layer4_out[3548];
    assign layer5_out[1525] = layer4_out[7908] & ~layer4_out[7909];
    assign layer5_out[1526] = layer4_out[7252] ^ layer4_out[7253];
    assign layer5_out[1527] = ~(layer4_out[6323] | layer4_out[6324]);
    assign layer5_out[1528] = ~(layer4_out[3065] | layer4_out[3066]);
    assign layer5_out[1529] = layer4_out[763] | layer4_out[764];
    assign layer5_out[1530] = layer4_out[4652] ^ layer4_out[4653];
    assign layer5_out[1531] = layer4_out[3787];
    assign layer5_out[1532] = layer4_out[1936] & layer4_out[1937];
    assign layer5_out[1533] = layer4_out[6006] & ~layer4_out[6007];
    assign layer5_out[1534] = 1'b0;
    assign layer5_out[1535] = layer4_out[5934] & ~layer4_out[5935];
    assign layer5_out[1536] = layer4_out[5094] ^ layer4_out[5095];
    assign layer5_out[1537] = layer4_out[5783];
    assign layer5_out[1538] = ~layer4_out[3271];
    assign layer5_out[1539] = ~(layer4_out[6736] ^ layer4_out[6737]);
    assign layer5_out[1540] = ~layer4_out[4923];
    assign layer5_out[1541] = layer4_out[1839] & layer4_out[1840];
    assign layer5_out[1542] = ~(layer4_out[669] & layer4_out[670]);
    assign layer5_out[1543] = ~layer4_out[3416] | layer4_out[3415];
    assign layer5_out[1544] = layer4_out[5586];
    assign layer5_out[1545] = ~(layer4_out[7406] | layer4_out[7407]);
    assign layer5_out[1546] = layer4_out[1644];
    assign layer5_out[1547] = layer4_out[2198] ^ layer4_out[2199];
    assign layer5_out[1548] = layer4_out[2659];
    assign layer5_out[1549] = ~(layer4_out[1458] ^ layer4_out[1459]);
    assign layer5_out[1550] = layer4_out[3421] ^ layer4_out[3422];
    assign layer5_out[1551] = ~(layer4_out[574] ^ layer4_out[575]);
    assign layer5_out[1552] = layer4_out[171] ^ layer4_out[172];
    assign layer5_out[1553] = ~(layer4_out[246] ^ layer4_out[247]);
    assign layer5_out[1554] = layer4_out[7700] ^ layer4_out[7701];
    assign layer5_out[1555] = ~layer4_out[5700];
    assign layer5_out[1556] = layer4_out[2936] & layer4_out[2937];
    assign layer5_out[1557] = ~(layer4_out[200] ^ layer4_out[201]);
    assign layer5_out[1558] = ~layer4_out[7273];
    assign layer5_out[1559] = layer4_out[1800];
    assign layer5_out[1560] = layer4_out[7333] ^ layer4_out[7334];
    assign layer5_out[1561] = ~(layer4_out[6353] | layer4_out[6354]);
    assign layer5_out[1562] = layer4_out[1982] & layer4_out[1983];
    assign layer5_out[1563] = ~layer4_out[1291];
    assign layer5_out[1564] = layer4_out[3154] & ~layer4_out[3155];
    assign layer5_out[1565] = layer4_out[1217];
    assign layer5_out[1566] = layer4_out[2964] ^ layer4_out[2965];
    assign layer5_out[1567] = layer4_out[2154];
    assign layer5_out[1568] = layer4_out[6471];
    assign layer5_out[1569] = layer4_out[1096];
    assign layer5_out[1570] = layer4_out[5350] & ~layer4_out[5351];
    assign layer5_out[1571] = layer4_out[3082];
    assign layer5_out[1572] = ~(layer4_out[7372] & layer4_out[7373]);
    assign layer5_out[1573] = ~(layer4_out[1967] ^ layer4_out[1968]);
    assign layer5_out[1574] = ~(layer4_out[2471] ^ layer4_out[2472]);
    assign layer5_out[1575] = ~layer4_out[1154];
    assign layer5_out[1576] = layer4_out[7838] & layer4_out[7839];
    assign layer5_out[1577] = ~(layer4_out[3952] ^ layer4_out[3953]);
    assign layer5_out[1578] = ~layer4_out[7080];
    assign layer5_out[1579] = layer4_out[6583];
    assign layer5_out[1580] = ~(layer4_out[4621] ^ layer4_out[4622]);
    assign layer5_out[1581] = layer4_out[2564] ^ layer4_out[2565];
    assign layer5_out[1582] = layer4_out[555] ^ layer4_out[556];
    assign layer5_out[1583] = layer4_out[1763] & ~layer4_out[1762];
    assign layer5_out[1584] = ~(layer4_out[4569] ^ layer4_out[4570]);
    assign layer5_out[1585] = ~layer4_out[3493] | layer4_out[3492];
    assign layer5_out[1586] = ~layer4_out[7131] | layer4_out[7132];
    assign layer5_out[1587] = ~layer4_out[400];
    assign layer5_out[1588] = layer4_out[3767] & ~layer4_out[3768];
    assign layer5_out[1589] = layer4_out[623];
    assign layer5_out[1590] = layer4_out[4866] ^ layer4_out[4867];
    assign layer5_out[1591] = layer4_out[5605] ^ layer4_out[5606];
    assign layer5_out[1592] = layer4_out[120];
    assign layer5_out[1593] = ~(layer4_out[4585] & layer4_out[4586]);
    assign layer5_out[1594] = layer4_out[3823] & ~layer4_out[3822];
    assign layer5_out[1595] = ~layer4_out[1598];
    assign layer5_out[1596] = layer4_out[2728] & layer4_out[2729];
    assign layer5_out[1597] = layer4_out[6368] ^ layer4_out[6369];
    assign layer5_out[1598] = ~layer4_out[3886] | layer4_out[3885];
    assign layer5_out[1599] = layer4_out[833] ^ layer4_out[834];
    assign layer5_out[1600] = layer4_out[7290] ^ layer4_out[7291];
    assign layer5_out[1601] = ~layer4_out[3161];
    assign layer5_out[1602] = ~(layer4_out[878] & layer4_out[879]);
    assign layer5_out[1603] = ~(layer4_out[2721] | layer4_out[2722]);
    assign layer5_out[1604] = layer4_out[2506] & layer4_out[2507];
    assign layer5_out[1605] = ~layer4_out[3191];
    assign layer5_out[1606] = ~(layer4_out[3623] & layer4_out[3624]);
    assign layer5_out[1607] = ~layer4_out[6867];
    assign layer5_out[1608] = ~layer4_out[2971];
    assign layer5_out[1609] = layer4_out[2943] & layer4_out[2944];
    assign layer5_out[1610] = layer4_out[3550] & layer4_out[3551];
    assign layer5_out[1611] = ~layer4_out[2319];
    assign layer5_out[1612] = ~(layer4_out[790] | layer4_out[791]);
    assign layer5_out[1613] = layer4_out[3289];
    assign layer5_out[1614] = layer4_out[5882] & layer4_out[5883];
    assign layer5_out[1615] = ~layer4_out[2867] | layer4_out[2868];
    assign layer5_out[1616] = ~layer4_out[7511];
    assign layer5_out[1617] = ~layer4_out[5028];
    assign layer5_out[1618] = layer4_out[5739];
    assign layer5_out[1619] = layer4_out[7040];
    assign layer5_out[1620] = layer4_out[3891];
    assign layer5_out[1621] = ~layer4_out[3555];
    assign layer5_out[1622] = layer4_out[4844] ^ layer4_out[4845];
    assign layer5_out[1623] = layer4_out[4563] ^ layer4_out[4564];
    assign layer5_out[1624] = layer4_out[5229] & layer4_out[5230];
    assign layer5_out[1625] = layer4_out[2306] ^ layer4_out[2307];
    assign layer5_out[1626] = layer4_out[7028] & ~layer4_out[7027];
    assign layer5_out[1627] = layer4_out[4832] & ~layer4_out[4833];
    assign layer5_out[1628] = layer4_out[3864] ^ layer4_out[3865];
    assign layer5_out[1629] = layer4_out[2274] & ~layer4_out[2275];
    assign layer5_out[1630] = layer4_out[3323];
    assign layer5_out[1631] = layer4_out[7409];
    assign layer5_out[1632] = layer4_out[3964] & layer4_out[3965];
    assign layer5_out[1633] = layer4_out[3153] | layer4_out[3154];
    assign layer5_out[1634] = layer4_out[5616];
    assign layer5_out[1635] = layer4_out[5950] ^ layer4_out[5951];
    assign layer5_out[1636] = ~layer4_out[6006];
    assign layer5_out[1637] = ~layer4_out[4634];
    assign layer5_out[1638] = layer4_out[4740] | layer4_out[4741];
    assign layer5_out[1639] = layer4_out[5065];
    assign layer5_out[1640] = layer4_out[3591] & ~layer4_out[3592];
    assign layer5_out[1641] = layer4_out[2599] & layer4_out[2600];
    assign layer5_out[1642] = layer4_out[4952];
    assign layer5_out[1643] = layer4_out[6260] & ~layer4_out[6259];
    assign layer5_out[1644] = layer4_out[7293] ^ layer4_out[7294];
    assign layer5_out[1645] = ~layer4_out[3951];
    assign layer5_out[1646] = ~layer4_out[985];
    assign layer5_out[1647] = layer4_out[7494];
    assign layer5_out[1648] = layer4_out[2199] & layer4_out[2200];
    assign layer5_out[1649] = ~(layer4_out[7361] ^ layer4_out[7362]);
    assign layer5_out[1650] = ~layer4_out[110];
    assign layer5_out[1651] = ~layer4_out[5653];
    assign layer5_out[1652] = layer4_out[4771] & ~layer4_out[4772];
    assign layer5_out[1653] = layer4_out[1079];
    assign layer5_out[1654] = layer4_out[3111];
    assign layer5_out[1655] = ~layer4_out[2652];
    assign layer5_out[1656] = ~layer4_out[2331];
    assign layer5_out[1657] = layer4_out[4135] & ~layer4_out[4136];
    assign layer5_out[1658] = ~(layer4_out[7639] ^ layer4_out[7640]);
    assign layer5_out[1659] = layer4_out[7777] | layer4_out[7778];
    assign layer5_out[1660] = ~(layer4_out[6003] ^ layer4_out[6004]);
    assign layer5_out[1661] = ~(layer4_out[1063] & layer4_out[1064]);
    assign layer5_out[1662] = layer4_out[3219] | layer4_out[3220];
    assign layer5_out[1663] = layer4_out[2271] & ~layer4_out[2270];
    assign layer5_out[1664] = layer4_out[739] | layer4_out[740];
    assign layer5_out[1665] = ~layer4_out[1934] | layer4_out[1933];
    assign layer5_out[1666] = ~(layer4_out[378] | layer4_out[379]);
    assign layer5_out[1667] = ~(layer4_out[741] ^ layer4_out[742]);
    assign layer5_out[1668] = layer4_out[5553] & ~layer4_out[5552];
    assign layer5_out[1669] = ~(layer4_out[679] ^ layer4_out[680]);
    assign layer5_out[1670] = layer4_out[1359];
    assign layer5_out[1671] = layer4_out[393] & ~layer4_out[392];
    assign layer5_out[1672] = layer4_out[6451] | layer4_out[6452];
    assign layer5_out[1673] = layer4_out[1471] ^ layer4_out[1472];
    assign layer5_out[1674] = layer4_out[1271];
    assign layer5_out[1675] = ~(layer4_out[4889] ^ layer4_out[4890]);
    assign layer5_out[1676] = layer4_out[7827];
    assign layer5_out[1677] = ~layer4_out[7429] | layer4_out[7430];
    assign layer5_out[1678] = ~(layer4_out[294] ^ layer4_out[295]);
    assign layer5_out[1679] = ~layer4_out[4306] | layer4_out[4305];
    assign layer5_out[1680] = layer4_out[7642] ^ layer4_out[7643];
    assign layer5_out[1681] = ~layer4_out[4533] | layer4_out[4534];
    assign layer5_out[1682] = layer4_out[5520] & layer4_out[5521];
    assign layer5_out[1683] = ~(layer4_out[5626] & layer4_out[5627]);
    assign layer5_out[1684] = ~layer4_out[3448] | layer4_out[3449];
    assign layer5_out[1685] = ~(layer4_out[5793] ^ layer4_out[5794]);
    assign layer5_out[1686] = layer4_out[723];
    assign layer5_out[1687] = ~layer4_out[5291];
    assign layer5_out[1688] = ~layer4_out[6473] | layer4_out[6474];
    assign layer5_out[1689] = layer4_out[3787] & layer4_out[3788];
    assign layer5_out[1690] = ~layer4_out[6223];
    assign layer5_out[1691] = layer4_out[2490];
    assign layer5_out[1692] = ~layer4_out[558];
    assign layer5_out[1693] = ~(layer4_out[4275] ^ layer4_out[4276]);
    assign layer5_out[1694] = ~layer4_out[5670];
    assign layer5_out[1695] = layer4_out[1935] ^ layer4_out[1936];
    assign layer5_out[1696] = layer4_out[260] | layer4_out[261];
    assign layer5_out[1697] = ~layer4_out[6400];
    assign layer5_out[1698] = layer4_out[2466] ^ layer4_out[2467];
    assign layer5_out[1699] = layer4_out[3564];
    assign layer5_out[1700] = ~layer4_out[2454] | layer4_out[2455];
    assign layer5_out[1701] = layer4_out[7599] ^ layer4_out[7600];
    assign layer5_out[1702] = ~(layer4_out[3698] ^ layer4_out[3699]);
    assign layer5_out[1703] = ~layer4_out[7915];
    assign layer5_out[1704] = ~layer4_out[6386] | layer4_out[6385];
    assign layer5_out[1705] = ~(layer4_out[3479] ^ layer4_out[3480]);
    assign layer5_out[1706] = layer4_out[1509] & ~layer4_out[1510];
    assign layer5_out[1707] = ~layer4_out[4972];
    assign layer5_out[1708] = ~layer4_out[4489];
    assign layer5_out[1709] = ~layer4_out[1580];
    assign layer5_out[1710] = ~layer4_out[413];
    assign layer5_out[1711] = ~(layer4_out[4355] ^ layer4_out[4356]);
    assign layer5_out[1712] = ~(layer4_out[4260] ^ layer4_out[4261]);
    assign layer5_out[1713] = layer4_out[2323] & ~layer4_out[2322];
    assign layer5_out[1714] = ~layer4_out[412];
    assign layer5_out[1715] = layer4_out[3726];
    assign layer5_out[1716] = layer4_out[7134] & ~layer4_out[7135];
    assign layer5_out[1717] = ~(layer4_out[3363] | layer4_out[3364]);
    assign layer5_out[1718] = layer4_out[7988];
    assign layer5_out[1719] = ~layer4_out[7715];
    assign layer5_out[1720] = ~(layer4_out[6263] ^ layer4_out[6264]);
    assign layer5_out[1721] = ~layer4_out[4274] | layer4_out[4275];
    assign layer5_out[1722] = layer4_out[6661];
    assign layer5_out[1723] = ~layer4_out[4991] | layer4_out[4992];
    assign layer5_out[1724] = ~layer4_out[3694];
    assign layer5_out[1725] = ~layer4_out[2335];
    assign layer5_out[1726] = ~(layer4_out[3062] & layer4_out[3063]);
    assign layer5_out[1727] = ~(layer4_out[5788] | layer4_out[5789]);
    assign layer5_out[1728] = ~layer4_out[6080];
    assign layer5_out[1729] = layer4_out[7719] & ~layer4_out[7720];
    assign layer5_out[1730] = ~layer4_out[1978] | layer4_out[1979];
    assign layer5_out[1731] = ~layer4_out[4024] | layer4_out[4023];
    assign layer5_out[1732] = ~layer4_out[3429];
    assign layer5_out[1733] = ~layer4_out[3636] | layer4_out[3635];
    assign layer5_out[1734] = ~layer4_out[6404] | layer4_out[6405];
    assign layer5_out[1735] = ~(layer4_out[4196] ^ layer4_out[4197]);
    assign layer5_out[1736] = layer4_out[4969];
    assign layer5_out[1737] = ~(layer4_out[1474] | layer4_out[1475]);
    assign layer5_out[1738] = layer4_out[610] & ~layer4_out[611];
    assign layer5_out[1739] = ~layer4_out[487];
    assign layer5_out[1740] = ~(layer4_out[4033] | layer4_out[4034]);
    assign layer5_out[1741] = ~layer4_out[424];
    assign layer5_out[1742] = ~layer4_out[1744] | layer4_out[1743];
    assign layer5_out[1743] = layer4_out[6601] & ~layer4_out[6602];
    assign layer5_out[1744] = layer4_out[4063];
    assign layer5_out[1745] = layer4_out[3845];
    assign layer5_out[1746] = ~layer4_out[396];
    assign layer5_out[1747] = layer4_out[5219] ^ layer4_out[5220];
    assign layer5_out[1748] = layer4_out[2603];
    assign layer5_out[1749] = layer4_out[1261];
    assign layer5_out[1750] = layer4_out[4334];
    assign layer5_out[1751] = ~(layer4_out[5126] & layer4_out[5127]);
    assign layer5_out[1752] = layer4_out[6172];
    assign layer5_out[1753] = layer4_out[7126] ^ layer4_out[7127];
    assign layer5_out[1754] = ~layer4_out[3765];
    assign layer5_out[1755] = ~(layer4_out[5123] | layer4_out[5124]);
    assign layer5_out[1756] = ~(layer4_out[6943] ^ layer4_out[6944]);
    assign layer5_out[1757] = ~layer4_out[6780];
    assign layer5_out[1758] = layer4_out[2139];
    assign layer5_out[1759] = layer4_out[2450] & ~layer4_out[2451];
    assign layer5_out[1760] = layer4_out[4870] & ~layer4_out[4871];
    assign layer5_out[1761] = layer4_out[1703];
    assign layer5_out[1762] = layer4_out[4942];
    assign layer5_out[1763] = ~layer4_out[6998] | layer4_out[6999];
    assign layer5_out[1764] = ~layer4_out[434];
    assign layer5_out[1765] = layer4_out[7680] ^ layer4_out[7681];
    assign layer5_out[1766] = ~layer4_out[3470];
    assign layer5_out[1767] = layer4_out[5565] & ~layer4_out[5566];
    assign layer5_out[1768] = ~layer4_out[1955] | layer4_out[1954];
    assign layer5_out[1769] = layer4_out[5674];
    assign layer5_out[1770] = layer4_out[2026] & layer4_out[2027];
    assign layer5_out[1771] = ~layer4_out[2661];
    assign layer5_out[1772] = layer4_out[1827] ^ layer4_out[1828];
    assign layer5_out[1773] = layer4_out[3984];
    assign layer5_out[1774] = ~layer4_out[3975];
    assign layer5_out[1775] = layer4_out[4953] ^ layer4_out[4954];
    assign layer5_out[1776] = ~layer4_out[2534] | layer4_out[2533];
    assign layer5_out[1777] = layer4_out[1866];
    assign layer5_out[1778] = layer4_out[3459];
    assign layer5_out[1779] = layer4_out[4268] ^ layer4_out[4269];
    assign layer5_out[1780] = layer4_out[2456] ^ layer4_out[2457];
    assign layer5_out[1781] = layer4_out[4353];
    assign layer5_out[1782] = layer4_out[6423] & layer4_out[6424];
    assign layer5_out[1783] = layer4_out[3589] | layer4_out[3590];
    assign layer5_out[1784] = ~layer4_out[4950] | layer4_out[4951];
    assign layer5_out[1785] = ~layer4_out[7278];
    assign layer5_out[1786] = ~(layer4_out[4142] ^ layer4_out[4143]);
    assign layer5_out[1787] = ~(layer4_out[1450] ^ layer4_out[1451]);
    assign layer5_out[1788] = layer4_out[75];
    assign layer5_out[1789] = ~layer4_out[7841];
    assign layer5_out[1790] = ~layer4_out[3822];
    assign layer5_out[1791] = layer4_out[1080];
    assign layer5_out[1792] = ~(layer4_out[3832] ^ layer4_out[3833]);
    assign layer5_out[1793] = ~layer4_out[5314];
    assign layer5_out[1794] = layer4_out[7568] & ~layer4_out[7567];
    assign layer5_out[1795] = layer4_out[360];
    assign layer5_out[1796] = layer4_out[4284];
    assign layer5_out[1797] = ~(layer4_out[4519] | layer4_out[4520]);
    assign layer5_out[1798] = ~(layer4_out[7637] | layer4_out[7638]);
    assign layer5_out[1799] = layer4_out[1568];
    assign layer5_out[1800] = layer4_out[2839] ^ layer4_out[2840];
    assign layer5_out[1801] = layer4_out[5564];
    assign layer5_out[1802] = ~layer4_out[3138];
    assign layer5_out[1803] = layer4_out[7164];
    assign layer5_out[1804] = ~(layer4_out[6549] | layer4_out[6550]);
    assign layer5_out[1805] = ~layer4_out[5478];
    assign layer5_out[1806] = layer4_out[889] & layer4_out[890];
    assign layer5_out[1807] = ~layer4_out[7092];
    assign layer5_out[1808] = ~(layer4_out[1975] ^ layer4_out[1976]);
    assign layer5_out[1809] = layer4_out[3212];
    assign layer5_out[1810] = ~(layer4_out[7720] | layer4_out[7721]);
    assign layer5_out[1811] = layer4_out[2697] & ~layer4_out[2698];
    assign layer5_out[1812] = ~layer4_out[5984];
    assign layer5_out[1813] = ~(layer4_out[2477] ^ layer4_out[2478]);
    assign layer5_out[1814] = ~layer4_out[4617];
    assign layer5_out[1815] = ~(layer4_out[4424] ^ layer4_out[4425]);
    assign layer5_out[1816] = layer4_out[2992] & ~layer4_out[2993];
    assign layer5_out[1817] = layer4_out[7502] & ~layer4_out[7501];
    assign layer5_out[1818] = layer4_out[3561] & ~layer4_out[3560];
    assign layer5_out[1819] = layer4_out[1553] | layer4_out[1554];
    assign layer5_out[1820] = layer4_out[1587];
    assign layer5_out[1821] = ~layer4_out[6016];
    assign layer5_out[1822] = layer4_out[5340] & layer4_out[5341];
    assign layer5_out[1823] = layer4_out[5518];
    assign layer5_out[1824] = layer4_out[2096] ^ layer4_out[2097];
    assign layer5_out[1825] = layer4_out[2889] ^ layer4_out[2890];
    assign layer5_out[1826] = layer4_out[3101] | layer4_out[3102];
    assign layer5_out[1827] = ~layer4_out[1694];
    assign layer5_out[1828] = layer4_out[4062] | layer4_out[4063];
    assign layer5_out[1829] = layer4_out[1718];
    assign layer5_out[1830] = layer4_out[4383];
    assign layer5_out[1831] = ~(layer4_out[1791] ^ layer4_out[1792]);
    assign layer5_out[1832] = ~layer4_out[3544];
    assign layer5_out[1833] = layer4_out[6728] ^ layer4_out[6729];
    assign layer5_out[1834] = ~(layer4_out[3035] ^ layer4_out[3036]);
    assign layer5_out[1835] = ~(layer4_out[2321] ^ layer4_out[2322]);
    assign layer5_out[1836] = layer4_out[7662] ^ layer4_out[7663];
    assign layer5_out[1837] = layer4_out[913] ^ layer4_out[914];
    assign layer5_out[1838] = ~(layer4_out[6655] ^ layer4_out[6656]);
    assign layer5_out[1839] = layer4_out[358];
    assign layer5_out[1840] = layer4_out[5245];
    assign layer5_out[1841] = layer4_out[5781] ^ layer4_out[5782];
    assign layer5_out[1842] = ~(layer4_out[3315] | layer4_out[3316]);
    assign layer5_out[1843] = ~(layer4_out[7592] ^ layer4_out[7593]);
    assign layer5_out[1844] = ~(layer4_out[6462] ^ layer4_out[6463]);
    assign layer5_out[1845] = ~(layer4_out[5847] | layer4_out[5848]);
    assign layer5_out[1846] = layer4_out[3739] ^ layer4_out[3740];
    assign layer5_out[1847] = layer4_out[5667] & ~layer4_out[5668];
    assign layer5_out[1848] = ~layer4_out[5411];
    assign layer5_out[1849] = layer4_out[1353] ^ layer4_out[1354];
    assign layer5_out[1850] = ~layer4_out[6941];
    assign layer5_out[1851] = layer4_out[5475] | layer4_out[5476];
    assign layer5_out[1852] = ~(layer4_out[7152] | layer4_out[7153]);
    assign layer5_out[1853] = ~layer4_out[7994];
    assign layer5_out[1854] = layer4_out[5386] & ~layer4_out[5385];
    assign layer5_out[1855] = layer4_out[6800];
    assign layer5_out[1856] = layer4_out[7507] | layer4_out[7508];
    assign layer5_out[1857] = ~(layer4_out[5215] & layer4_out[5216]);
    assign layer5_out[1858] = layer4_out[2795];
    assign layer5_out[1859] = ~(layer4_out[3705] ^ layer4_out[3706]);
    assign layer5_out[1860] = layer4_out[2268] & ~layer4_out[2269];
    assign layer5_out[1861] = layer4_out[1540] & ~layer4_out[1541];
    assign layer5_out[1862] = layer4_out[6331] & layer4_out[6332];
    assign layer5_out[1863] = layer4_out[1171] | layer4_out[1172];
    assign layer5_out[1864] = ~layer4_out[7795];
    assign layer5_out[1865] = ~(layer4_out[1883] ^ layer4_out[1884]);
    assign layer5_out[1866] = ~layer4_out[4276];
    assign layer5_out[1867] = layer4_out[5636] ^ layer4_out[5637];
    assign layer5_out[1868] = ~layer4_out[1087];
    assign layer5_out[1869] = ~layer4_out[7346] | layer4_out[7345];
    assign layer5_out[1870] = ~layer4_out[6457];
    assign layer5_out[1871] = layer4_out[7243] & ~layer4_out[7244];
    assign layer5_out[1872] = ~(layer4_out[4565] | layer4_out[4566]);
    assign layer5_out[1873] = layer4_out[5042];
    assign layer5_out[1874] = layer4_out[2275] ^ layer4_out[2276];
    assign layer5_out[1875] = layer4_out[7284] & layer4_out[7285];
    assign layer5_out[1876] = ~layer4_out[2366];
    assign layer5_out[1877] = ~(layer4_out[6890] ^ layer4_out[6891]);
    assign layer5_out[1878] = ~layer4_out[694] | layer4_out[693];
    assign layer5_out[1879] = ~(layer4_out[3510] ^ layer4_out[3511]);
    assign layer5_out[1880] = ~(layer4_out[938] ^ layer4_out[939]);
    assign layer5_out[1881] = ~(layer4_out[895] ^ layer4_out[896]);
    assign layer5_out[1882] = ~layer4_out[1663];
    assign layer5_out[1883] = ~(layer4_out[4041] ^ layer4_out[4042]);
    assign layer5_out[1884] = ~layer4_out[6442];
    assign layer5_out[1885] = ~(layer4_out[7330] ^ layer4_out[7331]);
    assign layer5_out[1886] = layer4_out[7618] & layer4_out[7619];
    assign layer5_out[1887] = ~(layer4_out[5069] | layer4_out[5070]);
    assign layer5_out[1888] = layer4_out[547];
    assign layer5_out[1889] = layer4_out[6786];
    assign layer5_out[1890] = ~(layer4_out[7259] ^ layer4_out[7260]);
    assign layer5_out[1891] = ~(layer4_out[3261] & layer4_out[3262]);
    assign layer5_out[1892] = ~layer4_out[1176];
    assign layer5_out[1893] = ~layer4_out[3037];
    assign layer5_out[1894] = ~layer4_out[2298];
    assign layer5_out[1895] = layer4_out[1115] & ~layer4_out[1116];
    assign layer5_out[1896] = layer4_out[5222];
    assign layer5_out[1897] = ~(layer4_out[5884] ^ layer4_out[5885]);
    assign layer5_out[1898] = ~layer4_out[5848];
    assign layer5_out[1899] = layer4_out[967];
    assign layer5_out[1900] = ~layer4_out[6291] | layer4_out[6292];
    assign layer5_out[1901] = layer4_out[1379];
    assign layer5_out[1902] = layer4_out[3483] & layer4_out[3484];
    assign layer5_out[1903] = ~layer4_out[1852] | layer4_out[1853];
    assign layer5_out[1904] = layer4_out[4151];
    assign layer5_out[1905] = ~layer4_out[6299];
    assign layer5_out[1906] = ~(layer4_out[4379] & layer4_out[4380]);
    assign layer5_out[1907] = layer4_out[5981];
    assign layer5_out[1908] = layer4_out[3369] | layer4_out[3370];
    assign layer5_out[1909] = ~layer4_out[6947] | layer4_out[6948];
    assign layer5_out[1910] = layer4_out[7618] & ~layer4_out[7617];
    assign layer5_out[1911] = ~(layer4_out[4778] ^ layer4_out[4779]);
    assign layer5_out[1912] = layer4_out[4877] & layer4_out[4878];
    assign layer5_out[1913] = layer4_out[3754];
    assign layer5_out[1914] = ~layer4_out[3978];
    assign layer5_out[1915] = ~(layer4_out[251] ^ layer4_out[252]);
    assign layer5_out[1916] = ~(layer4_out[268] | layer4_out[269]);
    assign layer5_out[1917] = ~layer4_out[5586];
    assign layer5_out[1918] = ~(layer4_out[2095] ^ layer4_out[2096]);
    assign layer5_out[1919] = layer4_out[1150];
    assign layer5_out[1920] = ~layer4_out[7652];
    assign layer5_out[1921] = ~(layer4_out[1285] ^ layer4_out[1286]);
    assign layer5_out[1922] = layer4_out[5505];
    assign layer5_out[1923] = layer4_out[778];
    assign layer5_out[1924] = ~layer4_out[3526] | layer4_out[3525];
    assign layer5_out[1925] = layer4_out[1957] & ~layer4_out[1958];
    assign layer5_out[1926] = layer4_out[3179];
    assign layer5_out[1927] = layer4_out[6480];
    assign layer5_out[1928] = layer4_out[7485] & layer4_out[7486];
    assign layer5_out[1929] = ~layer4_out[7811];
    assign layer5_out[1930] = layer4_out[2113] | layer4_out[2114];
    assign layer5_out[1931] = layer4_out[4482] & ~layer4_out[4483];
    assign layer5_out[1932] = layer4_out[6600];
    assign layer5_out[1933] = ~layer4_out[3159];
    assign layer5_out[1934] = layer4_out[7489] | layer4_out[7490];
    assign layer5_out[1935] = layer4_out[2337] & layer4_out[2338];
    assign layer5_out[1936] = layer4_out[3601] & ~layer4_out[3600];
    assign layer5_out[1937] = layer4_out[5745] ^ layer4_out[5746];
    assign layer5_out[1938] = ~(layer4_out[453] ^ layer4_out[454]);
    assign layer5_out[1939] = layer4_out[4283];
    assign layer5_out[1940] = layer4_out[2912] | layer4_out[2913];
    assign layer5_out[1941] = layer4_out[2610] ^ layer4_out[2611];
    assign layer5_out[1942] = layer4_out[5878];
    assign layer5_out[1943] = ~(layer4_out[7585] ^ layer4_out[7586]);
    assign layer5_out[1944] = layer4_out[7827];
    assign layer5_out[1945] = layer4_out[7775];
    assign layer5_out[1946] = ~layer4_out[7584];
    assign layer5_out[1947] = layer4_out[5017];
    assign layer5_out[1948] = layer4_out[1949];
    assign layer5_out[1949] = layer4_out[5463] | layer4_out[5464];
    assign layer5_out[1950] = ~layer4_out[5556] | layer4_out[5557];
    assign layer5_out[1951] = layer4_out[5151] ^ layer4_out[5152];
    assign layer5_out[1952] = layer4_out[54] | layer4_out[55];
    assign layer5_out[1953] = ~(layer4_out[2706] ^ layer4_out[2707]);
    assign layer5_out[1954] = layer4_out[7572] & ~layer4_out[7573];
    assign layer5_out[1955] = layer4_out[5002];
    assign layer5_out[1956] = ~(layer4_out[7352] & layer4_out[7353]);
    assign layer5_out[1957] = ~layer4_out[2035] | layer4_out[2034];
    assign layer5_out[1958] = ~(layer4_out[7105] & layer4_out[7106]);
    assign layer5_out[1959] = layer4_out[3602];
    assign layer5_out[1960] = ~(layer4_out[4871] ^ layer4_out[4872]);
    assign layer5_out[1961] = layer4_out[5352];
    assign layer5_out[1962] = layer4_out[882] & ~layer4_out[881];
    assign layer5_out[1963] = layer4_out[6659] & ~layer4_out[6658];
    assign layer5_out[1964] = layer4_out[2766];
    assign layer5_out[1965] = layer4_out[639] ^ layer4_out[640];
    assign layer5_out[1966] = layer4_out[1295];
    assign layer5_out[1967] = ~layer4_out[5120];
    assign layer5_out[1968] = ~layer4_out[1533];
    assign layer5_out[1969] = layer4_out[740] & ~layer4_out[741];
    assign layer5_out[1970] = ~(layer4_out[1191] & layer4_out[1192]);
    assign layer5_out[1971] = layer4_out[7890];
    assign layer5_out[1972] = layer4_out[815];
    assign layer5_out[1973] = ~(layer4_out[4667] | layer4_out[4668]);
    assign layer5_out[1974] = layer4_out[6698] & layer4_out[6699];
    assign layer5_out[1975] = ~layer4_out[4401];
    assign layer5_out[1976] = layer4_out[4811];
    assign layer5_out[1977] = layer4_out[6107];
    assign layer5_out[1978] = ~layer4_out[814];
    assign layer5_out[1979] = layer4_out[2580];
    assign layer5_out[1980] = ~layer4_out[3009];
    assign layer5_out[1981] = ~layer4_out[247];
    assign layer5_out[1982] = ~layer4_out[5144];
    assign layer5_out[1983] = ~layer4_out[5987] | layer4_out[5986];
    assign layer5_out[1984] = ~layer4_out[4242];
    assign layer5_out[1985] = ~(layer4_out[3966] ^ layer4_out[3967]);
    assign layer5_out[1986] = layer4_out[4407] & ~layer4_out[4408];
    assign layer5_out[1987] = layer4_out[1973] ^ layer4_out[1974];
    assign layer5_out[1988] = ~layer4_out[281];
    assign layer5_out[1989] = layer4_out[7098] & layer4_out[7099];
    assign layer5_out[1990] = layer4_out[6643] | layer4_out[6644];
    assign layer5_out[1991] = ~(layer4_out[2444] | layer4_out[2445]);
    assign layer5_out[1992] = ~(layer4_out[7783] ^ layer4_out[7784]);
    assign layer5_out[1993] = ~layer4_out[7580];
    assign layer5_out[1994] = layer4_out[6636] & ~layer4_out[6637];
    assign layer5_out[1995] = ~layer4_out[5326];
    assign layer5_out[1996] = ~(layer4_out[5338] ^ layer4_out[5339]);
    assign layer5_out[1997] = ~layer4_out[3166];
    assign layer5_out[1998] = ~layer4_out[103] | layer4_out[102];
    assign layer5_out[1999] = ~(layer4_out[5905] ^ layer4_out[5906]);
    assign layer5_out[2000] = layer4_out[1335] ^ layer4_out[1336];
    assign layer5_out[2001] = ~(layer4_out[4644] | layer4_out[4645]);
    assign layer5_out[2002] = layer4_out[4993] & ~layer4_out[4994];
    assign layer5_out[2003] = ~(layer4_out[3338] ^ layer4_out[3339]);
    assign layer5_out[2004] = ~(layer4_out[6665] ^ layer4_out[6666]);
    assign layer5_out[2005] = ~(layer4_out[265] & layer4_out[266]);
    assign layer5_out[2006] = layer4_out[1475] ^ layer4_out[1476];
    assign layer5_out[2007] = ~layer4_out[6907] | layer4_out[6906];
    assign layer5_out[2008] = ~(layer4_out[5762] & layer4_out[5763]);
    assign layer5_out[2009] = layer4_out[1455] ^ layer4_out[1456];
    assign layer5_out[2010] = ~layer4_out[5292];
    assign layer5_out[2011] = ~(layer4_out[7314] ^ layer4_out[7315]);
    assign layer5_out[2012] = layer4_out[1482];
    assign layer5_out[2013] = ~layer4_out[4145];
    assign layer5_out[2014] = ~(layer4_out[4104] | layer4_out[4105]);
    assign layer5_out[2015] = layer4_out[5878];
    assign layer5_out[2016] = layer4_out[324];
    assign layer5_out[2017] = layer4_out[7815];
    assign layer5_out[2018] = ~layer4_out[6219];
    assign layer5_out[2019] = ~layer4_out[2584];
    assign layer5_out[2020] = layer4_out[6327];
    assign layer5_out[2021] = ~layer4_out[5080];
    assign layer5_out[2022] = ~layer4_out[4506];
    assign layer5_out[2023] = layer4_out[2505] & ~layer4_out[2504];
    assign layer5_out[2024] = ~layer4_out[7483];
    assign layer5_out[2025] = layer4_out[1860] | layer4_out[1861];
    assign layer5_out[2026] = ~layer4_out[5091] | layer4_out[5092];
    assign layer5_out[2027] = ~layer4_out[476];
    assign layer5_out[2028] = ~(layer4_out[1048] ^ layer4_out[1049]);
    assign layer5_out[2029] = layer4_out[1110];
    assign layer5_out[2030] = layer4_out[448];
    assign layer5_out[2031] = ~layer4_out[6994];
    assign layer5_out[2032] = layer4_out[5717] & ~layer4_out[5718];
    assign layer5_out[2033] = ~layer4_out[3540] | layer4_out[3541];
    assign layer5_out[2034] = layer4_out[3064] | layer4_out[3065];
    assign layer5_out[2035] = ~(layer4_out[3805] ^ layer4_out[3806]);
    assign layer5_out[2036] = ~(layer4_out[4087] ^ layer4_out[4088]);
    assign layer5_out[2037] = ~layer4_out[7609];
    assign layer5_out[2038] = ~layer4_out[2111];
    assign layer5_out[2039] = ~(layer4_out[7300] ^ layer4_out[7301]);
    assign layer5_out[2040] = layer4_out[6132] & layer4_out[6133];
    assign layer5_out[2041] = layer4_out[197] & ~layer4_out[196];
    assign layer5_out[2042] = layer4_out[2988] & layer4_out[2989];
    assign layer5_out[2043] = layer4_out[6178] | layer4_out[6179];
    assign layer5_out[2044] = layer4_out[184];
    assign layer5_out[2045] = layer4_out[1410] & ~layer4_out[1409];
    assign layer5_out[2046] = ~layer4_out[649] | layer4_out[648];
    assign layer5_out[2047] = layer4_out[4387];
    assign layer5_out[2048] = ~layer4_out[1689] | layer4_out[1690];
    assign layer5_out[2049] = layer4_out[7477];
    assign layer5_out[2050] = ~layer4_out[3461];
    assign layer5_out[2051] = layer4_out[851];
    assign layer5_out[2052] = layer4_out[7798];
    assign layer5_out[2053] = ~layer4_out[2668];
    assign layer5_out[2054] = layer4_out[4129];
    assign layer5_out[2055] = ~layer4_out[5573];
    assign layer5_out[2056] = ~layer4_out[1976];
    assign layer5_out[2057] = ~layer4_out[7064];
    assign layer5_out[2058] = layer4_out[5005];
    assign layer5_out[2059] = layer4_out[2666];
    assign layer5_out[2060] = layer4_out[1487] & ~layer4_out[1486];
    assign layer5_out[2061] = ~(layer4_out[4112] ^ layer4_out[4113]);
    assign layer5_out[2062] = layer4_out[445];
    assign layer5_out[2063] = layer4_out[4660] ^ layer4_out[4661];
    assign layer5_out[2064] = ~(layer4_out[7957] ^ layer4_out[7958]);
    assign layer5_out[2065] = layer4_out[1411] ^ layer4_out[1412];
    assign layer5_out[2066] = layer4_out[7575];
    assign layer5_out[2067] = layer4_out[919];
    assign layer5_out[2068] = ~layer4_out[3986];
    assign layer5_out[2069] = layer4_out[4493] ^ layer4_out[4494];
    assign layer5_out[2070] = ~layer4_out[2656];
    assign layer5_out[2071] = ~layer4_out[2549];
    assign layer5_out[2072] = layer4_out[2882] ^ layer4_out[2883];
    assign layer5_out[2073] = layer4_out[2510] ^ layer4_out[2511];
    assign layer5_out[2074] = ~(layer4_out[1192] & layer4_out[1193]);
    assign layer5_out[2075] = layer4_out[6775] | layer4_out[6776];
    assign layer5_out[2076] = ~(layer4_out[2259] ^ layer4_out[2260]);
    assign layer5_out[2077] = layer4_out[98] ^ layer4_out[99];
    assign layer5_out[2078] = layer4_out[6722] & ~layer4_out[6721];
    assign layer5_out[2079] = ~(layer4_out[6666] ^ layer4_out[6667]);
    assign layer5_out[2080] = ~(layer4_out[7963] ^ layer4_out[7964]);
    assign layer5_out[2081] = ~layer4_out[6792];
    assign layer5_out[2082] = ~(layer4_out[4084] & layer4_out[4085]);
    assign layer5_out[2083] = ~(layer4_out[3950] | layer4_out[3951]);
    assign layer5_out[2084] = layer4_out[4987] ^ layer4_out[4988];
    assign layer5_out[2085] = layer4_out[1189];
    assign layer5_out[2086] = layer4_out[5116];
    assign layer5_out[2087] = ~layer4_out[2799];
    assign layer5_out[2088] = layer4_out[574];
    assign layer5_out[2089] = layer4_out[520] & layer4_out[521];
    assign layer5_out[2090] = ~layer4_out[6038] | layer4_out[6039];
    assign layer5_out[2091] = ~layer4_out[1834];
    assign layer5_out[2092] = ~layer4_out[3582];
    assign layer5_out[2093] = layer4_out[6961] ^ layer4_out[6962];
    assign layer5_out[2094] = layer4_out[5949] ^ layer4_out[5950];
    assign layer5_out[2095] = ~layer4_out[2172];
    assign layer5_out[2096] = ~layer4_out[1349];
    assign layer5_out[2097] = layer4_out[2930];
    assign layer5_out[2098] = layer4_out[2934] & layer4_out[2935];
    assign layer5_out[2099] = layer4_out[5829] | layer4_out[5830];
    assign layer5_out[2100] = ~(layer4_out[2628] ^ layer4_out[2629]);
    assign layer5_out[2101] = layer4_out[620];
    assign layer5_out[2102] = ~layer4_out[6044];
    assign layer5_out[2103] = ~layer4_out[3519];
    assign layer5_out[2104] = ~layer4_out[5530];
    assign layer5_out[2105] = layer4_out[2399] & layer4_out[2400];
    assign layer5_out[2106] = ~layer4_out[3158];
    assign layer5_out[2107] = ~(layer4_out[6874] ^ layer4_out[6875]);
    assign layer5_out[2108] = ~(layer4_out[6133] ^ layer4_out[6134]);
    assign layer5_out[2109] = layer4_out[1777];
    assign layer5_out[2110] = ~layer4_out[633] | layer4_out[632];
    assign layer5_out[2111] = ~layer4_out[1038] | layer4_out[1037];
    assign layer5_out[2112] = ~layer4_out[3461];
    assign layer5_out[2113] = ~layer4_out[4596];
    assign layer5_out[2114] = ~(layer4_out[5509] ^ layer4_out[5510]);
    assign layer5_out[2115] = layer4_out[7563] & layer4_out[7564];
    assign layer5_out[2116] = ~layer4_out[1057];
    assign layer5_out[2117] = layer4_out[1959] & ~layer4_out[1960];
    assign layer5_out[2118] = layer4_out[4179] ^ layer4_out[4180];
    assign layer5_out[2119] = ~(layer4_out[4371] & layer4_out[4372]);
    assign layer5_out[2120] = ~layer4_out[4238] | layer4_out[4239];
    assign layer5_out[2121] = layer4_out[626] & layer4_out[627];
    assign layer5_out[2122] = layer4_out[4857];
    assign layer5_out[2123] = layer4_out[6053] & layer4_out[6054];
    assign layer5_out[2124] = layer4_out[908] & layer4_out[909];
    assign layer5_out[2125] = layer4_out[5760] & layer4_out[5761];
    assign layer5_out[2126] = layer4_out[6217] ^ layer4_out[6218];
    assign layer5_out[2127] = ~layer4_out[4694] | layer4_out[4695];
    assign layer5_out[2128] = ~(layer4_out[6401] ^ layer4_out[6402]);
    assign layer5_out[2129] = ~layer4_out[3173] | layer4_out[3172];
    assign layer5_out[2130] = ~layer4_out[2954];
    assign layer5_out[2131] = layer4_out[1238];
    assign layer5_out[2132] = layer4_out[1290];
    assign layer5_out[2133] = ~layer4_out[1325] | layer4_out[1324];
    assign layer5_out[2134] = ~layer4_out[1435];
    assign layer5_out[2135] = layer4_out[3342] | layer4_out[3343];
    assign layer5_out[2136] = ~layer4_out[7184];
    assign layer5_out[2137] = ~(layer4_out[3087] ^ layer4_out[3088]);
    assign layer5_out[2138] = layer4_out[7191];
    assign layer5_out[2139] = layer4_out[5034] & ~layer4_out[5033];
    assign layer5_out[2140] = layer4_out[1070];
    assign layer5_out[2141] = ~layer4_out[5903];
    assign layer5_out[2142] = ~(layer4_out[4227] ^ layer4_out[4228]);
    assign layer5_out[2143] = ~(layer4_out[5592] ^ layer4_out[5593]);
    assign layer5_out[2144] = layer4_out[4472] ^ layer4_out[4473];
    assign layer5_out[2145] = layer4_out[3691] ^ layer4_out[3692];
    assign layer5_out[2146] = layer4_out[5805];
    assign layer5_out[2147] = layer4_out[7415] & ~layer4_out[7416];
    assign layer5_out[2148] = layer4_out[3549];
    assign layer5_out[2149] = ~layer4_out[4703];
    assign layer5_out[2150] = layer4_out[3408] ^ layer4_out[3409];
    assign layer5_out[2151] = ~layer4_out[4319] | layer4_out[4320];
    assign layer5_out[2152] = ~layer4_out[1481] | layer4_out[1482];
    assign layer5_out[2153] = layer4_out[7939];
    assign layer5_out[2154] = layer4_out[4326];
    assign layer5_out[2155] = ~(layer4_out[6993] & layer4_out[6994]);
    assign layer5_out[2156] = layer4_out[6340];
    assign layer5_out[2157] = ~(layer4_out[1655] | layer4_out[1656]);
    assign layer5_out[2158] = layer4_out[1084] & ~layer4_out[1083];
    assign layer5_out[2159] = layer4_out[2680] & ~layer4_out[2679];
    assign layer5_out[2160] = ~(layer4_out[34] | layer4_out[35]);
    assign layer5_out[2161] = layer4_out[225];
    assign layer5_out[2162] = ~(layer4_out[1184] ^ layer4_out[1185]);
    assign layer5_out[2163] = ~layer4_out[3538] | layer4_out[3539];
    assign layer5_out[2164] = layer4_out[6593] & layer4_out[6594];
    assign layer5_out[2165] = layer4_out[1605] & ~layer4_out[1604];
    assign layer5_out[2166] = ~(layer4_out[4406] ^ layer4_out[4407]);
    assign layer5_out[2167] = layer4_out[2146] & ~layer4_out[2145];
    assign layer5_out[2168] = ~(layer4_out[4358] ^ layer4_out[4359]);
    assign layer5_out[2169] = layer4_out[3715] & ~layer4_out[3716];
    assign layer5_out[2170] = ~layer4_out[6080];
    assign layer5_out[2171] = layer4_out[1453];
    assign layer5_out[2172] = ~layer4_out[7738];
    assign layer5_out[2173] = ~(layer4_out[1164] | layer4_out[1165]);
    assign layer5_out[2174] = ~(layer4_out[5574] ^ layer4_out[5575]);
    assign layer5_out[2175] = ~(layer4_out[1195] & layer4_out[1196]);
    assign layer5_out[2176] = layer4_out[3713] ^ layer4_out[3714];
    assign layer5_out[2177] = ~layer4_out[1490];
    assign layer5_out[2178] = ~layer4_out[1449];
    assign layer5_out[2179] = layer4_out[6364] ^ layer4_out[6365];
    assign layer5_out[2180] = ~layer4_out[4709];
    assign layer5_out[2181] = ~layer4_out[5336];
    assign layer5_out[2182] = layer4_out[1543] ^ layer4_out[1544];
    assign layer5_out[2183] = ~layer4_out[6486];
    assign layer5_out[2184] = ~layer4_out[3793];
    assign layer5_out[2185] = layer4_out[198] | layer4_out[199];
    assign layer5_out[2186] = ~layer4_out[6283];
    assign layer5_out[2187] = ~layer4_out[5213];
    assign layer5_out[2188] = ~layer4_out[3118];
    assign layer5_out[2189] = ~(layer4_out[1572] & layer4_out[1573]);
    assign layer5_out[2190] = ~(layer4_out[623] ^ layer4_out[624]);
    assign layer5_out[2191] = ~(layer4_out[2048] ^ layer4_out[2049]);
    assign layer5_out[2192] = layer4_out[61] & ~layer4_out[62];
    assign layer5_out[2193] = layer4_out[7193] ^ layer4_out[7194];
    assign layer5_out[2194] = layer4_out[2829];
    assign layer5_out[2195] = layer4_out[1338] ^ layer4_out[1339];
    assign layer5_out[2196] = layer4_out[6498] & ~layer4_out[6497];
    assign layer5_out[2197] = layer4_out[3854] & ~layer4_out[3853];
    assign layer5_out[2198] = layer4_out[669] & ~layer4_out[668];
    assign layer5_out[2199] = ~(layer4_out[89] ^ layer4_out[90]);
    assign layer5_out[2200] = layer4_out[6289] ^ layer4_out[6290];
    assign layer5_out[2201] = ~layer4_out[6663];
    assign layer5_out[2202] = layer4_out[99] & ~layer4_out[100];
    assign layer5_out[2203] = layer4_out[7405] ^ layer4_out[7406];
    assign layer5_out[2204] = layer4_out[577] ^ layer4_out[578];
    assign layer5_out[2205] = ~(layer4_out[470] ^ layer4_out[471]);
    assign layer5_out[2206] = layer4_out[3026] | layer4_out[3027];
    assign layer5_out[2207] = ~(layer4_out[5602] & layer4_out[5603]);
    assign layer5_out[2208] = layer4_out[3859];
    assign layer5_out[2209] = layer4_out[3387];
    assign layer5_out[2210] = ~(layer4_out[1385] | layer4_out[1386]);
    assign layer5_out[2211] = ~layer4_out[4194];
    assign layer5_out[2212] = layer4_out[5444];
    assign layer5_out[2213] = layer4_out[1054] ^ layer4_out[1055];
    assign layer5_out[2214] = layer4_out[6148];
    assign layer5_out[2215] = ~layer4_out[1417] | layer4_out[1418];
    assign layer5_out[2216] = ~layer4_out[4917];
    assign layer5_out[2217] = ~layer4_out[5090];
    assign layer5_out[2218] = layer4_out[5635];
    assign layer5_out[2219] = layer4_out[373];
    assign layer5_out[2220] = ~layer4_out[6544];
    assign layer5_out[2221] = layer4_out[5458] & ~layer4_out[5457];
    assign layer5_out[2222] = layer4_out[4633] & ~layer4_out[4634];
    assign layer5_out[2223] = ~(layer4_out[2080] ^ layer4_out[2081]);
    assign layer5_out[2224] = ~layer4_out[209];
    assign layer5_out[2225] = ~layer4_out[3255];
    assign layer5_out[2226] = ~layer4_out[2277] | layer4_out[2276];
    assign layer5_out[2227] = layer4_out[6099];
    assign layer5_out[2228] = layer4_out[521];
    assign layer5_out[2229] = ~(layer4_out[7199] | layer4_out[7200]);
    assign layer5_out[2230] = ~layer4_out[7963] | layer4_out[7962];
    assign layer5_out[2231] = layer4_out[3204];
    assign layer5_out[2232] = layer4_out[3226] & layer4_out[3227];
    assign layer5_out[2233] = layer4_out[510];
    assign layer5_out[2234] = ~(layer4_out[4924] ^ layer4_out[4925]);
    assign layer5_out[2235] = ~layer4_out[451] | layer4_out[452];
    assign layer5_out[2236] = ~layer4_out[1212];
    assign layer5_out[2237] = ~layer4_out[2209];
    assign layer5_out[2238] = layer4_out[7095];
    assign layer5_out[2239] = layer4_out[153] ^ layer4_out[154];
    assign layer5_out[2240] = ~layer4_out[2142];
    assign layer5_out[2241] = layer4_out[2473];
    assign layer5_out[2242] = layer4_out[1419];
    assign layer5_out[2243] = ~layer4_out[4032];
    assign layer5_out[2244] = layer4_out[7291] & ~layer4_out[7292];
    assign layer5_out[2245] = ~layer4_out[1262] | layer4_out[1261];
    assign layer5_out[2246] = layer4_out[1080];
    assign layer5_out[2247] = layer4_out[1626];
    assign layer5_out[2248] = ~(layer4_out[5466] ^ layer4_out[5467]);
    assign layer5_out[2249] = layer4_out[6245] & ~layer4_out[6246];
    assign layer5_out[2250] = layer4_out[5449] & layer4_out[5450];
    assign layer5_out[2251] = layer4_out[1394] & ~layer4_out[1393];
    assign layer5_out[2252] = ~(layer4_out[3520] & layer4_out[3521]);
    assign layer5_out[2253] = layer4_out[6822] ^ layer4_out[6823];
    assign layer5_out[2254] = layer4_out[6849];
    assign layer5_out[2255] = ~(layer4_out[3169] | layer4_out[3170]);
    assign layer5_out[2256] = layer4_out[1557] & ~layer4_out[1558];
    assign layer5_out[2257] = ~layer4_out[7609] | layer4_out[7610];
    assign layer5_out[2258] = layer4_out[745] ^ layer4_out[746];
    assign layer5_out[2259] = ~layer4_out[2254];
    assign layer5_out[2260] = layer4_out[4689];
    assign layer5_out[2261] = ~(layer4_out[4234] ^ layer4_out[4235]);
    assign layer5_out[2262] = layer4_out[510];
    assign layer5_out[2263] = ~layer4_out[3000] | layer4_out[2999];
    assign layer5_out[2264] = layer4_out[1892];
    assign layer5_out[2265] = layer4_out[1311];
    assign layer5_out[2266] = layer4_out[6856] ^ layer4_out[6857];
    assign layer5_out[2267] = layer4_out[5922] | layer4_out[5923];
    assign layer5_out[2268] = layer4_out[2580];
    assign layer5_out[2269] = ~(layer4_out[3668] | layer4_out[3669]);
    assign layer5_out[2270] = ~(layer4_out[3905] ^ layer4_out[3906]);
    assign layer5_out[2271] = ~(layer4_out[7456] | layer4_out[7457]);
    assign layer5_out[2272] = layer4_out[887] | layer4_out[888];
    assign layer5_out[2273] = ~layer4_out[1087];
    assign layer5_out[2274] = ~(layer4_out[7652] | layer4_out[7653]);
    assign layer5_out[2275] = layer4_out[2225] ^ layer4_out[2226];
    assign layer5_out[2276] = layer4_out[5859];
    assign layer5_out[2277] = ~layer4_out[5734];
    assign layer5_out[2278] = layer4_out[6397];
    assign layer5_out[2279] = ~layer4_out[7761];
    assign layer5_out[2280] = layer4_out[2];
    assign layer5_out[2281] = layer4_out[3789];
    assign layer5_out[2282] = layer4_out[5722];
    assign layer5_out[2283] = layer4_out[3484];
    assign layer5_out[2284] = ~(layer4_out[922] ^ layer4_out[923]);
    assign layer5_out[2285] = layer4_out[6812];
    assign layer5_out[2286] = ~layer4_out[2549];
    assign layer5_out[2287] = ~layer4_out[5668];
    assign layer5_out[2288] = layer4_out[5776];
    assign layer5_out[2289] = ~layer4_out[4555] | layer4_out[4556];
    assign layer5_out[2290] = ~layer4_out[7994];
    assign layer5_out[2291] = ~layer4_out[6685];
    assign layer5_out[2292] = ~(layer4_out[7215] ^ layer4_out[7216]);
    assign layer5_out[2293] = layer4_out[2572] | layer4_out[2573];
    assign layer5_out[2294] = ~(layer4_out[1769] ^ layer4_out[1770]);
    assign layer5_out[2295] = ~layer4_out[7159];
    assign layer5_out[2296] = layer4_out[291] & ~layer4_out[290];
    assign layer5_out[2297] = ~layer4_out[1726];
    assign layer5_out[2298] = layer4_out[2248] ^ layer4_out[2249];
    assign layer5_out[2299] = layer4_out[2691] & ~layer4_out[2690];
    assign layer5_out[2300] = layer4_out[1187] ^ layer4_out[1188];
    assign layer5_out[2301] = ~layer4_out[4863] | layer4_out[4864];
    assign layer5_out[2302] = layer4_out[7282];
    assign layer5_out[2303] = ~layer4_out[1039];
    assign layer5_out[2304] = ~(layer4_out[2044] ^ layer4_out[2045]);
    assign layer5_out[2305] = ~(layer4_out[1714] ^ layer4_out[1715]);
    assign layer5_out[2306] = ~(layer4_out[942] ^ layer4_out[943]);
    assign layer5_out[2307] = ~layer4_out[6489] | layer4_out[6490];
    assign layer5_out[2308] = ~layer4_out[415];
    assign layer5_out[2309] = layer4_out[5836];
    assign layer5_out[2310] = layer4_out[3420] ^ layer4_out[3421];
    assign layer5_out[2311] = layer4_out[5993] ^ layer4_out[5994];
    assign layer5_out[2312] = layer4_out[4978] ^ layer4_out[4979];
    assign layer5_out[2313] = layer4_out[2097] ^ layer4_out[2098];
    assign layer5_out[2314] = ~(layer4_out[692] ^ layer4_out[693]);
    assign layer5_out[2315] = ~layer4_out[1872];
    assign layer5_out[2316] = ~layer4_out[7580];
    assign layer5_out[2317] = ~layer4_out[2087];
    assign layer5_out[2318] = ~layer4_out[3037];
    assign layer5_out[2319] = layer4_out[2616] & ~layer4_out[2617];
    assign layer5_out[2320] = layer4_out[617];
    assign layer5_out[2321] = layer4_out[6679] & ~layer4_out[6678];
    assign layer5_out[2322] = layer4_out[1352] & ~layer4_out[1351];
    assign layer5_out[2323] = ~layer4_out[2540];
    assign layer5_out[2324] = layer4_out[4562] & ~layer4_out[4561];
    assign layer5_out[2325] = ~layer4_out[633];
    assign layer5_out[2326] = ~layer4_out[4914];
    assign layer5_out[2327] = ~layer4_out[3005];
    assign layer5_out[2328] = layer4_out[4762] ^ layer4_out[4763];
    assign layer5_out[2329] = layer4_out[664];
    assign layer5_out[2330] = ~layer4_out[2781];
    assign layer5_out[2331] = ~(layer4_out[2390] & layer4_out[2391]);
    assign layer5_out[2332] = ~(layer4_out[3384] ^ layer4_out[3385]);
    assign layer5_out[2333] = ~layer4_out[7576];
    assign layer5_out[2334] = ~layer4_out[6216];
    assign layer5_out[2335] = ~(layer4_out[398] & layer4_out[399]);
    assign layer5_out[2336] = ~layer4_out[5415];
    assign layer5_out[2337] = ~(layer4_out[742] ^ layer4_out[743]);
    assign layer5_out[2338] = ~layer4_out[6606];
    assign layer5_out[2339] = layer4_out[7516] & ~layer4_out[7517];
    assign layer5_out[2340] = layer4_out[3523];
    assign layer5_out[2341] = ~(layer4_out[3842] ^ layer4_out[3843]);
    assign layer5_out[2342] = layer4_out[1216];
    assign layer5_out[2343] = layer4_out[6564] ^ layer4_out[6565];
    assign layer5_out[2344] = layer4_out[941] & ~layer4_out[940];
    assign layer5_out[2345] = layer4_out[7775];
    assign layer5_out[2346] = ~(layer4_out[2678] ^ layer4_out[2679]);
    assign layer5_out[2347] = layer4_out[5484] ^ layer4_out[5485];
    assign layer5_out[2348] = ~(layer4_out[7016] ^ layer4_out[7017]);
    assign layer5_out[2349] = layer4_out[1932];
    assign layer5_out[2350] = layer4_out[7749] & ~layer4_out[7750];
    assign layer5_out[2351] = layer4_out[5940] ^ layer4_out[5941];
    assign layer5_out[2352] = layer4_out[6724] & ~layer4_out[6725];
    assign layer5_out[2353] = ~(layer4_out[6101] ^ layer4_out[6102]);
    assign layer5_out[2354] = ~layer4_out[579] | layer4_out[578];
    assign layer5_out[2355] = layer4_out[5105];
    assign layer5_out[2356] = ~layer4_out[4205];
    assign layer5_out[2357] = layer4_out[734] ^ layer4_out[735];
    assign layer5_out[2358] = layer4_out[5469] & ~layer4_out[5468];
    assign layer5_out[2359] = layer4_out[2632];
    assign layer5_out[2360] = layer4_out[3083] & ~layer4_out[3084];
    assign layer5_out[2361] = layer4_out[6754];
    assign layer5_out[2362] = layer4_out[7634];
    assign layer5_out[2363] = ~layer4_out[3667];
    assign layer5_out[2364] = ~layer4_out[1900] | layer4_out[1901];
    assign layer5_out[2365] = ~layer4_out[7934];
    assign layer5_out[2366] = ~(layer4_out[1044] ^ layer4_out[1045]);
    assign layer5_out[2367] = ~(layer4_out[2324] ^ layer4_out[2325]);
    assign layer5_out[2368] = layer4_out[4295];
    assign layer5_out[2369] = ~layer4_out[660];
    assign layer5_out[2370] = layer4_out[6917];
    assign layer5_out[2371] = ~layer4_out[514] | layer4_out[515];
    assign layer5_out[2372] = ~(layer4_out[4981] | layer4_out[4982]);
    assign layer5_out[2373] = layer4_out[3868];
    assign layer5_out[2374] = ~layer4_out[3020];
    assign layer5_out[2375] = layer4_out[1222] ^ layer4_out[1223];
    assign layer5_out[2376] = ~layer4_out[5446];
    assign layer5_out[2377] = ~layer4_out[396];
    assign layer5_out[2378] = ~(layer4_out[5175] | layer4_out[5176]);
    assign layer5_out[2379] = ~layer4_out[6789];
    assign layer5_out[2380] = ~(layer4_out[1120] ^ layer4_out[1121]);
    assign layer5_out[2381] = ~layer4_out[3683];
    assign layer5_out[2382] = layer4_out[6481] & layer4_out[6482];
    assign layer5_out[2383] = layer4_out[7074] & layer4_out[7075];
    assign layer5_out[2384] = ~layer4_out[5966];
    assign layer5_out[2385] = layer4_out[2165] & layer4_out[2166];
    assign layer5_out[2386] = ~(layer4_out[6135] ^ layer4_out[6136]);
    assign layer5_out[2387] = layer4_out[1534] & ~layer4_out[1535];
    assign layer5_out[2388] = layer4_out[2763];
    assign layer5_out[2389] = layer4_out[6917];
    assign layer5_out[2390] = layer4_out[4107];
    assign layer5_out[2391] = ~(layer4_out[7175] ^ layer4_out[7176]);
    assign layer5_out[2392] = ~(layer4_out[206] ^ layer4_out[207]);
    assign layer5_out[2393] = ~layer4_out[4919];
    assign layer5_out[2394] = layer4_out[1571] & ~layer4_out[1572];
    assign layer5_out[2395] = ~layer4_out[2046];
    assign layer5_out[2396] = layer4_out[5565];
    assign layer5_out[2397] = ~layer4_out[1473] | layer4_out[1472];
    assign layer5_out[2398] = ~layer4_out[2351] | layer4_out[2350];
    assign layer5_out[2399] = layer4_out[4236];
    assign layer5_out[2400] = layer4_out[6014] & ~layer4_out[6013];
    assign layer5_out[2401] = ~(layer4_out[4108] ^ layer4_out[4109]);
    assign layer5_out[2402] = ~layer4_out[2324];
    assign layer5_out[2403] = ~(layer4_out[5715] ^ layer4_out[5716]);
    assign layer5_out[2404] = ~layer4_out[1897] | layer4_out[1898];
    assign layer5_out[2405] = ~layer4_out[5162];
    assign layer5_out[2406] = layer4_out[4252] ^ layer4_out[4253];
    assign layer5_out[2407] = ~(layer4_out[7275] ^ layer4_out[7276]);
    assign layer5_out[2408] = layer4_out[2735] | layer4_out[2736];
    assign layer5_out[2409] = layer4_out[5191] ^ layer4_out[5192];
    assign layer5_out[2410] = layer4_out[6508] ^ layer4_out[6509];
    assign layer5_out[2411] = layer4_out[5355] & layer4_out[5356];
    assign layer5_out[2412] = layer4_out[2518] | layer4_out[2519];
    assign layer5_out[2413] = layer4_out[2257] ^ layer4_out[2258];
    assign layer5_out[2414] = ~(layer4_out[4894] ^ layer4_out[4895]);
    assign layer5_out[2415] = layer4_out[6853] & ~layer4_out[6852];
    assign layer5_out[2416] = layer4_out[7842];
    assign layer5_out[2417] = ~layer4_out[6914];
    assign layer5_out[2418] = layer4_out[5844] & ~layer4_out[5845];
    assign layer5_out[2419] = layer4_out[7419] & layer4_out[7420];
    assign layer5_out[2420] = layer4_out[5750] ^ layer4_out[5751];
    assign layer5_out[2421] = ~(layer4_out[2152] ^ layer4_out[2153]);
    assign layer5_out[2422] = ~layer4_out[1909];
    assign layer5_out[2423] = ~layer4_out[7332] | layer4_out[7331];
    assign layer5_out[2424] = layer4_out[7093] ^ layer4_out[7094];
    assign layer5_out[2425] = layer4_out[7052] ^ layer4_out[7053];
    assign layer5_out[2426] = ~(layer4_out[3719] | layer4_out[3720]);
    assign layer5_out[2427] = ~(layer4_out[3641] & layer4_out[3642]);
    assign layer5_out[2428] = layer4_out[4930] ^ layer4_out[4931];
    assign layer5_out[2429] = layer4_out[386] & layer4_out[387];
    assign layer5_out[2430] = ~(layer4_out[4053] ^ layer4_out[4054]);
    assign layer5_out[2431] = layer4_out[1929] | layer4_out[1930];
    assign layer5_out[2432] = ~(layer4_out[1392] ^ layer4_out[1393]);
    assign layer5_out[2433] = ~(layer4_out[7570] | layer4_out[7571]);
    assign layer5_out[2434] = layer4_out[7535];
    assign layer5_out[2435] = layer4_out[5826] ^ layer4_out[5827];
    assign layer5_out[2436] = layer4_out[5460] & ~layer4_out[5459];
    assign layer5_out[2437] = layer4_out[4712] & ~layer4_out[4711];
    assign layer5_out[2438] = layer4_out[1369];
    assign layer5_out[2439] = layer4_out[3410];
    assign layer5_out[2440] = ~layer4_out[6426];
    assign layer5_out[2441] = layer4_out[310];
    assign layer5_out[2442] = layer4_out[1929];
    assign layer5_out[2443] = layer4_out[5168] ^ layer4_out[5169];
    assign layer5_out[2444] = layer4_out[7709];
    assign layer5_out[2445] = layer4_out[6992] & ~layer4_out[6993];
    assign layer5_out[2446] = layer4_out[6762] & layer4_out[6763];
    assign layer5_out[2447] = ~layer4_out[5931] | layer4_out[5932];
    assign layer5_out[2448] = layer4_out[6996] ^ layer4_out[6997];
    assign layer5_out[2449] = ~(layer4_out[3670] | layer4_out[3671]);
    assign layer5_out[2450] = ~layer4_out[1099];
    assign layer5_out[2451] = ~(layer4_out[4542] | layer4_out[4543]);
    assign layer5_out[2452] = layer4_out[58] & ~layer4_out[57];
    assign layer5_out[2453] = ~(layer4_out[5845] | layer4_out[5846]);
    assign layer5_out[2454] = ~(layer4_out[4974] | layer4_out[4975]);
    assign layer5_out[2455] = layer4_out[4380] ^ layer4_out[4381];
    assign layer5_out[2456] = ~layer4_out[6372];
    assign layer5_out[2457] = ~layer4_out[3743];
    assign layer5_out[2458] = ~layer4_out[7654] | layer4_out[7653];
    assign layer5_out[2459] = ~layer4_out[5027];
    assign layer5_out[2460] = ~(layer4_out[6299] ^ layer4_out[6300]);
    assign layer5_out[2461] = ~(layer4_out[2103] ^ layer4_out[2104]);
    assign layer5_out[2462] = ~(layer4_out[3638] & layer4_out[3639]);
    assign layer5_out[2463] = ~(layer4_out[3808] ^ layer4_out[3809]);
    assign layer5_out[2464] = layer4_out[381] | layer4_out[382];
    assign layer5_out[2465] = layer4_out[6409] & ~layer4_out[6408];
    assign layer5_out[2466] = layer4_out[6781];
    assign layer5_out[2467] = layer4_out[4432] ^ layer4_out[4433];
    assign layer5_out[2468] = ~(layer4_out[4143] | layer4_out[4144]);
    assign layer5_out[2469] = ~layer4_out[7986] | layer4_out[7985];
    assign layer5_out[2470] = ~(layer4_out[4884] & layer4_out[4885]);
    assign layer5_out[2471] = layer4_out[1213] ^ layer4_out[1214];
    assign layer5_out[2472] = ~(layer4_out[7625] ^ layer4_out[7626]);
    assign layer5_out[2473] = ~(layer4_out[7795] ^ layer4_out[7796]);
    assign layer5_out[2474] = ~layer4_out[6970];
    assign layer5_out[2475] = layer4_out[3376] & ~layer4_out[3375];
    assign layer5_out[2476] = layer4_out[4110];
    assign layer5_out[2477] = ~layer4_out[4682];
    assign layer5_out[2478] = layer4_out[2512] & layer4_out[2513];
    assign layer5_out[2479] = layer4_out[4] & ~layer4_out[5];
    assign layer5_out[2480] = layer4_out[2227] & layer4_out[2228];
    assign layer5_out[2481] = layer4_out[4081] | layer4_out[4082];
    assign layer5_out[2482] = ~layer4_out[5139] | layer4_out[5138];
    assign layer5_out[2483] = layer4_out[4443];
    assign layer5_out[2484] = ~(layer4_out[3497] ^ layer4_out[3498]);
    assign layer5_out[2485] = ~(layer4_out[6776] ^ layer4_out[6777]);
    assign layer5_out[2486] = ~layer4_out[3780];
    assign layer5_out[2487] = ~layer4_out[2529];
    assign layer5_out[2488] = layer4_out[3452] & layer4_out[3453];
    assign layer5_out[2489] = layer4_out[642];
    assign layer5_out[2490] = ~(layer4_out[7192] | layer4_out[7193]);
    assign layer5_out[2491] = layer4_out[3950];
    assign layer5_out[2492] = layer4_out[3235];
    assign layer5_out[2493] = layer4_out[4410];
    assign layer5_out[2494] = layer4_out[3816] & ~layer4_out[3817];
    assign layer5_out[2495] = ~layer4_out[2567] | layer4_out[2568];
    assign layer5_out[2496] = layer4_out[5758] ^ layer4_out[5759];
    assign layer5_out[2497] = layer4_out[5265] ^ layer4_out[5266];
    assign layer5_out[2498] = ~layer4_out[1343];
    assign layer5_out[2499] = ~(layer4_out[3976] ^ layer4_out[3977]);
    assign layer5_out[2500] = layer4_out[1570] & ~layer4_out[1571];
    assign layer5_out[2501] = layer4_out[3124] & ~layer4_out[3125];
    assign layer5_out[2502] = layer4_out[4025] ^ layer4_out[4026];
    assign layer5_out[2503] = layer4_out[5875] ^ layer4_out[5876];
    assign layer5_out[2504] = ~layer4_out[3786];
    assign layer5_out[2505] = ~layer4_out[5308];
    assign layer5_out[2506] = ~(layer4_out[1828] ^ layer4_out[1829]);
    assign layer5_out[2507] = ~layer4_out[6859];
    assign layer5_out[2508] = ~(layer4_out[1106] | layer4_out[1107]);
    assign layer5_out[2509] = ~layer4_out[335];
    assign layer5_out[2510] = layer4_out[840];
    assign layer5_out[2511] = ~layer4_out[7938];
    assign layer5_out[2512] = layer4_out[1765] & ~layer4_out[1766];
    assign layer5_out[2513] = ~layer4_out[4822];
    assign layer5_out[2514] = layer4_out[6276] & ~layer4_out[6277];
    assign layer5_out[2515] = ~(layer4_out[1767] | layer4_out[1768]);
    assign layer5_out[2516] = layer4_out[4396] ^ layer4_out[4397];
    assign layer5_out[2517] = layer4_out[6963];
    assign layer5_out[2518] = layer4_out[7095] ^ layer4_out[7096];
    assign layer5_out[2519] = layer4_out[7919];
    assign layer5_out[2520] = layer4_out[2495] ^ layer4_out[2496];
    assign layer5_out[2521] = ~(layer4_out[3702] ^ layer4_out[3703]);
    assign layer5_out[2522] = ~layer4_out[3532];
    assign layer5_out[2523] = layer4_out[3716] ^ layer4_out[3717];
    assign layer5_out[2524] = ~layer4_out[4590];
    assign layer5_out[2525] = layer4_out[5649] | layer4_out[5650];
    assign layer5_out[2526] = layer4_out[7065] ^ layer4_out[7066];
    assign layer5_out[2527] = layer4_out[277] & ~layer4_out[278];
    assign layer5_out[2528] = ~layer4_out[238];
    assign layer5_out[2529] = ~layer4_out[4722] | layer4_out[4721];
    assign layer5_out[2530] = ~layer4_out[1530];
    assign layer5_out[2531] = ~layer4_out[4056];
    assign layer5_out[2532] = ~layer4_out[2929];
    assign layer5_out[2533] = layer4_out[3908];
    assign layer5_out[2534] = layer4_out[6409] & ~layer4_out[6410];
    assign layer5_out[2535] = ~layer4_out[818] | layer4_out[817];
    assign layer5_out[2536] = layer4_out[5774] & layer4_out[5775];
    assign layer5_out[2537] = ~layer4_out[7213] | layer4_out[7214];
    assign layer5_out[2538] = ~layer4_out[1806];
    assign layer5_out[2539] = ~layer4_out[585];
    assign layer5_out[2540] = layer4_out[6611];
    assign layer5_out[2541] = layer4_out[5166] & ~layer4_out[5167];
    assign layer5_out[2542] = ~(layer4_out[12] ^ layer4_out[13]);
    assign layer5_out[2543] = ~layer4_out[7955];
    assign layer5_out[2544] = ~(layer4_out[5361] ^ layer4_out[5362]);
    assign layer5_out[2545] = layer4_out[6337];
    assign layer5_out[2546] = layer4_out[2738] & ~layer4_out[2739];
    assign layer5_out[2547] = layer4_out[6551] ^ layer4_out[6552];
    assign layer5_out[2548] = layer4_out[2993] & ~layer4_out[2994];
    assign layer5_out[2549] = ~(layer4_out[4814] ^ layer4_out[4815]);
    assign layer5_out[2550] = ~layer4_out[5908];
    assign layer5_out[2551] = layer4_out[1526];
    assign layer5_out[2552] = ~layer4_out[7965];
    assign layer5_out[2553] = layer4_out[2823];
    assign layer5_out[2554] = layer4_out[3415];
    assign layer5_out[2555] = ~(layer4_out[6472] & layer4_out[6473]);
    assign layer5_out[2556] = ~layer4_out[3139];
    assign layer5_out[2557] = ~layer4_out[5278];
    assign layer5_out[2558] = layer4_out[6897] & ~layer4_out[6898];
    assign layer5_out[2559] = layer4_out[476];
    assign layer5_out[2560] = layer4_out[3450];
    assign layer5_out[2561] = ~layer4_out[2010];
    assign layer5_out[2562] = ~layer4_out[4021];
    assign layer5_out[2563] = layer4_out[4200] ^ layer4_out[4201];
    assign layer5_out[2564] = ~(layer4_out[2602] ^ layer4_out[2603]);
    assign layer5_out[2565] = layer4_out[2469];
    assign layer5_out[2566] = ~(layer4_out[6319] ^ layer4_out[6320]);
    assign layer5_out[2567] = ~layer4_out[4272] | layer4_out[4271];
    assign layer5_out[2568] = ~(layer4_out[5544] | layer4_out[5545]);
    assign layer5_out[2569] = layer4_out[1160] ^ layer4_out[1161];
    assign layer5_out[2570] = layer4_out[4846] & layer4_out[4847];
    assign layer5_out[2571] = ~layer4_out[6627];
    assign layer5_out[2572] = ~(layer4_out[1399] & layer4_out[1400]);
    assign layer5_out[2573] = ~layer4_out[963] | layer4_out[962];
    assign layer5_out[2574] = layer4_out[6110] & ~layer4_out[6109];
    assign layer5_out[2575] = layer4_out[6877] & layer4_out[6878];
    assign layer5_out[2576] = layer4_out[2284];
    assign layer5_out[2577] = layer4_out[1869];
    assign layer5_out[2578] = ~(layer4_out[6474] ^ layer4_out[6475]);
    assign layer5_out[2579] = layer4_out[7126];
    assign layer5_out[2580] = ~layer4_out[3997];
    assign layer5_out[2581] = layer4_out[177] & ~layer4_out[176];
    assign layer5_out[2582] = layer4_out[1069];
    assign layer5_out[2583] = layer4_out[5767];
    assign layer5_out[2584] = layer4_out[5141];
    assign layer5_out[2585] = layer4_out[6390] & ~layer4_out[6391];
    assign layer5_out[2586] = ~layer4_out[4068];
    assign layer5_out[2587] = layer4_out[2408];
    assign layer5_out[2588] = layer4_out[1549];
    assign layer5_out[2589] = ~(layer4_out[1033] ^ layer4_out[1034]);
    assign layer5_out[2590] = ~layer4_out[5730] | layer4_out[5729];
    assign layer5_out[2591] = ~layer4_out[3941];
    assign layer5_out[2592] = ~(layer4_out[4503] & layer4_out[4504]);
    assign layer5_out[2593] = layer4_out[444] ^ layer4_out[445];
    assign layer5_out[2594] = layer4_out[7360];
    assign layer5_out[2595] = ~layer4_out[6415];
    assign layer5_out[2596] = ~(layer4_out[3935] ^ layer4_out[3936]);
    assign layer5_out[2597] = ~(layer4_out[524] | layer4_out[525]);
    assign layer5_out[2598] = ~layer4_out[6523] | layer4_out[6524];
    assign layer5_out[2599] = layer4_out[6292];
    assign layer5_out[2600] = layer4_out[2622];
    assign layer5_out[2601] = layer4_out[1251] & layer4_out[1252];
    assign layer5_out[2602] = ~layer4_out[760] | layer4_out[761];
    assign layer5_out[2603] = layer4_out[5391] ^ layer4_out[5392];
    assign layer5_out[2604] = ~(layer4_out[3168] | layer4_out[3169]);
    assign layer5_out[2605] = ~layer4_out[1885] | layer4_out[1884];
    assign layer5_out[2606] = layer4_out[505];
    assign layer5_out[2607] = ~layer4_out[4619];
    assign layer5_out[2608] = layer4_out[7364];
    assign layer5_out[2609] = ~layer4_out[2461];
    assign layer5_out[2610] = ~layer4_out[2575];
    assign layer5_out[2611] = layer4_out[7188] ^ layer4_out[7189];
    assign layer5_out[2612] = ~(layer4_out[131] ^ layer4_out[132]);
    assign layer5_out[2613] = ~(layer4_out[5239] | layer4_out[5240]);
    assign layer5_out[2614] = layer4_out[5625] & ~layer4_out[5624];
    assign layer5_out[2615] = layer4_out[342] | layer4_out[343];
    assign layer5_out[2616] = layer4_out[3557];
    assign layer5_out[2617] = ~layer4_out[2382];
    assign layer5_out[2618] = ~(layer4_out[7734] ^ layer4_out[7735]);
    assign layer5_out[2619] = ~(layer4_out[5081] ^ layer4_out[5082]);
    assign layer5_out[2620] = ~(layer4_out[7208] | layer4_out[7209]);
    assign layer5_out[2621] = ~(layer4_out[278] | layer4_out[279]);
    assign layer5_out[2622] = ~layer4_out[3038];
    assign layer5_out[2623] = ~layer4_out[765];
    assign layer5_out[2624] = ~(layer4_out[4354] ^ layer4_out[4355]);
    assign layer5_out[2625] = layer4_out[4707] & layer4_out[4708];
    assign layer5_out[2626] = ~layer4_out[5821];
    assign layer5_out[2627] = layer4_out[5860] ^ layer4_out[5861];
    assign layer5_out[2628] = ~(layer4_out[1947] | layer4_out[1948]);
    assign layer5_out[2629] = layer4_out[1638];
    assign layer5_out[2630] = ~layer4_out[2295] | layer4_out[2296];
    assign layer5_out[2631] = layer4_out[3532] ^ layer4_out[3533];
    assign layer5_out[2632] = ~layer4_out[5240];
    assign layer5_out[2633] = ~layer4_out[7157];
    assign layer5_out[2634] = layer4_out[7770] & layer4_out[7771];
    assign layer5_out[2635] = ~(layer4_out[5963] ^ layer4_out[5964]);
    assign layer5_out[2636] = ~layer4_out[7857];
    assign layer5_out[2637] = layer4_out[6097] ^ layer4_out[6098];
    assign layer5_out[2638] = layer4_out[2699] & ~layer4_out[2700];
    assign layer5_out[2639] = ~layer4_out[3766];
    assign layer5_out[2640] = layer4_out[500] & layer4_out[501];
    assign layer5_out[2641] = ~(layer4_out[1754] ^ layer4_out[1755]);
    assign layer5_out[2642] = layer4_out[3980] ^ layer4_out[3981];
    assign layer5_out[2643] = layer4_out[31] & ~layer4_out[30];
    assign layer5_out[2644] = layer4_out[713] ^ layer4_out[714];
    assign layer5_out[2645] = ~layer4_out[3241] | layer4_out[3242];
    assign layer5_out[2646] = ~(layer4_out[6348] ^ layer4_out[6349]);
    assign layer5_out[2647] = layer4_out[6688];
    assign layer5_out[2648] = layer4_out[6476];
    assign layer5_out[2649] = layer4_out[1465];
    assign layer5_out[2650] = ~(layer4_out[5190] ^ layer4_out[5191]);
    assign layer5_out[2651] = ~layer4_out[7550];
    assign layer5_out[2652] = layer4_out[5061] & ~layer4_out[5062];
    assign layer5_out[2653] = ~(layer4_out[417] ^ layer4_out[418]);
    assign layer5_out[2654] = layer4_out[7417];
    assign layer5_out[2655] = layer4_out[3339] ^ layer4_out[3340];
    assign layer5_out[2656] = ~layer4_out[1759];
    assign layer5_out[2657] = layer4_out[4819];
    assign layer5_out[2658] = ~layer4_out[2367];
    assign layer5_out[2659] = layer4_out[2415];
    assign layer5_out[2660] = layer4_out[7124];
    assign layer5_out[2661] = ~(layer4_out[711] & layer4_out[712]);
    assign layer5_out[2662] = ~layer4_out[5595];
    assign layer5_out[2663] = layer4_out[2155] & ~layer4_out[2156];
    assign layer5_out[2664] = ~layer4_out[6819] | layer4_out[6818];
    assign layer5_out[2665] = layer4_out[4089];
    assign layer5_out[2666] = layer4_out[5813] & ~layer4_out[5814];
    assign layer5_out[2667] = layer4_out[2544] ^ layer4_out[2545];
    assign layer5_out[2668] = ~layer4_out[6330];
    assign layer5_out[2669] = layer4_out[7222] ^ layer4_out[7223];
    assign layer5_out[2670] = ~(layer4_out[5633] | layer4_out[5634]);
    assign layer5_out[2671] = ~layer4_out[784] | layer4_out[785];
    assign layer5_out[2672] = layer4_out[3305];
    assign layer5_out[2673] = layer4_out[18] ^ layer4_out[19];
    assign layer5_out[2674] = ~(layer4_out[4277] ^ layer4_out[4278]);
    assign layer5_out[2675] = ~layer4_out[7032];
    assign layer5_out[2676] = ~(layer4_out[7554] | layer4_out[7555]);
    assign layer5_out[2677] = layer4_out[5942];
    assign layer5_out[2678] = ~(layer4_out[3458] & layer4_out[3459]);
    assign layer5_out[2679] = ~(layer4_out[4726] & layer4_out[4727]);
    assign layer5_out[2680] = layer4_out[4000] & layer4_out[4001];
    assign layer5_out[2681] = layer4_out[1824];
    assign layer5_out[2682] = ~(layer4_out[6224] | layer4_out[6225]);
    assign layer5_out[2683] = layer4_out[5924] & ~layer4_out[5923];
    assign layer5_out[2684] = ~(layer4_out[5487] ^ layer4_out[5488]);
    assign layer5_out[2685] = ~(layer4_out[3077] ^ layer4_out[3078]);
    assign layer5_out[2686] = layer4_out[2908] ^ layer4_out[2909];
    assign layer5_out[2687] = ~layer4_out[3023] | layer4_out[3024];
    assign layer5_out[2688] = ~(layer4_out[2051] | layer4_out[2052]);
    assign layer5_out[2689] = ~layer4_out[524] | layer4_out[523];
    assign layer5_out[2690] = ~(layer4_out[1389] ^ layer4_out[1390]);
    assign layer5_out[2691] = layer4_out[862];
    assign layer5_out[2692] = ~(layer4_out[1364] | layer4_out[1365]);
    assign layer5_out[2693] = layer4_out[2914];
    assign layer5_out[2694] = ~layer4_out[4625];
    assign layer5_out[2695] = layer4_out[4799] & layer4_out[4800];
    assign layer5_out[2696] = ~layer4_out[1022];
    assign layer5_out[2697] = layer4_out[3683] & layer4_out[3684];
    assign layer5_out[2698] = layer4_out[5236] ^ layer4_out[5237];
    assign layer5_out[2699] = layer4_out[5792] | layer4_out[5793];
    assign layer5_out[2700] = ~layer4_out[5480];
    assign layer5_out[2701] = layer4_out[1550] ^ layer4_out[1551];
    assign layer5_out[2702] = ~(layer4_out[1000] | layer4_out[1001]);
    assign layer5_out[2703] = ~(layer4_out[165] | layer4_out[166]);
    assign layer5_out[2704] = layer4_out[138] & ~layer4_out[139];
    assign layer5_out[2705] = layer4_out[6901];
    assign layer5_out[2706] = layer4_out[2569] ^ layer4_out[2570];
    assign layer5_out[2707] = ~layer4_out[1095];
    assign layer5_out[2708] = layer4_out[1524];
    assign layer5_out[2709] = ~(layer4_out[5422] ^ layer4_out[5423]);
    assign layer5_out[2710] = ~(layer4_out[7136] ^ layer4_out[7137]);
    assign layer5_out[2711] = ~layer4_out[5580];
    assign layer5_out[2712] = ~layer4_out[3420] | layer4_out[3419];
    assign layer5_out[2713] = layer4_out[4684] & ~layer4_out[4683];
    assign layer5_out[2714] = layer4_out[2359];
    assign layer5_out[2715] = layer4_out[1678] | layer4_out[1679];
    assign layer5_out[2716] = layer4_out[5478];
    assign layer5_out[2717] = layer4_out[1659];
    assign layer5_out[2718] = layer4_out[7349] & layer4_out[7350];
    assign layer5_out[2719] = ~(layer4_out[2344] ^ layer4_out[2345]);
    assign layer5_out[2720] = ~layer4_out[4626] | layer4_out[4627];
    assign layer5_out[2721] = layer4_out[7576] ^ layer4_out[7577];
    assign layer5_out[2722] = ~layer4_out[4461];
    assign layer5_out[2723] = ~layer4_out[796];
    assign layer5_out[2724] = layer4_out[2434] & layer4_out[2435];
    assign layer5_out[2725] = ~(layer4_out[4281] ^ layer4_out[4282]);
    assign layer5_out[2726] = layer4_out[6];
    assign layer5_out[2727] = ~(layer4_out[5444] ^ layer4_out[5445]);
    assign layer5_out[2728] = ~layer4_out[6078];
    assign layer5_out[2729] = layer4_out[1642] ^ layer4_out[1643];
    assign layer5_out[2730] = layer4_out[4935] & ~layer4_out[4934];
    assign layer5_out[2731] = layer4_out[2265] & layer4_out[2266];
    assign layer5_out[2732] = ~layer4_out[3306];
    assign layer5_out[2733] = ~layer4_out[4342];
    assign layer5_out[2734] = ~layer4_out[4697];
    assign layer5_out[2735] = ~(layer4_out[7167] ^ layer4_out[7168]);
    assign layer5_out[2736] = layer4_out[103] & ~layer4_out[104];
    assign layer5_out[2737] = layer4_out[1287];
    assign layer5_out[2738] = layer4_out[4545] & layer4_out[4546];
    assign layer5_out[2739] = ~layer4_out[5771] | layer4_out[5772];
    assign layer5_out[2740] = layer4_out[7048];
    assign layer5_out[2741] = layer4_out[6861];
    assign layer5_out[2742] = layer4_out[3931];
    assign layer5_out[2743] = layer4_out[7464] & layer4_out[7465];
    assign layer5_out[2744] = layer4_out[7111];
    assign layer5_out[2745] = layer4_out[7707];
    assign layer5_out[2746] = ~layer4_out[5728];
    assign layer5_out[2747] = layer4_out[4136] ^ layer4_out[4137];
    assign layer5_out[2748] = layer4_out[5460];
    assign layer5_out[2749] = layer4_out[5787];
    assign layer5_out[2750] = layer4_out[156] ^ layer4_out[157];
    assign layer5_out[2751] = layer4_out[182] ^ layer4_out[183];
    assign layer5_out[2752] = layer4_out[3627] | layer4_out[3628];
    assign layer5_out[2753] = ~layer4_out[634] | layer4_out[635];
    assign layer5_out[2754] = ~layer4_out[2197];
    assign layer5_out[2755] = layer4_out[2946] ^ layer4_out[2947];
    assign layer5_out[2756] = layer4_out[6316];
    assign layer5_out[2757] = layer4_out[7630] ^ layer4_out[7631];
    assign layer5_out[2758] = layer4_out[6468] | layer4_out[6469];
    assign layer5_out[2759] = ~layer4_out[6641];
    assign layer5_out[2760] = layer4_out[3944];
    assign layer5_out[2761] = ~layer4_out[1402];
    assign layer5_out[2762] = layer4_out[5326] ^ layer4_out[5327];
    assign layer5_out[2763] = layer4_out[2892];
    assign layer5_out[2764] = layer4_out[3856];
    assign layer5_out[2765] = layer4_out[6964] ^ layer4_out[6965];
    assign layer5_out[2766] = layer4_out[5194] | layer4_out[5195];
    assign layer5_out[2767] = layer4_out[1442];
    assign layer5_out[2768] = layer4_out[7199] & ~layer4_out[7198];
    assign layer5_out[2769] = ~layer4_out[1490];
    assign layer5_out[2770] = layer4_out[1082];
    assign layer5_out[2771] = layer4_out[5372];
    assign layer5_out[2772] = layer4_out[3717] ^ layer4_out[3718];
    assign layer5_out[2773] = ~layer4_out[4038];
    assign layer5_out[2774] = ~layer4_out[356];
    assign layer5_out[2775] = ~(layer4_out[35] ^ layer4_out[36]);
    assign layer5_out[2776] = layer4_out[2093] ^ layer4_out[2094];
    assign layer5_out[2777] = layer4_out[6715] ^ layer4_out[6716];
    assign layer5_out[2778] = layer4_out[2734];
    assign layer5_out[2779] = layer4_out[230];
    assign layer5_out[2780] = layer4_out[4130] ^ layer4_out[4131];
    assign layer5_out[2781] = ~(layer4_out[3663] ^ layer4_out[3664]);
    assign layer5_out[2782] = ~(layer4_out[3494] ^ layer4_out[3495]);
    assign layer5_out[2783] = ~(layer4_out[5827] ^ layer4_out[5828]);
    assign layer5_out[2784] = ~(layer4_out[207] ^ layer4_out[208]);
    assign layer5_out[2785] = ~(layer4_out[2809] ^ layer4_out[2810]);
    assign layer5_out[2786] = layer4_out[5926] & ~layer4_out[5927];
    assign layer5_out[2787] = ~(layer4_out[7358] & layer4_out[7359]);
    assign layer5_out[2788] = ~(layer4_out[4434] | layer4_out[4435]);
    assign layer5_out[2789] = ~layer4_out[3361];
    assign layer5_out[2790] = layer4_out[6246] ^ layer4_out[6247];
    assign layer5_out[2791] = layer4_out[5719];
    assign layer5_out[2792] = layer4_out[2194] & layer4_out[2195];
    assign layer5_out[2793] = layer4_out[41] ^ layer4_out[42];
    assign layer5_out[2794] = layer4_out[7325] ^ layer4_out[7326];
    assign layer5_out[2795] = ~layer4_out[2147];
    assign layer5_out[2796] = ~layer4_out[7333];
    assign layer5_out[2797] = layer4_out[5287] & layer4_out[5288];
    assign layer5_out[2798] = layer4_out[2245] & ~layer4_out[2246];
    assign layer5_out[2799] = layer4_out[7746] ^ layer4_out[7747];
    assign layer5_out[2800] = ~layer4_out[5665];
    assign layer5_out[2801] = layer4_out[5928] ^ layer4_out[5929];
    assign layer5_out[2802] = layer4_out[3566] & ~layer4_out[3565];
    assign layer5_out[2803] = ~layer4_out[2966];
    assign layer5_out[2804] = layer4_out[7156];
    assign layer5_out[2805] = ~layer4_out[7846];
    assign layer5_out[2806] = ~(layer4_out[4004] ^ layer4_out[4005]);
    assign layer5_out[2807] = layer4_out[1804] ^ layer4_out[1805];
    assign layer5_out[2808] = ~layer4_out[5229];
    assign layer5_out[2809] = ~(layer4_out[469] ^ layer4_out[470]);
    assign layer5_out[2810] = layer4_out[7010] ^ layer4_out[7011];
    assign layer5_out[2811] = ~layer4_out[6256];
    assign layer5_out[2812] = ~(layer4_out[6683] | layer4_out[6684]);
    assign layer5_out[2813] = layer4_out[1893] & ~layer4_out[1892];
    assign layer5_out[2814] = layer4_out[4851] | layer4_out[4852];
    assign layer5_out[2815] = layer4_out[49] & ~layer4_out[48];
    assign layer5_out[2816] = layer4_out[7989] & layer4_out[7990];
    assign layer5_out[2817] = layer4_out[1972] & ~layer4_out[1973];
    assign layer5_out[2818] = ~layer4_out[4985];
    assign layer5_out[2819] = ~(layer4_out[5685] ^ layer4_out[5686]);
    assign layer5_out[2820] = ~layer4_out[1838];
    assign layer5_out[2821] = ~(layer4_out[7998] ^ layer4_out[7999]);
    assign layer5_out[2822] = layer4_out[2359] & ~layer4_out[2358];
    assign layer5_out[2823] = ~layer4_out[7487];
    assign layer5_out[2824] = layer4_out[248];
    assign layer5_out[2825] = layer4_out[5121] & layer4_out[5122];
    assign layer5_out[2826] = layer4_out[1887] & layer4_out[1888];
    assign layer5_out[2827] = ~layer4_out[5959];
    assign layer5_out[2828] = ~(layer4_out[1996] ^ layer4_out[1997]);
    assign layer5_out[2829] = layer4_out[244];
    assign layer5_out[2830] = ~(layer4_out[4296] & layer4_out[4297]);
    assign layer5_out[2831] = ~layer4_out[6132] | layer4_out[6131];
    assign layer5_out[2832] = ~(layer4_out[2590] ^ layer4_out[2591]);
    assign layer5_out[2833] = ~(layer4_out[3658] | layer4_out[3659]);
    assign layer5_out[2834] = layer4_out[2233];
    assign layer5_out[2835] = layer4_out[6320];
    assign layer5_out[2836] = ~(layer4_out[4589] | layer4_out[4590]);
    assign layer5_out[2837] = ~(layer4_out[3400] ^ layer4_out[3401]);
    assign layer5_out[2838] = ~layer4_out[3265];
    assign layer5_out[2839] = layer4_out[6550] & layer4_out[6551];
    assign layer5_out[2840] = ~layer4_out[6607];
    assign layer5_out[2841] = ~(layer4_out[1185] ^ layer4_out[1186]);
    assign layer5_out[2842] = layer4_out[4893];
    assign layer5_out[2843] = layer4_out[1925] & ~layer4_out[1924];
    assign layer5_out[2844] = layer4_out[5270];
    assign layer5_out[2845] = layer4_out[4780] ^ layer4_out[4781];
    assign layer5_out[2846] = layer4_out[6050] & layer4_out[6051];
    assign layer5_out[2847] = ~(layer4_out[1691] ^ layer4_out[1692]);
    assign layer5_out[2848] = ~layer4_out[4891];
    assign layer5_out[2849] = ~layer4_out[5302];
    assign layer5_out[2850] = ~layer4_out[5434] | layer4_out[5433];
    assign layer5_out[2851] = ~(layer4_out[4504] ^ layer4_out[4505]);
    assign layer5_out[2852] = ~layer4_out[6934];
    assign layer5_out[2853] = ~layer4_out[112];
    assign layer5_out[2854] = layer4_out[6190] & layer4_out[6191];
    assign layer5_out[2855] = ~layer4_out[1631];
    assign layer5_out[2856] = ~layer4_out[1806];
    assign layer5_out[2857] = layer4_out[680] ^ layer4_out[681];
    assign layer5_out[2858] = ~layer4_out[3308];
    assign layer5_out[2859] = ~layer4_out[651] | layer4_out[652];
    assign layer5_out[2860] = layer4_out[6203] | layer4_out[6204];
    assign layer5_out[2861] = ~layer4_out[6672] | layer4_out[6671];
    assign layer5_out[2862] = layer4_out[6611];
    assign layer5_out[2863] = ~layer4_out[6228];
    assign layer5_out[2864] = ~layer4_out[5756];
    assign layer5_out[2865] = layer4_out[2951] ^ layer4_out[2952];
    assign layer5_out[2866] = layer4_out[6543];
    assign layer5_out[2867] = ~layer4_out[3028];
    assign layer5_out[2868] = ~layer4_out[1048];
    assign layer5_out[2869] = ~(layer4_out[4016] ^ layer4_out[4017]);
    assign layer5_out[2870] = ~layer4_out[1728];
    assign layer5_out[2871] = layer4_out[1594] & ~layer4_out[1593];
    assign layer5_out[2872] = ~(layer4_out[6234] ^ layer4_out[6235]);
    assign layer5_out[2873] = ~(layer4_out[1629] ^ layer4_out[1630]);
    assign layer5_out[2874] = layer4_out[1439];
    assign layer5_out[2875] = layer4_out[600] & ~layer4_out[599];
    assign layer5_out[2876] = layer4_out[7343];
    assign layer5_out[2877] = ~layer4_out[7594];
    assign layer5_out[2878] = ~layer4_out[2481] | layer4_out[2482];
    assign layer5_out[2879] = layer4_out[4715] ^ layer4_out[4716];
    assign layer5_out[2880] = layer4_out[930] & ~layer4_out[929];
    assign layer5_out[2881] = layer4_out[2409];
    assign layer5_out[2882] = layer4_out[3412];
    assign layer5_out[2883] = layer4_out[4121] ^ layer4_out[4122];
    assign layer5_out[2884] = layer4_out[1800] ^ layer4_out[1801];
    assign layer5_out[2885] = ~layer4_out[7648];
    assign layer5_out[2886] = ~layer4_out[7228];
    assign layer5_out[2887] = layer4_out[1972];
    assign layer5_out[2888] = ~layer4_out[3611];
    assign layer5_out[2889] = ~(layer4_out[2033] ^ layer4_out[2034]);
    assign layer5_out[2890] = layer4_out[110];
    assign layer5_out[2891] = ~(layer4_out[494] ^ layer4_out[495]);
    assign layer5_out[2892] = ~layer4_out[2874];
    assign layer5_out[2893] = ~layer4_out[7278];
    assign layer5_out[2894] = layer4_out[5748] & ~layer4_out[5749];
    assign layer5_out[2895] = ~layer4_out[5069];
    assign layer5_out[2896] = ~layer4_out[3780] | layer4_out[3781];
    assign layer5_out[2897] = ~layer4_out[3639] | layer4_out[3640];
    assign layer5_out[2898] = ~layer4_out[1578] | layer4_out[1579];
    assign layer5_out[2899] = ~(layer4_out[4847] ^ layer4_out[4848]);
    assign layer5_out[2900] = ~layer4_out[6520];
    assign layer5_out[2901] = ~layer4_out[7824] | layer4_out[7825];
    assign layer5_out[2902] = ~layer4_out[7426] | layer4_out[7427];
    assign layer5_out[2903] = ~layer4_out[2058] | layer4_out[2059];
    assign layer5_out[2904] = ~layer4_out[4870] | layer4_out[4869];
    assign layer5_out[2905] = ~(layer4_out[1168] ^ layer4_out[1169]);
    assign layer5_out[2906] = layer4_out[5397];
    assign layer5_out[2907] = layer4_out[3771] & ~layer4_out[3770];
    assign layer5_out[2908] = ~(layer4_out[2804] | layer4_out[2805]);
    assign layer5_out[2909] = layer4_out[2716] & ~layer4_out[2717];
    assign layer5_out[2910] = layer4_out[171];
    assign layer5_out[2911] = layer4_out[4406];
    assign layer5_out[2912] = ~layer4_out[4087];
    assign layer5_out[2913] = layer4_out[7091];
    assign layer5_out[2914] = ~layer4_out[4720] | layer4_out[4721];
    assign layer5_out[2915] = ~(layer4_out[3009] ^ layer4_out[3010]);
    assign layer5_out[2916] = ~(layer4_out[7377] ^ layer4_out[7378]);
    assign layer5_out[2917] = layer4_out[777] & ~layer4_out[776];
    assign layer5_out[2918] = layer4_out[3860] | layer4_out[3861];
    assign layer5_out[2919] = ~layer4_out[2537];
    assign layer5_out[2920] = ~layer4_out[5462] | layer4_out[5461];
    assign layer5_out[2921] = layer4_out[3955];
    assign layer5_out[2922] = ~layer4_out[909];
    assign layer5_out[2923] = ~layer4_out[1740];
    assign layer5_out[2924] = ~layer4_out[6431];
    assign layer5_out[2925] = ~layer4_out[6933] | layer4_out[6932];
    assign layer5_out[2926] = ~layer4_out[6988];
    assign layer5_out[2927] = layer4_out[1584] & ~layer4_out[1583];
    assign layer5_out[2928] = ~layer4_out[4736];
    assign layer5_out[2929] = ~(layer4_out[3270] ^ layer4_out[3271]);
    assign layer5_out[2930] = layer4_out[1076];
    assign layer5_out[2931] = layer4_out[5255];
    assign layer5_out[2932] = ~(layer4_out[3979] ^ layer4_out[3980]);
    assign layer5_out[2933] = layer4_out[7463];
    assign layer5_out[2934] = layer4_out[496] & ~layer4_out[497];
    assign layer5_out[2935] = ~layer4_out[1873];
    assign layer5_out[2936] = layer4_out[7586] & layer4_out[7587];
    assign layer5_out[2937] = ~layer4_out[7399];
    assign layer5_out[2938] = ~layer4_out[2831] | layer4_out[2830];
    assign layer5_out[2939] = layer4_out[7845] & ~layer4_out[7844];
    assign layer5_out[2940] = ~layer4_out[2131] | layer4_out[2130];
    assign layer5_out[2941] = layer4_out[7943] & layer4_out[7944];
    assign layer5_out[2942] = layer4_out[5081];
    assign layer5_out[2943] = layer4_out[522] ^ layer4_out[523];
    assign layer5_out[2944] = ~layer4_out[4865];
    assign layer5_out[2945] = ~layer4_out[4392];
    assign layer5_out[2946] = layer4_out[3208];
    assign layer5_out[2947] = ~layer4_out[1504] | layer4_out[1505];
    assign layer5_out[2948] = ~layer4_out[2955];
    assign layer5_out[2949] = ~(layer4_out[4607] ^ layer4_out[4608]);
    assign layer5_out[2950] = layer4_out[4074] ^ layer4_out[4075];
    assign layer5_out[2951] = layer4_out[7058];
    assign layer5_out[2952] = layer4_out[6460] & ~layer4_out[6459];
    assign layer5_out[2953] = layer4_out[3114] & layer4_out[3115];
    assign layer5_out[2954] = layer4_out[5149] & ~layer4_out[5150];
    assign layer5_out[2955] = layer4_out[5424] ^ layer4_out[5425];
    assign layer5_out[2956] = layer4_out[7181];
    assign layer5_out[2957] = ~layer4_out[5618];
    assign layer5_out[2958] = ~layer4_out[7166];
    assign layer5_out[2959] = ~(layer4_out[293] | layer4_out[294]);
    assign layer5_out[2960] = ~(layer4_out[323] ^ layer4_out[324]);
    assign layer5_out[2961] = ~layer4_out[3846];
    assign layer5_out[2962] = ~layer4_out[3966];
    assign layer5_out[2963] = layer4_out[5680] ^ layer4_out[5681];
    assign layer5_out[2964] = layer4_out[5641] & ~layer4_out[5642];
    assign layer5_out[2965] = ~layer4_out[4019] | layer4_out[4020];
    assign layer5_out[2966] = ~layer4_out[6882];
    assign layer5_out[2967] = layer4_out[3889];
    assign layer5_out[2968] = layer4_out[7906] ^ layer4_out[7907];
    assign layer5_out[2969] = ~layer4_out[6478] | layer4_out[6477];
    assign layer5_out[2970] = ~(layer4_out[6032] | layer4_out[6033]);
    assign layer5_out[2971] = layer4_out[6573] ^ layer4_out[6574];
    assign layer5_out[2972] = ~layer4_out[3286] | layer4_out[3285];
    assign layer5_out[2973] = ~layer4_out[5302];
    assign layer5_out[2974] = ~layer4_out[1866];
    assign layer5_out[2975] = ~layer4_out[1832];
    assign layer5_out[2976] = layer4_out[5014] & ~layer4_out[5013];
    assign layer5_out[2977] = ~(layer4_out[4588] ^ layer4_out[4589]);
    assign layer5_out[2978] = ~layer4_out[6738];
    assign layer5_out[2979] = layer4_out[2315];
    assign layer5_out[2980] = ~layer4_out[2399];
    assign layer5_out[2981] = layer4_out[602];
    assign layer5_out[2982] = ~(layer4_out[7756] | layer4_out[7757]);
    assign layer5_out[2983] = ~(layer4_out[6112] ^ layer4_out[6113]);
    assign layer5_out[2984] = ~layer4_out[1276];
    assign layer5_out[2985] = layer4_out[4017] ^ layer4_out[4018];
    assign layer5_out[2986] = ~layer4_out[7538] | layer4_out[7537];
    assign layer5_out[2987] = ~(layer4_out[6903] | layer4_out[6904]);
    assign layer5_out[2988] = ~layer4_out[6347];
    assign layer5_out[2989] = ~(layer4_out[1581] ^ layer4_out[1582]);
    assign layer5_out[2990] = layer4_out[7713] & layer4_out[7714];
    assign layer5_out[2991] = layer4_out[7376] ^ layer4_out[7377];
    assign layer5_out[2992] = ~layer4_out[238];
    assign layer5_out[2993] = layer4_out[4332] ^ layer4_out[4333];
    assign layer5_out[2994] = ~layer4_out[7873];
    assign layer5_out[2995] = layer4_out[2396] & ~layer4_out[2395];
    assign layer5_out[2996] = ~layer4_out[5315] | layer4_out[5316];
    assign layer5_out[2997] = ~layer4_out[2727];
    assign layer5_out[2998] = layer4_out[719] ^ layer4_out[720];
    assign layer5_out[2999] = layer4_out[5178] & ~layer4_out[5179];
    assign layer5_out[3000] = layer4_out[6851] & ~layer4_out[6852];
    assign layer5_out[3001] = layer4_out[5421] ^ layer4_out[5422];
    assign layer5_out[3002] = layer4_out[5214] ^ layer4_out[5215];
    assign layer5_out[3003] = ~layer4_out[3390] | layer4_out[3391];
    assign layer5_out[3004] = ~(layer4_out[4536] & layer4_out[4537]);
    assign layer5_out[3005] = ~(layer4_out[3645] ^ layer4_out[3646]);
    assign layer5_out[3006] = ~layer4_out[5031];
    assign layer5_out[3007] = layer4_out[677] & layer4_out[678];
    assign layer5_out[3008] = layer4_out[2840] & ~layer4_out[2841];
    assign layer5_out[3009] = ~(layer4_out[1040] | layer4_out[1041]);
    assign layer5_out[3010] = layer4_out[7544];
    assign layer5_out[3011] = layer4_out[7525] ^ layer4_out[7526];
    assign layer5_out[3012] = layer4_out[7764] & ~layer4_out[7765];
    assign layer5_out[3013] = layer4_out[1799] & ~layer4_out[1798];
    assign layer5_out[3014] = ~(layer4_out[4944] | layer4_out[4945]);
    assign layer5_out[3015] = layer4_out[3052] ^ layer4_out[3053];
    assign layer5_out[3016] = layer4_out[3279] ^ layer4_out[3280];
    assign layer5_out[3017] = ~layer4_out[169];
    assign layer5_out[3018] = layer4_out[7760];
    assign layer5_out[3019] = layer4_out[2703] & ~layer4_out[2702];
    assign layer5_out[3020] = layer4_out[172];
    assign layer5_out[3021] = ~(layer4_out[4836] ^ layer4_out[4837]);
    assign layer5_out[3022] = layer4_out[2170] ^ layer4_out[2171];
    assign layer5_out[3023] = ~(layer4_out[1413] ^ layer4_out[1414]);
    assign layer5_out[3024] = layer4_out[7731];
    assign layer5_out[3025] = ~layer4_out[5482] | layer4_out[5481];
    assign layer5_out[3026] = ~(layer4_out[4593] ^ layer4_out[4594]);
    assign layer5_out[3027] = layer4_out[5723];
    assign layer5_out[3028] = layer4_out[1573] & layer4_out[1574];
    assign layer5_out[3029] = ~(layer4_out[5503] | layer4_out[5504]);
    assign layer5_out[3030] = layer4_out[2121];
    assign layer5_out[3031] = layer4_out[4501];
    assign layer5_out[3032] = layer4_out[2906] & ~layer4_out[2907];
    assign layer5_out[3033] = ~(layer4_out[3473] ^ layer4_out[3474]);
    assign layer5_out[3034] = layer4_out[6159];
    assign layer5_out[3035] = ~layer4_out[2382];
    assign layer5_out[3036] = layer4_out[5437];
    assign layer5_out[3037] = layer4_out[1995] & ~layer4_out[1996];
    assign layer5_out[3038] = ~layer4_out[5739];
    assign layer5_out[3039] = layer4_out[7590];
    assign layer5_out[3040] = ~(layer4_out[4534] ^ layer4_out[4535]);
    assign layer5_out[3041] = ~layer4_out[7224];
    assign layer5_out[3042] = ~layer4_out[4018];
    assign layer5_out[3043] = ~(layer4_out[2566] & layer4_out[2567]);
    assign layer5_out[3044] = layer4_out[6258];
    assign layer5_out[3045] = layer4_out[2286];
    assign layer5_out[3046] = ~layer4_out[1326] | layer4_out[1327];
    assign layer5_out[3047] = ~layer4_out[547];
    assign layer5_out[3048] = layer4_out[6589] & layer4_out[6590];
    assign layer5_out[3049] = ~(layer4_out[2347] & layer4_out[2348]);
    assign layer5_out[3050] = layer4_out[2878];
    assign layer5_out[3051] = layer4_out[931];
    assign layer5_out[3052] = layer4_out[5362] & ~layer4_out[5363];
    assign layer5_out[3053] = layer4_out[5681];
    assign layer5_out[3054] = layer4_out[2996] ^ layer4_out[2997];
    assign layer5_out[3055] = ~(layer4_out[1204] ^ layer4_out[1205]);
    assign layer5_out[3056] = layer4_out[933] & layer4_out[934];
    assign layer5_out[3057] = layer4_out[3940] & ~layer4_out[3939];
    assign layer5_out[3058] = ~(layer4_out[7235] ^ layer4_out[7236]);
    assign layer5_out[3059] = layer4_out[1432] ^ layer4_out[1433];
    assign layer5_out[3060] = layer4_out[4636] & layer4_out[4637];
    assign layer5_out[3061] = layer4_out[4729];
    assign layer5_out[3062] = layer4_out[1333] ^ layer4_out[1334];
    assign layer5_out[3063] = ~(layer4_out[3102] ^ layer4_out[3103]);
    assign layer5_out[3064] = ~(layer4_out[533] | layer4_out[534]);
    assign layer5_out[3065] = layer4_out[2463] ^ layer4_out[2464];
    assign layer5_out[3066] = layer4_out[2312] & layer4_out[2313];
    assign layer5_out[3067] = ~layer4_out[7565];
    assign layer5_out[3068] = layer4_out[6880];
    assign layer5_out[3069] = ~layer4_out[1991] | layer4_out[1990];
    assign layer5_out[3070] = ~layer4_out[2884];
    assign layer5_out[3071] = ~(layer4_out[7006] ^ layer4_out[7007]);
    assign layer5_out[3072] = layer4_out[4030] & ~layer4_out[4029];
    assign layer5_out[3073] = ~(layer4_out[1280] ^ layer4_out[1281]);
    assign layer5_out[3074] = ~layer4_out[7025];
    assign layer5_out[3075] = ~layer4_out[1278];
    assign layer5_out[3076] = ~(layer4_out[6597] | layer4_out[6598]);
    assign layer5_out[3077] = layer4_out[4647];
    assign layer5_out[3078] = layer4_out[6561] & ~layer4_out[6562];
    assign layer5_out[3079] = ~layer4_out[811];
    assign layer5_out[3080] = layer4_out[7702];
    assign layer5_out[3081] = layer4_out[552];
    assign layer5_out[3082] = ~layer4_out[6399];
    assign layer5_out[3083] = ~(layer4_out[1991] ^ layer4_out[1992]);
    assign layer5_out[3084] = layer4_out[6726] & layer4_out[6727];
    assign layer5_out[3085] = layer4_out[4752];
    assign layer5_out[3086] = layer4_out[6137] | layer4_out[6138];
    assign layer5_out[3087] = ~layer4_out[1954];
    assign layer5_out[3088] = ~(layer4_out[7066] ^ layer4_out[7067]);
    assign layer5_out[3089] = ~layer4_out[2211];
    assign layer5_out[3090] = ~(layer4_out[1701] ^ layer4_out[1702]);
    assign layer5_out[3091] = layer4_out[3094] & layer4_out[3095];
    assign layer5_out[3092] = layer4_out[4318] ^ layer4_out[4319];
    assign layer5_out[3093] = layer4_out[4901] | layer4_out[4902];
    assign layer5_out[3094] = ~layer4_out[5611];
    assign layer5_out[3095] = layer4_out[3180];
    assign layer5_out[3096] = ~layer4_out[7864];
    assign layer5_out[3097] = layer4_out[3034] & ~layer4_out[3033];
    assign layer5_out[3098] = layer4_out[728] & layer4_out[729];
    assign layer5_out[3099] = layer4_out[2426] | layer4_out[2427];
    assign layer5_out[3100] = layer4_out[2879] ^ layer4_out[2880];
    assign layer5_out[3101] = layer4_out[5495];
    assign layer5_out[3102] = ~(layer4_out[6504] | layer4_out[6505]);
    assign layer5_out[3103] = layer4_out[3824];
    assign layer5_out[3104] = ~(layer4_out[6908] | layer4_out[6909]);
    assign layer5_out[3105] = ~(layer4_out[5130] | layer4_out[5131]);
    assign layer5_out[3106] = ~(layer4_out[7982] | layer4_out[7983]);
    assign layer5_out[3107] = layer4_out[2924] ^ layer4_out[2925];
    assign layer5_out[3108] = ~layer4_out[3537];
    assign layer5_out[3109] = ~layer4_out[6812];
    assign layer5_out[3110] = ~(layer4_out[4805] ^ layer4_out[4806]);
    assign layer5_out[3111] = ~(layer4_out[7267] ^ layer4_out[7268]);
    assign layer5_out[3112] = layer4_out[4501];
    assign layer5_out[3113] = ~layer4_out[2559];
    assign layer5_out[3114] = ~layer4_out[6091];
    assign layer5_out[3115] = layer4_out[2074];
    assign layer5_out[3116] = ~layer4_out[3568] | layer4_out[3567];
    assign layer5_out[3117] = layer4_out[4635] | layer4_out[4636];
    assign layer5_out[3118] = ~layer4_out[6091];
    assign layer5_out[3119] = ~layer4_out[4841];
    assign layer5_out[3120] = ~(layer4_out[2136] | layer4_out[2137]);
    assign layer5_out[3121] = ~(layer4_out[1854] ^ layer4_out[1855]);
    assign layer5_out[3122] = ~layer4_out[5918];
    assign layer5_out[3123] = layer4_out[3274];
    assign layer5_out[3124] = layer4_out[3280] & ~layer4_out[3281];
    assign layer5_out[3125] = layer4_out[5144] ^ layer4_out[5145];
    assign layer5_out[3126] = layer4_out[6426] ^ layer4_out[6427];
    assign layer5_out[3127] = ~(layer4_out[3760] & layer4_out[3761]);
    assign layer5_out[3128] = layer4_out[7587] ^ layer4_out[7588];
    assign layer5_out[3129] = layer4_out[4750];
    assign layer5_out[3130] = layer4_out[2807] | layer4_out[2808];
    assign layer5_out[3131] = layer4_out[6152] | layer4_out[6153];
    assign layer5_out[3132] = layer4_out[4502];
    assign layer5_out[3133] = ~(layer4_out[7347] ^ layer4_out[7348]);
    assign layer5_out[3134] = ~(layer4_out[6084] ^ layer4_out[6085]);
    assign layer5_out[3135] = layer4_out[6773] ^ layer4_out[6774];
    assign layer5_out[3136] = ~(layer4_out[7187] | layer4_out[7188]);
    assign layer5_out[3137] = layer4_out[5389] & ~layer4_out[5390];
    assign layer5_out[3138] = layer4_out[7079] & ~layer4_out[7078];
    assign layer5_out[3139] = layer4_out[2663] ^ layer4_out[2664];
    assign layer5_out[3140] = layer4_out[2881] ^ layer4_out[2882];
    assign layer5_out[3141] = ~layer4_out[503];
    assign layer5_out[3142] = ~(layer4_out[3286] ^ layer4_out[3287]);
    assign layer5_out[3143] = ~layer4_out[423];
    assign layer5_out[3144] = layer4_out[7623] & ~layer4_out[7622];
    assign layer5_out[3145] = layer4_out[3248] ^ layer4_out[3249];
    assign layer5_out[3146] = ~layer4_out[6157];
    assign layer5_out[3147] = layer4_out[1063] & ~layer4_out[1062];
    assign layer5_out[3148] = ~layer4_out[5810];
    assign layer5_out[3149] = layer4_out[6178];
    assign layer5_out[3150] = ~layer4_out[5881];
    assign layer5_out[3151] = layer4_out[4255];
    assign layer5_out[3152] = ~layer4_out[888];
    assign layer5_out[3153] = layer4_out[1345];
    assign layer5_out[3154] = layer4_out[7197] & ~layer4_out[7198];
    assign layer5_out[3155] = layer4_out[7491];
    assign layer5_out[3156] = ~layer4_out[5106];
    assign layer5_out[3157] = ~layer4_out[6095];
    assign layer5_out[3158] = ~layer4_out[2498];
    assign layer5_out[3159] = layer4_out[2135] ^ layer4_out[2136];
    assign layer5_out[3160] = layer4_out[1826];
    assign layer5_out[3161] = layer4_out[2705];
    assign layer5_out[3162] = ~layer4_out[6576];
    assign layer5_out[3163] = ~layer4_out[4106];
    assign layer5_out[3164] = ~(layer4_out[6193] ^ layer4_out[6194]);
    assign layer5_out[3165] = layer4_out[1676] & ~layer4_out[1675];
    assign layer5_out[3166] = ~layer4_out[289];
    assign layer5_out[3167] = layer4_out[387] & layer4_out[388];
    assign layer5_out[3168] = layer4_out[2792] ^ layer4_out[2793];
    assign layer5_out[3169] = layer4_out[7974] & layer4_out[7975];
    assign layer5_out[3170] = layer4_out[5038];
    assign layer5_out[3171] = ~layer4_out[5978];
    assign layer5_out[3172] = layer4_out[14];
    assign layer5_out[3173] = layer4_out[1025];
    assign layer5_out[3174] = ~layer4_out[916];
    assign layer5_out[3175] = layer4_out[6841] | layer4_out[6842];
    assign layer5_out[3176] = layer4_out[5932] & layer4_out[5933];
    assign layer5_out[3177] = ~(layer4_out[2707] ^ layer4_out[2708]);
    assign layer5_out[3178] = ~layer4_out[2520] | layer4_out[2519];
    assign layer5_out[3179] = ~(layer4_out[5678] & layer4_out[5679]);
    assign layer5_out[3180] = layer4_out[4573] & ~layer4_out[4572];
    assign layer5_out[3181] = ~layer4_out[2523] | layer4_out[2522];
    assign layer5_out[3182] = layer4_out[1267];
    assign layer5_out[3183] = layer4_out[4664];
    assign layer5_out[3184] = layer4_out[5119] ^ layer4_out[5120];
    assign layer5_out[3185] = ~layer4_out[4998];
    assign layer5_out[3186] = ~layer4_out[344];
    assign layer5_out[3187] = layer4_out[724];
    assign layer5_out[3188] = ~(layer4_out[3478] ^ layer4_out[3479]);
    assign layer5_out[3189] = ~layer4_out[2520];
    assign layer5_out[3190] = layer4_out[2871];
    assign layer5_out[3191] = layer4_out[4610] | layer4_out[4611];
    assign layer5_out[3192] = ~layer4_out[7219] | layer4_out[7220];
    assign layer5_out[3193] = layer4_out[4584];
    assign layer5_out[3194] = layer4_out[4351];
    assign layer5_out[3195] = layer4_out[7432];
    assign layer5_out[3196] = ~layer4_out[7396];
    assign layer5_out[3197] = ~(layer4_out[7547] ^ layer4_out[7548]);
    assign layer5_out[3198] = ~layer4_out[6379];
    assign layer5_out[3199] = layer4_out[4069];
    assign layer5_out[3200] = layer4_out[4376] & ~layer4_out[4375];
    assign layer5_out[3201] = ~layer4_out[4951];
    assign layer5_out[3202] = layer4_out[4138];
    assign layer5_out[3203] = ~layer4_out[6363];
    assign layer5_out[3204] = ~layer4_out[1460];
    assign layer5_out[3205] = layer4_out[5528];
    assign layer5_out[3206] = ~(layer4_out[0] ^ layer4_out[1]);
    assign layer5_out[3207] = ~layer4_out[587];
    assign layer5_out[3208] = layer4_out[6631] & ~layer4_out[6632];
    assign layer5_out[3209] = layer4_out[6727] ^ layer4_out[6728];
    assign layer5_out[3210] = ~(layer4_out[7916] ^ layer4_out[7917]);
    assign layer5_out[3211] = ~(layer4_out[2919] | layer4_out[2920]);
    assign layer5_out[3212] = ~layer4_out[3502];
    assign layer5_out[3213] = layer4_out[4622] | layer4_out[4623];
    assign layer5_out[3214] = layer4_out[4949] ^ layer4_out[4950];
    assign layer5_out[3215] = ~layer4_out[4598] | layer4_out[4599];
    assign layer5_out[3216] = ~layer4_out[3990];
    assign layer5_out[3217] = ~(layer4_out[4083] ^ layer4_out[4084]);
    assign layer5_out[3218] = layer4_out[4827] & layer4_out[4828];
    assign layer5_out[3219] = layer4_out[6075] ^ layer4_out[6076];
    assign layer5_out[3220] = ~layer4_out[7739] | layer4_out[7740];
    assign layer5_out[3221] = layer4_out[2425] & ~layer4_out[2424];
    assign layer5_out[3222] = ~(layer4_out[1101] | layer4_out[1102]);
    assign layer5_out[3223] = ~layer4_out[5152];
    assign layer5_out[3224] = layer4_out[4173] ^ layer4_out[4174];
    assign layer5_out[3225] = layer4_out[1803] & ~layer4_out[1804];
    assign layer5_out[3226] = layer4_out[121] & layer4_out[122];
    assign layer5_out[3227] = layer4_out[2815] ^ layer4_out[2816];
    assign layer5_out[3228] = layer4_out[6576] & ~layer4_out[6577];
    assign layer5_out[3229] = ~(layer4_out[6256] ^ layer4_out[6257]);
    assign layer5_out[3230] = ~layer4_out[4400];
    assign layer5_out[3231] = layer4_out[4111] & ~layer4_out[4110];
    assign layer5_out[3232] = ~(layer4_out[6752] ^ layer4_out[6753]);
    assign layer5_out[3233] = layer4_out[2152];
    assign layer5_out[3234] = ~(layer4_out[205] | layer4_out[206]);
    assign layer5_out[3235] = ~layer4_out[2227] | layer4_out[2226];
    assign layer5_out[3236] = ~layer4_out[1576];
    assign layer5_out[3237] = layer4_out[7553];
    assign layer5_out[3238] = ~(layer4_out[1520] | layer4_out[1521]);
    assign layer5_out[3239] = layer4_out[450];
    assign layer5_out[3240] = layer4_out[3489];
    assign layer5_out[3241] = ~(layer4_out[3333] ^ layer4_out[3334]);
    assign layer5_out[3242] = ~(layer4_out[6434] ^ layer4_out[6435]);
    assign layer5_out[3243] = layer4_out[2656];
    assign layer5_out[3244] = layer4_out[5648];
    assign layer5_out[3245] = layer4_out[4612];
    assign layer5_out[3246] = layer4_out[4685];
    assign layer5_out[3247] = ~layer4_out[2886] | layer4_out[2885];
    assign layer5_out[3248] = ~(layer4_out[1357] | layer4_out[1358]);
    assign layer5_out[3249] = layer4_out[7977] & ~layer4_out[7976];
    assign layer5_out[3250] = layer4_out[6599] & ~layer4_out[6598];
    assign layer5_out[3251] = ~(layer4_out[2561] ^ layer4_out[2562]);
    assign layer5_out[3252] = layer4_out[4656];
    assign layer5_out[3253] = ~(layer4_out[4760] & layer4_out[4761]);
    assign layer5_out[3254] = layer4_out[1879] ^ layer4_out[1880];
    assign layer5_out[3255] = ~layer4_out[6053] | layer4_out[6052];
    assign layer5_out[3256] = layer4_out[152];
    assign layer5_out[3257] = ~(layer4_out[2843] ^ layer4_out[2844]);
    assign layer5_out[3258] = layer4_out[1847] & ~layer4_out[1846];
    assign layer5_out[3259] = layer4_out[3293] & ~layer4_out[3294];
    assign layer5_out[3260] = ~layer4_out[892];
    assign layer5_out[3261] = layer4_out[2143];
    assign layer5_out[3262] = layer4_out[2606] & layer4_out[2607];
    assign layer5_out[3263] = ~(layer4_out[365] ^ layer4_out[366]);
    assign layer5_out[3264] = layer4_out[1591] & ~layer4_out[1590];
    assign layer5_out[3265] = ~layer4_out[1771];
    assign layer5_out[3266] = ~layer4_out[7525];
    assign layer5_out[3267] = ~layer4_out[3205] | layer4_out[3204];
    assign layer5_out[3268] = layer4_out[3434] ^ layer4_out[3435];
    assign layer5_out[3269] = layer4_out[6270] & ~layer4_out[6271];
    assign layer5_out[3270] = ~layer4_out[7355];
    assign layer5_out[3271] = ~layer4_out[2105];
    assign layer5_out[3272] = layer4_out[6072] & layer4_out[6073];
    assign layer5_out[3273] = layer4_out[646] & layer4_out[647];
    assign layer5_out[3274] = ~layer4_out[4348];
    assign layer5_out[3275] = layer4_out[7313];
    assign layer5_out[3276] = layer4_out[5057] ^ layer4_out[5058];
    assign layer5_out[3277] = ~(layer4_out[1479] | layer4_out[1480]);
    assign layer5_out[3278] = ~layer4_out[328];
    assign layer5_out[3279] = ~(layer4_out[6744] ^ layer4_out[6745]);
    assign layer5_out[3280] = layer4_out[7605];
    assign layer5_out[3281] = ~layer4_out[3183];
    assign layer5_out[3282] = ~layer4_out[3080];
    assign layer5_out[3283] = layer4_out[2581] ^ layer4_out[2582];
    assign layer5_out[3284] = ~layer4_out[4990];
    assign layer5_out[3285] = layer4_out[2278] ^ layer4_out[2279];
    assign layer5_out[3286] = layer4_out[6157];
    assign layer5_out[3287] = ~layer4_out[2037];
    assign layer5_out[3288] = layer4_out[2092];
    assign layer5_out[3289] = layer4_out[1016];
    assign layer5_out[3290] = ~(layer4_out[6475] | layer4_out[6476]);
    assign layer5_out[3291] = layer4_out[5145] & layer4_out[5146];
    assign layer5_out[3292] = layer4_out[1141] ^ layer4_out[1142];
    assign layer5_out[3293] = layer4_out[4027] | layer4_out[4028];
    assign layer5_out[3294] = ~layer4_out[5189];
    assign layer5_out[3295] = ~layer4_out[7889];
    assign layer5_out[3296] = ~layer4_out[6788] | layer4_out[6787];
    assign layer5_out[3297] = layer4_out[1011] & ~layer4_out[1010];
    assign layer5_out[3298] = ~(layer4_out[4692] ^ layer4_out[4693]);
    assign layer5_out[3299] = ~layer4_out[6240] | layer4_out[6241];
    assign layer5_out[3300] = layer4_out[5084];
    assign layer5_out[3301] = ~(layer4_out[2725] ^ layer4_out[2726]);
    assign layer5_out[3302] = ~layer4_out[366];
    assign layer5_out[3303] = ~layer4_out[614];
    assign layer5_out[3304] = layer4_out[4423] | layer4_out[4424];
    assign layer5_out[3305] = ~layer4_out[2007];
    assign layer5_out[3306] = layer4_out[7650];
    assign layer5_out[3307] = ~(layer4_out[5476] | layer4_out[5477]);
    assign layer5_out[3308] = layer4_out[1872];
    assign layer5_out[3309] = layer4_out[5661] | layer4_out[5662];
    assign layer5_out[3310] = ~layer4_out[5164];
    assign layer5_out[3311] = layer4_out[2176] & ~layer4_out[2175];
    assign layer5_out[3312] = ~layer4_out[6333];
    assign layer5_out[3313] = layer4_out[6904] ^ layer4_out[6905];
    assign layer5_out[3314] = layer4_out[6723];
    assign layer5_out[3315] = layer4_out[4264];
    assign layer5_out[3316] = layer4_out[5915];
    assign layer5_out[3317] = layer4_out[3732];
    assign layer5_out[3318] = layer4_out[7009] | layer4_out[7010];
    assign layer5_out[3319] = layer4_out[7767];
    assign layer5_out[3320] = ~(layer4_out[4992] & layer4_out[4993]);
    assign layer5_out[3321] = layer4_out[7892];
    assign layer5_out[3322] = ~(layer4_out[2403] ^ layer4_out[2404]);
    assign layer5_out[3323] = ~(layer4_out[1715] ^ layer4_out[1716]);
    assign layer5_out[3324] = ~(layer4_out[5818] ^ layer4_out[5819]);
    assign layer5_out[3325] = layer4_out[3729];
    assign layer5_out[3326] = layer4_out[3200];
    assign layer5_out[3327] = layer4_out[6186] ^ layer4_out[6187];
    assign layer5_out[3328] = ~layer4_out[1723];
    assign layer5_out[3329] = ~layer4_out[2697];
    assign layer5_out[3330] = layer4_out[6023];
    assign layer5_out[3331] = layer4_out[2563] & layer4_out[2564];
    assign layer5_out[3332] = layer4_out[7857];
    assign layer5_out[3333] = layer4_out[2841];
    assign layer5_out[3334] = ~layer4_out[151];
    assign layer5_out[3335] = ~(layer4_out[1912] ^ layer4_out[1913]);
    assign layer5_out[3336] = layer4_out[5019] ^ layer4_out[5020];
    assign layer5_out[3337] = layer4_out[292] | layer4_out[293];
    assign layer5_out[3338] = layer4_out[5403] & layer4_out[5404];
    assign layer5_out[3339] = layer4_out[4357] & ~layer4_out[4358];
    assign layer5_out[3340] = layer4_out[501] ^ layer4_out[502];
    assign layer5_out[3341] = ~layer4_out[1163];
    assign layer5_out[3342] = ~layer4_out[5113] | layer4_out[5112];
    assign layer5_out[3343] = layer4_out[3872] ^ layer4_out[3873];
    assign layer5_out[3344] = layer4_out[3619] ^ layer4_out[3620];
    assign layer5_out[3345] = layer4_out[517];
    assign layer5_out[3346] = ~(layer4_out[6805] ^ layer4_out[6806]);
    assign layer5_out[3347] = ~(layer4_out[3855] & layer4_out[3856]);
    assign layer5_out[3348] = ~(layer4_out[4801] ^ layer4_out[4802]);
    assign layer5_out[3349] = ~layer4_out[4560];
    assign layer5_out[3350] = layer4_out[5060] ^ layer4_out[5061];
    assign layer5_out[3351] = layer4_out[7176] | layer4_out[7177];
    assign layer5_out[3352] = layer4_out[5378] & ~layer4_out[5377];
    assign layer5_out[3353] = ~layer4_out[605];
    assign layer5_out[3354] = layer4_out[5024] & layer4_out[5025];
    assign layer5_out[3355] = layer4_out[1263];
    assign layer5_out[3356] = ~layer4_out[2880] | layer4_out[2881];
    assign layer5_out[3357] = layer4_out[254];
    assign layer5_out[3358] = ~layer4_out[1066];
    assign layer5_out[3359] = layer4_out[7528];
    assign layer5_out[3360] = ~layer4_out[3323] | layer4_out[3322];
    assign layer5_out[3361] = ~(layer4_out[6175] ^ layer4_out[6176]);
    assign layer5_out[3362] = layer4_out[4372] ^ layer4_out[4373];
    assign layer5_out[3363] = ~layer4_out[3502];
    assign layer5_out[3364] = ~(layer4_out[4240] ^ layer4_out[4241]);
    assign layer5_out[3365] = ~layer4_out[5274];
    assign layer5_out[3366] = ~layer4_out[500] | layer4_out[499];
    assign layer5_out[3367] = ~layer4_out[6152];
    assign layer5_out[3368] = ~layer4_out[85] | layer4_out[86];
    assign layer5_out[3369] = layer4_out[7887];
    assign layer5_out[3370] = layer4_out[202] ^ layer4_out[203];
    assign layer5_out[3371] = layer4_out[7226] & ~layer4_out[7227];
    assign layer5_out[3372] = ~(layer4_out[6957] | layer4_out[6958]);
    assign layer5_out[3373] = ~(layer4_out[3269] ^ layer4_out[3270]);
    assign layer5_out[3374] = ~layer4_out[4455];
    assign layer5_out[3375] = ~(layer4_out[946] ^ layer4_out[947]);
    assign layer5_out[3376] = layer4_out[1908] ^ layer4_out[1909];
    assign layer5_out[3377] = layer4_out[2338] ^ layer4_out[2339];
    assign layer5_out[3378] = layer4_out[5387];
    assign layer5_out[3379] = layer4_out[7362];
    assign layer5_out[3380] = layer4_out[6855];
    assign layer5_out[3381] = layer4_out[782];
    assign layer5_out[3382] = layer4_out[1732];
    assign layer5_out[3383] = layer4_out[4434];
    assign layer5_out[3384] = ~layer4_out[4624] | layer4_out[4623];
    assign layer5_out[3385] = ~layer4_out[5272];
    assign layer5_out[3386] = ~(layer4_out[4049] ^ layer4_out[4050]);
    assign layer5_out[3387] = ~layer4_out[869];
    assign layer5_out[3388] = layer4_out[1270];
    assign layer5_out[3389] = layer4_out[647];
    assign layer5_out[3390] = layer4_out[6341];
    assign layer5_out[3391] = layer4_out[4725];
    assign layer5_out[3392] = ~layer4_out[6969];
    assign layer5_out[3393] = ~layer4_out[5383];
    assign layer5_out[3394] = layer4_out[6071] & layer4_out[6072];
    assign layer5_out[3395] = ~layer4_out[850];
    assign layer5_out[3396] = ~layer4_out[4704];
    assign layer5_out[3397] = ~layer4_out[1723];
    assign layer5_out[3398] = ~(layer4_out[3111] | layer4_out[3112]);
    assign layer5_out[3399] = layer4_out[7881] ^ layer4_out[7882];
    assign layer5_out[3400] = layer4_out[6302] ^ layer4_out[6303];
    assign layer5_out[3401] = layer4_out[988];
    assign layer5_out[3402] = ~(layer4_out[5542] ^ layer4_out[5543]);
    assign layer5_out[3403] = ~layer4_out[1608] | layer4_out[1607];
    assign layer5_out[3404] = ~layer4_out[3300];
    assign layer5_out[3405] = ~(layer4_out[3659] ^ layer4_out[3660]);
    assign layer5_out[3406] = ~(layer4_out[1147] | layer4_out[1148]);
    assign layer5_out[3407] = ~layer4_out[5981] | layer4_out[5980];
    assign layer5_out[3408] = ~layer4_out[3697];
    assign layer5_out[3409] = ~layer4_out[1848];
    assign layer5_out[3410] = ~(layer4_out[2960] & layer4_out[2961]);
    assign layer5_out[3411] = ~layer4_out[2936] | layer4_out[2935];
    assign layer5_out[3412] = ~(layer4_out[490] | layer4_out[491]);
    assign layer5_out[3413] = ~(layer4_out[1176] | layer4_out[1177]);
    assign layer5_out[3414] = layer4_out[5160] ^ layer4_out[5161];
    assign layer5_out[3415] = ~layer4_out[7608];
    assign layer5_out[3416] = ~layer4_out[750];
    assign layer5_out[3417] = layer4_out[1354] ^ layer4_out[1355];
    assign layer5_out[3418] = ~(layer4_out[3194] ^ layer4_out[3195]);
    assign layer5_out[3419] = layer4_out[5021];
    assign layer5_out[3420] = ~(layer4_out[1927] ^ layer4_out[1928]);
    assign layer5_out[3421] = ~layer4_out[6593];
    assign layer5_out[3422] = ~layer4_out[7214] | layer4_out[7215];
    assign layer5_out[3423] = layer4_out[537];
    assign layer5_out[3424] = ~layer4_out[5136];
    assign layer5_out[3425] = layer4_out[6114];
    assign layer5_out[3426] = ~(layer4_out[3103] ^ layer4_out[3104]);
    assign layer5_out[3427] = ~layer4_out[3785];
    assign layer5_out[3428] = ~layer4_out[4097];
    assign layer5_out[3429] = layer4_out[2386];
    assign layer5_out[3430] = ~layer4_out[6169] | layer4_out[6168];
    assign layer5_out[3431] = ~layer4_out[3886];
    assign layer5_out[3432] = layer4_out[6580] & ~layer4_out[6579];
    assign layer5_out[3433] = ~(layer4_out[1424] ^ layer4_out[1425]);
    assign layer5_out[3434] = ~layer4_out[1946];
    assign layer5_out[3435] = layer4_out[4549];
    assign layer5_out[3436] = ~layer4_out[4331];
    assign layer5_out[3437] = ~(layer4_out[1156] | layer4_out[1157]);
    assign layer5_out[3438] = ~layer4_out[1492];
    assign layer5_out[3439] = layer4_out[6103] ^ layer4_out[6104];
    assign layer5_out[3440] = ~(layer4_out[4713] | layer4_out[4714]);
    assign layer5_out[3441] = layer4_out[6266] & ~layer4_out[6267];
    assign layer5_out[3442] = ~(layer4_out[937] ^ layer4_out[938]);
    assign layer5_out[3443] = ~layer4_out[6866];
    assign layer5_out[3444] = layer4_out[2033];
    assign layer5_out[3445] = ~layer4_out[7879];
    assign layer5_out[3446] = ~layer4_out[3661];
    assign layer5_out[3447] = ~(layer4_out[2508] ^ layer4_out[2509]);
    assign layer5_out[3448] = layer4_out[4727] & ~layer4_out[4728];
    assign layer5_out[3449] = layer4_out[2468];
    assign layer5_out[3450] = ~layer4_out[2272] | layer4_out[2273];
    assign layer5_out[3451] = ~(layer4_out[214] & layer4_out[215]);
    assign layer5_out[3452] = ~layer4_out[6363];
    assign layer5_out[3453] = ~layer4_out[607];
    assign layer5_out[3454] = layer4_out[2933];
    assign layer5_out[3455] = ~layer4_out[1055];
    assign layer5_out[3456] = ~layer4_out[5304];
    assign layer5_out[3457] = ~(layer4_out[5938] | layer4_out[5939]);
    assign layer5_out[3458] = ~(layer4_out[5695] ^ layer4_out[5696]);
    assign layer5_out[3459] = layer4_out[2431];
    assign layer5_out[3460] = layer4_out[6778];
    assign layer5_out[3461] = ~(layer4_out[1206] ^ layer4_out[1207]);
    assign layer5_out[3462] = ~layer4_out[460];
    assign layer5_out[3463] = layer4_out[6790];
    assign layer5_out[3464] = layer4_out[7021];
    assign layer5_out[3465] = layer4_out[2973] ^ layer4_out[2974];
    assign layer5_out[3466] = layer4_out[5102];
    assign layer5_out[3467] = layer4_out[3499] | layer4_out[3500];
    assign layer5_out[3468] = ~layer4_out[5244];
    assign layer5_out[3469] = layer4_out[7969] ^ layer4_out[7970];
    assign layer5_out[3470] = layer4_out[904] | layer4_out[905];
    assign layer5_out[3471] = ~layer4_out[306];
    assign layer5_out[3472] = layer4_out[453];
    assign layer5_out[3473] = layer4_out[6272];
    assign layer5_out[3474] = layer4_out[1955] | layer4_out[1956];
    assign layer5_out[3475] = layer4_out[488] & layer4_out[489];
    assign layer5_out[3476] = ~layer4_out[7679];
    assign layer5_out[3477] = layer4_out[4300] ^ layer4_out[4301];
    assign layer5_out[3478] = ~(layer4_out[4735] ^ layer4_out[4736]);
    assign layer5_out[3479] = ~layer4_out[2878];
    assign layer5_out[3480] = layer4_out[6893];
    assign layer5_out[3481] = layer4_out[3078] & layer4_out[3079];
    assign layer5_out[3482] = ~layer4_out[2985];
    assign layer5_out[3483] = layer4_out[6925];
    assign layer5_out[3484] = layer4_out[7440];
    assign layer5_out[3485] = layer4_out[1123] & layer4_out[1124];
    assign layer5_out[3486] = ~layer4_out[5597];
    assign layer5_out[3487] = layer4_out[5359] ^ layer4_out[5360];
    assign layer5_out[3488] = ~(layer4_out[5791] ^ layer4_out[5792]);
    assign layer5_out[3489] = layer4_out[3376] & ~layer4_out[3377];
    assign layer5_out[3490] = ~layer4_out[6138];
    assign layer5_out[3491] = ~layer4_out[4614];
    assign layer5_out[3492] = layer4_out[5534];
    assign layer5_out[3493] = layer4_out[612] ^ layer4_out[613];
    assign layer5_out[3494] = layer4_out[3853];
    assign layer5_out[3495] = ~layer4_out[4512];
    assign layer5_out[3496] = layer4_out[2492] ^ layer4_out[2493];
    assign layer5_out[3497] = ~(layer4_out[6622] | layer4_out[6623]);
    assign layer5_out[3498] = ~(layer4_out[3582] ^ layer4_out[3583]);
    assign layer5_out[3499] = ~layer4_out[5750];
    assign layer5_out[3500] = layer4_out[6159] & ~layer4_out[6160];
    assign layer5_out[3501] = layer4_out[5659] ^ layer4_out[5660];
    assign layer5_out[3502] = layer4_out[225] ^ layer4_out[226];
    assign layer5_out[3503] = layer4_out[33] & ~layer4_out[32];
    assign layer5_out[3504] = ~layer4_out[5170];
    assign layer5_out[3505] = layer4_out[74] ^ layer4_out[75];
    assign layer5_out[3506] = ~(layer4_out[6873] ^ layer4_out[6874]);
    assign layer5_out[3507] = layer4_out[7390] & layer4_out[7391];
    assign layer5_out[3508] = ~layer4_out[2751];
    assign layer5_out[3509] = layer4_out[7542] ^ layer4_out[7543];
    assign layer5_out[3510] = ~(layer4_out[5773] & layer4_out[5774]);
    assign layer5_out[3511] = ~layer4_out[7321] | layer4_out[7322];
    assign layer5_out[3512] = ~(layer4_out[1684] ^ layer4_out[1685]);
    assign layer5_out[3513] = layer4_out[621] & layer4_out[622];
    assign layer5_out[3514] = ~layer4_out[7551];
    assign layer5_out[3515] = ~layer4_out[5656];
    assign layer5_out[3516] = layer4_out[7631] ^ layer4_out[7632];
    assign layer5_out[3517] = layer4_out[1284];
    assign layer5_out[3518] = ~layer4_out[2598];
    assign layer5_out[3519] = layer4_out[468];
    assign layer5_out[3520] = ~(layer4_out[6609] ^ layer4_out[6610]);
    assign layer5_out[3521] = ~(layer4_out[7160] ^ layer4_out[7161]);
    assign layer5_out[3522] = layer4_out[4629];
    assign layer5_out[3523] = layer4_out[2420];
    assign layer5_out[3524] = ~(layer4_out[7638] | layer4_out[7639]);
    assign layer5_out[3525] = ~layer4_out[6063] | layer4_out[6064];
    assign layer5_out[3526] = ~(layer4_out[2131] ^ layer4_out[2132]);
    assign layer5_out[3527] = layer4_out[7313];
    assign layer5_out[3528] = layer4_out[5311] ^ layer4_out[5312];
    assign layer5_out[3529] = layer4_out[876] & ~layer4_out[875];
    assign layer5_out[3530] = ~layer4_out[4460];
    assign layer5_out[3531] = ~(layer4_out[5432] | layer4_out[5433]);
    assign layer5_out[3532] = layer4_out[7745] & layer4_out[7746];
    assign layer5_out[3533] = layer4_out[4686] & layer4_out[4687];
    assign layer5_out[3534] = layer4_out[5551];
    assign layer5_out[3535] = ~layer4_out[2244] | layer4_out[2243];
    assign layer5_out[3536] = ~layer4_out[3205];
    assign layer5_out[3537] = ~layer4_out[7000];
    assign layer5_out[3538] = ~layer4_out[1957] | layer4_out[1956];
    assign layer5_out[3539] = layer4_out[7039];
    assign layer5_out[3540] = ~(layer4_out[4429] ^ layer4_out[4430]);
    assign layer5_out[3541] = layer4_out[3267];
    assign layer5_out[3542] = layer4_out[1712] ^ layer4_out[1713];
    assign layer5_out[3543] = layer4_out[4232];
    assign layer5_out[3544] = ~layer4_out[1510];
    assign layer5_out[3545] = ~layer4_out[992];
    assign layer5_out[3546] = ~layer4_out[6099] | layer4_out[6100];
    assign layer5_out[3547] = ~layer4_out[6404];
    assign layer5_out[3548] = layer4_out[3468] ^ layer4_out[3469];
    assign layer5_out[3549] = ~layer4_out[1749];
    assign layer5_out[3550] = ~layer4_out[3885];
    assign layer5_out[3551] = layer4_out[1159] & layer4_out[1160];
    assign layer5_out[3552] = ~layer4_out[869];
    assign layer5_out[3553] = ~layer4_out[3721] | layer4_out[3720];
    assign layer5_out[3554] = layer4_out[4134];
    assign layer5_out[3555] = ~layer4_out[5173];
    assign layer5_out[3556] = layer4_out[3609] ^ layer4_out[3610];
    assign layer5_out[3557] = layer4_out[4259] ^ layer4_out[4260];
    assign layer5_out[3558] = layer4_out[6130];
    assign layer5_out[3559] = ~(layer4_out[7315] | layer4_out[7316]);
    assign layer5_out[3560] = ~layer4_out[5075] | layer4_out[5074];
    assign layer5_out[3561] = ~layer4_out[2452] | layer4_out[2451];
    assign layer5_out[3562] = layer4_out[6046] ^ layer4_out[6047];
    assign layer5_out[3563] = layer4_out[2867] & ~layer4_out[2866];
    assign layer5_out[3564] = layer4_out[1486];
    assign layer5_out[3565] = layer4_out[6243] ^ layer4_out[6244];
    assign layer5_out[3566] = layer4_out[7458] ^ layer4_out[7459];
    assign layer5_out[3567] = layer4_out[5011] & ~layer4_out[5010];
    assign layer5_out[3568] = layer4_out[611] ^ layer4_out[612];
    assign layer5_out[3569] = ~layer4_out[4664] | layer4_out[4665];
    assign layer5_out[3570] = layer4_out[3050] ^ layer4_out[3051];
    assign layer5_out[3571] = ~(layer4_out[3143] | layer4_out[3144]);
    assign layer5_out[3572] = layer4_out[7669];
    assign layer5_out[3573] = ~(layer4_out[4153] | layer4_out[4154]);
    assign layer5_out[3574] = layer4_out[543];
    assign layer5_out[3575] = layer4_out[1210] & ~layer4_out[1211];
    assign layer5_out[3576] = layer4_out[53] & ~layer4_out[54];
    assign layer5_out[3577] = ~layer4_out[4990];
    assign layer5_out[3578] = ~layer4_out[1851];
    assign layer5_out[3579] = ~layer4_out[3551];
    assign layer5_out[3580] = layer4_out[4756] | layer4_out[4757];
    assign layer5_out[3581] = layer4_out[6511];
    assign layer5_out[3582] = layer4_out[1481] & ~layer4_out[1480];
    assign layer5_out[3583] = ~(layer4_out[441] ^ layer4_out[442]);
    assign layer5_out[3584] = layer4_out[7414];
    assign layer5_out[3585] = layer4_out[6093];
    assign layer5_out[3586] = layer4_out[7261];
    assign layer5_out[3587] = layer4_out[4302] ^ layer4_out[4303];
    assign layer5_out[3588] = ~layer4_out[87];
    assign layer5_out[3589] = ~(layer4_out[7303] ^ layer4_out[7304]);
    assign layer5_out[3590] = ~(layer4_out[5312] ^ layer4_out[5313]);
    assign layer5_out[3591] = layer4_out[6440];
    assign layer5_out[3592] = ~(layer4_out[7975] | layer4_out[7976]);
    assign layer5_out[3593] = layer4_out[2440] ^ layer4_out[2441];
    assign layer5_out[3594] = layer4_out[6885];
    assign layer5_out[3595] = ~layer4_out[959];
    assign layer5_out[3596] = ~layer4_out[4930];
    assign layer5_out[3597] = ~(layer4_out[2279] ^ layer4_out[2280]);
    assign layer5_out[3598] = layer4_out[3571] ^ layer4_out[3572];
    assign layer5_out[3599] = layer4_out[7443];
    assign layer5_out[3600] = ~(layer4_out[952] & layer4_out[953]);
    assign layer5_out[3601] = ~layer4_out[3066];
    assign layer5_out[3602] = layer4_out[1623] ^ layer4_out[1624];
    assign layer5_out[3603] = ~layer4_out[538];
    assign layer5_out[3604] = layer4_out[235];
    assign layer5_out[3605] = layer4_out[2069] ^ layer4_out[2070];
    assign layer5_out[3606] = layer4_out[1728];
    assign layer5_out[3607] = layer4_out[4757] | layer4_out[4758];
    assign layer5_out[3608] = ~layer4_out[5758];
    assign layer5_out[3609] = ~layer4_out[3992];
    assign layer5_out[3610] = layer4_out[2018] | layer4_out[2019];
    assign layer5_out[3611] = layer4_out[2062];
    assign layer5_out[3612] = layer4_out[5944] ^ layer4_out[5945];
    assign layer5_out[3613] = layer4_out[583] | layer4_out[584];
    assign layer5_out[3614] = ~(layer4_out[1200] ^ layer4_out[1201]);
    assign layer5_out[3615] = layer4_out[6373] & ~layer4_out[6374];
    assign layer5_out[3616] = layer4_out[7460];
    assign layer5_out[3617] = layer4_out[7861] & ~layer4_out[7860];
    assign layer5_out[3618] = ~(layer4_out[4703] | layer4_out[4704]);
    assign layer5_out[3619] = layer4_out[7481] & ~layer4_out[7480];
    assign layer5_out[3620] = ~layer4_out[3892];
    assign layer5_out[3621] = layer4_out[6111] ^ layer4_out[6112];
    assign layer5_out[3622] = ~(layer4_out[1716] ^ layer4_out[1717]);
    assign layer5_out[3623] = ~layer4_out[3585];
    assign layer5_out[3624] = layer4_out[3228] | layer4_out[3229];
    assign layer5_out[3625] = ~layer4_out[91];
    assign layer5_out[3626] = ~layer4_out[608];
    assign layer5_out[3627] = layer4_out[525] ^ layer4_out[526];
    assign layer5_out[3628] = layer4_out[5423] | layer4_out[5424];
    assign layer5_out[3629] = layer4_out[1416] & ~layer4_out[1417];
    assign layer5_out[3630] = layer4_out[5569] ^ layer4_out[5570];
    assign layer5_out[3631] = ~layer4_out[3057] | layer4_out[3056];
    assign layer5_out[3632] = layer4_out[7071] & ~layer4_out[7072];
    assign layer5_out[3633] = layer4_out[3850];
    assign layer5_out[3634] = layer4_out[395];
    assign layer5_out[3635] = layer4_out[4995] & ~layer4_out[4996];
    assign layer5_out[3636] = ~layer4_out[5237] | layer4_out[5238];
    assign layer5_out[3637] = ~layer4_out[3799];
    assign layer5_out[3638] = layer4_out[6326];
    assign layer5_out[3639] = layer4_out[6531];
    assign layer5_out[3640] = layer4_out[811];
    assign layer5_out[3641] = ~(layer4_out[1786] & layer4_out[1787]);
    assign layer5_out[3642] = layer4_out[3148];
    assign layer5_out[3643] = layer4_out[245];
    assign layer5_out[3644] = ~(layer4_out[4389] ^ layer4_out[4390]);
    assign layer5_out[3645] = layer4_out[4826] | layer4_out[4827];
    assign layer5_out[3646] = ~(layer4_out[361] & layer4_out[362]);
    assign layer5_out[3647] = ~layer4_out[3313];
    assign layer5_out[3648] = ~layer4_out[7703];
    assign layer5_out[3649] = layer4_out[5871] & ~layer4_out[5872];
    assign layer5_out[3650] = ~layer4_out[3427];
    assign layer5_out[3651] = layer4_out[7446] & layer4_out[7447];
    assign layer5_out[3652] = ~layer4_out[123] | layer4_out[122];
    assign layer5_out[3653] = ~layer4_out[3635];
    assign layer5_out[3654] = layer4_out[691];
    assign layer5_out[3655] = ~layer4_out[3553];
    assign layer5_out[3656] = ~(layer4_out[4559] & layer4_out[4560]);
    assign layer5_out[3657] = layer4_out[3291];
    assign layer5_out[3658] = ~layer4_out[4023];
    assign layer5_out[3659] = layer4_out[4175];
    assign layer5_out[3660] = layer4_out[1500];
    assign layer5_out[3661] = layer4_out[2109];
    assign layer5_out[3662] = layer4_out[2208] & ~layer4_out[2207];
    assign layer5_out[3663] = layer4_out[1454];
    assign layer5_out[3664] = ~(layer4_out[129] ^ layer4_out[130]);
    assign layer5_out[3665] = layer4_out[5192] | layer4_out[5193];
    assign layer5_out[3666] = layer4_out[926] & ~layer4_out[925];
    assign layer5_out[3667] = layer4_out[842];
    assign layer5_out[3668] = layer4_out[6584];
    assign layer5_out[3669] = layer4_out[1697] & ~layer4_out[1696];
    assign layer5_out[3670] = layer4_out[5953];
    assign layer5_out[3671] = ~layer4_out[1797] | layer4_out[1798];
    assign layer5_out[3672] = layer4_out[6682];
    assign layer5_out[3673] = layer4_out[2209] ^ layer4_out[2210];
    assign layer5_out[3674] = ~layer4_out[4630];
    assign layer5_out[3675] = layer4_out[5434] & layer4_out[5435];
    assign layer5_out[3676] = layer4_out[3107];
    assign layer5_out[3677] = layer4_out[6073];
    assign layer5_out[3678] = layer4_out[4241] ^ layer4_out[4242];
    assign layer5_out[3679] = ~layer4_out[6560];
    assign layer5_out[3680] = ~layer4_out[5183];
    assign layer5_out[3681] = ~(layer4_out[7177] ^ layer4_out[7178]);
    assign layer5_out[3682] = ~layer4_out[7430];
    assign layer5_out[3683] = layer4_out[1542] & ~layer4_out[1543];
    assign layer5_out[3684] = layer4_out[450];
    assign layer5_out[3685] = layer4_out[6377];
    assign layer5_out[3686] = layer4_out[3641];
    assign layer5_out[3687] = ~layer4_out[4559] | layer4_out[4558];
    assign layer5_out[3688] = ~layer4_out[4764];
    assign layer5_out[3689] = ~layer4_out[2134];
    assign layer5_out[3690] = ~layer4_out[850];
    assign layer5_out[3691] = ~layer4_out[1813];
    assign layer5_out[3692] = layer4_out[5492] ^ layer4_out[5493];
    assign layer5_out[3693] = layer4_out[4583];
    assign layer5_out[3694] = layer4_out[6352] & ~layer4_out[6353];
    assign layer5_out[3695] = ~layer4_out[3943];
    assign layer5_out[3696] = ~(layer4_out[6505] ^ layer4_out[6506]);
    assign layer5_out[3697] = ~(layer4_out[3330] & layer4_out[3331]);
    assign layer5_out[3698] = layer4_out[4385] ^ layer4_out[4386];
    assign layer5_out[3699] = layer4_out[7014] | layer4_out[7015];
    assign layer5_out[3700] = layer4_out[5911] | layer4_out[5912];
    assign layer5_out[3701] = ~layer4_out[5298];
    assign layer5_out[3702] = layer4_out[535] | layer4_out[536];
    assign layer5_out[3703] = ~(layer4_out[4879] ^ layer4_out[4880]);
    assign layer5_out[3704] = ~layer4_out[7853];
    assign layer5_out[3705] = ~layer4_out[959] | layer4_out[960];
    assign layer5_out[3706] = ~(layer4_out[5282] | layer4_out[5283]);
    assign layer5_out[3707] = ~layer4_out[3436];
    assign layer5_out[3708] = ~(layer4_out[698] ^ layer4_out[699]);
    assign layer5_out[3709] = layer4_out[7195];
    assign layer5_out[3710] = layer4_out[7565];
    assign layer5_out[3711] = layer4_out[906] & ~layer4_out[907];
    assign layer5_out[3712] = layer4_out[5225] ^ layer4_out[5226];
    assign layer5_out[3713] = layer4_out[1309] & layer4_out[1310];
    assign layer5_out[3714] = layer4_out[3871];
    assign layer5_out[3715] = ~(layer4_out[3654] & layer4_out[3655]);
    assign layer5_out[3716] = ~(layer4_out[934] & layer4_out[935]);
    assign layer5_out[3717] = ~(layer4_out[116] & layer4_out[117]);
    assign layer5_out[3718] = ~layer4_out[3406];
    assign layer5_out[3719] = ~layer4_out[7155];
    assign layer5_out[3720] = ~(layer4_out[3305] ^ layer4_out[3306]);
    assign layer5_out[3721] = layer4_out[95] ^ layer4_out[96];
    assign layer5_out[3722] = layer4_out[7104] & ~layer4_out[7105];
    assign layer5_out[3723] = layer4_out[5915] & layer4_out[5916];
    assign layer5_out[3724] = ~layer4_out[5558];
    assign layer5_out[3725] = ~(layer4_out[3837] ^ layer4_out[3838]);
    assign layer5_out[3726] = ~(layer4_out[587] & layer4_out[588]);
    assign layer5_out[3727] = ~layer4_out[3920];
    assign layer5_out[3728] = layer4_out[4524] | layer4_out[4525];
    assign layer5_out[3729] = ~layer4_out[1580];
    assign layer5_out[3730] = layer4_out[1817];
    assign layer5_out[3731] = ~layer4_out[4688];
    assign layer5_out[3732] = ~layer4_out[5095];
    assign layer5_out[3733] = ~(layer4_out[3686] ^ layer4_out[3687]);
    assign layer5_out[3734] = ~layer4_out[173];
    assign layer5_out[3735] = layer4_out[3924] & ~layer4_out[3925];
    assign layer5_out[3736] = layer4_out[2457] ^ layer4_out[2458];
    assign layer5_out[3737] = layer4_out[3470];
    assign layer5_out[3738] = layer4_out[2377] & ~layer4_out[2376];
    assign layer5_out[3739] = layer4_out[563] ^ layer4_out[564];
    assign layer5_out[3740] = ~layer4_out[6659];
    assign layer5_out[3741] = layer4_out[817];
    assign layer5_out[3742] = layer4_out[3700];
    assign layer5_out[3743] = layer4_out[6312];
    assign layer5_out[3744] = ~(layer4_out[437] | layer4_out[438]);
    assign layer5_out[3745] = ~(layer4_out[3672] ^ layer4_out[3673]);
    assign layer5_out[3746] = ~layer4_out[632];
    assign layer5_out[3747] = layer4_out[1149] ^ layer4_out[1150];
    assign layer5_out[3748] = layer4_out[3801] ^ layer4_out[3802];
    assign layer5_out[3749] = layer4_out[3316];
    assign layer5_out[3750] = ~(layer4_out[7329] & layer4_out[7330]);
    assign layer5_out[3751] = layer4_out[1232] & layer4_out[1233];
    assign layer5_out[3752] = ~layer4_out[1932];
    assign layer5_out[3753] = ~layer4_out[3949];
    assign layer5_out[3754] = layer4_out[6706] ^ layer4_out[6707];
    assign layer5_out[3755] = ~layer4_out[3015];
    assign layer5_out[3756] = ~layer4_out[3085];
    assign layer5_out[3757] = ~layer4_out[3524];
    assign layer5_out[3758] = ~(layer4_out[5000] | layer4_out[5001]);
    assign layer5_out[3759] = ~layer4_out[375];
    assign layer5_out[3760] = layer4_out[493];
    assign layer5_out[3761] = ~(layer4_out[4301] ^ layer4_out[4302]);
    assign layer5_out[3762] = layer4_out[3744];
    assign layer5_out[3763] = ~(layer4_out[5970] ^ layer4_out[5971]);
    assign layer5_out[3764] = layer4_out[4292] & ~layer4_out[4291];
    assign layer5_out[3765] = ~(layer4_out[6350] ^ layer4_out[6351]);
    assign layer5_out[3766] = ~(layer4_out[47] & layer4_out[48]);
    assign layer5_out[3767] = ~layer4_out[2127];
    assign layer5_out[3768] = ~(layer4_out[1496] ^ layer4_out[1497]);
    assign layer5_out[3769] = ~layer4_out[409];
    assign layer5_out[3770] = layer4_out[7923] & ~layer4_out[7924];
    assign layer5_out[3771] = ~(layer4_out[6279] & layer4_out[6280]);
    assign layer5_out[3772] = ~layer4_out[3319];
    assign layer5_out[3773] = ~layer4_out[6693];
    assign layer5_out[3774] = ~layer4_out[5826];
    assign layer5_out[3775] = layer4_out[5820];
    assign layer5_out[3776] = layer4_out[7953] & ~layer4_out[7952];
    assign layer5_out[3777] = layer4_out[1613] ^ layer4_out[1614];
    assign layer5_out[3778] = layer4_out[4679];
    assign layer5_out[3779] = ~layer4_out[3820];
    assign layer5_out[3780] = layer4_out[7133];
    assign layer5_out[3781] = layer4_out[7656] & ~layer4_out[7655];
    assign layer5_out[3782] = ~layer4_out[4825] | layer4_out[4826];
    assign layer5_out[3783] = layer4_out[1671] | layer4_out[1672];
    assign layer5_out[3784] = layer4_out[7397] | layer4_out[7398];
    assign layer5_out[3785] = layer4_out[5840] ^ layer4_out[5841];
    assign layer5_out[3786] = layer4_out[263] ^ layer4_out[264];
    assign layer5_out[3787] = ~layer4_out[3943];
    assign layer5_out[3788] = layer4_out[4066];
    assign layer5_out[3789] = ~layer4_out[306];
    assign layer5_out[3790] = layer4_out[592];
    assign layer5_out[3791] = ~(layer4_out[6745] ^ layer4_out[6746]);
    assign layer5_out[3792] = layer4_out[1500];
    assign layer5_out[3793] = layer4_out[3516];
    assign layer5_out[3794] = ~layer4_out[2812];
    assign layer5_out[3795] = layer4_out[2214] ^ layer4_out[2215];
    assign layer5_out[3796] = layer4_out[1270];
    assign layer5_out[3797] = layer4_out[736] | layer4_out[737];
    assign layer5_out[3798] = layer4_out[6008];
    assign layer5_out[3799] = layer4_out[7715] & ~layer4_out[7716];
    assign layer5_out[3800] = layer4_out[3141] & ~layer4_out[3140];
    assign layer5_out[3801] = layer4_out[3028];
    assign layer5_out[3802] = layer4_out[1790];
    assign layer5_out[3803] = layer4_out[7902];
    assign layer5_out[3804] = layer4_out[3674];
    assign layer5_out[3805] = layer4_out[2211] & ~layer4_out[2210];
    assign layer5_out[3806] = layer4_out[4631];
    assign layer5_out[3807] = layer4_out[6452] | layer4_out[6453];
    assign layer5_out[3808] = ~(layer4_out[5868] ^ layer4_out[5869]);
    assign layer5_out[3809] = layer4_out[5367];
    assign layer5_out[3810] = ~layer4_out[328];
    assign layer5_out[3811] = ~layer4_out[4326];
    assign layer5_out[3812] = ~(layer4_out[6793] ^ layer4_out[6794]);
    assign layer5_out[3813] = ~layer4_out[5804];
    assign layer5_out[3814] = layer4_out[5224];
    assign layer5_out[3815] = ~(layer4_out[2869] & layer4_out[2870]);
    assign layer5_out[3816] = layer4_out[359];
    assign layer5_out[3817] = layer4_out[567];
    assign layer5_out[3818] = ~layer4_out[6927];
    assign layer5_out[3819] = layer4_out[5157] & layer4_out[5158];
    assign layer5_out[3820] = ~layer4_out[550];
    assign layer5_out[3821] = layer4_out[4754];
    assign layer5_out[3822] = ~layer4_out[1039] | layer4_out[1040];
    assign layer5_out[3823] = layer4_out[6068] | layer4_out[6069];
    assign layer5_out[3824] = layer4_out[6008] & ~layer4_out[6009];
    assign layer5_out[3825] = ~(layer4_out[4725] ^ layer4_out[4726]);
    assign layer5_out[3826] = ~(layer4_out[7457] ^ layer4_out[7458]);
    assign layer5_out[3827] = layer4_out[6902] ^ layer4_out[6903];
    assign layer5_out[3828] = layer4_out[686];
    assign layer5_out[3829] = ~layer4_out[5629];
    assign layer5_out[3830] = layer4_out[1381] & ~layer4_out[1382];
    assign layer5_out[3831] = ~layer4_out[509];
    assign layer5_out[3832] = layer4_out[2573] ^ layer4_out[2574];
    assign layer5_out[3833] = layer4_out[4048];
    assign layer5_out[3834] = layer4_out[1253] | layer4_out[1254];
    assign layer5_out[3835] = ~layer4_out[7788] | layer4_out[7787];
    assign layer5_out[3836] = ~layer4_out[3300];
    assign layer5_out[3837] = layer4_out[7548] & layer4_out[7549];
    assign layer5_out[3838] = ~layer4_out[4496];
    assign layer5_out[3839] = ~(layer4_out[146] ^ layer4_out[147]);
    assign layer5_out[3840] = layer4_out[4042] & layer4_out[4043];
    assign layer5_out[3841] = ~layer4_out[4346];
    assign layer5_out[3842] = layer4_out[1609] ^ layer4_out[1610];
    assign layer5_out[3843] = layer4_out[1937] & ~layer4_out[1938];
    assign layer5_out[3844] = ~layer4_out[2998];
    assign layer5_out[3845] = layer4_out[5055] ^ layer4_out[5056];
    assign layer5_out[3846] = ~layer4_out[1893];
    assign layer5_out[3847] = ~(layer4_out[4994] ^ layer4_out[4995]);
    assign layer5_out[3848] = ~layer4_out[2430] | layer4_out[2431];
    assign layer5_out[3849] = ~layer4_out[3468];
    assign layer5_out[3850] = ~layer4_out[3074];
    assign layer5_out[3851] = ~layer4_out[550];
    assign layer5_out[3852] = ~layer4_out[7401];
    assign layer5_out[3853] = ~layer4_out[3189];
    assign layer5_out[3854] = ~layer4_out[3832] | layer4_out[3831];
    assign layer5_out[3855] = layer4_out[7097];
    assign layer5_out[3856] = ~(layer4_out[6969] | layer4_out[6970]);
    assign layer5_out[3857] = layer4_out[5746];
    assign layer5_out[3858] = ~(layer4_out[6760] ^ layer4_out[6761]);
    assign layer5_out[3859] = ~layer4_out[5483] | layer4_out[5482];
    assign layer5_out[3860] = ~layer4_out[3485];
    assign layer5_out[3861] = ~layer4_out[6279] | layer4_out[6278];
    assign layer5_out[3862] = layer4_out[1711] ^ layer4_out[1712];
    assign layer5_out[3863] = layer4_out[7820] & ~layer4_out[7819];
    assign layer5_out[3864] = layer4_out[7288] ^ layer4_out[7289];
    assign layer5_out[3865] = ~layer4_out[1585];
    assign layer5_out[3866] = layer4_out[3345];
    assign layer5_out[3867] = layer4_out[5414];
    assign layer5_out[3868] = layer4_out[3817] ^ layer4_out[3818];
    assign layer5_out[3869] = ~layer4_out[6214] | layer4_out[6215];
    assign layer5_out[3870] = layer4_out[5068];
    assign layer5_out[3871] = ~(layer4_out[752] ^ layer4_out[753]);
    assign layer5_out[3872] = layer4_out[2904];
    assign layer5_out[3873] = layer4_out[7147] ^ layer4_out[7148];
    assign layer5_out[3874] = layer4_out[7151];
    assign layer5_out[3875] = layer4_out[717] ^ layer4_out[718];
    assign layer5_out[3876] = layer4_out[2303] & ~layer4_out[2304];
    assign layer5_out[3877] = ~layer4_out[2689];
    assign layer5_out[3878] = ~layer4_out[68] | layer4_out[67];
    assign layer5_out[3879] = ~layer4_out[2304];
    assign layer5_out[3880] = layer4_out[3];
    assign layer5_out[3881] = layer4_out[6756] ^ layer4_out[6757];
    assign layer5_out[3882] = ~(layer4_out[5694] ^ layer4_out[5695]);
    assign layer5_out[3883] = ~layer4_out[5658];
    assign layer5_out[3884] = layer4_out[873] ^ layer4_out[874];
    assign layer5_out[3885] = layer4_out[2076] ^ layer4_out[2077];
    assign layer5_out[3886] = layer4_out[6570] ^ layer4_out[6571];
    assign layer5_out[3887] = ~(layer4_out[4040] ^ layer4_out[4041]);
    assign layer5_out[3888] = ~layer4_out[5043] | layer4_out[5044];
    assign layer5_out[3889] = ~(layer4_out[658] ^ layer4_out[659]);
    assign layer5_out[3890] = layer4_out[7460];
    assign layer5_out[3891] = layer4_out[5903];
    assign layer5_out[3892] = ~layer4_out[3313];
    assign layer5_out[3893] = layer4_out[4157];
    assign layer5_out[3894] = layer4_out[7953] & ~layer4_out[7954];
    assign layer5_out[3895] = ~(layer4_out[4880] ^ layer4_out[4881]);
    assign layer5_out[3896] = ~(layer4_out[1886] & layer4_out[1887]);
    assign layer5_out[3897] = layer4_out[3013];
    assign layer5_out[3898] = ~(layer4_out[5380] ^ layer4_out[5381]);
    assign layer5_out[3899] = ~(layer4_out[1652] & layer4_out[1653]);
    assign layer5_out[3900] = layer4_out[3311];
    assign layer5_out[3901] = ~layer4_out[5717];
    assign layer5_out[3902] = layer4_out[6037] ^ layer4_out[6038];
    assign layer5_out[3903] = layer4_out[5479];
    assign layer5_out[3904] = layer4_out[4576] & ~layer4_out[4575];
    assign layer5_out[3905] = layer4_out[5426];
    assign layer5_out[3906] = ~(layer4_out[3044] ^ layer4_out[3045]);
    assign layer5_out[3907] = layer4_out[3314] ^ layer4_out[3315];
    assign layer5_out[3908] = layer4_out[7205];
    assign layer5_out[3909] = ~(layer4_out[7469] ^ layer4_out[7470]);
    assign layer5_out[3910] = layer4_out[1463];
    assign layer5_out[3911] = layer4_out[1560];
    assign layer5_out[3912] = layer4_out[5714] | layer4_out[5715];
    assign layer5_out[3913] = ~layer4_out[2219];
    assign layer5_out[3914] = ~(layer4_out[1084] | layer4_out[1085]);
    assign layer5_out[3915] = ~(layer4_out[2784] & layer4_out[2785]);
    assign layer5_out[3916] = layer4_out[4781];
    assign layer5_out[3917] = layer4_out[3489];
    assign layer5_out[3918] = ~layer4_out[1121];
    assign layer5_out[3919] = ~(layer4_out[7885] & layer4_out[7886]);
    assign layer5_out[3920] = layer4_out[1221] ^ layer4_out[1222];
    assign layer5_out[3921] = ~layer4_out[4548];
    assign layer5_out[3922] = layer4_out[2015];
    assign layer5_out[3923] = ~layer4_out[6484];
    assign layer5_out[3924] = layer4_out[6537];
    assign layer5_out[3925] = layer4_out[863] & layer4_out[864];
    assign layer5_out[3926] = layer4_out[1560] ^ layer4_out[1561];
    assign layer5_out[3927] = layer4_out[7405];
    assign layer5_out[3928] = ~layer4_out[4216];
    assign layer5_out[3929] = layer4_out[6224];
    assign layer5_out[3930] = ~(layer4_out[7920] ^ layer4_out[7921]);
    assign layer5_out[3931] = ~(layer4_out[397] ^ layer4_out[398]);
    assign layer5_out[3932] = ~layer4_out[1218];
    assign layer5_out[3933] = layer4_out[4795] | layer4_out[4796];
    assign layer5_out[3934] = layer4_out[1355] ^ layer4_out[1356];
    assign layer5_out[3935] = layer4_out[7621] & layer4_out[7622];
    assign layer5_out[3936] = ~layer4_out[7385];
    assign layer5_out[3937] = ~layer4_out[6240];
    assign layer5_out[3938] = layer4_out[3700];
    assign layer5_out[3939] = ~(layer4_out[5471] & layer4_out[5472]);
    assign layer5_out[3940] = ~(layer4_out[3655] & layer4_out[3656]);
    assign layer5_out[3941] = layer4_out[5894];
    assign layer5_out[3942] = layer4_out[161] ^ layer4_out[162];
    assign layer5_out[3943] = layer4_out[3863];
    assign layer5_out[3944] = layer4_out[3750];
    assign layer5_out[3945] = layer4_out[5357] & layer4_out[5358];
    assign layer5_out[3946] = ~layer4_out[3834];
    assign layer5_out[3947] = ~layer4_out[2815];
    assign layer5_out[3948] = ~(layer4_out[330] | layer4_out[331]);
    assign layer5_out[3949] = layer4_out[4541] | layer4_out[4542];
    assign layer5_out[3950] = layer4_out[2541] & layer4_out[2542];
    assign layer5_out[3951] = ~layer4_out[6950];
    assign layer5_out[3952] = layer4_out[5022] | layer4_out[5023];
    assign layer5_out[3953] = ~layer4_out[3278];
    assign layer5_out[3954] = layer4_out[5083] & layer4_out[5084];
    assign layer5_out[3955] = layer4_out[2884];
    assign layer5_out[3956] = layer4_out[7122] ^ layer4_out[7123];
    assign layer5_out[3957] = layer4_out[7594] & layer4_out[7595];
    assign layer5_out[3958] = layer4_out[2356];
    assign layer5_out[3959] = ~layer4_out[4001] | layer4_out[4002];
    assign layer5_out[3960] = ~layer4_out[5505];
    assign layer5_out[3961] = ~layer4_out[1570];
    assign layer5_out[3962] = layer4_out[921] & ~layer4_out[922];
    assign layer5_out[3963] = layer4_out[6758] & ~layer4_out[6759];
    assign layer5_out[3964] = ~(layer4_out[2658] ^ layer4_out[2659]);
    assign layer5_out[3965] = layer4_out[3070];
    assign layer5_out[3966] = ~layer4_out[6920];
    assign layer5_out[3967] = ~layer4_out[3426];
    assign layer5_out[3968] = ~layer4_out[4103];
    assign layer5_out[3969] = layer4_out[1320] & ~layer4_out[1321];
    assign layer5_out[3970] = layer4_out[5412] ^ layer4_out[5413];
    assign layer5_out[3971] = ~layer4_out[5811];
    assign layer5_out[3972] = layer4_out[6844];
    assign layer5_out[3973] = layer4_out[5015];
    assign layer5_out[3974] = ~layer4_out[5418];
    assign layer5_out[3975] = layer4_out[1385];
    assign layer5_out[3976] = ~(layer4_out[1507] ^ layer4_out[1508]);
    assign layer5_out[3977] = layer4_out[4226];
    assign layer5_out[3978] = ~(layer4_out[6487] ^ layer4_out[6488]);
    assign layer5_out[3979] = layer4_out[1421] & layer4_out[1422];
    assign layer5_out[3980] = layer4_out[7146];
    assign layer5_out[3981] = layer4_out[5611] & ~layer4_out[5612];
    assign layer5_out[3982] = ~layer4_out[3172];
    assign layer5_out[3983] = layer4_out[6394] & ~layer4_out[6395];
    assign layer5_out[3984] = ~layer4_out[1208];
    assign layer5_out[3985] = layer4_out[3818] ^ layer4_out[3819];
    assign layer5_out[3986] = layer4_out[7173];
    assign layer5_out[3987] = ~layer4_out[7468];
    assign layer5_out[3988] = layer4_out[1272];
    assign layer5_out[3989] = layer4_out[6980];
    assign layer5_out[3990] = ~layer4_out[4512];
    assign layer5_out[3991] = layer4_out[6525] ^ layer4_out[6526];
    assign layer5_out[3992] = layer4_out[6162];
    assign layer5_out[3993] = ~(layer4_out[6795] | layer4_out[6796]);
    assign layer5_out[3994] = ~(layer4_out[5640] ^ layer4_out[5641]);
    assign layer5_out[3995] = layer4_out[4088];
    assign layer5_out[3996] = layer4_out[2966];
    assign layer5_out[3997] = layer4_out[6705];
    assign layer5_out[3998] = layer4_out[5628];
    assign layer5_out[3999] = layer4_out[2592];
    assign layer5_out[4000] = layer4_out[5772] ^ layer4_out[5773];
    assign layer5_out[4001] = layer4_out[3025];
    assign layer5_out[4002] = layer4_out[1529] & layer4_out[1530];
    assign layer5_out[4003] = layer4_out[1682];
    assign layer5_out[4004] = ~layer4_out[1484];
    assign layer5_out[4005] = layer4_out[3768] | layer4_out[3769];
    assign layer5_out[4006] = ~layer4_out[911];
    assign layer5_out[4007] = ~(layer4_out[1807] | layer4_out[1808]);
    assign layer5_out[4008] = ~layer4_out[3289];
    assign layer5_out[4009] = layer4_out[7151];
    assign layer5_out[4010] = layer4_out[6318] & ~layer4_out[6317];
    assign layer5_out[4011] = layer4_out[5517] & ~layer4_out[5518];
    assign layer5_out[4012] = ~layer4_out[1372];
    assign layer5_out[4013] = layer4_out[1501] ^ layer4_out[1502];
    assign layer5_out[4014] = ~layer4_out[2432] | layer4_out[2433];
    assign layer5_out[4015] = layer4_out[7504] & layer4_out[7505];
    assign layer5_out[4016] = ~(layer4_out[4330] ^ layer4_out[4331]);
    assign layer5_out[4017] = ~(layer4_out[4306] ^ layer4_out[4307]);
    assign layer5_out[4018] = ~layer4_out[6708];
    assign layer5_out[4019] = ~(layer4_out[7239] ^ layer4_out[7240]);
    assign layer5_out[4020] = ~layer4_out[5651];
    assign layer5_out[4021] = ~(layer4_out[6953] ^ layer4_out[6954]);
    assign layer5_out[4022] = ~layer4_out[3106];
    assign layer5_out[4023] = ~(layer4_out[6705] | layer4_out[6706]);
    assign layer5_out[4024] = layer4_out[7871];
    assign layer5_out[4025] = ~layer4_out[404];
    assign layer5_out[4026] = layer4_out[2947] & layer4_out[2948];
    assign layer5_out[4027] = ~layer4_out[638];
    assign layer5_out[4028] = ~layer4_out[1030];
    assign layer5_out[4029] = layer4_out[6590] & ~layer4_out[6591];
    assign layer5_out[4030] = ~layer4_out[2471] | layer4_out[2470];
    assign layer5_out[4031] = layer4_out[3676] & ~layer4_out[3677];
    assign layer5_out[4032] = layer4_out[7645] ^ layer4_out[7646];
    assign layer5_out[4033] = ~(layer4_out[6181] ^ layer4_out[6182]);
    assign layer5_out[4034] = ~(layer4_out[1676] ^ layer4_out[1677]);
    assign layer5_out[4035] = ~layer4_out[7443] | layer4_out[7442];
    assign layer5_out[4036] = layer4_out[1059];
    assign layer5_out[4037] = layer4_out[7287] & ~layer4_out[7288];
    assign layer5_out[4038] = layer4_out[673] & ~layer4_out[674];
    assign layer5_out[4039] = layer4_out[5163];
    assign layer5_out[4040] = layer4_out[2437];
    assign layer5_out[4041] = layer4_out[1746] & ~layer4_out[1745];
    assign layer5_out[4042] = layer4_out[185];
    assign layer5_out[4043] = layer4_out[44] & ~layer4_out[45];
    assign layer5_out[4044] = layer4_out[7792];
    assign layer5_out[4045] = layer4_out[4829] & ~layer4_out[4830];
    assign layer5_out[4046] = ~(layer4_out[5886] ^ layer4_out[5887]);
    assign layer5_out[4047] = layer4_out[2978] | layer4_out[2979];
    assign layer5_out[4048] = layer4_out[7045];
    assign layer5_out[4049] = layer4_out[5560];
    assign layer5_out[4050] = layer4_out[898] | layer4_out[899];
    assign layer5_out[4051] = ~layer4_out[7936];
    assign layer5_out[4052] = layer4_out[7319];
    assign layer5_out[4053] = ~(layer4_out[5962] ^ layer4_out[5963]);
    assign layer5_out[4054] = ~(layer4_out[4412] ^ layer4_out[4413]);
    assign layer5_out[4055] = ~layer4_out[5719];
    assign layer5_out[4056] = ~(layer4_out[7002] ^ layer4_out[7003]);
    assign layer5_out[4057] = ~(layer4_out[2290] ^ layer4_out[2291]);
    assign layer5_out[4058] = layer4_out[6526] ^ layer4_out[6527];
    assign layer5_out[4059] = layer4_out[6763] & layer4_out[6764];
    assign layer5_out[4060] = layer4_out[6586];
    assign layer5_out[4061] = ~layer4_out[2251] | layer4_out[2252];
    assign layer5_out[4062] = layer4_out[7829] & layer4_out[7830];
    assign layer5_out[4063] = ~layer4_out[620];
    assign layer5_out[4064] = layer4_out[7672];
    assign layer5_out[4065] = layer4_out[6956];
    assign layer5_out[4066] = ~layer4_out[6062] | layer4_out[6061];
    assign layer5_out[4067] = ~layer4_out[1299];
    assign layer5_out[4068] = ~layer4_out[3399] | layer4_out[3398];
    assign layer5_out[4069] = ~(layer4_out[6419] ^ layer4_out[6420]);
    assign layer5_out[4070] = layer4_out[4932];
    assign layer5_out[4071] = layer4_out[4669];
    assign layer5_out[4072] = ~(layer4_out[2406] ^ layer4_out[2407]);
    assign layer5_out[4073] = ~layer4_out[1590];
    assign layer5_out[4074] = ~(layer4_out[1547] ^ layer4_out[1548]);
    assign layer5_out[4075] = layer4_out[1245] ^ layer4_out[1246];
    assign layer5_out[4076] = ~layer4_out[7753] | layer4_out[7754];
    assign layer5_out[4077] = layer4_out[2718];
    assign layer5_out[4078] = layer4_out[7321];
    assign layer5_out[4079] = ~layer4_out[3126];
    assign layer5_out[4080] = layer4_out[597];
    assign layer5_out[4081] = layer4_out[2665] ^ layer4_out[2666];
    assign layer5_out[4082] = ~layer4_out[5265];
    assign layer5_out[4083] = layer4_out[2600] ^ layer4_out[2601];
    assign layer5_out[4084] = ~layer4_out[5450] | layer4_out[5451];
    assign layer5_out[4085] = ~(layer4_out[7623] & layer4_out[7624]);
    assign layer5_out[4086] = ~layer4_out[655] | layer4_out[656];
    assign layer5_out[4087] = layer4_out[6813] ^ layer4_out[6814];
    assign layer5_out[4088] = ~layer4_out[6082] | layer4_out[6083];
    assign layer5_out[4089] = ~layer4_out[1577] | layer4_out[1578];
    assign layer5_out[4090] = ~layer4_out[4466];
    assign layer5_out[4091] = ~layer4_out[3488];
    assign layer5_out[4092] = layer4_out[4948] & ~layer4_out[4947];
    assign layer5_out[4093] = layer4_out[435];
    assign layer5_out[4094] = ~(layer4_out[2637] & layer4_out[2638]);
    assign layer5_out[4095] = layer4_out[1072];
    assign layer5_out[4096] = layer4_out[7683] & ~layer4_out[7682];
    assign layer5_out[4097] = layer4_out[5185] ^ layer4_out[5186];
    assign layer5_out[4098] = layer4_out[2939] & layer4_out[2940];
    assign layer5_out[4099] = layer4_out[6771] & layer4_out[6772];
    assign layer5_out[4100] = layer4_out[1994] ^ layer4_out[1995];
    assign layer5_out[4101] = ~layer4_out[7868];
    assign layer5_out[4102] = layer4_out[7843] ^ layer4_out[7844];
    assign layer5_out[4103] = ~(layer4_out[5114] & layer4_out[5115]);
    assign layer5_out[4104] = ~(layer4_out[5696] & layer4_out[5697]);
    assign layer5_out[4105] = layer4_out[1603] & ~layer4_out[1604];
    assign layer5_out[4106] = layer4_out[2392] | layer4_out[2393];
    assign layer5_out[4107] = layer4_out[7917] ^ layer4_out[7918];
    assign layer5_out[4108] = layer4_out[5751] & ~layer4_out[5752];
    assign layer5_out[4109] = layer4_out[6134] ^ layer4_out[6135];
    assign layer5_out[4110] = layer4_out[4426];
    assign layer5_out[4111] = layer4_out[1182];
    assign layer5_out[4112] = ~layer4_out[2141];
    assign layer5_out[4113] = ~(layer4_out[7207] ^ layer4_out[7208]);
    assign layer5_out[4114] = layer4_out[879] ^ layer4_out[880];
    assign layer5_out[4115] = ~layer4_out[6690];
    assign layer5_out[4116] = layer4_out[3424] & ~layer4_out[3425];
    assign layer5_out[4117] = ~layer4_out[3772];
    assign layer5_out[4118] = ~layer4_out[6309];
    assign layer5_out[4119] = layer4_out[3046];
    assign layer5_out[4120] = layer4_out[6273] & ~layer4_out[6274];
    assign layer5_out[4121] = layer4_out[7004] ^ layer4_out[7005];
    assign layer5_out[4122] = ~(layer4_out[769] | layer4_out[770]);
    assign layer5_out[4123] = layer4_out[4927] & ~layer4_out[4928];
    assign layer5_out[4124] = ~layer4_out[6872];
    assign layer5_out[4125] = layer4_out[1696];
    assign layer5_out[4126] = layer4_out[7352] & ~layer4_out[7351];
    assign layer5_out[4127] = ~layer4_out[3068];
    assign layer5_out[4128] = layer4_out[3395];
    assign layer5_out[4129] = ~(layer4_out[3302] & layer4_out[3303]);
    assign layer5_out[4130] = layer4_out[7141] | layer4_out[7142];
    assign layer5_out[4131] = ~layer4_out[2982] | layer4_out[2981];
    assign layer5_out[4132] = layer4_out[1782];
    assign layer5_out[4133] = ~layer4_out[1007];
    assign layer5_out[4134] = layer4_out[7107];
    assign layer5_out[4135] = ~(layer4_out[6030] ^ layer4_out[6031]);
    assign layer5_out[4136] = layer4_out[7424] & layer4_out[7425];
    assign layer5_out[4137] = layer4_out[6166] ^ layer4_out[6167];
    assign layer5_out[4138] = ~layer4_out[4616];
    assign layer5_out[4139] = layer4_out[2802] & ~layer4_out[2801];
    assign layer5_out[4140] = ~(layer4_out[2277] ^ layer4_out[2278]);
    assign layer5_out[4141] = layer4_out[3947];
    assign layer5_out[4142] = ~(layer4_out[3706] ^ layer4_out[3707]);
    assign layer5_out[4143] = layer4_out[4280];
    assign layer5_out[4144] = ~layer4_out[2372];
    assign layer5_out[4145] = ~layer4_out[4674];
    assign layer5_out[4146] = ~layer4_out[2858] | layer4_out[2859];
    assign layer5_out[4147] = ~(layer4_out[953] ^ layer4_out[954]);
    assign layer5_out[4148] = layer4_out[2825] & ~layer4_out[2824];
    assign layer5_out[4149] = layer4_out[1645] & ~layer4_out[1646];
    assign layer5_out[4150] = layer4_out[169];
    assign layer5_out[4151] = layer4_out[2739] & ~layer4_out[2740];
    assign layer5_out[4152] = layer4_out[93] & ~layer4_out[92];
    assign layer5_out[4153] = ~(layer4_out[1653] | layer4_out[1654]);
    assign layer5_out[4154] = ~(layer4_out[213] ^ layer4_out[214]);
    assign layer5_out[4155] = ~(layer4_out[544] | layer4_out[545]);
    assign layer5_out[4156] = layer4_out[1562];
    assign layer5_out[4157] = layer4_out[3186] & ~layer4_out[3185];
    assign layer5_out[4158] = layer4_out[3762];
    assign layer5_out[4159] = layer4_out[5947];
    assign layer5_out[4160] = ~layer4_out[2535];
    assign layer5_out[4161] = ~layer4_out[6441];
    assign layer5_out[4162] = layer4_out[4194] & ~layer4_out[4195];
    assign layer5_out[4163] = ~layer4_out[6128];
    assign layer5_out[4164] = layer4_out[1426] & layer4_out[1427];
    assign layer5_out[4165] = ~(layer4_out[1513] ^ layer4_out[1514]);
    assign layer5_out[4166] = ~layer4_out[2732];
    assign layer5_out[4167] = layer4_out[113];
    assign layer5_out[4168] = ~layer4_out[813];
    assign layer5_out[4169] = layer4_out[7113] ^ layer4_out[7114];
    assign layer5_out[4170] = layer4_out[3350] & layer4_out[3351];
    assign layer5_out[4171] = ~layer4_out[4295];
    assign layer5_out[4172] = layer4_out[533];
    assign layer5_out[4173] = ~layer4_out[4514];
    assign layer5_out[4174] = layer4_out[6580] ^ layer4_out[6581];
    assign layer5_out[4175] = ~(layer4_out[7007] & layer4_out[7008]);
    assign layer5_out[4176] = layer4_out[4640];
    assign layer5_out[4177] = ~layer4_out[7557];
    assign layer5_out[4178] = layer4_out[2514] & ~layer4_out[2515];
    assign layer5_out[4179] = layer4_out[919] ^ layer4_out[920];
    assign layer5_out[4180] = ~layer4_out[1986];
    assign layer5_out[4181] = ~(layer4_out[5295] ^ layer4_out[5296]);
    assign layer5_out[4182] = layer4_out[2404] ^ layer4_out[2405];
    assign layer5_out[4183] = layer4_out[1819];
    assign layer5_out[4184] = layer4_out[2671] & layer4_out[2672];
    assign layer5_out[4185] = layer4_out[5101];
    assign layer5_out[4186] = layer4_out[3235];
    assign layer5_out[4187] = layer4_out[1783];
    assign layer5_out[4188] = layer4_out[3336] & ~layer4_out[3335];
    assign layer5_out[4189] = ~(layer4_out[5519] ^ layer4_out[5520]);
    assign layer5_out[4190] = ~layer4_out[5063];
    assign layer5_out[4191] = layer4_out[4014] & layer4_out[4015];
    assign layer5_out[4192] = layer4_out[418];
    assign layer5_out[4193] = ~(layer4_out[3643] ^ layer4_out[3644]);
    assign layer5_out[4194] = layer4_out[3404] & ~layer4_out[3403];
    assign layer5_out[4195] = ~(layer4_out[6422] ^ layer4_out[6423]);
    assign layer5_out[4196] = layer4_out[2316] ^ layer4_out[2317];
    assign layer5_out[4197] = layer4_out[7637];
    assign layer5_out[4198] = ~(layer4_out[6067] ^ layer4_out[6068]);
    assign layer5_out[4199] = layer4_out[440] ^ layer4_out[441];
    assign layer5_out[4200] = layer4_out[3685];
    assign layer5_out[4201] = ~layer4_out[3798];
    assign layer5_out[4202] = layer4_out[3957] & ~layer4_out[3958];
    assign layer5_out[4203] = layer4_out[2168];
    assign layer5_out[4204] = ~(layer4_out[7897] & layer4_out[7898]);
    assign layer5_out[4205] = ~layer4_out[2078];
    assign layer5_out[4206] = layer4_out[4059];
    assign layer5_out[4207] = ~(layer4_out[4835] | layer4_out[4836]);
    assign layer5_out[4208] = ~layer4_out[1748];
    assign layer5_out[4209] = ~(layer4_out[4594] | layer4_out[4595]);
    assign layer5_out[4210] = layer4_out[7590] & ~layer4_out[7591];
    assign layer5_out[4211] = layer4_out[7115];
    assign layer5_out[4212] = ~(layer4_out[2750] ^ layer4_out[2751]);
    assign layer5_out[4213] = ~(layer4_out[6262] & layer4_out[6263]);
    assign layer5_out[4214] = layer4_out[5670] ^ layer4_out[5671];
    assign layer5_out[4215] = layer4_out[3835] | layer4_out[3836];
    assign layer5_out[4216] = layer4_out[4247];
    assign layer5_out[4217] = layer4_out[1193] & layer4_out[1194];
    assign layer5_out[4218] = ~layer4_out[7366];
    assign layer5_out[4219] = layer4_out[5346] & ~layer4_out[5347];
    assign layer5_out[4220] = layer4_out[6049];
    assign layer5_out[4221] = layer4_out[2027] & layer4_out[2028];
    assign layer5_out[4222] = layer4_out[3191];
    assign layer5_out[4223] = ~(layer4_out[2183] ^ layer4_out[2184]);
    assign layer5_out[4224] = layer4_out[135];
    assign layer5_out[4225] = layer4_out[2677] | layer4_out[2678];
    assign layer5_out[4226] = ~layer4_out[4604];
    assign layer5_out[4227] = layer4_out[588];
    assign layer5_out[4228] = ~layer4_out[2539];
    assign layer5_out[4229] = ~(layer4_out[4115] | layer4_out[4116]);
    assign layer5_out[4230] = ~layer4_out[3237];
    assign layer5_out[4231] = layer4_out[307] & ~layer4_out[308];
    assign layer5_out[4232] = ~(layer4_out[2386] ^ layer4_out[2387]);
    assign layer5_out[4233] = ~layer4_out[1345] | layer4_out[1344];
    assign layer5_out[4234] = ~layer4_out[4685];
    assign layer5_out[4235] = layer4_out[7435];
    assign layer5_out[4236] = layer4_out[6833] ^ layer4_out[6834];
    assign layer5_out[4237] = layer4_out[5556] & ~layer4_out[5555];
    assign layer5_out[4238] = ~layer4_out[2759];
    assign layer5_out[4239] = ~layer4_out[3646];
    assign layer5_out[4240] = ~layer4_out[483];
    assign layer5_out[4241] = ~(layer4_out[5857] ^ layer4_out[5858]);
    assign layer5_out[4242] = ~layer4_out[74];
    assign layer5_out[4243] = ~layer4_out[4405];
    assign layer5_out[4244] = ~layer4_out[731];
    assign layer5_out[4245] = layer4_out[2230] | layer4_out[2231];
    assign layer5_out[4246] = ~layer4_out[1103];
    assign layer5_out[4247] = layer4_out[2187];
    assign layer5_out[4248] = layer4_out[1257];
    assign layer5_out[4249] = layer4_out[1895];
    assign layer5_out[4250] = ~layer4_out[432];
    assign layer5_out[4251] = layer4_out[7722] | layer4_out[7723];
    assign layer5_out[4252] = layer4_out[462] & ~layer4_out[463];
    assign layer5_out[4253] = layer4_out[7491] ^ layer4_out[7492];
    assign layer5_out[4254] = layer4_out[4507];
    assign layer5_out[4255] = layer4_out[6095];
    assign layer5_out[4256] = layer4_out[6815] | layer4_out[6816];
    assign layer5_out[4257] = layer4_out[7724] ^ layer4_out[7725];
    assign layer5_out[4258] = layer4_out[2055] & layer4_out[2056];
    assign layer5_out[4259] = ~layer4_out[6371] | layer4_out[6370];
    assign layer5_out[4260] = layer4_out[4224] & layer4_out[4225];
    assign layer5_out[4261] = layer4_out[1098] ^ layer4_out[1099];
    assign layer5_out[4262] = ~(layer4_out[3150] ^ layer4_out[3151]);
    assign layer5_out[4263] = layer4_out[4892];
    assign layer5_out[4264] = ~layer4_out[6847];
    assign layer5_out[4265] = layer4_out[6304];
    assign layer5_out[4266] = ~layer4_out[6840];
    assign layer5_out[4267] = ~(layer4_out[6735] ^ layer4_out[6736]);
    assign layer5_out[4268] = ~(layer4_out[2296] | layer4_out[2297]);
    assign layer5_out[4269] = ~(layer4_out[755] ^ layer4_out[756]);
    assign layer5_out[4270] = layer4_out[4520] | layer4_out[4521];
    assign layer5_out[4271] = ~(layer4_out[967] | layer4_out[968]);
    assign layer5_out[4272] = layer4_out[5672] & ~layer4_out[5671];
    assign layer5_out[4273] = layer4_out[2061] & ~layer4_out[2060];
    assign layer5_out[4274] = layer4_out[3577] & ~layer4_out[3578];
    assign layer5_out[4275] = layer4_out[5045];
    assign layer5_out[4276] = layer4_out[7582] & ~layer4_out[7583];
    assign layer5_out[4277] = ~(layer4_out[3430] | layer4_out[3431]);
    assign layer5_out[4278] = layer4_out[7045];
    assign layer5_out[4279] = layer4_out[3072] ^ layer4_out[3073];
    assign layer5_out[4280] = ~layer4_out[3439];
    assign layer5_out[4281] = ~layer4_out[3862];
    assign layer5_out[4282] = ~layer4_out[3607];
    assign layer5_out[4283] = ~layer4_out[3439];
    assign layer5_out[4284] = ~(layer4_out[4945] | layer4_out[4946]);
    assign layer5_out[4285] = ~(layer4_out[7663] | layer4_out[7664]);
    assign layer5_out[4286] = layer4_out[4690] & layer4_out[4691];
    assign layer5_out[4287] = ~layer4_out[802];
    assign layer5_out[4288] = ~(layer4_out[6322] & layer4_out[6323]);
    assign layer5_out[4289] = layer4_out[1730];
    assign layer5_out[4290] = ~layer4_out[4485];
    assign layer5_out[4291] = layer4_out[5576];
    assign layer5_out[4292] = layer4_out[4309];
    assign layer5_out[4293] = ~layer4_out[2762];
    assign layer5_out[4294] = ~layer4_out[7172];
    assign layer5_out[4295] = ~(layer4_out[2636] ^ layer4_out[2637]);
    assign layer5_out[4296] = ~(layer4_out[1117] ^ layer4_out[1118]);
    assign layer5_out[4297] = layer4_out[3255] ^ layer4_out[3256];
    assign layer5_out[4298] = ~(layer4_out[2740] ^ layer4_out[2741]);
    assign layer5_out[4299] = layer4_out[7371] & layer4_out[7372];
    assign layer5_out[4300] = layer4_out[2850] & ~layer4_out[2851];
    assign layer5_out[4301] = ~layer4_out[3755];
    assign layer5_out[4302] = ~layer4_out[65];
    assign layer5_out[4303] = layer4_out[2933] ^ layer4_out[2934];
    assign layer5_out[4304] = layer4_out[5239];
    assign layer5_out[4305] = layer4_out[2126] | layer4_out[2127];
    assign layer5_out[4306] = ~layer4_out[228];
    assign layer5_out[4307] = ~(layer4_out[1634] | layer4_out[1635]);
    assign layer5_out[4308] = ~layer4_out[5680];
    assign layer5_out[4309] = layer4_out[3085] & ~layer4_out[3086];
    assign layer5_out[4310] = ~layer4_out[2777] | layer4_out[2776];
    assign layer5_out[4311] = ~(layer4_out[4671] ^ layer4_out[4672]);
    assign layer5_out[4312] = layer4_out[2309];
    assign layer5_out[4313] = ~(layer4_out[3462] ^ layer4_out[3463]);
    assign layer5_out[4314] = ~layer4_out[6770];
    assign layer5_out[4315] = ~layer4_out[272];
    assign layer5_out[4316] = layer4_out[1870];
    assign layer5_out[4317] = ~(layer4_out[4213] ^ layer4_out[4214]);
    assign layer5_out[4318] = ~layer4_out[5456];
    assign layer5_out[4319] = layer4_out[2055] & ~layer4_out[2054];
    assign layer5_out[4320] = layer4_out[6235];
    assign layer5_out[4321] = ~layer4_out[5074] | layer4_out[5073];
    assign layer5_out[4322] = layer4_out[2088];
    assign layer5_out[4323] = layer4_out[4549];
    assign layer5_out[4324] = ~(layer4_out[1343] ^ layer4_out[1344]);
    assign layer5_out[4325] = layer4_out[2081] & layer4_out[2082];
    assign layer5_out[4326] = layer4_out[4298];
    assign layer5_out[4327] = layer4_out[7728];
    assign layer5_out[4328] = layer4_out[7924];
    assign layer5_out[4329] = layer4_out[4439] | layer4_out[4440];
    assign layer5_out[4330] = layer4_out[3396] & ~layer4_out[3397];
    assign layer5_out[4331] = ~layer4_out[6108];
    assign layer5_out[4332] = ~layer4_out[7397];
    assign layer5_out[4333] = ~(layer4_out[3926] ^ layer4_out[3927]);
    assign layer5_out[4334] = ~(layer4_out[4364] | layer4_out[4365]);
    assign layer5_out[4335] = layer4_out[370];
    assign layer5_out[4336] = ~(layer4_out[917] ^ layer4_out[918]);
    assign layer5_out[4337] = layer4_out[2555] & layer4_out[2556];
    assign layer5_out[4338] = ~(layer4_out[7793] ^ layer4_out[7794]);
    assign layer5_out[4339] = layer4_out[4640] ^ layer4_out[4641];
    assign layer5_out[4340] = layer4_out[840];
    assign layer5_out[4341] = ~layer4_out[2638];
    assign layer5_out[4342] = ~layer4_out[2963];
    assign layer5_out[4343] = ~(layer4_out[986] ^ layer4_out[987]);
    assign layer5_out[4344] = ~layer4_out[6119];
    assign layer5_out[4345] = ~(layer4_out[5554] | layer4_out[5555]);
    assign layer5_out[4346] = layer4_out[6673] | layer4_out[6674];
    assign layer5_out[4347] = layer4_out[6988];
    assign layer5_out[4348] = ~layer4_out[6388];
    assign layer5_out[4349] = layer4_out[3008];
    assign layer5_out[4350] = ~layer4_out[5320];
    assign layer5_out[4351] = ~layer4_out[927];
    assign layer5_out[4352] = ~layer4_out[936] | layer4_out[935];
    assign layer5_out[4353] = layer4_out[7886];
    assign layer5_out[4354] = ~(layer4_out[5801] ^ layer4_out[5802]);
    assign layer5_out[4355] = layer4_out[5578];
    assign layer5_out[4356] = ~(layer4_out[7931] & layer4_out[7932]);
    assign layer5_out[4357] = layer4_out[164] ^ layer4_out[165];
    assign layer5_out[4358] = layer4_out[4732];
    assign layer5_out[4359] = layer4_out[5778] & ~layer4_out[5779];
    assign layer5_out[4360] = ~layer4_out[7203];
    assign layer5_out[4361] = layer4_out[115] | layer4_out[116];
    assign layer5_out[4362] = ~layer4_out[1239];
    assign layer5_out[4363] = ~(layer4_out[1508] & layer4_out[1509]);
    assign layer5_out[4364] = ~(layer4_out[4174] ^ layer4_out[4175]);
    assign layer5_out[4365] = ~(layer4_out[6019] ^ layer4_out[6020]);
    assign layer5_out[4366] = layer4_out[1821] & ~layer4_out[1820];
    assign layer5_out[4367] = layer4_out[2636] & ~layer4_out[2635];
    assign layer5_out[4368] = layer4_out[132];
    assign layer5_out[4369] = layer4_out[2162] ^ layer4_out[2163];
    assign layer5_out[4370] = layer4_out[3017] | layer4_out[3018];
    assign layer5_out[4371] = layer4_out[2724];
    assign layer5_out[4372] = ~(layer4_out[3825] & layer4_out[3826]);
    assign layer5_out[4373] = ~layer4_out[7020] | layer4_out[7019];
    assign layer5_out[4374] = ~(layer4_out[1899] ^ layer4_out[1900]);
    assign layer5_out[4375] = ~layer4_out[2811] | layer4_out[2810];
    assign layer5_out[4376] = layer4_out[7688] & ~layer4_out[7689];
    assign layer5_out[4377] = layer4_out[6959] ^ layer4_out[6960];
    assign layer5_out[4378] = layer4_out[6624];
    assign layer5_out[4379] = layer4_out[5373];
    assign layer5_out[4380] = ~layer4_out[7873];
    assign layer5_out[4381] = layer4_out[1346];
    assign layer5_out[4382] = layer4_out[2621] ^ layer4_out[2622];
    assign layer5_out[4383] = layer4_out[4979] & ~layer4_out[4980];
    assign layer5_out[4384] = layer4_out[5271];
    assign layer5_out[4385] = ~(layer4_out[645] | layer4_out[646]);
    assign layer5_out[4386] = layer4_out[3355];
    assign layer5_out[4387] = ~layer4_out[7711];
    assign layer5_out[4388] = layer4_out[143];
    assign layer5_out[4389] = layer4_out[6185];
    assign layer5_out[4390] = layer4_out[6457] & ~layer4_out[6456];
    assign layer5_out[4391] = layer4_out[6458];
    assign layer5_out[4392] = layer4_out[629] & layer4_out[630];
    assign layer5_out[4393] = ~(layer4_out[3381] ^ layer4_out[3382]);
    assign layer5_out[4394] = layer4_out[7956];
    assign layer5_out[4395] = ~(layer4_out[4336] ^ layer4_out[4337]);
    assign layer5_out[4396] = layer4_out[6618] | layer4_out[6619];
    assign layer5_out[4397] = layer4_out[4480] ^ layer4_out[4481];
    assign layer5_out[4398] = ~layer4_out[3206];
    assign layer5_out[4399] = layer4_out[3777] & ~layer4_out[3778];
    assign layer5_out[4400] = layer4_out[1409];
    assign layer5_out[4401] = layer4_out[2687];
    assign layer5_out[4402] = ~layer4_out[5975];
    assign layer5_out[4403] = layer4_out[4300] & ~layer4_out[4299];
    assign layer5_out[4404] = layer4_out[6729] ^ layer4_out[6730];
    assign layer5_out[4405] = layer4_out[3881];
    assign layer5_out[4406] = layer4_out[3095];
    assign layer5_out[4407] = ~layer4_out[6090] | layer4_out[6089];
    assign layer5_out[4408] = layer4_out[4486] ^ layer4_out[4487];
    assign layer5_out[4409] = layer4_out[77] & ~layer4_out[78];
    assign layer5_out[4410] = ~(layer4_out[526] ^ layer4_out[527]);
    assign layer5_out[4411] = ~layer4_out[6711];
    assign layer5_out[4412] = layer4_out[2647] ^ layer4_out[2648];
    assign layer5_out[4413] = layer4_out[4812];
    assign layer5_out[4414] = ~(layer4_out[1303] ^ layer4_out[1304]);
    assign layer5_out[4415] = layer4_out[430] & layer4_out[431];
    assign layer5_out[4416] = layer4_out[1921];
    assign layer5_out[4417] = layer4_out[1626] ^ layer4_out[1627];
    assign layer5_out[4418] = ~(layer4_out[3548] ^ layer4_out[3549]);
    assign layer5_out[4419] = ~(layer4_out[1118] ^ layer4_out[1119]);
    assign layer5_out[4420] = ~layer4_out[6972] | layer4_out[6973];
    assign layer5_out[4421] = ~layer4_out[7251];
    assign layer5_out[4422] = layer4_out[3215];
    assign layer5_out[4423] = ~(layer4_out[192] & layer4_out[193]);
    assign layer5_out[4424] = layer4_out[3340] & layer4_out[3341];
    assign layer5_out[4425] = layer4_out[580] ^ layer4_out[581];
    assign layer5_out[4426] = layer4_out[4360];
    assign layer5_out[4427] = ~layer4_out[6516];
    assign layer5_out[4428] = ~layer4_out[3878];
    assign layer5_out[4429] = ~layer4_out[7809];
    assign layer5_out[4430] = ~(layer4_out[3851] ^ layer4_out[3852]);
    assign layer5_out[4431] = ~layer4_out[2385];
    assign layer5_out[4432] = layer4_out[2144];
    assign layer5_out[4433] = ~layer4_out[5408];
    assign layer5_out[4434] = ~layer4_out[1086];
    assign layer5_out[4435] = ~(layer4_out[6711] | layer4_out[6712]);
    assign layer5_out[4436] = layer4_out[7732] & ~layer4_out[7733];
    assign layer5_out[4437] = layer4_out[4528] & layer4_out[4529];
    assign layer5_out[4438] = layer4_out[55] ^ layer4_out[56];
    assign layer5_out[4439] = ~layer4_out[5131];
    assign layer5_out[4440] = layer4_out[2589] | layer4_out[2590];
    assign layer5_out[4441] = layer4_out[6668] ^ layer4_out[6669];
    assign layer5_out[4442] = layer4_out[5127];
    assign layer5_out[4443] = ~layer4_out[4605];
    assign layer5_out[4444] = layer4_out[6189];
    assign layer5_out[4445] = layer4_out[4144];
    assign layer5_out[4446] = layer4_out[2743] ^ layer4_out[2744];
    assign layer5_out[4447] = ~(layer4_out[6982] ^ layer4_out[6983]);
    assign layer5_out[4448] = layer4_out[4525] ^ layer4_out[4526];
    assign layer5_out[4449] = layer4_out[3938];
    assign layer5_out[4450] = layer4_out[6981];
    assign layer5_out[4451] = layer4_out[287];
    assign layer5_out[4452] = ~layer4_out[1588];
    assign layer5_out[4453] = layer4_out[4708] & layer4_out[4709];
    assign layer5_out[4454] = ~layer4_out[3750];
    assign layer5_out[4455] = layer4_out[914] & layer4_out[915];
    assign layer5_out[4456] = ~layer4_out[3934];
    assign layer5_out[4457] = layer4_out[7550];
    assign layer5_out[4458] = ~layer4_out[1093];
    assign layer5_out[4459] = layer4_out[6565] ^ layer4_out[6566];
    assign layer5_out[4460] = layer4_out[3988] & layer4_out[3989];
    assign layer5_out[4461] = ~(layer4_out[2692] | layer4_out[2693]);
    assign layer5_out[4462] = layer4_out[5212] ^ layer4_out[5213];
    assign layer5_out[4463] = layer4_out[7118];
    assign layer5_out[4464] = layer4_out[1874] & layer4_out[1875];
    assign layer5_out[4465] = ~layer4_out[1299];
    assign layer5_out[4466] = ~(layer4_out[6858] | layer4_out[6859]);
    assign layer5_out[4467] = layer4_out[4813] ^ layer4_out[4814];
    assign layer5_out[4468] = layer4_out[4803];
    assign layer5_out[4469] = layer4_out[3834] | layer4_out[3835];
    assign layer5_out[4470] = ~(layer4_out[1906] & layer4_out[1907]);
    assign layer5_out[4471] = ~(layer4_out[1460] | layer4_out[1461]);
    assign layer5_out[4472] = layer4_out[6639] ^ layer4_out[6640];
    assign layer5_out[4473] = ~layer4_out[7201] | layer4_out[7200];
    assign layer5_out[4474] = layer4_out[2050];
    assign layer5_out[4475] = ~layer4_out[4188];
    assign layer5_out[4476] = layer4_out[7226];
    assign layer5_out[4477] = layer4_out[4156];
    assign layer5_out[4478] = layer4_out[3400] & ~layer4_out[3399];
    assign layer5_out[4479] = layer4_out[6481] & ~layer4_out[6480];
    assign layer5_out[4480] = ~(layer4_out[1017] ^ layer4_out[1018]);
    assign layer5_out[4481] = ~layer4_out[4776] | layer4_out[4775];
    assign layer5_out[4482] = ~(layer4_out[1155] ^ layer4_out[1156]);
    assign layer5_out[4483] = layer4_out[5516];
    assign layer5_out[4484] = layer4_out[2400] ^ layer4_out[2401];
    assign layer5_out[4485] = layer4_out[1466];
    assign layer5_out[4486] = layer4_out[6333];
    assign layer5_out[4487] = layer4_out[5966];
    assign layer5_out[4488] = layer4_out[4768] ^ layer4_out[4769];
    assign layer5_out[4489] = layer4_out[6748] & layer4_out[6749];
    assign layer5_out[4490] = ~layer4_out[71];
    assign layer5_out[4491] = ~layer4_out[7666];
    assign layer5_out[4492] = ~layer4_out[7521];
    assign layer5_out[4493] = layer4_out[7119] ^ layer4_out[7120];
    assign layer5_out[4494] = layer4_out[7240] & ~layer4_out[7241];
    assign layer5_out[4495] = layer4_out[3277] & layer4_out[3278];
    assign layer5_out[4496] = ~layer4_out[1030];
    assign layer5_out[4497] = layer4_out[6254] & layer4_out[6255];
    assign layer5_out[4498] = layer4_out[915];
    assign layer5_out[4499] = ~layer4_out[220];
    assign layer5_out[4500] = ~layer4_out[2630];
    assign layer5_out[4501] = layer4_out[2797];
    assign layer5_out[4502] = layer4_out[5570];
    assign layer5_out[4503] = ~layer4_out[5813];
    assign layer5_out[4504] = layer4_out[5232] & ~layer4_out[5233];
    assign layer5_out[4505] = ~layer4_out[6578];
    assign layer5_out[4506] = layer4_out[5330] & layer4_out[5331];
    assign layer5_out[4507] = layer4_out[2709];
    assign layer5_out[4508] = layer4_out[3021];
    assign layer5_out[4509] = layer4_out[6556] & ~layer4_out[6555];
    assign layer5_out[4510] = ~layer4_out[722];
    assign layer5_out[4511] = ~layer4_out[2826];
    assign layer5_out[4512] = ~(layer4_out[5453] ^ layer4_out[5454]);
    assign layer5_out[4513] = layer4_out[7422];
    assign layer5_out[4514] = ~layer4_out[2318];
    assign layer5_out[4515] = ~layer4_out[275];
    assign layer5_out[4516] = ~layer4_out[4443];
    assign layer5_out[4517] = ~(layer4_out[5207] ^ layer4_out[5208]);
    assign layer5_out[4518] = ~layer4_out[4569];
    assign layer5_out[4519] = layer4_out[4658] ^ layer4_out[4659];
    assign layer5_out[4520] = layer4_out[3129] & ~layer4_out[3130];
    assign layer5_out[4521] = ~(layer4_out[7676] | layer4_out[7677]);
    assign layer5_out[4522] = layer4_out[4452] & layer4_out[4453];
    assign layer5_out[4523] = layer4_out[2374];
    assign layer5_out[4524] = layer4_out[7037] ^ layer4_out[7038];
    assign layer5_out[4525] = layer4_out[1692] & ~layer4_out[1693];
    assign layer5_out[4526] = ~layer4_out[460];
    assign layer5_out[4527] = layer4_out[5638];
    assign layer5_out[4528] = ~(layer4_out[897] ^ layer4_out[898]);
    assign layer5_out[4529] = ~(layer4_out[1669] ^ layer4_out[1670]);
    assign layer5_out[4530] = ~(layer4_out[45] | layer4_out[46]);
    assign layer5_out[4531] = ~(layer4_out[3893] ^ layer4_out[3894]);
    assign layer5_out[4532] = ~layer4_out[4537];
    assign layer5_out[4533] = layer4_out[5049] ^ layer4_out[5050];
    assign layer5_out[4534] = ~layer4_out[5697];
    assign layer5_out[4535] = ~layer4_out[1026];
    assign layer5_out[4536] = layer4_out[4782];
    assign layer5_out[4537] = ~layer4_out[4760] | layer4_out[4759];
    assign layer5_out[4538] = ~layer4_out[1953] | layer4_out[1952];
    assign layer5_out[4539] = layer4_out[528] ^ layer4_out[529];
    assign layer5_out[4540] = ~layer4_out[3068];
    assign layer5_out[4541] = ~(layer4_out[7519] ^ layer4_out[7520]);
    assign layer5_out[4542] = ~layer4_out[5736] | layer4_out[5735];
    assign layer5_out[4543] = layer4_out[6153];
    assign layer5_out[4544] = ~(layer4_out[2164] & layer4_out[2165]);
    assign layer5_out[4545] = ~layer4_out[3791];
    assign layer5_out[4546] = ~layer4_out[3674] | layer4_out[3675];
    assign layer5_out[4547] = layer4_out[6504];
    assign layer5_out[4548] = layer4_out[6672];
    assign layer5_out[4549] = ~(layer4_out[3630] | layer4_out[3631]);
    assign layer5_out[4550] = layer4_out[1034] & layer4_out[1035];
    assign layer5_out[4551] = layer4_out[3722] ^ layer4_out[3723];
    assign layer5_out[4552] = layer4_out[3545] & ~layer4_out[3546];
    assign layer5_out[4553] = ~layer4_out[67];
    assign layer5_out[4554] = ~(layer4_out[6616] ^ layer4_out[6617]);
    assign layer5_out[4555] = layer4_out[1845] ^ layer4_out[1846];
    assign layer5_out[4556] = layer4_out[1319] & ~layer4_out[1320];
    assign layer5_out[4557] = ~layer4_out[568];
    assign layer5_out[4558] = ~layer4_out[7603];
    assign layer5_out[4559] = ~layer4_out[4189];
    assign layer5_out[4560] = ~layer4_out[5862];
    assign layer5_out[4561] = layer4_out[405] ^ layer4_out[406];
    assign layer5_out[4562] = layer4_out[1843] & ~layer4_out[1842];
    assign layer5_out[4563] = layer4_out[3631] ^ layer4_out[3632];
    assign layer5_out[4564] = ~layer4_out[5378];
    assign layer5_out[4565] = layer4_out[3759];
    assign layer5_out[4566] = layer4_out[2718];
    assign layer5_out[4567] = layer4_out[7968] ^ layer4_out[7969];
    assign layer5_out[4568] = ~(layer4_out[4172] ^ layer4_out[4173]);
    assign layer5_out[4569] = layer4_out[6501] & ~layer4_out[6502];
    assign layer5_out[4570] = ~layer4_out[1734];
    assign layer5_out[4571] = ~(layer4_out[454] | layer4_out[455]);
    assign layer5_out[4572] = ~layer4_out[7477];
    assign layer5_out[4573] = layer4_out[3515];
    assign layer5_out[4574] = ~(layer4_out[6810] ^ layer4_out[6811]);
    assign layer5_out[4575] = layer4_out[1697];
    assign layer5_out[4576] = ~layer4_out[1939];
    assign layer5_out[4577] = layer4_out[2988] & ~layer4_out[2987];
    assign layer5_out[4578] = layer4_out[2876];
    assign layer5_out[4579] = layer4_out[2369] ^ layer4_out[2370];
    assign layer5_out[4580] = layer4_out[3394] ^ layer4_out[3395];
    assign layer5_out[4581] = layer4_out[7977] & ~layer4_out[7978];
    assign layer5_out[4582] = ~layer4_out[7206];
    assign layer5_out[4583] = ~(layer4_out[2532] | layer4_out[2533]);
    assign layer5_out[4584] = layer4_out[5007] & ~layer4_out[5006];
    assign layer5_out[4585] = ~layer4_out[739];
    assign layer5_out[4586] = layer4_out[4179] & ~layer4_out[4178];
    assign layer5_out[4587] = ~(layer4_out[858] ^ layer4_out[859]);
    assign layer5_out[4588] = ~layer4_out[604];
    assign layer5_out[4589] = layer4_out[5635] ^ layer4_out[5636];
    assign layer5_out[4590] = layer4_out[7547] & ~layer4_out[7546];
    assign layer5_out[4591] = ~layer4_out[5486];
    assign layer5_out[4592] = ~layer4_out[3998];
    assign layer5_out[4593] = ~layer4_out[5309] | layer4_out[5310];
    assign layer5_out[4594] = layer4_out[6494] ^ layer4_out[6495];
    assign layer5_out[4595] = ~(layer4_out[1740] & layer4_out[1741]);
    assign layer5_out[4596] = ~layer4_out[4797] | layer4_out[4796];
    assign layer5_out[4597] = layer4_out[1201] ^ layer4_out[1202];
    assign layer5_out[4598] = layer4_out[5283];
    assign layer5_out[4599] = layer4_out[2768] & ~layer4_out[2767];
    assign layer5_out[4600] = ~layer4_out[3741];
    assign layer5_out[4601] = layer4_out[6372];
    assign layer5_out[4602] = layer4_out[2357];
    assign layer5_out[4603] = layer4_out[6113] & ~layer4_out[6114];
    assign layer5_out[4604] = layer4_out[3854] & layer4_out[3855];
    assign layer5_out[4605] = ~(layer4_out[5687] ^ layer4_out[5688]);
    assign layer5_out[4606] = ~(layer4_out[7182] ^ layer4_out[7183]);
    assign layer5_out[4607] = layer4_out[5924];
    assign layer5_out[4608] = ~layer4_out[1734];
    assign layer5_out[4609] = layer4_out[266];
    assign layer5_out[4610] = ~layer4_out[1780];
    assign layer5_out[4611] = layer4_out[6143] ^ layer4_out[6144];
    assign layer5_out[4612] = ~(layer4_out[6066] ^ layer4_out[6067]);
    assign layer5_out[4613] = ~layer4_out[2911];
    assign layer5_out[4614] = ~layer4_out[489];
    assign layer5_out[4615] = ~layer4_out[493] | layer4_out[492];
    assign layer5_out[4616] = ~layer4_out[1657];
    assign layer5_out[4617] = ~(layer4_out[7189] | layer4_out[7190]);
    assign layer5_out[4618] = ~layer4_out[6491] | layer4_out[6492];
    assign layer5_out[4619] = layer4_out[7738] | layer4_out[7739];
    assign layer5_out[4620] = layer4_out[6974] ^ layer4_out[6975];
    assign layer5_out[4621] = ~layer4_out[972];
    assign layer5_out[4622] = layer4_out[167] ^ layer4_out[168];
    assign layer5_out[4623] = ~layer4_out[7709];
    assign layer5_out[4624] = layer4_out[3937] & ~layer4_out[3936];
    assign layer5_out[4625] = layer4_out[2112] & layer4_out[2113];
    assign layer5_out[4626] = ~layer4_out[5483];
    assign layer5_out[4627] = ~layer4_out[5682];
    assign layer5_out[4628] = ~layer4_out[280];
    assign layer5_out[4629] = layer4_out[1818] & ~layer4_out[1817];
    assign layer5_out[4630] = layer4_out[4716] | layer4_out[4717];
    assign layer5_out[4631] = layer4_out[1602] & layer4_out[1603];
    assign layer5_out[4632] = layer4_out[2970] & ~layer4_out[2971];
    assign layer5_out[4633] = layer4_out[3781] ^ layer4_out[3782];
    assign layer5_out[4634] = ~layer4_out[439];
    assign layer5_out[4635] = ~layer4_out[7513] | layer4_out[7514];
    assign layer5_out[4636] = layer4_out[7080] & ~layer4_out[7081];
    assign layer5_out[4637] = layer4_out[1136] & ~layer4_out[1137];
    assign layer5_out[4638] = layer4_out[6545] ^ layer4_out[6546];
    assign layer5_out[4639] = ~layer4_out[3397] | layer4_out[3398];
    assign layer5_out[4640] = ~layer4_out[2158];
    assign layer5_out[4641] = layer4_out[7422];
    assign layer5_out[4642] = ~(layer4_out[7111] & layer4_out[7112]);
    assign layer5_out[4643] = ~layer4_out[562];
    assign layer5_out[4644] = ~layer4_out[6120];
    assign layer5_out[4645] = ~(layer4_out[2972] ^ layer4_out[2973]);
    assign layer5_out[4646] = layer4_out[5982] & layer4_out[5983];
    assign layer5_out[4647] = layer4_out[7078];
    assign layer5_out[4648] = ~layer4_out[6405];
    assign layer5_out[4649] = ~(layer4_out[5202] ^ layer4_out[5203]);
    assign layer5_out[4650] = layer4_out[26] ^ layer4_out[27];
    assign layer5_out[4651] = ~(layer4_out[7195] | layer4_out[7196]);
    assign layer5_out[4652] = ~layer4_out[3739];
    assign layer5_out[4653] = layer4_out[3840];
    assign layer5_out[4654] = layer4_out[7071];
    assign layer5_out[4655] = ~layer4_out[6058];
    assign layer5_out[4656] = layer4_out[3883] & layer4_out[3884];
    assign layer5_out[4657] = ~(layer4_out[3268] ^ layer4_out[3269]);
    assign layer5_out[4658] = ~layer4_out[5285];
    assign layer5_out[4659] = layer4_out[2576] & layer4_out[2577];
    assign layer5_out[4660] = ~layer4_out[7725];
    assign layer5_out[4661] = layer4_out[1950];
    assign layer5_out[4662] = layer4_out[2412] & layer4_out[2413];
    assign layer5_out[4663] = ~layer4_out[6597];
    assign layer5_out[4664] = ~layer4_out[3162];
    assign layer5_out[4665] = layer4_out[1943] ^ layer4_out[1944];
    assign layer5_out[4666] = ~(layer4_out[3217] ^ layer4_out[3218]);
    assign layer5_out[4667] = ~layer4_out[7081] | layer4_out[7082];
    assign layer5_out[4668] = layer4_out[2571] | layer4_out[2572];
    assign layer5_out[4669] = layer4_out[4250] | layer4_out[4251];
    assign layer5_out[4670] = ~(layer4_out[862] | layer4_out[863]);
    assign layer5_out[4671] = layer4_out[1648];
    assign layer5_out[4672] = layer4_out[145];
    assign layer5_out[4673] = ~(layer4_out[481] ^ layer4_out[482]);
    assign layer5_out[4674] = layer4_out[6166] & ~layer4_out[6165];
    assign layer5_out[4675] = layer4_out[3960];
    assign layer5_out[4676] = ~layer4_out[4218];
    assign layer5_out[4677] = ~layer4_out[1767] | layer4_out[1766];
    assign layer5_out[4678] = ~layer4_out[5042] | layer4_out[5041];
    assign layer5_out[4679] = layer4_out[391] | layer4_out[392];
    assign layer5_out[4680] = ~(layer4_out[2084] | layer4_out[2085]);
    assign layer5_out[4681] = layer4_out[7545] & ~layer4_out[7546];
    assign layer5_out[4682] = ~(layer4_out[7768] ^ layer4_out[7769]);
    assign layer5_out[4683] = ~layer4_out[3919];
    assign layer5_out[4684] = layer4_out[7661];
    assign layer5_out[4685] = ~layer4_out[16];
    assign layer5_out[4686] = ~layer4_out[780];
    assign layer5_out[4687] = ~(layer4_out[1259] ^ layer4_out[1260]);
    assign layer5_out[4688] = ~layer4_out[3734];
    assign layer5_out[4689] = ~layer4_out[3651];
    assign layer5_out[4690] = ~(layer4_out[399] ^ layer4_out[400]);
    assign layer5_out[4691] = layer4_out[885] ^ layer4_out[886];
    assign layer5_out[4692] = layer4_out[2513] & layer4_out[2514];
    assign layer5_out[4693] = ~layer4_out[3903];
    assign layer5_out[4694] = ~layer4_out[3772];
    assign layer5_out[4695] = ~layer4_out[3919] | layer4_out[3920];
    assign layer5_out[4696] = layer4_out[7054];
    assign layer5_out[4697] = ~(layer4_out[7850] ^ layer4_out[7851]);
    assign layer5_out[4698] = layer4_out[3320];
    assign layer5_out[4699] = layer4_out[5597];
    assign layer5_out[4700] = ~layer4_out[3220];
    assign layer5_out[4701] = ~layer4_out[2421];
    assign layer5_out[4702] = layer4_out[4030];
    assign layer5_out[4703] = ~layer4_out[5036];
    assign layer5_out[4704] = layer4_out[6301] & ~layer4_out[6300];
    assign layer5_out[4705] = ~layer4_out[3976];
    assign layer5_out[4706] = ~(layer4_out[372] | layer4_out[373]);
    assign layer5_out[4707] = ~layer4_out[6818];
    assign layer5_out[4708] = ~(layer4_out[7863] ^ layer4_out[7864]);
    assign layer5_out[4709] = layer4_out[2608] ^ layer4_out[2609];
    assign layer5_out[4710] = layer4_out[6140];
    assign layer5_out[4711] = ~layer4_out[4317];
    assign layer5_out[4712] = layer4_out[5844] & ~layer4_out[5843];
    assign layer5_out[4713] = layer4_out[4858] ^ layer4_out[4859];
    assign layer5_out[4714] = layer4_out[4258];
    assign layer5_out[4715] = ~layer4_out[1617];
    assign layer5_out[4716] = layer4_out[7972] & layer4_out[7973];
    assign layer5_out[4717] = ~layer4_out[14];
    assign layer5_out[4718] = ~layer4_out[175];
    assign layer5_out[4719] = ~layer4_out[535];
    assign layer5_out[4720] = ~layer4_out[1282];
    assign layer5_out[4721] = layer4_out[7544] ^ layer4_out[7545];
    assign layer5_out[4722] = layer4_out[3312] & ~layer4_out[3311];
    assign layer5_out[4723] = layer4_out[4377] ^ layer4_out[4378];
    assign layer5_out[4724] = layer4_out[5568];
    assign layer5_out[4725] = ~layer4_out[5038] | layer4_out[5039];
    assign layer5_out[4726] = layer4_out[4345];
    assign layer5_out[4727] = layer4_out[787];
    assign layer5_out[4728] = ~layer4_out[5588];
    assign layer5_out[4729] = ~layer4_out[5019];
    assign layer5_out[4730] = ~(layer4_out[6863] & layer4_out[6864]);
    assign layer5_out[4731] = ~layer4_out[4530];
    assign layer5_out[4732] = layer4_out[7648];
    assign layer5_out[4733] = ~layer4_out[1061];
    assign layer5_out[4734] = layer4_out[5769] | layer4_out[5770];
    assign layer5_out[4735] = ~layer4_out[5580];
    assign layer5_out[4736] = layer4_out[1327] ^ layer4_out[1328];
    assign layer5_out[4737] = ~layer4_out[4734] | layer4_out[4735];
    assign layer5_out[4738] = layer4_out[7306] ^ layer4_out[7307];
    assign layer5_out[4739] = ~layer4_out[3367];
    assign layer5_out[4740] = layer4_out[5838] | layer4_out[5839];
    assign layer5_out[4741] = layer4_out[1713];
    assign layer5_out[4742] = layer4_out[6800] ^ layer4_out[6801];
    assign layer5_out[4743] = layer4_out[2366] & ~layer4_out[2367];
    assign layer5_out[4744] = ~layer4_out[3581];
    assign layer5_out[4745] = layer4_out[7086];
    assign layer5_out[4746] = layer4_out[3002] & ~layer4_out[3003];
    assign layer5_out[4747] = ~layer4_out[6120];
    assign layer5_out[4748] = ~(layer4_out[1656] ^ layer4_out[1657]);
    assign layer5_out[4749] = ~(layer4_out[6369] ^ layer4_out[6370]);
    assign layer5_out[4750] = layer4_out[4456] ^ layer4_out[4457];
    assign layer5_out[4751] = layer4_out[6125];
    assign layer5_out[4752] = layer4_out[5517];
    assign layer5_out[4753] = ~layer4_out[6701];
    assign layer5_out[4754] = ~(layer4_out[2077] | layer4_out[2078]);
    assign layer5_out[4755] = layer4_out[3605] ^ layer4_out[3606];
    assign layer5_out[4756] = layer4_out[3662] & layer4_out[3663];
    assign layer5_out[4757] = ~(layer4_out[4100] | layer4_out[4101]);
    assign layer5_out[4758] = layer4_out[6855];
    assign layer5_out[4759] = layer4_out[4310] ^ layer4_out[4311];
    assign layer5_out[4760] = ~layer4_out[1546];
    assign layer5_out[4761] = layer4_out[5990];
    assign layer5_out[4762] = layer4_out[3177];
    assign layer5_out[4763] = ~layer4_out[2080];
    assign layer5_out[4764] = layer4_out[142];
    assign layer5_out[4765] = layer4_out[7346];
    assign layer5_out[4766] = layer4_out[2819] ^ layer4_out[2820];
    assign layer5_out[4767] = layer4_out[2461] & layer4_out[2462];
    assign layer5_out[4768] = layer4_out[5300] & ~layer4_out[5299];
    assign layer5_out[4769] = ~layer4_out[5957];
    assign layer5_out[4770] = layer4_out[6911] & ~layer4_out[6912];
    assign layer5_out[4771] = layer4_out[6772];
    assign layer5_out[4772] = ~(layer4_out[5960] | layer4_out[5961]);
    assign layer5_out[4773] = ~(layer4_out[1628] | layer4_out[1629]);
    assign layer5_out[4774] = layer4_out[3806] & layer4_out[3807];
    assign layer5_out[4775] = layer4_out[4521];
    assign layer5_out[4776] = layer4_out[1166];
    assign layer5_out[4777] = ~(layer4_out[7227] ^ layer4_out[7228]);
    assign layer5_out[4778] = layer4_out[7047] ^ layer4_out[7048];
    assign layer5_out[4779] = layer4_out[1202] ^ layer4_out[1203];
    assign layer5_out[4780] = ~layer4_out[5816];
    assign layer5_out[4781] = layer4_out[7971];
    assign layer5_out[4782] = ~layer4_out[2190] | layer4_out[2189];
    assign layer5_out[4783] = layer4_out[4921];
    assign layer5_out[4784] = ~layer4_out[6165];
    assign layer5_out[4785] = layer4_out[2778] & ~layer4_out[2779];
    assign layer5_out[4786] = layer4_out[5452] ^ layer4_out[5453];
    assign layer5_out[4787] = ~layer4_out[4771];
    assign layer5_out[4788] = ~layer4_out[3240] | layer4_out[3241];
    assign layer5_out[4789] = ~layer4_out[1737] | layer4_out[1736];
    assign layer5_out[4790] = layer4_out[2601] | layer4_out[2602];
    assign layer5_out[4791] = layer4_out[4007] ^ layer4_out[4008];
    assign layer5_out[4792] = ~(layer4_out[5608] ^ layer4_out[5609]);
    assign layer5_out[4793] = layer4_out[1146];
    assign layer5_out[4794] = ~(layer4_out[4478] ^ layer4_out[4479]);
    assign layer5_out[4795] = layer4_out[3937] & layer4_out[3938];
    assign layer5_out[4796] = ~(layer4_out[1810] ^ layer4_out[1811]);
    assign layer5_out[4797] = ~layer4_out[2040] | layer4_out[2041];
    assign layer5_out[4798] = layer4_out[694] ^ layer4_out[695];
    assign layer5_out[4799] = ~layer4_out[3862];
    assign layer5_out[4800] = ~(layer4_out[6241] | layer4_out[6242]);
    assign layer5_out[4801] = ~layer4_out[3215];
    assign layer5_out[4802] = layer4_out[6206];
    assign layer5_out[4803] = layer4_out[5064];
    assign layer5_out[4804] = ~(layer4_out[2891] ^ layer4_out[2892]);
    assign layer5_out[4805] = layer4_out[5021] ^ layer4_out[5022];
    assign layer5_out[4806] = ~(layer4_out[6899] | layer4_out[6900]);
    assign layer5_out[4807] = layer4_out[5980];
    assign layer5_out[4808] = ~layer4_out[6036];
    assign layer5_out[4809] = layer4_out[3304];
    assign layer5_out[4810] = ~(layer4_out[320] | layer4_out[321]);
    assign layer5_out[4811] = layer4_out[2352];
    assign layer5_out[4812] = layer4_out[6059] ^ layer4_out[6060];
    assign layer5_out[4813] = ~layer4_out[7561];
    assign layer5_out[4814] = ~layer4_out[6048];
    assign layer5_out[4815] = layer4_out[5545] ^ layer4_out[5546];
    assign layer5_out[4816] = ~(layer4_out[412] & layer4_out[413]);
    assign layer5_out[4817] = ~layer4_out[7242];
    assign layer5_out[4818] = ~layer4_out[4366];
    assign layer5_out[4819] = layer4_out[561] & layer4_out[562];
    assign layer5_out[4820] = layer4_out[1611] | layer4_out[1612];
    assign layer5_out[4821] = ~layer4_out[5997];
    assign layer5_out[4822] = layer4_out[3298] ^ layer4_out[3299];
    assign layer5_out[4823] = layer4_out[5047];
    assign layer5_out[4824] = layer4_out[3624] ^ layer4_out[3625];
    assign layer5_out[4825] = layer4_out[2937];
    assign layer5_out[4826] = ~(layer4_out[4468] ^ layer4_out[4469]);
    assign layer5_out[4827] = layer4_out[4314];
    assign layer5_out[4828] = ~layer4_out[4117];
    assign layer5_out[4829] = ~(layer4_out[5889] ^ layer4_out[5890]);
    assign layer5_out[4830] = layer4_out[1915] & ~layer4_out[1914];
    assign layer5_out[4831] = ~layer4_out[4170];
    assign layer5_out[4832] = layer4_out[7210] & ~layer4_out[7211];
    assign layer5_out[4833] = layer4_out[4997];
    assign layer5_out[4834] = layer4_out[1112] & ~layer4_out[1113];
    assign layer5_out[4835] = layer4_out[1843];
    assign layer5_out[4836] = layer4_out[1548];
    assign layer5_out[4837] = ~layer4_out[459] | layer4_out[458];
    assign layer5_out[4838] = layer4_out[4718];
    assign layer5_out[4839] = ~(layer4_out[7901] ^ layer4_out[7902]);
    assign layer5_out[4840] = layer4_out[3375] & ~layer4_out[3374];
    assign layer5_out[4841] = layer4_out[3016] | layer4_out[3017];
    assign layer5_out[4842] = ~(layer4_out[2160] ^ layer4_out[2161]);
    assign layer5_out[4843] = layer4_out[3252];
    assign layer5_out[4844] = ~(layer4_out[3866] | layer4_out[3867]);
    assign layer5_out[4845] = layer4_out[5475];
    assign layer5_out[4846] = ~layer4_out[641];
    assign layer5_out[4847] = ~layer4_out[4316];
    assign layer5_out[4848] = ~(layer4_out[4475] ^ layer4_out[4476]);
    assign layer5_out[4849] = ~layer4_out[793];
    assign layer5_out[4850] = ~layer4_out[1890];
    assign layer5_out[4851] = ~layer4_out[2771] | layer4_out[2772];
    assign layer5_out[4852] = ~layer4_out[5818];
    assign layer5_out[4853] = layer4_out[7717];
    assign layer5_out[4854] = layer4_out[4734];
    assign layer5_out[4855] = ~layer4_out[4044];
    assign layer5_out[4856] = ~layer4_out[7442];
    assign layer5_out[4857] = ~layer4_out[7540] | layer4_out[7539];
    assign layer5_out[4858] = ~layer4_out[860];
    assign layer5_out[4859] = layer4_out[6587] & ~layer4_out[6588];
    assign layer5_out[4860] = layer4_out[4008] ^ layer4_out[4009];
    assign layer5_out[4861] = layer4_out[1131] & ~layer4_out[1132];
    assign layer5_out[4862] = ~layer4_out[3678];
    assign layer5_out[4863] = layer4_out[6849];
    assign layer5_out[4864] = ~(layer4_out[2640] ^ layer4_out[2641]);
    assign layer5_out[4865] = ~(layer4_out[5538] ^ layer4_out[5539]);
    assign layer5_out[4866] = layer4_out[2118];
    assign layer5_out[4867] = layer4_out[3618];
    assign layer5_out[4868] = ~layer4_out[3364];
    assign layer5_out[4869] = layer4_out[7473] ^ layer4_out[7474];
    assign layer5_out[4870] = ~(layer4_out[1558] ^ layer4_out[1559]);
    assign layer5_out[4871] = layer4_out[1498] & layer4_out[1499];
    assign layer5_out[4872] = ~layer4_out[2821];
    assign layer5_out[4873] = ~layer4_out[2766];
    assign layer5_out[4874] = ~(layer4_out[133] ^ layer4_out[134]);
    assign layer5_out[4875] = layer4_out[2862] & ~layer4_out[2861];
    assign layer5_out[4876] = ~(layer4_out[3404] & layer4_out[3405]);
    assign layer5_out[4877] = layer4_out[5890] & layer4_out[5891];
    assign layer5_out[4878] = ~layer4_out[4964] | layer4_out[4963];
    assign layer5_out[4879] = layer4_out[1977] & ~layer4_out[1978];
    assign layer5_out[4880] = ~layer4_out[6140] | layer4_out[6141];
    assign layer5_out[4881] = layer4_out[4747];
    assign layer5_out[4882] = layer4_out[7323] & ~layer4_out[7324];
    assign layer5_out[4883] = layer4_out[2300];
    assign layer5_out[4884] = layer4_out[117] ^ layer4_out[118];
    assign layer5_out[4885] = ~(layer4_out[3259] ^ layer4_out[3260]);
    assign layer5_out[4886] = layer4_out[4903] & ~layer4_out[4902];
    assign layer5_out[4887] = layer4_out[7432];
    assign layer5_out[4888] = ~layer4_out[6621];
    assign layer5_out[4889] = layer4_out[2030];
    assign layer5_out[4890] = ~layer4_out[7162];
    assign layer5_out[4891] = ~(layer4_out[5056] ^ layer4_out[5057]);
    assign layer5_out[4892] = ~(layer4_out[2859] | layer4_out[2860]);
    assign layer5_out[4893] = ~layer4_out[5306];
    assign layer5_out[4894] = ~(layer4_out[2239] | layer4_out[2240]);
    assign layer5_out[4895] = layer4_out[2852] & ~layer4_out[2853];
    assign layer5_out[4896] = ~(layer4_out[3059] ^ layer4_out[3060]);
    assign layer5_out[4897] = layer4_out[7767] ^ layer4_out[7768];
    assign layer5_out[4898] = layer4_out[5687];
    assign layer5_out[4899] = ~layer4_out[3735] | layer4_out[3736];
    assign layer5_out[4900] = layer4_out[2554];
    assign layer5_out[4901] = layer4_out[3941];
    assign layer5_out[4902] = layer4_out[2023] ^ layer4_out[2024];
    assign layer5_out[4903] = ~(layer4_out[3108] | layer4_out[3109]);
    assign layer5_out[4904] = layer4_out[7248] & ~layer4_out[7249];
    assign layer5_out[4905] = layer4_out[1519];
    assign layer5_out[4906] = layer4_out[421] ^ layer4_out[422];
    assign layer5_out[4907] = ~(layer4_out[6650] ^ layer4_out[6651]);
    assign layer5_out[4908] = layer4_out[576];
    assign layer5_out[4909] = layer4_out[1895];
    assign layer5_out[4910] = layer4_out[5253];
    assign layer5_out[4911] = ~layer4_out[1852] | layer4_out[1851];
    assign layer5_out[4912] = layer4_out[604];
    assign layer5_out[4913] = layer4_out[1511] | layer4_out[1512];
    assign layer5_out[4914] = ~(layer4_out[6248] ^ layer4_out[6249]);
    assign layer5_out[4915] = ~layer4_out[4362];
    assign layer5_out[4916] = layer4_out[1612];
    assign layer5_out[4917] = layer4_out[2281];
    assign layer5_out[4918] = ~layer4_out[2205] | layer4_out[2204];
    assign layer5_out[4919] = layer4_out[2360];
    assign layer5_out[4920] = ~layer4_out[2982] | layer4_out[2983];
    assign layer5_out[4921] = layer4_out[2266] ^ layer4_out[2267];
    assign layer5_out[4922] = layer4_out[735] | layer4_out[736];
    assign layer5_out[4923] = layer4_out[2475] ^ layer4_out[2476];
    assign layer5_out[4924] = ~layer4_out[442];
    assign layer5_out[4925] = ~(layer4_out[978] ^ layer4_out[979]);
    assign layer5_out[4926] = ~layer4_out[3649];
    assign layer5_out[4927] = ~layer4_out[1340];
    assign layer5_out[4928] = ~layer4_out[5183];
    assign layer5_out[4929] = ~layer4_out[1132] | layer4_out[1133];
    assign layer5_out[4930] = layer4_out[3564] & ~layer4_out[3565];
    assign layer5_out[4931] = layer4_out[367];
    assign layer5_out[4932] = ~layer4_out[7635];
    assign layer5_out[4933] = ~layer4_out[3857];
    assign layer5_out[4934] = ~(layer4_out[6161] | layer4_out[6162]);
    assign layer5_out[4935] = ~layer4_out[4824];
    assign layer5_out[4936] = ~layer4_out[7224];
    assign layer5_out[4937] = ~layer4_out[4567] | layer4_out[4566];
    assign layer5_out[4938] = layer4_out[82];
    assign layer5_out[4939] = layer4_out[7804] ^ layer4_out[7805];
    assign layer5_out[4940] = layer4_out[1133] | layer4_out[1134];
    assign layer5_out[4941] = layer4_out[7987];
    assign layer5_out[4942] = layer4_out[5023] ^ layer4_out[5024];
    assign layer5_out[4943] = ~layer4_out[1141];
    assign layer5_out[4944] = layer4_out[7023] & layer4_out[7024];
    assign layer5_out[4945] = layer4_out[189];
    assign layer5_out[4946] = layer4_out[1234];
    assign layer5_out[4947] = layer4_out[7125] & ~layer4_out[7124];
    assign layer5_out[4948] = layer4_out[972];
    assign layer5_out[4949] = layer4_out[7382];
    assign layer5_out[4950] = ~layer4_out[270];
    assign layer5_out[4951] = layer4_out[2737] ^ layer4_out[2738];
    assign layer5_out[4952] = layer4_out[1073] ^ layer4_out[1074];
    assign layer5_out[4953] = layer4_out[5994];
    assign layer5_out[4954] = layer4_out[2395] & ~layer4_out[2394];
    assign layer5_out[4955] = ~layer4_out[3503];
    assign layer5_out[4956] = layer4_out[3511] | layer4_out[3512];
    assign layer5_out[4957] = ~layer4_out[4141];
    assign layer5_out[4958] = layer4_out[7462];
    assign layer5_out[4959] = layer4_out[1275] | layer4_out[1276];
    assign layer5_out[4960] = layer4_out[1595];
    assign layer5_out[4961] = ~layer4_out[767];
    assign layer5_out[4962] = layer4_out[7247] & layer4_out[7248];
    assign layer5_out[4963] = layer4_out[6351] ^ layer4_out[6352];
    assign layer5_out[4964] = ~layer4_out[4168];
    assign layer5_out[4965] = layer4_out[4449];
    assign layer5_out[4966] = layer4_out[3887];
    assign layer5_out[4967] = ~layer4_out[2428];
    assign layer5_out[4968] = layer4_out[7452] ^ layer4_out[7453];
    assign layer5_out[4969] = layer4_out[6109];
    assign layer5_out[4970] = ~layer4_out[4526] | layer4_out[4527];
    assign layer5_out[4971] = layer4_out[285];
    assign layer5_out[4972] = layer4_out[2302];
    assign layer5_out[4973] = layer4_out[195] ^ layer4_out[196];
    assign layer5_out[4974] = layer4_out[1811];
    assign layer5_out[4975] = ~layer4_out[3107];
    assign layer5_out[4976] = ~layer4_out[3097];
    assign layer5_out[4977] = ~(layer4_out[3648] & layer4_out[3649]);
    assign layer5_out[4978] = layer4_out[6025];
    assign layer5_out[4979] = layer4_out[6285] & ~layer4_out[6284];
    assign layer5_out[4980] = ~(layer4_out[326] | layer4_out[327]);
    assign layer5_out[4981] = layer4_out[7559] ^ layer4_out[7560];
    assign layer5_out[4982] = layer4_out[22] & ~layer4_out[21];
    assign layer5_out[4983] = layer4_out[4497];
    assign layer5_out[4984] = layer4_out[405] & ~layer4_out[404];
    assign layer5_out[4985] = ~layer4_out[7566];
    assign layer5_out[4986] = layer4_out[2219];
    assign layer5_out[4987] = ~(layer4_out[2428] | layer4_out[2429]);
    assign layer5_out[4988] = ~layer4_out[4129] | layer4_out[4128];
    assign layer5_out[4989] = layer4_out[6039] & ~layer4_out[6040];
    assign layer5_out[4990] = layer4_out[3599] & ~layer4_out[3600];
    assign layer5_out[4991] = layer4_out[845] & layer4_out[846];
    assign layer5_out[4992] = ~layer4_out[580];
    assign layer5_out[4993] = ~layer4_out[4588];
    assign layer5_out[4994] = ~(layer4_out[6615] ^ layer4_out[6616]);
    assign layer5_out[4995] = ~layer4_out[5975] | layer4_out[5974];
    assign layer5_out[4996] = ~layer4_out[1317];
    assign layer5_out[4997] = ~layer4_out[5897];
    assign layer5_out[4998] = ~(layer4_out[234] ^ layer4_out[235]);
    assign layer5_out[4999] = ~(layer4_out[5156] | layer4_out[5157]);
    assign layer5_out[5000] = ~layer4_out[5945];
    assign layer5_out[5001] = ~layer4_out[5825];
    assign layer5_out[5002] = layer4_out[5313] & layer4_out[5314];
    assign layer5_out[5003] = ~layer4_out[2064] | layer4_out[2065];
    assign layer5_out[5004] = ~layer4_out[4621] | layer4_out[4620];
    assign layer5_out[5005] = layer4_out[6967] | layer4_out[6968];
    assign layer5_out[5006] = ~layer4_out[4562];
    assign layer5_out[5007] = layer4_out[6501];
    assign layer5_out[5008] = ~(layer4_out[2827] | layer4_out[2828]);
    assign layer5_out[5009] = ~(layer4_out[4245] ^ layer4_out[4246]);
    assign layer5_out[5010] = ~layer4_out[280];
    assign layer5_out[5011] = layer4_out[5691] & ~layer4_out[5690];
    assign layer5_out[5012] = layer4_out[6764] & layer4_out[6765];
    assign layer5_out[5013] = layer4_out[653];
    assign layer5_out[5014] = layer4_out[3928] & layer4_out[3929];
    assign layer5_out[5015] = ~(layer4_out[3418] & layer4_out[3419]);
    assign layer5_out[5016] = layer4_out[6832];
    assign layer5_out[5017] = ~layer4_out[2229];
    assign layer5_out[5018] = ~(layer4_out[2897] | layer4_out[2898]);
    assign layer5_out[5019] = layer4_out[5317];
    assign layer5_out[5020] = ~layer4_out[5264];
    assign layer5_out[5021] = ~layer4_out[6569];
    assign layer5_out[5022] = layer4_out[3015] | layer4_out[3016];
    assign layer5_out[5023] = layer4_out[1677];
    assign layer5_out[5024] = layer4_out[4550] | layer4_out[4551];
    assign layer5_out[5025] = ~layer4_out[1566];
    assign layer5_out[5026] = layer4_out[6028] & ~layer4_out[6027];
    assign layer5_out[5027] = ~layer4_out[6388];
    assign layer5_out[5028] = layer4_out[2040];
    assign layer5_out[5029] = ~layer4_out[4783] | layer4_out[4784];
    assign layer5_out[5030] = layer4_out[957] ^ layer4_out[958];
    assign layer5_out[5031] = layer4_out[7058];
    assign layer5_out[5032] = ~layer4_out[212] | layer4_out[211];
    assign layer5_out[5033] = ~layer4_out[1784];
    assign layer5_out[5034] = ~layer4_out[1729];
    assign layer5_out[5035] = ~layer4_out[6802] | layer4_out[6801];
    assign layer5_out[5036] = ~(layer4_out[6288] ^ layer4_out[6289]);
    assign layer5_out[5037] = ~(layer4_out[2177] | layer4_out[2178]);
    assign layer5_out[5038] = ~(layer4_out[3346] | layer4_out[3347]);
    assign layer5_out[5039] = layer4_out[5154] & ~layer4_out[5155];
    assign layer5_out[5040] = layer4_out[2995] & ~layer4_out[2994];
    assign layer5_out[5041] = ~layer4_out[4666];
    assign layer5_out[5042] = ~layer4_out[7220];
    assign layer5_out[5043] = ~layer4_out[6582];
    assign layer5_out[5044] = ~layer4_out[7695];
    assign layer5_out[5045] = layer4_out[3910] ^ layer4_out[3911];
    assign layer5_out[5046] = ~layer4_out[6946] | layer4_out[6945];
    assign layer5_out[5047] = ~layer4_out[1324];
    assign layer5_out[5048] = ~layer4_out[1669];
    assign layer5_out[5049] = layer4_out[6642];
    assign layer5_out[5050] = ~(layer4_out[428] ^ layer4_out[429]);
    assign layer5_out[5051] = layer4_out[5539] ^ layer4_out[5540];
    assign layer5_out[5052] = layer4_out[313] ^ layer4_out[314];
    assign layer5_out[5053] = ~layer4_out[7450];
    assign layer5_out[5054] = ~layer4_out[5149];
    assign layer5_out[5055] = ~layer4_out[3914];
    assign layer5_out[5056] = layer4_out[448] & ~layer4_out[447];
    assign layer5_out[5057] = layer4_out[6559] & ~layer4_out[6558];
    assign layer5_out[5058] = layer4_out[2045] ^ layer4_out[2046];
    assign layer5_out[5059] = layer4_out[6417];
    assign layer5_out[5060] = layer4_out[1304] ^ layer4_out[1305];
    assign layer5_out[5061] = ~layer4_out[4366];
    assign layer5_out[5062] = layer4_out[1983] ^ layer4_out[1984];
    assign layer5_out[5063] = ~layer4_out[4269];
    assign layer5_out[5064] = ~layer4_out[5437];
    assign layer5_out[5065] = ~layer4_out[1841];
    assign layer5_out[5066] = layer4_out[7698];
    assign layer5_out[5067] = ~(layer4_out[6085] | layer4_out[6086]);
    assign layer5_out[5068] = layer4_out[6522] & ~layer4_out[6523];
    assign layer5_out[5069] = ~layer4_out[1428];
    assign layer5_out[5070] = ~(layer4_out[4920] ^ layer4_out[4921]);
    assign layer5_out[5071] = ~layer4_out[5706];
    assign layer5_out[5072] = ~layer4_out[2652];
    assign layer5_out[5073] = layer4_out[2596];
    assign layer5_out[5074] = layer4_out[2607] & layer4_out[2608];
    assign layer5_out[5075] = layer4_out[4312] & ~layer4_out[4311];
    assign layer5_out[5076] = ~layer4_out[7391] | layer4_out[7392];
    assign layer5_out[5077] = ~layer4_out[7068] | layer4_out[7069];
    assign layer5_out[5078] = layer4_out[4006] ^ layer4_out[4007];
    assign layer5_out[5079] = layer4_out[4162] & ~layer4_out[4161];
    assign layer5_out[5080] = ~layer4_out[6553];
    assign layer5_out[5081] = ~layer4_out[2423];
    assign layer5_out[5082] = layer4_out[6375];
    assign layer5_out[5083] = ~(layer4_out[7137] | layer4_out[7138]);
    assign layer5_out[5084] = ~layer4_out[6554];
    assign layer5_out[5085] = ~layer4_out[2800] | layer4_out[2799];
    assign layer5_out[5086] = ~layer4_out[4337];
    assign layer5_out[5087] = layer4_out[4266] & ~layer4_out[4265];
    assign layer5_out[5088] = ~layer4_out[1414] | layer4_out[1415];
    assign layer5_out[5089] = ~(layer4_out[5430] ^ layer4_out[5431]);
    assign layer5_out[5090] = ~(layer4_out[872] ^ layer4_out[873]);
    assign layer5_out[5091] = layer4_out[1858];
    assign layer5_out[5092] = ~layer4_out[1841];
    assign layer5_out[5093] = layer4_out[7666] ^ layer4_out[7667];
    assign layer5_out[5094] = ~(layer4_out[1752] | layer4_out[1753]);
    assign layer5_out[5095] = ~layer4_out[4955];
    assign layer5_out[5096] = ~layer4_out[7950];
    assign layer5_out[5097] = layer4_out[6998];
    assign layer5_out[5098] = layer4_out[6681] ^ layer4_out[6682];
    assign layer5_out[5099] = ~layer4_out[3898];
    assign layer5_out[5100] = ~layer4_out[1284];
    assign layer5_out[5101] = layer4_out[7051] & layer4_out[7052];
    assign layer5_out[5102] = layer4_out[464];
    assign layer5_out[5103] = ~(layer4_out[436] ^ layer4_out[437]);
    assign layer5_out[5104] = layer4_out[4789];
    assign layer5_out[5105] = layer4_out[1661] & ~layer4_out[1660];
    assign layer5_out[5106] = ~layer4_out[1999];
    assign layer5_out[5107] = layer4_out[4906];
    assign layer5_out[5108] = layer4_out[4164] ^ layer4_out[4165];
    assign layer5_out[5109] = ~layer4_out[7042];
    assign layer5_out[5110] = ~layer4_out[1555];
    assign layer5_out[5111] = ~(layer4_out[7526] ^ layer4_out[7527]);
    assign layer5_out[5112] = layer4_out[3543] ^ layer4_out[3544];
    assign layer5_out[5113] = ~layer4_out[3237];
    assign layer5_out[5114] = ~layer4_out[243];
    assign layer5_out[5115] = ~(layer4_out[3657] | layer4_out[3658]);
    assign layer5_out[5116] = ~(layer4_out[94] ^ layer4_out[95]);
    assign layer5_out[5117] = ~layer4_out[1935] | layer4_out[1934];
    assign layer5_out[5118] = layer4_out[7613];
    assign layer5_out[5119] = ~layer4_out[3374];
    assign layer5_out[5120] = ~layer4_out[7497];
    assign layer5_out[5121] = layer4_out[845] & ~layer4_out[844];
    assign layer5_out[5122] = layer4_out[2742];
    assign layer5_out[5123] = layer4_out[5181];
    assign layer5_out[5124] = layer4_out[4312];
    assign layer5_out[5125] = layer4_out[1620];
    assign layer5_out[5126] = ~(layer4_out[5925] ^ layer4_out[5926]);
    assign layer5_out[5127] = layer4_out[5442] ^ layer4_out[5443];
    assign layer5_out[5128] = ~layer4_out[3041] | layer4_out[3040];
    assign layer5_out[5129] = ~(layer4_out[19] | layer4_out[20]);
    assign layer5_out[5130] = layer4_out[7369];
    assign layer5_out[5131] = ~(layer4_out[1986] & layer4_out[1987]);
    assign layer5_out[5132] = layer4_out[3774] & layer4_out[3775];
    assign layer5_out[5133] = layer4_out[376];
    assign layer5_out[5134] = layer4_out[2223] ^ layer4_out[2224];
    assign layer5_out[5135] = layer4_out[6002];
    assign layer5_out[5136] = layer4_out[2118];
    assign layer5_out[5137] = layer4_out[866];
    assign layer5_out[5138] = layer4_out[4352] & layer4_out[4353];
    assign layer5_out[5139] = ~(layer4_out[5946] ^ layer4_out[5947]);
    assign layer5_out[5140] = layer4_out[4592] | layer4_out[4593];
    assign layer5_out[5141] = layer4_out[6750];
    assign layer5_out[5142] = layer4_out[5985] | layer4_out[5986];
    assign layer5_out[5143] = layer4_out[617] | layer4_out[618];
    assign layer5_out[5144] = layer4_out[1011] ^ layer4_out[1012];
    assign layer5_out[5145] = layer4_out[3498];
    assign layer5_out[5146] = layer4_out[2761];
    assign layer5_out[5147] = ~(layer4_out[6324] ^ layer4_out[6325]);
    assign layer5_out[5148] = layer4_out[85];
    assign layer5_out[5149] = layer4_out[296] & ~layer4_out[297];
    assign layer5_out[5150] = layer4_out[6867];
    assign layer5_out[5151] = ~(layer4_out[5919] ^ layer4_out[5920]);
    assign layer5_out[5152] = ~layer4_out[7560];
    assign layer5_out[5153] = ~(layer4_out[5230] ^ layer4_out[5231]);
    assign layer5_out[5154] = layer4_out[2499] & layer4_out[2500];
    assign layer5_out[5155] = ~layer4_out[2990];
    assign layer5_out[5156] = ~layer4_out[4580];
    assign layer5_out[5157] = ~layer4_out[6231];
    assign layer5_out[5158] = ~(layer4_out[368] ^ layer4_out[369]);
    assign layer5_out[5159] = layer4_out[809];
    assign layer5_out[5160] = layer4_out[7374] & ~layer4_out[7373];
    assign layer5_out[5161] = ~layer4_out[4699] | layer4_out[4698];
    assign layer5_out[5162] = layer4_out[7915];
    assign layer5_out[5163] = layer4_out[3776];
    assign layer5_out[5164] = layer4_out[2166];
    assign layer5_out[5165] = ~(layer4_out[4251] | layer4_out[4252]);
    assign layer5_out[5166] = layer4_out[4060];
    assign layer5_out[5167] = layer4_out[4450] ^ layer4_out[4451];
    assign layer5_out[5168] = ~(layer4_out[1788] ^ layer4_out[1789]);
    assign layer5_out[5169] = layer4_out[5934];
    assign layer5_out[5170] = layer4_out[5322] ^ layer4_out[5323];
    assign layer5_out[5171] = ~layer4_out[7184] | layer4_out[7185];
    assign layer5_out[5172] = layer4_out[4233] ^ layer4_out[4234];
    assign layer5_out[5173] = layer4_out[1719] & ~layer4_out[1720];
    assign layer5_out[5174] = ~(layer4_out[1404] & layer4_out[1405]);
    assign layer5_out[5175] = layer4_out[667];
    assign layer5_out[5176] = layer4_out[2271] ^ layer4_out[2272];
    assign layer5_out[5177] = layer4_out[6909];
    assign layer5_out[5178] = layer4_out[2787] & layer4_out[2788];
    assign layer5_out[5179] = ~(layer4_out[1987] & layer4_out[1988]);
    assign layer5_out[5180] = layer4_out[3653] & ~layer4_out[3652];
    assign layer5_out[5181] = layer4_out[65];
    assign layer5_out[5182] = layer4_out[2122] ^ layer4_out[2123];
    assign layer5_out[5183] = layer4_out[5991];
    assign layer5_out[5184] = ~(layer4_out[3379] | layer4_out[3380]);
    assign layer5_out[5185] = layer4_out[6019];
    assign layer5_out[5186] = ~(layer4_out[6056] & layer4_out[6057]);
    assign layer5_out[5187] = ~(layer4_out[1708] ^ layer4_out[1709]);
    assign layer5_out[5188] = ~layer4_out[6827];
    assign layer5_out[5189] = layer4_out[7121] & layer4_out[7122];
    assign layer5_out[5190] = layer4_out[3618];
    assign layer5_out[5191] = ~layer4_out[6440];
    assign layer5_out[5192] = layer4_out[5883] ^ layer4_out[5884];
    assign layer5_out[5193] = ~(layer4_out[150] | layer4_out[151]);
    assign layer5_out[5194] = ~layer4_out[6608];
    assign layer5_out[5195] = ~layer4_out[2202] | layer4_out[2201];
    assign layer5_out[5196] = ~layer4_out[6097];
    assign layer5_out[5197] = layer4_out[1211];
    assign layer5_out[5198] = layer4_out[6564];
    assign layer5_out[5199] = ~layer4_out[2256];
    assign layer5_out[5200] = ~(layer4_out[4498] & layer4_out[4499]);
    assign layer5_out[5201] = layer4_out[4970];
    assign layer5_out[5202] = ~layer4_out[3660];
    assign layer5_out[5203] = ~layer4_out[31];
    assign layer5_out[5204] = layer4_out[3764] & ~layer4_out[3763];
    assign layer5_out[5205] = ~layer4_out[843];
    assign layer5_out[5206] = layer4_out[6306] & layer4_out[6307];
    assign layer5_out[5207] = ~(layer4_out[7677] ^ layer4_out[7678]);
    assign layer5_out[5208] = ~(layer4_out[6251] ^ layer4_out[6252]);
    assign layer5_out[5209] = layer4_out[6220] ^ layer4_out[6221];
    assign layer5_out[5210] = ~layer4_out[4094] | layer4_out[4095];
    assign layer5_out[5211] = ~layer4_out[930];
    assign layer5_out[5212] = ~(layer4_out[4943] | layer4_out[4944]);
    assign layer5_out[5213] = ~layer4_out[830];
    assign layer5_out[5214] = layer4_out[6449] ^ layer4_out[6450];
    assign layer5_out[5215] = ~layer4_out[2233];
    assign layer5_out[5216] = ~layer4_out[7807];
    assign layer5_out[5217] = ~layer4_out[2261];
    assign layer5_out[5218] = ~(layer4_out[7369] ^ layer4_out[7370]);
    assign layer5_out[5219] = ~(layer4_out[4068] | layer4_out[4069]);
    assign layer5_out[5220] = layer4_out[7762] & layer4_out[7763];
    assign layer5_out[5221] = layer4_out[3978] & ~layer4_out[3979];
    assign layer5_out[5222] = layer4_out[7668] & ~layer4_out[7669];
    assign layer5_out[5223] = layer4_out[6934];
    assign layer5_out[5224] = layer4_out[3243] ^ layer4_out[3244];
    assign layer5_out[5225] = layer4_out[4655];
    assign layer5_out[5226] = ~layer4_out[5446];
    assign layer5_out[5227] = ~(layer4_out[7675] ^ layer4_out[7676]);
    assign layer5_out[5228] = ~(layer4_out[2774] | layer4_out[2775]);
    assign layer5_out[5229] = ~(layer4_out[4075] ^ layer4_out[4076]);
    assign layer5_out[5230] = ~(layer4_out[7299] ^ layer4_out[7300]);
    assign layer5_out[5231] = ~layer4_out[7245];
    assign layer5_out[5232] = ~layer4_out[7805];
    assign layer5_out[5233] = layer4_out[837] & ~layer4_out[836];
    assign layer5_out[5234] = ~layer4_out[3518];
    assign layer5_out[5235] = layer4_out[3247] ^ layer4_out[3248];
    assign layer5_out[5236] = layer4_out[4906];
    assign layer5_out[5237] = layer4_out[2486] & ~layer4_out[2487];
    assign layer5_out[5238] = ~(layer4_out[154] | layer4_out[155]);
    assign layer5_out[5239] = layer4_out[4292];
    assign layer5_out[5240] = ~(layer4_out[5998] & layer4_out[5999]);
    assign layer5_out[5241] = layer4_out[1107] ^ layer4_out[1108];
    assign layer5_out[5242] = layer4_out[7510];
    assign layer5_out[5243] = layer4_out[4819] ^ layer4_out[4820];
    assign layer5_out[5244] = ~layer4_out[5561];
    assign layer5_out[5245] = layer4_out[899];
    assign layer5_out[5246] = layer4_out[1834];
    assign layer5_out[5247] = layer4_out[3751];
    assign layer5_out[5248] = layer4_out[2983] & ~layer4_out[2984];
    assign layer5_out[5249] = layer4_out[4530] & ~layer4_out[4529];
    assign layer5_out[5250] = layer4_out[1142] | layer4_out[1143];
    assign layer5_out[5251] = layer4_out[2242];
    assign layer5_out[5252] = ~layer4_out[1966];
    assign layer5_out[5253] = ~(layer4_out[4567] ^ layer4_out[4568]);
    assign layer5_out[5254] = layer4_out[5709] & ~layer4_out[5710];
    assign layer5_out[5255] = ~(layer4_out[1302] ^ layer4_out[1303]);
    assign layer5_out[5256] = ~(layer4_out[8] | layer4_out[9]);
    assign layer5_out[5257] = layer4_out[69];
    assign layer5_out[5258] = ~layer4_out[1308] | layer4_out[1309];
    assign layer5_out[5259] = ~layer4_out[5603];
    assign layer5_out[5260] = ~layer4_out[2057];
    assign layer5_out[5261] = layer4_out[5524] & ~layer4_out[5525];
    assign layer5_out[5262] = ~(layer4_out[5117] | layer4_out[5118]);
    assign layer5_out[5263] = ~layer4_out[3293];
    assign layer5_out[5264] = layer4_out[194];
    assign layer5_out[5265] = ~(layer4_out[2896] | layer4_out[2897]);
    assign layer5_out[5266] = layer4_out[6467];
    assign layer5_out[5267] = layer4_out[2825] & layer4_out[2826];
    assign layer5_out[5268] = ~layer4_out[6926];
    assign layer5_out[5269] = ~(layer4_out[2836] ^ layer4_out[2837]);
    assign layer5_out[5270] = layer4_out[1186];
    assign layer5_out[5271] = layer4_out[2207] & ~layer4_out[2206];
    assign layer5_out[5272] = ~layer4_out[4893];
    assign layer5_out[5273] = layer4_out[1288];
    assign layer5_out[5274] = layer4_out[7115] & layer4_out[7116];
    assign layer5_out[5275] = ~(layer4_out[1045] ^ layer4_out[1046]);
    assign layer5_out[5276] = layer4_out[1648] ^ layer4_out[1649];
    assign layer5_out[5277] = layer4_out[5612];
    assign layer5_out[5278] = layer4_out[2794];
    assign layer5_out[5279] = layer4_out[7865] | layer4_out[7866];
    assign layer5_out[5280] = ~(layer4_out[2525] & layer4_out[2526]);
    assign layer5_out[5281] = layer4_out[1837];
    assign layer5_out[5282] = layer4_out[7069] | layer4_out[7070];
    assign layer5_out[5283] = ~layer4_out[3335] | layer4_out[3334];
    assign layer5_out[5284] = ~layer4_out[7438];
    assign layer5_out[5285] = ~(layer4_out[5353] & layer4_out[5354]);
    assign layer5_out[5286] = layer4_out[1144] & layer4_out[1145];
    assign layer5_out[5287] = ~layer4_out[4793];
    assign layer5_out[5288] = layer4_out[886] & ~layer4_out[887];
    assign layer5_out[5289] = layer4_out[2857] & ~layer4_out[2858];
    assign layer5_out[5290] = ~layer4_out[4357];
    assign layer5_out[5291] = layer4_out[1293];
    assign layer5_out[5292] = layer4_out[7830] ^ layer4_out[7831];
    assign layer5_out[5293] = layer4_out[3586] | layer4_out[3587];
    assign layer5_out[5294] = ~(layer4_out[4838] | layer4_out[4839]);
    assign layer5_out[5295] = layer4_out[2645] ^ layer4_out[2646];
    assign layer5_out[5296] = layer4_out[7470] & layer4_out[7471];
    assign layer5_out[5297] = layer4_out[3167] & layer4_out[3168];
    assign layer5_out[5298] = ~(layer4_out[3152] ^ layer4_out[3153]);
    assign layer5_out[5299] = ~layer4_out[4874];
    assign layer5_out[5300] = layer4_out[7633] & ~layer4_out[7632];
    assign layer5_out[5301] = ~layer4_out[5498];
    assign layer5_out[5302] = layer4_out[1068] ^ layer4_out[1069];
    assign layer5_out[5303] = layer4_out[4148] ^ layer4_out[4149];
    assign layer5_out[5304] = ~layer4_out[3726];
    assign layer5_out[5305] = layer4_out[5494] & layer4_out[5495];
    assign layer5_out[5306] = ~(layer4_out[2583] | layer4_out[2584]);
    assign layer5_out[5307] = layer4_out[1323];
    assign layer5_out[5308] = layer4_out[7686];
    assign layer5_out[5309] = ~layer4_out[4189];
    assign layer5_out[5310] = ~layer4_out[2263];
    assign layer5_out[5311] = layer4_out[6521];
    assign layer5_out[5312] = layer4_out[6286] & layer4_out[6287];
    assign layer5_out[5313] = layer4_out[2405] & layer4_out[2406];
    assign layer5_out[5314] = layer4_out[375] | layer4_out[376];
    assign layer5_out[5315] = ~(layer4_out[793] ^ layer4_out[794]);
    assign layer5_out[5316] = ~layer4_out[5338];
    assign layer5_out[5317] = layer4_out[6270] & ~layer4_out[6269];
    assign layer5_out[5318] = layer4_out[5725] ^ layer4_out[5726];
    assign layer5_out[5319] = ~layer4_out[275];
    assign layer5_out[5320] = layer4_out[1488] & ~layer4_out[1487];
    assign layer5_out[5321] = layer4_out[464];
    assign layer5_out[5322] = layer4_out[7130];
    assign layer5_out[5323] = layer4_out[178] ^ layer4_out[179];
    assign layer5_out[5324] = ~(layer4_out[3250] ^ layer4_out[3251]);
    assign layer5_out[5325] = layer4_out[4436] | layer4_out[4437];
    assign layer5_out[5326] = ~layer4_out[1773];
    assign layer5_out[5327] = ~layer4_out[3145];
    assign layer5_out[5328] = layer4_out[7425];
    assign layer5_out[5329] = layer4_out[6614] ^ layer4_out[6615];
    assign layer5_out[5330] = ~(layer4_out[2676] ^ layer4_out[2677]);
    assign layer5_out[5331] = layer4_out[7921];
    assign layer5_out[5332] = ~layer4_out[600] | layer4_out[601];
    assign layer5_out[5333] = layer4_out[2523] ^ layer4_out[2524];
    assign layer5_out[5334] = layer4_out[1363];
    assign layer5_out[5335] = layer4_out[6670] ^ layer4_out[6671];
    assign layer5_out[5336] = ~layer4_out[2229];
    assign layer5_out[5337] = layer4_out[6453] & layer4_out[6454];
    assign layer5_out[5338] = ~layer4_out[4081] | layer4_out[4080];
    assign layer5_out[5339] = ~(layer4_out[1427] ^ layer4_out[1428]);
    assign layer5_out[5340] = ~(layer4_out[1058] & layer4_out[1059]);
    assign layer5_out[5341] = ~layer4_out[1965];
    assign layer5_out[5342] = ~layer4_out[347] | layer4_out[346];
    assign layer5_out[5343] = ~(layer4_out[6534] ^ layer4_out[6535]);
    assign layer5_out[5344] = ~layer4_out[4447];
    assign layer5_out[5345] = layer4_out[5110] & ~layer4_out[5111];
    assign layer5_out[5346] = layer4_out[7682];
    assign layer5_out[5347] = ~layer4_out[1005];
    assign layer5_out[5348] = layer4_out[382] ^ layer4_out[383];
    assign layer5_out[5349] = ~layer4_out[939];
    assign layer5_out[5350] = layer4_out[5900];
    assign layer5_out[5351] = ~layer4_out[2038];
    assign layer5_out[5352] = layer4_out[5833];
    assign layer5_out[5353] = ~layer4_out[7118] | layer4_out[7117];
    assign layer5_out[5354] = ~layer4_out[3145] | layer4_out[3144];
    assign layer5_out[5355] = layer4_out[3946];
    assign layer5_out[5356] = layer4_out[218] & layer4_out[219];
    assign layer5_out[5357] = ~layer4_out[6844];
    assign layer5_out[5358] = ~layer4_out[836];
    assign layer5_out[5359] = layer4_out[2462] ^ layer4_out[2463];
    assign layer5_out[5360] = ~layer4_out[4609];
    assign layer5_out[5361] = ~layer4_out[5492];
    assign layer5_out[5362] = ~layer4_out[6708];
    assign layer5_out[5363] = ~(layer4_out[6850] & layer4_out[6851]);
    assign layer5_out[5364] = layer4_out[3946];
    assign layer5_out[5365] = layer4_out[98];
    assign layer5_out[5366] = layer4_out[3615];
    assign layer5_out[5367] = ~(layer4_out[5071] | layer4_out[5072]);
    assign layer5_out[5368] = ~layer4_out[6470];
    assign layer5_out[5369] = layer4_out[2102];
    assign layer5_out[5370] = layer4_out[846];
    assign layer5_out[5371] = ~(layer4_out[5600] & layer4_out[5601]);
    assign layer5_out[5372] = ~(layer4_out[118] & layer4_out[119]);
    assign layer5_out[5373] = layer4_out[5106];
    assign layer5_out[5374] = ~layer4_out[6446];
    assign layer5_out[5375] = layer4_out[5623];
    assign layer5_out[5376] = ~(layer4_out[1516] ^ layer4_out[1517]);
    assign layer5_out[5377] = ~layer4_out[6982];
    assign layer5_out[5378] = ~(layer4_out[2670] ^ layer4_out[2671]);
    assign layer5_out[5379] = ~(layer4_out[6201] | layer4_out[6202]);
    assign layer5_out[5380] = ~(layer4_out[2476] ^ layer4_out[2477]);
    assign layer5_out[5381] = layer4_out[7230] ^ layer4_out[7231];
    assign layer5_out[5382] = layer4_out[5562] ^ layer4_out[5563];
    assign layer5_out[5383] = layer4_out[6548] & ~layer4_out[6549];
    assign layer5_out[5384] = ~(layer4_out[2291] | layer4_out[2292]);
    assign layer5_out[5385] = layer4_out[2775] ^ layer4_out[2776];
    assign layer5_out[5386] = layer4_out[1224];
    assign layer5_out[5387] = ~layer4_out[2181];
    assign layer5_out[5388] = layer4_out[5753] & layer4_out[5754];
    assign layer5_out[5389] = layer4_out[2627] ^ layer4_out[2628];
    assign layer5_out[5390] = layer4_out[7607];
    assign layer5_out[5391] = layer4_out[1049] ^ layer4_out[1050];
    assign layer5_out[5392] = layer4_out[37];
    assign layer5_out[5393] = layer4_out[4744];
    assign layer5_out[5394] = layer4_out[5777];
    assign layer5_out[5395] = layer4_out[424];
    assign layer5_out[5396] = layer4_out[6595] & ~layer4_out[6594];
    assign layer5_out[5397] = ~(layer4_out[1151] ^ layer4_out[1152]);
    assign layer5_out[5398] = layer4_out[6431];
    assign layer5_out[5399] = ~layer4_out[6543];
    assign layer5_out[5400] = layer4_out[613] ^ layer4_out[614];
    assign layer5_out[5401] = ~layer4_out[1888];
    assign layer5_out[5402] = layer4_out[4050];
    assign layer5_out[5403] = layer4_out[7408];
    assign layer5_out[5404] = ~layer4_out[5416] | layer4_out[5415];
    assign layer5_out[5405] = layer4_out[4913];
    assign layer5_out[5406] = layer4_out[3588];
    assign layer5_out[5407] = layer4_out[3934];
    assign layer5_out[5408] = ~layer4_out[2894] | layer4_out[2895];
    assign layer5_out[5409] = layer4_out[996];
    assign layer5_out[5410] = ~layer4_out[3101];
    assign layer5_out[5411] = ~(layer4_out[6402] ^ layer4_out[6403]);
    assign layer5_out[5412] = layer4_out[3050];
    assign layer5_out[5413] = ~layer4_out[678];
    assign layer5_out[5414] = layer4_out[4038];
    assign layer5_out[5415] = layer4_out[7386] & layer4_out[7387];
    assign layer5_out[5416] = ~layer4_out[6605] | layer4_out[6606];
    assign layer5_out[5417] = layer4_out[5662];
    assign layer5_out[5418] = ~layer4_out[2053];
    assign layer5_out[5419] = layer4_out[5965];
    assign layer5_out[5420] = layer4_out[5159];
    assign layer5_out[5421] = layer4_out[3290];
    assign layer5_out[5422] = ~layer4_out[4037];
    assign layer5_out[5423] = layer4_out[4519];
    assign layer5_out[5424] = layer4_out[3961] ^ layer4_out[3962];
    assign layer5_out[5425] = layer4_out[3733];
    assign layer5_out[5426] = ~layer4_out[2850] | layer4_out[2849];
    assign layer5_out[5427] = ~layer4_out[6379];
    assign layer5_out[5428] = ~(layer4_out[1756] ^ layer4_out[1757]);
    assign layer5_out[5429] = layer4_out[420] ^ layer4_out[421];
    assign layer5_out[5430] = layer4_out[5276];
    assign layer5_out[5431] = ~layer4_out[257];
    assign layer5_out[5432] = ~layer4_out[5490];
    assign layer5_out[5433] = layer4_out[7281];
    assign layer5_out[5434] = layer4_out[4658] & ~layer4_out[4657];
    assign layer5_out[5435] = layer4_out[4831] & ~layer4_out[4830];
    assign layer5_out[5436] = layer4_out[6034];
    assign layer5_out[5437] = layer4_out[6924];
    assign layer5_out[5438] = layer4_out[3727] & ~layer4_out[3728];
    assign layer5_out[5439] = layer4_out[481];
    assign layer5_out[5440] = ~layer4_out[3389];
    assign layer5_out[5441] = layer4_out[5055];
    assign layer5_out[5442] = ~(layer4_out[3454] | layer4_out[3455]);
    assign layer5_out[5443] = ~layer4_out[3198];
    assign layer5_out[5444] = layer4_out[1312] ^ layer4_out[1313];
    assign layer5_out[5445] = layer4_out[6358];
    assign layer5_out[5446] = layer4_out[923] ^ layer4_out[924];
    assign layer5_out[5447] = ~layer4_out[6752];
    assign layer5_out[5448] = ~(layer4_out[2958] | layer4_out[2959]);
    assign layer5_out[5449] = layer4_out[4882];
    assign layer5_out[5450] = layer4_out[2551] & ~layer4_out[2552];
    assign layer5_out[5451] = ~(layer4_out[364] | layer4_out[365]);
    assign layer5_out[5452] = layer4_out[637] | layer4_out[638];
    assign layer5_out[5453] = ~(layer4_out[1984] | layer4_out[1985]);
    assign layer5_out[5454] = ~(layer4_out[2014] ^ layer4_out[2015]);
    assign layer5_out[5455] = layer4_out[7991] ^ layer4_out[7992];
    assign layer5_out[5456] = ~layer4_out[4127] | layer4_out[4128];
    assign layer5_out[5457] = layer4_out[363];
    assign layer5_out[5458] = ~layer4_out[4291];
    assign layer5_out[5459] = ~layer4_out[5344];
    assign layer5_out[5460] = layer4_out[3035];
    assign layer5_out[5461] = layer4_out[4415];
    assign layer5_out[5462] = ~layer4_out[312] | layer4_out[311];
    assign layer5_out[5463] = ~(layer4_out[1265] | layer4_out[1266]);
    assign layer5_out[5464] = layer4_out[2339] ^ layer4_out[2340];
    assign layer5_out[5465] = ~(layer4_out[1614] & layer4_out[1615]);
    assign layer5_out[5466] = ~(layer4_out[4149] & layer4_out[4150]);
    assign layer5_out[5467] = ~(layer4_out[843] ^ layer4_out[844]);
    assign layer5_out[5468] = ~layer4_out[5319] | layer4_out[5318];
    assign layer5_out[5469] = ~layer4_out[6718];
    assign layer5_out[5470] = layer4_out[2959] ^ layer4_out[2960];
    assign layer5_out[5471] = ~layer4_out[7264];
    assign layer5_out[5472] = ~(layer4_out[744] & layer4_out[745]);
    assign layer5_out[5473] = ~layer4_out[3393] | layer4_out[3394];
    assign layer5_out[5474] = layer4_out[3223] ^ layer4_out[3224];
    assign layer5_out[5475] = ~(layer4_out[2247] ^ layer4_out[2248]);
    assign layer5_out[5476] = layer4_out[3245];
    assign layer5_out[5477] = layer4_out[4317] & ~layer4_out[4316];
    assign layer5_out[5478] = ~layer4_out[4391];
    assign layer5_out[5479] = layer4_out[40];
    assign layer5_out[5480] = layer4_out[1134] | layer4_out[1135];
    assign layer5_out[5481] = ~layer4_out[4258] | layer4_out[4257];
    assign layer5_out[5482] = layer4_out[2669] & ~layer4_out[2670];
    assign layer5_out[5483] = layer4_out[6105];
    assign layer5_out[5484] = ~layer4_out[5599];
    assign layer5_out[5485] = layer4_out[4403];
    assign layer5_out[5486] = layer4_out[6424] ^ layer4_out[6425];
    assign layer5_out[5487] = layer4_out[3770];
    assign layer5_out[5488] = layer4_out[4842] | layer4_out[4843];
    assign layer5_out[5489] = ~layer4_out[6303];
    assign layer5_out[5490] = layer4_out[6200] ^ layer4_out[6201];
    assign layer5_out[5491] = ~layer4_out[2860];
    assign layer5_out[5492] = ~(layer4_out[6020] | layer4_out[6021]);
    assign layer5_out[5493] = ~layer4_out[6150] | layer4_out[6149];
    assign layer5_out[5494] = ~(layer4_out[5743] ^ layer4_out[5744]);
    assign layer5_out[5495] = layer4_out[1379] | layer4_out[1380];
    assign layer5_out[5496] = layer4_out[5523];
    assign layer5_out[5497] = ~(layer4_out[2193] | layer4_out[2194]);
    assign layer5_out[5498] = ~(layer4_out[3898] | layer4_out[3899]);
    assign layer5_out[5499] = layer4_out[3791];
    assign layer5_out[5500] = layer4_out[6105] & ~layer4_out[6106];
    assign layer5_out[5501] = ~layer4_out[962];
    assign layer5_out[5502] = ~layer4_out[1494];
    assign layer5_out[5503] = layer4_out[7968] & ~layer4_out[7967];
    assign layer5_out[5504] = layer4_out[636] | layer4_out[637];
    assign layer5_out[5505] = layer4_out[652] ^ layer4_out[653];
    assign layer5_out[5506] = layer4_out[1994] & ~layer4_out[1993];
    assign layer5_out[5507] = layer4_out[2315];
    assign layer5_out[5508] = layer4_out[2632] & ~layer4_out[2631];
    assign layer5_out[5509] = ~(layer4_out[4850] ^ layer4_out[4851]);
    assign layer5_out[5510] = ~(layer4_out[5363] ^ layer4_out[5364]);
    assign layer5_out[5511] = ~layer4_out[5779];
    assign layer5_out[5512] = layer4_out[561];
    assign layer5_out[5513] = layer4_out[7671];
    assign layer5_out[5514] = ~layer4_out[4853] | layer4_out[4852];
    assign layer5_out[5515] = layer4_out[6910] ^ layer4_out[6911];
    assign layer5_out[5516] = ~(layer4_out[4313] ^ layer4_out[4314]);
    assign layer5_out[5517] = layer4_out[3282] ^ layer4_out[3283];
    assign layer5_out[5518] = layer4_out[705] & ~layer4_out[706];
    assign layer5_out[5519] = layer4_out[7847] ^ layer4_out[7848];
    assign layer5_out[5520] = ~layer4_out[357];
    assign layer5_out[5521] = layer4_out[2099] & ~layer4_out[2098];
    assign layer5_out[5522] = ~layer4_out[6603];
    assign layer5_out[5523] = layer4_out[2259];
    assign layer5_out[5524] = ~layer4_out[5936];
    assign layer5_out[5525] = ~(layer4_out[2391] ^ layer4_out[2392]);
    assign layer5_out[5526] = layer4_out[1673] & ~layer4_out[1674];
    assign layer5_out[5527] = layer4_out[4308] & ~layer4_out[4307];
    assign layer5_out[5528] = ~(layer4_out[5842] ^ layer4_out[5843]);
    assign layer5_out[5529] = layer4_out[7673] ^ layer4_out[7674];
    assign layer5_out[5530] = ~layer4_out[4960];
    assign layer5_out[5531] = layer4_out[4458];
    assign layer5_out[5532] = layer4_out[377] & layer4_out[378];
    assign layer5_out[5533] = layer4_out[78] ^ layer4_out[79];
    assign layer5_out[5534] = ~(layer4_out[3882] & layer4_out[3883]);
    assign layer5_out[5535] = layer4_out[2956] & ~layer4_out[2957];
    assign layer5_out[5536] = layer4_out[2146] ^ layer4_out[2147];
    assign layer5_out[5537] = ~(layer4_out[5619] & layer4_out[5620]);
    assign layer5_out[5538] = ~(layer4_out[7266] ^ layer4_out[7267]);
    assign layer5_out[5539] = layer4_out[4786] & layer4_out[4787];
    assign layer5_out[5540] = layer4_out[128];
    assign layer5_out[5541] = layer4_out[702];
    assign layer5_out[5542] = layer4_out[2169] & ~layer4_out[2170];
    assign layer5_out[5543] = ~layer4_out[2509];
    assign layer5_out[5544] = ~(layer4_out[7900] | layer4_out[7901]);
    assign layer5_out[5545] = ~(layer4_out[5268] ^ layer4_out[5269]);
    assign layer5_out[5546] = layer4_out[6991] & layer4_out[6992];
    assign layer5_out[5547] = ~layer4_out[6238];
    assign layer5_out[5548] = ~layer4_out[2979];
    assign layer5_out[5549] = layer4_out[72];
    assign layer5_out[5550] = ~layer4_out[3505];
    assign layer5_out[5551] = layer4_out[5011];
    assign layer5_out[5552] = ~layer4_out[7851];
    assign layer5_out[5553] = ~layer4_out[4127];
    assign layer5_out[5554] = layer4_out[1437];
    assign layer5_out[5555] = layer4_out[6212];
    assign layer5_out[5556] = ~(layer4_out[2148] & layer4_out[2149]);
    assign layer5_out[5557] = ~layer4_out[6961];
    assign layer5_out[5558] = ~(layer4_out[5410] | layer4_out[5411]);
    assign layer5_out[5559] = layer4_out[3756] ^ layer4_out[3757];
    assign layer5_out[5560] = layer4_out[2904];
    assign layer5_out[5561] = layer4_out[6175];
    assign layer5_out[5562] = ~(layer4_out[773] ^ layer4_out[774]);
    assign layer5_out[5563] = layer4_out[3535] & ~layer4_out[3536];
    assign layer5_out[5564] = layer4_out[3091];
    assign layer5_out[5565] = layer4_out[4100];
    assign layer5_out[5566] = layer4_out[130] & layer4_out[131];
    assign layer5_out[5567] = layer4_out[2570] | layer4_out[2571];
    assign layer5_out[5568] = layer4_out[6816] | layer4_out[6817];
    assign layer5_out[5569] = layer4_out[3332];
    assign layer5_out[5570] = layer4_out[527] | layer4_out[528];
    assign layer5_out[5571] = ~(layer4_out[7495] & layer4_out[7496]);
    assign layer5_out[5572] = layer4_out[7046];
    assign layer5_out[5573] = layer4_out[7338] & ~layer4_out[7337];
    assign layer5_out[5574] = ~layer4_out[3401] | layer4_out[3402];
    assign layer5_out[5575] = layer4_out[2761];
    assign layer5_out[5576] = ~(layer4_out[3233] ^ layer4_out[3234]);
    assign layer5_out[5577] = layer4_out[3187];
    assign layer5_out[5578] = ~layer4_out[2415];
    assign layer5_out[5579] = ~layer4_out[3124];
    assign layer5_out[5580] = layer4_out[7323] & ~layer4_out[7322];
    assign layer5_out[5581] = ~layer4_out[7948] | layer4_out[7949];
    assign layer5_out[5582] = ~layer4_out[3871];
    assign layer5_out[5583] = ~layer4_out[1926];
    assign layer5_out[5584] = layer4_out[6967];
    assign layer5_out[5585] = layer4_out[6362];
    assign layer5_out[5586] = ~(layer4_out[3820] ^ layer4_out[3821]);
    assign layer5_out[5587] = layer4_out[7582] & ~layer4_out[7581];
    assign layer5_out[5588] = layer4_out[2866];
    assign layer5_out[5589] = ~layer4_out[1396];
    assign layer5_out[5590] = layer4_out[7693];
    assign layer5_out[5591] = layer4_out[6061] & ~layer4_out[6060];
    assign layer5_out[5592] = layer4_out[4254] & ~layer4_out[4253];
    assign layer5_out[5593] = layer4_out[82];
    assign layer5_out[5594] = layer4_out[6412] & ~layer4_out[6411];
    assign layer5_out[5595] = ~layer4_out[3612];
    assign layer5_out[5596] = layer4_out[5688] ^ layer4_out[5689];
    assign layer5_out[5597] = layer4_out[6384] & ~layer4_out[6385];
    assign layer5_out[5598] = ~layer4_out[3583];
    assign layer5_out[5599] = layer4_out[6838];
    assign layer5_out[5600] = ~layer4_out[4651] | layer4_out[4652];
    assign layer5_out[5601] = ~layer4_out[6310];
    assign layer5_out[5602] = layer4_out[7706] ^ layer4_out[7707];
    assign layer5_out[5603] = ~layer4_out[4091];
    assign layer5_out[5604] = layer4_out[2796] & ~layer4_out[2797];
    assign layer5_out[5605] = layer4_out[6759];
    assign layer5_out[5606] = layer4_out[1347] | layer4_out[1348];
    assign layer5_out[5607] = layer4_out[4266] ^ layer4_out[4267];
    assign layer5_out[5608] = ~(layer4_out[6667] & layer4_out[6668]);
    assign layer5_out[5609] = ~(layer4_out[2813] ^ layer4_out[2814]);
    assign layer5_out[5610] = layer4_out[542] & ~layer4_out[543];
    assign layer5_out[5611] = ~(layer4_out[1681] | layer4_out[1682]);
    assign layer5_out[5612] = layer4_out[4926] & layer4_out[4927];
    assign layer5_out[5613] = ~layer4_out[1096];
    assign layer5_out[5614] = ~layer4_out[3616];
    assign layer5_out[5615] = layer4_out[6464] ^ layer4_out[6465];
    assign layer5_out[5616] = layer4_out[3958] | layer4_out[3959];
    assign layer5_out[5617] = layer4_out[5370];
    assign layer5_out[5618] = layer4_out[6918] | layer4_out[6919];
    assign layer5_out[5619] = ~(layer4_out[7891] ^ layer4_out[7892]);
    assign layer5_out[5620] = ~layer4_out[6925];
    assign layer5_out[5621] = ~(layer4_out[4668] & layer4_out[4669]);
    assign layer5_out[5622] = ~layer4_out[5440];
    assign layer5_out[5623] = layer4_out[1839] & ~layer4_out[1838];
    assign layer5_out[5624] = ~layer4_out[5073];
    assign layer5_out[5625] = ~(layer4_out[1139] | layer4_out[1140]);
    assign layer5_out[5626] = layer4_out[4898] | layer4_out[4899];
    assign layer5_out[5627] = ~layer4_out[7840];
    assign layer5_out[5628] = layer4_out[6946] ^ layer4_out[6947];
    assign layer5_out[5629] = layer4_out[6819] & ~layer4_out[6820];
    assign layer5_out[5630] = ~layer4_out[91] | layer4_out[92];
    assign layer5_out[5631] = layer4_out[4895] & ~layer4_out[4896];
    assign layer5_out[5632] = layer4_out[6730] & layer4_out[6731];
    assign layer5_out[5633] = layer4_out[6794] ^ layer4_out[6795];
    assign layer5_out[5634] = ~layer4_out[319] | layer4_out[320];
    assign layer5_out[5635] = layer4_out[2488] & layer4_out[2489];
    assign layer5_out[5636] = layer4_out[5548] | layer4_out[5549];
    assign layer5_out[5637] = layer4_out[5449] & ~layer4_out[5448];
    assign layer5_out[5638] = ~(layer4_out[5888] ^ layer4_out[5889]);
    assign layer5_out[5639] = ~layer4_out[2474];
    assign layer5_out[5640] = layer4_out[6115] & ~layer4_out[6116];
    assign layer5_out[5641] = layer4_out[7611] | layer4_out[7612];
    assign layer5_out[5642] = ~(layer4_out[7817] & layer4_out[7818]);
    assign layer5_out[5643] = layer4_out[4574] & ~layer4_out[4575];
    assign layer5_out[5644] = ~(layer4_out[5632] ^ layer4_out[5633]);
    assign layer5_out[5645] = layer4_out[270];
    assign layer5_out[5646] = layer4_out[1952];
    assign layer5_out[5647] = layer4_out[3971] | layer4_out[3972];
    assign layer5_out[5648] = layer4_out[7937] ^ layer4_out[7938];
    assign layer5_out[5649] = layer4_out[7836];
    assign layer5_out[5650] = layer4_out[3981];
    assign layer5_out[5651] = layer4_out[4544] ^ layer4_out[4545];
    assign layer5_out[5652] = ~layer4_out[6768];
    assign layer5_out[5653] = layer4_out[7062] | layer4_out[7063];
    assign layer5_out[5654] = layer4_out[6625];
    assign layer5_out[5655] = layer4_out[5690];
    assign layer5_out[5656] = ~(layer4_out[4009] ^ layer4_out[4010]);
    assign layer5_out[5657] = layer4_out[871];
    assign layer5_out[5658] = ~layer4_out[4824] | layer4_out[4823];
    assign layer5_out[5659] = ~layer4_out[2690];
    assign layer5_out[5660] = layer4_out[6205] & layer4_out[6206];
    assign layer5_out[5661] = layer4_out[5014] ^ layer4_out[5015];
    assign layer5_out[5662] = layer4_out[1406] & ~layer4_out[1407];
    assign layer5_out[5663] = layer4_out[3429];
    assign layer5_out[5664] = layer4_out[7167];
    assign layer5_out[5665] = layer4_out[7536];
    assign layer5_out[5666] = layer4_out[104];
    assign layer5_out[5667] = ~layer4_out[4376];
    assign layer5_out[5668] = layer4_out[2086];
    assign layer5_out[5669] = layer4_out[6647];
    assign layer5_out[5670] = ~layer4_out[3040];
    assign layer5_out[5671] = ~layer4_out[2745] | layer4_out[2744];
    assign layer5_out[5672] = ~layer4_out[5721];
    assign layer5_out[5673] = ~layer4_out[7169];
    assign layer5_out[5674] = layer4_out[3802] | layer4_out[3803];
    assign layer5_out[5675] = ~layer4_out[1790] | layer4_out[1789];
    assign layer5_out[5676] = layer4_out[4898];
    assign layer5_out[5677] = layer4_out[7624] ^ layer4_out[7625];
    assign layer5_out[5678] = layer4_out[2124] ^ layer4_out[2125];
    assign layer5_out[5679] = layer4_out[1721];
    assign layer5_out[5680] = ~(layer4_out[4705] & layer4_out[4706]);
    assign layer5_out[5681] = layer4_out[514];
    assign layer5_out[5682] = ~(layer4_out[7385] ^ layer4_out[7386]);
    assign layer5_out[5683] = ~layer4_out[6767] | layer4_out[6766];
    assign layer5_out[5684] = layer4_out[4212] ^ layer4_out[4213];
    assign layer5_out[5685] = layer4_out[1822] ^ layer4_out[1823];
    assign layer5_out[5686] = ~(layer4_out[4369] ^ layer4_out[4370]);
    assign layer5_out[5687] = layer4_out[6876] ^ layer4_out[6877];
    assign layer5_out[5688] = ~layer4_out[5291];
    assign layer5_out[5689] = layer4_out[4226] & ~layer4_out[4227];
    assign layer5_out[5690] = ~(layer4_out[4097] & layer4_out[4098]);
    assign layer5_out[5691] = ~(layer4_out[4896] ^ layer4_out[4897]);
    assign layer5_out[5692] = layer4_out[990];
    assign layer5_out[5693] = ~layer4_out[2232];
    assign layer5_out[5694] = layer4_out[1890];
    assign layer5_out[5695] = layer4_out[5457];
    assign layer5_out[5696] = layer4_out[1375] ^ layer4_out[1376];
    assign layer5_out[5697] = ~layer4_out[6170];
    assign layer5_out[5698] = ~layer4_out[7912];
    assign layer5_out[5699] = layer4_out[3609] & ~layer4_out[3608];
    assign layer5_out[5700] = layer4_out[2612];
    assign layer5_out[5701] = layer4_out[7854];
    assign layer5_out[5702] = layer4_out[7218] & ~layer4_out[7217];
    assign layer5_out[5703] = ~(layer4_out[4446] ^ layer4_out[4447]);
    assign layer5_out[5704] = layer4_out[3917];
    assign layer5_out[5705] = layer4_out[3202];
    assign layer5_out[5706] = ~(layer4_out[548] ^ layer4_out[549]);
    assign layer5_out[5707] = ~layer4_out[5721];
    assign layer5_out[5708] = ~layer4_out[1006] | layer4_out[1005];
    assign layer5_out[5709] = ~layer4_out[6747];
    assign layer5_out[5710] = ~layer4_out[2484];
    assign layer5_out[5711] = layer4_out[5324] | layer4_out[5325];
    assign layer5_out[5712] = ~layer4_out[5181];
    assign layer5_out[5713] = layer4_out[3135] & layer4_out[3136];
    assign layer5_out[5714] = ~(layer4_out[1362] | layer4_out[1363]);
    assign layer5_out[5715] = layer4_out[7474] | layer4_out[7475];
    assign layer5_out[5716] = layer4_out[111];
    assign layer5_out[5717] = layer4_out[3724] ^ layer4_out[3725];
    assign layer5_out[5718] = ~layer4_out[3913];
    assign layer5_out[5719] = layer4_out[781];
    assign layer5_out[5720] = ~layer4_out[4288];
    assign layer5_out[5721] = layer4_out[567];
    assign layer5_out[5722] = ~(layer4_out[5800] & layer4_out[5801]);
    assign layer5_out[5723] = layer4_out[4374] & ~layer4_out[4375];
    assign layer5_out[5724] = layer4_out[5187] | layer4_out[5188];
    assign layer5_out[5725] = ~(layer4_out[7108] | layer4_out[7109]);
    assign layer5_out[5726] = ~layer4_out[7272] | layer4_out[7273];
    assign layer5_out[5727] = ~(layer4_out[6354] ^ layer4_out[6355]);
    assign layer5_out[5728] = ~(layer4_out[4395] ^ layer4_out[4396]);
    assign layer5_out[5729] = ~layer4_out[2673];
    assign layer5_out[5730] = ~(layer4_out[4695] | layer4_out[4696]);
    assign layer5_out[5731] = ~(layer4_out[4415] ^ layer4_out[4416]);
    assign layer5_out[5732] = ~layer4_out[2436];
    assign layer5_out[5733] = ~(layer4_out[564] & layer4_out[565]);
    assign layer5_out[5734] = layer4_out[3445] ^ layer4_out[3446];
    assign layer5_out[5735] = layer4_out[511];
    assign layer5_out[5736] = layer4_out[276] & layer4_out[277];
    assign layer5_out[5737] = layer4_out[2609] ^ layer4_out[2610];
    assign layer5_out[5738] = layer4_out[251];
    assign layer5_out[5739] = layer4_out[4630];
    assign layer5_out[5740] = ~(layer4_out[4828] ^ layer4_out[4829]);
    assign layer5_out[5741] = ~layer4_out[5474] | layer4_out[5473];
    assign layer5_out[5742] = ~layer4_out[1403];
    assign layer5_out[5743] = layer4_out[2156] | layer4_out[2157];
    assign layer5_out[5744] = layer4_out[2962];
    assign layer5_out[5745] = layer4_out[4230];
    assign layer5_out[5746] = layer4_out[3198] & ~layer4_out[3197];
    assign layer5_out[5747] = layer4_out[2691];
    assign layer5_out[5748] = layer4_out[1181];
    assign layer5_out[5749] = layer4_out[3830] ^ layer4_out[3831];
    assign layer5_out[5750] = ~layer4_out[1556];
    assign layer5_out[5751] = ~(layer4_out[2524] ^ layer4_out[2525]);
    assign layer5_out[5752] = layer4_out[3680];
    assign layer5_out[5753] = ~layer4_out[7135];
    assign layer5_out[5754] = layer4_out[120] & layer4_out[121];
    assign layer5_out[5755] = ~(layer4_out[7073] ^ layer4_out[7074]);
    assign layer5_out[5756] = layer4_out[5763];
    assign layer5_out[5757] = layer4_out[5345];
    assign layer5_out[5758] = ~layer4_out[2186];
    assign layer5_out[5759] = layer4_out[2047] | layer4_out[2048];
    assign layer5_out[5760] = ~(layer4_out[743] ^ layer4_out[744]);
    assign layer5_out[5761] = layer4_out[5401];
    assign layer5_out[5762] = ~layer4_out[5350] | layer4_out[5349];
    assign layer5_out[5763] = ~layer4_out[503];
    assign layer5_out[5764] = ~(layer4_out[5536] | layer4_out[5537]);
    assign layer5_out[5765] = ~layer4_out[3061];
    assign layer5_out[5766] = ~layer4_out[7748];
    assign layer5_out[5767] = layer4_out[300] & layer4_out[301];
    assign layer5_out[5768] = layer4_out[2112];
    assign layer5_out[5769] = layer4_out[1625];
    assign layer5_out[5770] = layer4_out[1969] ^ layer4_out[1970];
    assign layer5_out[5771] = layer4_out[3839] ^ layer4_out[3840];
    assign layer5_out[5772] = ~layer4_out[3238];
    assign layer5_out[5773] = layer4_out[5403];
    assign layer5_out[5774] = ~(layer4_out[1050] | layer4_out[1051]);
    assign layer5_out[5775] = ~(layer4_out[3692] | layer4_out[3693]);
    assign layer5_out[5776] = ~layer4_out[1431];
    assign layer5_out[5777] = layer4_out[950];
    assign layer5_out[5778] = layer4_out[4707] & ~layer4_out[4706];
    assign layer5_out[5779] = layer4_out[1457];
    assign layer5_out[5780] = ~layer4_out[4403];
    assign layer5_out[5781] = layer4_out[1823] ^ layer4_out[1824];
    assign layer5_out[5782] = layer4_out[2597] & ~layer4_out[2596];
    assign layer5_out[5783] = ~(layer4_out[5012] | layer4_out[5013]);
    assign layer5_out[5784] = layer4_out[7295];
    assign layer5_out[5785] = ~layer4_out[5732];
    assign layer5_out[5786] = ~(layer4_out[1885] ^ layer4_out[1886]);
    assign layer5_out[5787] = ~(layer4_out[1627] ^ layer4_out[1628]);
    assign layer5_out[5788] = layer4_out[7246] ^ layer4_out[7247];
    assign layer5_out[5789] = ~layer4_out[5092];
    assign layer5_out[5790] = layer4_out[5406] ^ layer4_out[5407];
    assign layer5_out[5791] = ~layer4_out[1423] | layer4_out[1424];
    assign layer5_out[5792] = layer4_out[4051];
    assign layer5_out[5793] = layer4_out[1522];
    assign layer5_out[5794] = ~layer4_out[2343] | layer4_out[2342];
    assign layer5_out[5795] = layer4_out[5134] & ~layer4_out[5133];
    assign layer5_out[5796] = ~layer4_out[2502];
    assign layer5_out[5797] = layer4_out[315] ^ layer4_out[316];
    assign layer5_out[5798] = ~layer4_out[5171] | layer4_out[5172];
    assign layer5_out[5799] = ~layer4_out[1442];
    assign layer5_out[5800] = ~layer4_out[3813];
    assign layer5_out[5801] = layer4_out[3442] & ~layer4_out[3443];
    assign layer5_out[5802] = ~(layer4_out[1443] & layer4_out[1444]);
    assign layer5_out[5803] = layer4_out[4077];
    assign layer5_out[5804] = layer4_out[1170] & ~layer4_out[1171];
    assign layer5_out[5805] = layer4_out[3141] & layer4_out[3142];
    assign layer5_out[5806] = layer4_out[3455];
    assign layer5_out[5807] = layer4_out[553];
    assign layer5_out[5808] = ~layer4_out[6245];
    assign layer5_out[5809] = layer4_out[715];
    assign layer5_out[5810] = ~layer4_out[6339] | layer4_out[6340];
    assign layer5_out[5811] = ~(layer4_out[4552] | layer4_out[4553]);
    assign layer5_out[5812] = ~layer4_out[1242] | layer4_out[1243];
    assign layer5_out[5813] = ~(layer4_out[6337] ^ layer4_out[6338]);
    assign layer5_out[5814] = layer4_out[4868];
    assign layer5_out[5815] = layer4_out[7644] & layer4_out[7645];
    assign layer5_out[5816] = layer4_out[6571] ^ layer4_out[6572];
    assign layer5_out[5817] = layer4_out[7699];
    assign layer5_out[5818] = ~(layer4_out[6894] & layer4_out[6895]);
    assign layer5_out[5819] = layer4_out[4792] | layer4_out[4793];
    assign layer5_out[5820] = ~layer4_out[6460] | layer4_out[6461];
    assign layer5_out[5821] = ~(layer4_out[4093] | layer4_out[4094]);
    assign layer5_out[5822] = layer4_out[7672];
    assign layer5_out[5823] = layer4_out[15] | layer4_out[16];
    assign layer5_out[5824] = layer4_out[5973] & ~layer4_out[5974];
    assign layer5_out[5825] = ~(layer4_out[1832] ^ layer4_out[1833]);
    assign layer5_out[5826] = ~layer4_out[5128];
    assign layer5_out[5827] = layer4_out[7088] ^ layer4_out[7089];
    assign layer5_out[5828] = layer4_out[5747];
    assign layer5_out[5829] = ~layer4_out[883] | layer4_out[884];
    assign layer5_out[5830] = layer4_out[4489];
    assign layer5_out[5831] = ~layer4_out[3543];
    assign layer5_out[5832] = layer4_out[7821];
    assign layer5_out[5833] = layer4_out[140] ^ layer4_out[141];
    assign layer5_out[5834] = layer4_out[1911] ^ layer4_out[1912];
    assign layer5_out[5835] = ~layer4_out[2117] | layer4_out[2116];
    assign layer5_out[5836] = ~layer4_out[4027];
    assign layer5_out[5837] = ~(layer4_out[1380] ^ layer4_out[1381]);
    assign layer5_out[5838] = layer4_out[5390];
    assign layer5_out[5839] = layer4_out[3138] & layer4_out[3139];
    assign layer5_out[5840] = layer4_out[5607] & layer4_out[5608];
    assign layer5_out[5841] = ~layer4_out[3556];
    assign layer5_out[5842] = ~layer4_out[5294];
    assign layer5_out[5843] = layer4_out[2910] ^ layer4_out[2911];
    assign layer5_out[5844] = ~(layer4_out[7834] | layer4_out[7835]);
    assign layer5_out[5845] = ~layer4_out[4942];
    assign layer5_out[5846] = layer4_out[3441] | layer4_out[3442];
    assign layer5_out[5847] = ~(layer4_out[5374] ^ layer4_out[5375]);
    assign layer5_out[5848] = ~(layer4_out[5642] & layer4_out[5643]);
    assign layer5_out[5849] = layer4_out[4900];
    assign layer5_out[5850] = layer4_out[5852] & layer4_out[5853];
    assign layer5_out[5851] = layer4_out[429];
    assign layer5_out[5852] = layer4_out[1940];
    assign layer5_out[5853] = ~(layer4_out[5582] | layer4_out[5583]);
    assign layer5_out[5854] = ~(layer4_out[3327] & layer4_out[3328]);
    assign layer5_out[5855] = layer4_out[688];
    assign layer5_out[5856] = layer4_out[199] & layer4_out[200];
    assign layer5_out[5857] = layer4_out[3707] & layer4_out[3708];
    assign layer5_out[5858] = layer4_out[3664];
    assign layer5_out[5859] = layer4_out[4961] ^ layer4_out[4962];
    assign layer5_out[5860] = layer4_out[7882] | layer4_out[7883];
    assign layer5_out[5861] = layer4_out[6975] & layer4_out[6976];
    assign layer5_out[5862] = ~layer4_out[1812];
    assign layer5_out[5863] = layer4_out[7856];
    assign layer5_out[5864] = ~layer4_out[6122] | layer4_out[6123];
    assign layer5_out[5865] = layer4_out[2754] & ~layer4_out[2753];
    assign layer5_out[5866] = layer4_out[5356];
    assign layer5_out[5867] = layer4_out[2624] & ~layer4_out[2623];
    assign layer5_out[5868] = layer4_out[5266] | layer4_out[5267];
    assign layer5_out[5869] = ~layer4_out[1597];
    assign layer5_out[5870] = ~layer4_out[5742] | layer4_out[5743];
    assign layer5_out[5871] = ~(layer4_out[4932] | layer4_out[4933]);
    assign layer5_out[5872] = ~(layer4_out[262] & layer4_out[263]);
    assign layer5_out[5873] = layer4_out[3294] & layer4_out[3295];
    assign layer5_out[5874] = ~(layer4_out[7532] ^ layer4_out[7533]);
    assign layer5_out[5875] = layer4_out[1194] ^ layer4_out[1195];
    assign layer5_out[5876] = layer4_out[4745];
    assign layer5_out[5877] = ~(layer4_out[4600] ^ layer4_out[4601]);
    assign layer5_out[5878] = ~layer4_out[4350];
    assign layer5_out[5879] = ~layer4_out[1746];
    assign layer5_out[5880] = layer4_out[7757];
    assign layer5_out[5881] = layer4_out[4077];
    assign layer5_out[5882] = ~layer4_out[2301];
    assign layer5_out[5883] = layer4_out[715];
    assign layer5_out[5884] = layer4_out[3626] ^ layer4_out[3627];
    assign layer5_out[5885] = layer4_out[3637];
    assign layer5_out[5886] = layer4_out[6749] & ~layer4_out[6750];
    assign layer5_out[5887] = ~layer4_out[7572];
    assign layer5_out[5888] = ~layer4_out[1856];
    assign layer5_out[5889] = ~(layer4_out[6740] ^ layer4_out[6741]);
    assign layer5_out[5890] = ~(layer4_out[1506] | layer4_out[1507]);
    assign layer5_out[5891] = layer4_out[7506] ^ layer4_out[7507];
    assign layer5_out[5892] = layer4_out[6024] & ~layer4_out[6025];
    assign layer5_out[5893] = layer4_out[5252] & layer4_out[5253];
    assign layer5_out[5894] = ~layer4_out[1250];
    assign layer5_out[5895] = layer4_out[2001] | layer4_out[2002];
    assign layer5_out[5896] = ~layer4_out[4198];
    assign layer5_out[5897] = ~layer4_out[1724];
    assign layer5_out[5898] = ~layer4_out[7100];
    assign layer5_out[5899] = ~(layer4_out[3721] | layer4_out[3722]);
    assign layer5_out[5900] = ~layer4_out[804];
    assign layer5_out[5901] = layer4_out[1043];
    assign layer5_out[5902] = layer4_out[573] & ~layer4_out[572];
    assign layer5_out[5903] = layer4_out[956];
    assign layer5_out[5904] = ~(layer4_out[7540] ^ layer4_out[7541]);
    assign layer5_out[5905] = ~(layer4_out[7946] & layer4_out[7947]);
    assign layer5_out[5906] = layer4_out[3603] & ~layer4_out[3604];
    assign layer5_out[5907] = ~(layer4_out[5704] | layer4_out[5705]);
    assign layer5_out[5908] = ~layer4_out[3350];
    assign layer5_out[5909] = ~(layer4_out[7816] ^ layer4_out[7817]);
    assign layer5_out[5910] = ~(layer4_out[5297] ^ layer4_out[5298]);
    assign layer5_out[5911] = ~layer4_out[824];
    assign layer5_out[5912] = ~layer4_out[2876];
    assign layer5_out[5913] = ~(layer4_out[6199] ^ layer4_out[6200]);
    assign layer5_out[5914] = layer4_out[1844] & ~layer4_out[1845];
    assign layer5_out[5915] = layer4_out[598] | layer4_out[599];
    assign layer5_out[5916] = layer4_out[5610];
    assign layer5_out[5917] = layer4_out[1793];
    assign layer5_out[5918] = layer4_out[370] ^ layer4_out[371];
    assign layer5_out[5919] = ~layer4_out[7941];
    assign layer5_out[5920] = layer4_out[3453] & layer4_out[3454];
    assign layer5_out[5921] = layer4_out[81];
    assign layer5_out[5922] = ~layer4_out[7818];
    assign layer5_out[5923] = layer4_out[6291] & ~layer4_out[6290];
    assign layer5_out[5924] = layer4_out[4410] & layer4_out[4411];
    assign layer5_out[5925] = layer4_out[6078] & ~layer4_out[6077];
    assign layer5_out[5926] = layer4_out[419] | layer4_out[420];
    assign layer5_out[5927] = layer4_out[7022] & layer4_out[7023];
    assign layer5_out[5928] = layer4_out[308] | layer4_out[309];
    assign layer5_out[5929] = layer4_out[2357] & layer4_out[2358];
    assign layer5_out[5930] = layer4_out[2070] ^ layer4_out[2071];
    assign layer5_out[5931] = layer4_out[3874];
    assign layer5_out[5932] = ~layer4_out[5909] | layer4_out[5910];
    assign layer5_out[5933] = layer4_out[3850] & ~layer4_out[3851];
    assign layer5_out[5934] = ~(layer4_out[6657] | layer4_out[6658]);
    assign layer5_out[5935] = ~layer4_out[1130];
    assign layer5_out[5936] = layer4_out[7875];
    assign layer5_out[5937] = ~(layer4_out[2847] ^ layer4_out[2848]);
    assign layer5_out[5938] = ~layer4_out[834];
    assign layer5_out[5939] = ~(layer4_out[877] ^ layer4_out[878]);
    assign layer5_out[5940] = ~(layer4_out[6634] ^ layer4_out[6635]);
    assign layer5_out[5941] = ~layer4_out[156];
    assign layer5_out[5942] = layer4_out[5122] & ~layer4_out[5123];
    assign layer5_out[5943] = layer4_out[1905] & layer4_out[1906];
    assign layer5_out[5944] = ~layer4_out[4940];
    assign layer5_out[5945] = ~(layer4_out[7436] ^ layer4_out[7437]);
    assign layer5_out[5946] = layer4_out[7503];
    assign layer5_out[5947] = ~layer4_out[1821];
    assign layer5_out[5948] = layer4_out[6051] | layer4_out[6052];
    assign layer5_out[5949] = ~(layer4_out[2842] | layer4_out[2843]);
    assign layer5_out[5950] = layer4_out[515] ^ layer4_out[516];
    assign layer5_out[5951] = layer4_out[6128] ^ layer4_out[6129];
    assign layer5_out[5952] = ~layer4_out[6846] | layer4_out[6845];
    assign layer5_out[5953] = layer4_out[7950];
    assign layer5_out[5954] = layer4_out[3151] & layer4_out[3152];
    assign layer5_out[5955] = layer4_out[6633] & layer4_out[6634];
    assign layer5_out[5956] = layer4_out[5832] & ~layer4_out[5831];
    assign layer5_out[5957] = layer4_out[1615];
    assign layer5_out[5958] = ~(layer4_out[6420] & layer4_out[6421]);
    assign layer5_out[5959] = layer4_out[975] & ~layer4_out[974];
    assign layer5_out[5960] = ~(layer4_out[6141] ^ layer4_out[6142]);
    assign layer5_out[5961] = ~layer4_out[5426];
    assign layer5_out[5962] = layer4_out[4981];
    assign layer5_out[5963] = layer4_out[4491] & layer4_out[4492];
    assign layer5_out[5964] = ~(layer4_out[7379] & layer4_out[7380]);
    assign layer5_out[5965] = layer4_out[5554] & ~layer4_out[5553];
    assign layer5_out[5966] = layer4_out[2190] ^ layer4_out[2191];
    assign layer5_out[5967] = layer4_out[3447] ^ layer4_out[3448];
    assign layer5_out[5968] = layer4_out[6168];
    assign layer5_out[5969] = ~(layer4_out[6529] & layer4_out[6530]);
    assign layer5_out[5970] = layer4_out[6057];
    assign layer5_out[5971] = layer4_out[7480];
    assign layer5_out[5972] = layer4_out[6437] ^ layer4_out[6438];
    assign layer5_out[5973] = layer4_out[6010];
    assign layer5_out[5974] = layer4_out[2614];
    assign layer5_out[5975] = ~(layer4_out[477] ^ layer4_out[478]);
    assign layer5_out[5976] = ~(layer4_out[5198] | layer4_out[5199]);
    assign layer5_out[5977] = layer4_out[6792] ^ layer4_out[6793];
    assign layer5_out[5978] = layer4_out[1759];
    assign layer5_out[5979] = ~layer4_out[5583];
    assign layer5_out[5980] = layer4_out[6625] | layer4_out[6626];
    assign layer5_out[5981] = layer4_out[488] & ~layer4_out[487];
    assign layer5_out[5982] = layer4_out[1173];
    assign layer5_out[5983] = ~layer4_out[4279];
    assign layer5_out[5984] = layer4_out[2332] ^ layer4_out[2333];
    assign layer5_out[5985] = ~layer4_out[2236];
    assign layer5_out[5986] = ~layer4_out[4031] | layer4_out[4032];
    assign layer5_out[5987] = layer4_out[3906] ^ layer4_out[3907];
    assign layer5_out[5988] = layer4_out[7627];
    assign layer5_out[5989] = layer4_out[7338] ^ layer4_out[7339];
    assign layer5_out[5990] = layer4_out[7229];
    assign layer5_out[5991] = ~(layer4_out[5531] ^ layer4_out[5532]);
    assign layer5_out[5992] = ~(layer4_out[3385] | layer4_out[3386]);
    assign layer5_out[5993] = ~layer4_out[7380];
    assign layer5_out[5994] = ~layer4_out[261];
    assign layer5_out[5995] = layer4_out[3388] ^ layer4_out[3389];
    assign layer5_out[5996] = layer4_out[5098];
    assign layer5_out[5997] = layer4_out[1528];
    assign layer5_out[5998] = layer4_out[5954] & ~layer4_out[5955];
    assign layer5_out[5999] = ~layer4_out[6802] | layer4_out[6803];
    assign layer5_out[6000] = layer4_out[1599] & ~layer4_out[1600];
    assign layer5_out[6001] = layer4_out[5550] & ~layer4_out[5551];
    assign layer5_out[6002] = layer4_out[1144];
    assign layer5_out[6003] = ~layer4_out[6146] | layer4_out[6147];
    assign layer5_out[6004] = ~layer4_out[7862] | layer4_out[7861];
    assign layer5_out[6005] = ~(layer4_out[6219] ^ layer4_out[6220]);
    assign layer5_out[6006] = ~(layer4_out[2949] ^ layer4_out[2950]);
    assign layer5_out[6007] = ~(layer4_out[2768] ^ layer4_out[2769]);
    assign layer5_out[6008] = layer4_out[4973];
    assign layer5_out[6009] = ~layer4_out[2534];
    assign layer5_out[6010] = ~layer4_out[1865];
    assign layer5_out[6011] = layer4_out[977] ^ layer4_out[978];
    assign layer5_out[6012] = layer4_out[4722] ^ layer4_out[4723];
    assign layer5_out[6013] = layer4_out[4925] | layer4_out[4926];
    assign layer5_out[6014] = ~layer4_out[6176];
    assign layer5_out[6015] = ~(layer4_out[4808] | layer4_out[4809]);
    assign layer5_out[6016] = layer4_out[1316];
    assign layer5_out[6017] = layer4_out[6591] ^ layer4_out[6592];
    assign layer5_out[6018] = ~layer4_out[3326] | layer4_out[3325];
    assign layer5_out[6019] = layer4_out[7527] & ~layer4_out[7528];
    assign layer5_out[6020] = layer4_out[2803] ^ layer4_out[2804];
    assign layer5_out[6021] = layer4_out[3996];
    assign layer5_out[6022] = ~layer4_out[2926];
    assign layer5_out[6023] = ~(layer4_out[571] | layer4_out[572]);
    assign layer5_out[6024] = layer4_out[7316];
    assign layer5_out[6025] = layer4_out[7658] ^ layer4_out[7659];
    assign layer5_out[6026] = ~(layer4_out[6983] ^ layer4_out[6984]);
    assign layer5_out[6027] = ~layer4_out[3810];
    assign layer5_out[6028] = layer4_out[1502] | layer4_out[1503];
    assign layer5_out[6029] = ~(layer4_out[2200] | layer4_out[2201]);
    assign layer5_out[6030] = ~layer4_out[2484];
    assign layer5_out[6031] = layer4_out[4176] | layer4_out[4177];
    assign layer5_out[6032] = layer4_out[4111];
    assign layer5_out[6033] = ~(layer4_out[0] ^ layer4_out[2]);
    assign layer5_out[6034] = layer4_out[1153] & ~layer4_out[1154];
    assign layer5_out[6035] = layer4_out[4160];
    assign layer5_out[6036] = ~layer4_out[2072] | layer4_out[2071];
    assign layer5_out[6037] = layer4_out[5111] ^ layer4_out[5112];
    assign layer5_out[6038] = ~layer4_out[1398];
    assign layer5_out[6039] = layer4_out[3225] & ~layer4_out[3224];
    assign layer5_out[6040] = layer4_out[2795];
    assign layer5_out[6041] = layer4_out[6806];
    assign layer5_out[6042] = layer4_out[7034] | layer4_out[7035];
    assign layer5_out[6043] = ~(layer4_out[2340] ^ layer4_out[2341]);
    assign layer5_out[6044] = layer4_out[1877] & layer4_out[1878];
    assign layer5_out[6045] = layer4_out[3273] & ~layer4_out[3272];
    assign layer5_out[6046] = ~(layer4_out[5576] ^ layer4_out[5577]);
    assign layer5_out[6047] = ~layer4_out[7232];
    assign layer5_out[6048] = ~layer4_out[5151];
    assign layer5_out[6049] = layer4_out[6366];
    assign layer5_out[6050] = ~layer4_out[427];
    assign layer5_out[6051] = layer4_out[7831] & layer4_out[7832];
    assign layer5_out[6052] = layer4_out[3491];
    assign layer5_out[6053] = layer4_out[2060];
    assign layer5_out[6054] = layer4_out[2917] & ~layer4_out[2918];
    assign layer5_out[6055] = layer4_out[3505] & ~layer4_out[3506];
    assign layer5_out[6056] = layer4_out[6995];
    assign layer5_out[6057] = ~layer4_out[2091] | layer4_out[2090];
    assign layer5_out[6058] = layer4_out[2620];
    assign layer5_out[6059] = layer4_out[2928];
    assign layer5_out[6060] = layer4_out[825];
    assign layer5_out[6061] = layer4_out[507];
    assign layer5_out[6062] = layer4_out[6150] ^ layer4_out[6151];
    assign layer5_out[6063] = ~layer4_out[2657];
    assign layer5_out[6064] = ~layer4_out[7181];
    assign layer5_out[6065] = layer4_out[1089] & layer4_out[1090];
    assign layer5_out[6066] = ~layer4_out[3715];
    assign layer5_out[6067] = layer4_out[3478];
    assign layer5_out[6068] = ~(layer4_out[7271] & layer4_out[7272]);
    assign layer5_out[6069] = ~(layer4_out[2698] ^ layer4_out[2699]);
    assign layer5_out[6070] = ~(layer4_out[6015] ^ layer4_out[6016]);
    assign layer5_out[6071] = ~(layer4_out[746] | layer4_out[747]);
    assign layer5_out[6072] = layer4_out[304] & ~layer4_out[305];
    assign layer5_out[6073] = layer4_out[1700];
    assign layer5_out[6074] = ~(layer4_out[6912] ^ layer4_out[6913]);
    assign layer5_out[6075] = ~layer4_out[6547];
    assign layer5_out[6076] = layer4_out[1546];
    assign layer5_out[6077] = layer4_out[4183];
    assign layer5_out[6078] = layer4_out[530] ^ layer4_out[531];
    assign layer5_out[6079] = layer4_out[4160] & layer4_out[4161];
    assign layer5_out[6080] = layer4_out[6360] ^ layer4_out[6361];
    assign layer5_out[6081] = ~(layer4_out[5644] ^ layer4_out[5645]);
    assign layer5_out[6082] = layer4_out[3678];
    assign layer5_out[6083] = layer4_out[3379];
    assign layer5_out[6084] = layer4_out[4340];
    assign layer5_out[6085] = ~layer4_out[2282] | layer4_out[2283];
    assign layer5_out[6086] = layer4_out[4391];
    assign layer5_out[6087] = ~(layer4_out[4919] ^ layer4_out[4920]);
    assign layer5_out[6088] = ~layer4_out[4384];
    assign layer5_out[6089] = ~layer4_out[4064];
    assign layer5_out[6090] = ~(layer4_out[7909] | layer4_out[7910]);
    assign layer5_out[6091] = layer4_out[2816] & layer4_out[2817];
    assign layer5_out[6092] = ~layer4_out[258];
    assign layer5_out[6093] = layer4_out[4599];
    assign layer5_out[6094] = ~layer4_out[5952];
    assign layer5_out[6095] = layer4_out[434] & ~layer4_out[433];
    assign layer5_out[6096] = layer4_out[7591] & ~layer4_out[7592];
    assign layer5_out[6097] = layer4_out[2052] ^ layer4_out[2053];
    assign layer5_out[6098] = ~(layer4_out[4506] ^ layer4_out[4507]);
    assign layer5_out[6099] = ~(layer4_out[2969] ^ layer4_out[2970]);
    assign layer5_out[6100] = ~(layer4_out[7116] | layer4_out[7117]);
    assign layer5_out[6101] = layer4_out[7836] ^ layer4_out[7837];
    assign layer5_out[6102] = layer4_out[3847];
    assign layer5_out[6103] = ~(layer4_out[4368] | layer4_out[4369]);
    assign layer5_out[6104] = ~(layer4_out[3326] & layer4_out[3327]);
    assign layer5_out[6105] = layer4_out[3463] & ~layer4_out[3464];
    assign layer5_out[6106] = ~layer4_out[1032];
    assign layer5_out[6107] = layer4_out[3287];
    assign layer5_out[6108] = ~layer4_out[7599];
    assign layer5_out[6109] = ~(layer4_out[1214] ^ layer4_out[1215]);
    assign layer5_out[6110] = layer4_out[4693] ^ layer4_out[4694];
    assign layer5_out[6111] = layer4_out[1630] & layer4_out[1631];
    assign layer5_out[6112] = layer4_out[1227] | layer4_out[1228];
    assign layer5_out[6113] = layer4_out[7494];
    assign layer5_out[6114] = ~layer4_out[2176] | layer4_out[2177];
    assign layer5_out[6115] = layer4_out[4441];
    assign layer5_out[6116] = ~layer4_out[1623];
    assign layer5_out[6117] = layer4_out[7284] & ~layer4_out[7283];
    assign layer5_out[6118] = layer4_out[1127];
    assign layer5_out[6119] = ~(layer4_out[2789] ^ layer4_out[2790]);
    assign layer5_out[6120] = layer4_out[1876] ^ layer4_out[1877];
    assign layer5_out[6121] = ~(layer4_out[4675] ^ layer4_out[4676]);
    assign layer5_out[6122] = ~(layer4_out[2530] ^ layer4_out[2531]);
    assign layer5_out[6123] = ~(layer4_out[7568] & layer4_out[7569]);
    assign layer5_out[6124] = layer4_out[5296];
    assign layer5_out[6125] = ~(layer4_out[6511] | layer4_out[6512]);
    assign layer5_out[6126] = layer4_out[5607];
    assign layer5_out[6127] = layer4_out[187] & layer4_out[188];
    assign layer5_out[6128] = ~(layer4_out[5521] | layer4_out[5522]);
    assign layer5_out[6129] = ~(layer4_out[7728] ^ layer4_out[7729]);
    assign layer5_out[6130] = ~layer4_out[1539];
    assign layer5_out[6131] = layer4_out[3347] ^ layer4_out[3348];
    assign layer5_out[6132] = layer4_out[3732] & ~layer4_out[3731];
    assign layer5_out[6133] = layer4_out[2887];
    assign layer5_out[6134] = ~layer4_out[7773];
    assign layer5_out[6135] = layer4_out[1360] ^ layer4_out[1361];
    assign layer5_out[6136] = layer4_out[4168] ^ layer4_out[4169];
    assign layer5_out[6137] = ~(layer4_out[1741] ^ layer4_out[1742]);
    assign layer5_out[6138] = ~(layer4_out[1989] | layer4_out[1990]);
    assign layer5_out[6139] = layer4_out[1745];
    assign layer5_out[6140] = ~(layer4_out[2757] | layer4_out[2758]);
    assign layer5_out[6141] = layer4_out[4002];
    assign layer5_out[6142] = layer4_out[2035] ^ layer4_out[2036];
    assign layer5_out[6143] = ~(layer4_out[6447] ^ layer4_out[6448]);
    assign layer5_out[6144] = ~layer4_out[630];
    assign layer5_out[6145] = ~(layer4_out[7262] ^ layer4_out[7263]);
    assign layer5_out[6146] = ~layer4_out[7863];
    assign layer5_out[6147] = ~layer4_out[5836] | layer4_out[5835];
    assign layer5_out[6148] = ~(layer4_out[3744] ^ layer4_out[3745]);
    assign layer5_out[6149] = ~layer4_out[2213] | layer4_out[2212];
    assign layer5_out[6150] = layer4_out[7782] & ~layer4_out[7781];
    assign layer5_out[6151] = layer4_out[1237] & ~layer4_out[1238];
    assign layer5_out[6152] = ~layer4_out[33];
    assign layer5_out[6153] = ~(layer4_out[3568] ^ layer4_out[3569]);
    assign layer5_out[6154] = layer4_out[287] & layer4_out[288];
    assign layer5_out[6155] = ~layer4_out[1569];
    assign layer5_out[6156] = ~(layer4_out[4323] & layer4_out[4324]);
    assign layer5_out[6157] = layer4_out[3930] & ~layer4_out[3931];
    assign layer5_out[6158] = ~layer4_out[229];
    assign layer5_out[6159] = ~(layer4_out[2401] ^ layer4_out[2402]);
    assign layer5_out[6160] = layer4_out[1913];
    assign layer5_out[6161] = layer4_out[2726] | layer4_out[2727];
    assign layer5_out[6162] = layer4_out[6700] & layer4_out[6701];
    assign layer5_out[6163] = ~layer4_out[7339];
    assign layer5_out[6164] = layer4_out[2770] | layer4_out[2771];
    assign layer5_out[6165] = ~(layer4_out[333] ^ layer4_out[334]);
    assign layer5_out[6166] = layer4_out[1830] & ~layer4_out[1829];
    assign layer5_out[6167] = ~layer4_out[951];
    assign layer5_out[6168] = ~layer4_out[5009];
    assign layer5_out[6169] = ~layer4_out[2522];
    assign layer5_out[6170] = ~layer4_out[3320];
    assign layer5_out[6171] = layer4_out[6238] ^ layer4_out[6239];
    assign layer5_out[6172] = ~layer4_out[7569] | layer4_out[7570];
    assign layer5_out[6173] = layer4_out[4272] ^ layer4_out[4273];
    assign layer5_out[6174] = ~layer4_out[7387];
    assign layer5_out[6175] = ~layer4_out[3604];
    assign layer5_out[6176] = ~layer4_out[2905];
    assign layer5_out[6177] = ~layer4_out[3691];
    assign layer5_out[6178] = ~layer4_out[4057];
    assign layer5_out[6179] = ~layer4_out[2282];
    assign layer5_out[6180] = ~layer4_out[2370];
    assign layer5_out[6181] = ~layer4_out[2713] | layer4_out[2712];
    assign layer5_out[6182] = layer4_out[4765];
    assign layer5_out[6183] = layer4_out[5089];
    assign layer5_out[6184] = ~(layer4_out[4948] ^ layer4_out[4949]);
    assign layer5_out[6185] = ~layer4_out[5398];
    assign layer5_out[6186] = ~layer4_out[6496] | layer4_out[6497];
    assign layer5_out[6187] = ~(layer4_out[6305] ^ layer4_out[6306]);
    assign layer5_out[6188] = ~layer4_out[4766] | layer4_out[4767];
    assign layer5_out[6189] = layer4_out[1868];
    assign layer5_out[6190] = ~layer4_out[4544] | layer4_out[4543];
    assign layer5_out[6191] = ~layer4_out[532];
    assign layer5_out[6192] = layer4_out[6250] & ~layer4_out[6249];
    assign layer5_out[6193] = ~(layer4_out[4219] ^ layer4_out[4220]);
    assign layer5_out[6194] = layer4_out[2832];
    assign layer5_out[6195] = ~layer4_out[4209];
    assign layer5_out[6196] = layer4_out[7796] ^ layer4_out[7797];
    assign layer5_out[6197] = layer4_out[796] ^ layer4_out[797];
    assign layer5_out[6198] = ~layer4_out[675];
    assign layer5_out[6199] = ~layer4_out[1477];
    assign layer5_out[6200] = layer4_out[6062];
    assign layer5_out[6201] = layer4_out[6123];
    assign layer5_out[6202] = layer4_out[1753];
    assign layer5_out[6203] = layer4_out[698];
    assign layer5_out[6204] = layer4_out[2447] ^ layer4_out[2448];
    assign layer5_out[6205] = layer4_out[6436] | layer4_out[6437];
    assign layer5_out[6206] = ~layer4_out[3962] | layer4_out[3963];
    assign layer5_out[6207] = ~(layer4_out[6160] ^ layer4_out[6161]);
    assign layer5_out[6208] = layer4_out[3329] & ~layer4_out[3328];
    assign layer5_out[6209] = layer4_out[738] & ~layer4_out[737];
    assign layer5_out[6210] = layer4_out[1027];
    assign layer5_out[6211] = ~(layer4_out[7806] ^ layer4_out[7807]);
    assign layer5_out[6212] = layer4_out[7871] ^ layer4_out[7872];
    assign layer5_out[6213] = layer4_out[3134] & ~layer4_out[3133];
    assign layer5_out[6214] = ~(layer4_out[389] | layer4_out[390]);
    assign layer5_out[6215] = layer4_out[763];
    assign layer5_out[6216] = ~(layer4_out[5153] & layer4_out[5154]);
    assign layer5_out[6217] = layer4_out[5547] | layer4_out[5548];
    assign layer5_out[6218] = layer4_out[6307] ^ layer4_out[6308];
    assign layer5_out[6219] = layer4_out[5786] & ~layer4_out[5785];
    assign layer5_out[6220] = layer4_out[7417] | layer4_out[7418];
    assign layer5_out[6221] = layer4_out[5304];
    assign layer5_out[6222] = ~(layer4_out[3246] ^ layer4_out[3247]);
    assign layer5_out[6223] = ~(layer4_out[2037] ^ layer4_out[2038]);
    assign layer5_out[6224] = layer4_out[4492];
    assign layer5_out[6225] = layer4_out[83] & layer4_out[84];
    assign layer5_out[6226] = layer4_out[4285] ^ layer4_out[4286];
    assign layer5_out[6227] = ~layer4_out[6517];
    assign layer5_out[6228] = layer4_out[518] ^ layer4_out[519];
    assign layer5_out[6229] = ~layer4_out[474];
    assign layer5_out[6230] = layer4_out[4459];
    assign layer5_out[6231] = layer4_out[2832];
    assign layer5_out[6232] = layer4_out[685] ^ layer4_out[686];
    assign layer5_out[6233] = layer4_out[1760];
    assign layer5_out[6234] = layer4_out[6513] & ~layer4_out[6512];
    assign layer5_out[6235] = ~layer4_out[7499];
    assign layer5_out[6236] = layer4_out[1110];
    assign layer5_out[6237] = layer4_out[6227];
    assign layer5_out[6238] = layer4_out[3757] ^ layer4_out[3758];
    assign layer5_out[6239] = layer4_out[7799] ^ layer4_out[7800];
    assign layer5_out[6240] = ~layer4_out[2220];
    assign layer5_out[6241] = ~(layer4_out[7922] & layer4_out[7923]);
    assign layer5_out[6242] = ~(layer4_out[756] & layer4_out[757]);
    assign layer5_out[6243] = ~(layer4_out[6898] ^ layer4_out[6899]);
    assign layer5_out[6244] = ~layer4_out[2968] | layer4_out[2967];
    assign layer5_out[6245] = layer4_out[3120] & layer4_out[3121];
    assign layer5_out[6246] = layer4_out[2445] | layer4_out[2446];
    assign layer5_out[6247] = layer4_out[4073];
    assign layer5_out[6248] = layer4_out[6928] & layer4_out[6929];
    assign layer5_out[6249] = layer4_out[2791] & layer4_out[2792];
    assign layer5_out[6250] = ~layer4_out[1126] | layer4_out[1127];
    assign layer5_out[6251] = ~(layer4_out[5526] & layer4_out[5527]);
    assign layer5_out[6252] = layer4_out[3694] & ~layer4_out[3695];
    assign layer5_out[6253] = layer4_out[7747] ^ layer4_out[7748];
    assign layer5_out[6254] = layer4_out[4603];
    assign layer5_out[6255] = layer4_out[5571] ^ layer4_out[5572];
    assign layer5_out[6256] = ~(layer4_out[7947] ^ layer4_out[7948]);
    assign layer5_out[6257] = layer4_out[1356] ^ layer4_out[1357];
    assign layer5_out[6258] = ~(layer4_out[5581] | layer4_out[5582]);
    assign layer5_out[6259] = ~layer4_out[5071] | layer4_out[5070];
    assign layer5_out[6260] = layer4_out[942];
    assign layer5_out[6261] = ~layer4_out[2709] | layer4_out[2710];
    assign layer5_out[6262] = layer4_out[3109];
    assign layer5_out[6263] = layer4_out[4514] | layer4_out[4515];
    assign layer5_out[6264] = ~(layer4_out[4056] & layer4_out[4057]);
    assign layer5_out[6265] = ~layer4_out[713] | layer4_out[712];
    assign layer5_out[6266] = layer4_out[1961];
    assign layer5_out[6267] = ~(layer4_out[1220] ^ layer4_out[1221]);
    assign layer5_out[6268] = ~layer4_out[2061] | layer4_out[2062];
    assign layer5_out[6269] = layer4_out[2246] & layer4_out[2247];
    assign layer5_out[6270] = ~(layer4_out[2806] | layer4_out[2807]);
    assign layer5_out[6271] = layer4_out[5790] & layer4_out[5791];
    assign layer5_out[6272] = layer4_out[5808];
    assign layer5_out[6273] = layer4_out[1248];
    assign layer5_out[6274] = ~layer4_out[260];
    assign layer5_out[6275] = ~layer4_out[1430] | layer4_out[1429];
    assign layer5_out[6276] = ~(layer4_out[3348] ^ layer4_out[3349]);
    assign layer5_out[6277] = layer4_out[6651];
    assign layer5_out[6278] = ~layer4_out[3573];
    assign layer5_out[6279] = ~layer4_out[4381];
    assign layer5_out[6280] = layer4_out[6432] & layer4_out[6433];
    assign layer5_out[6281] = ~layer4_out[2396];
    assign layer5_out[6282] = layer4_out[295] ^ layer4_out[296];
    assign layer5_out[6283] = layer4_out[3336];
    assign layer5_out[6284] = ~layer4_out[5676] | layer4_out[5677];
    assign layer5_out[6285] = layer4_out[190] & ~layer4_out[189];
    assign layer5_out[6286] = ~layer4_out[560];
    assign layer5_out[6287] = layer4_out[1721];
    assign layer5_out[6288] = layer4_out[5113] ^ layer4_out[5114];
    assign layer5_out[6289] = layer4_out[2661];
    assign layer5_out[6290] = layer4_out[1735];
    assign layer5_out[6291] = layer4_out[7930] ^ layer4_out[7931];
    assign layer5_out[6292] = layer4_out[1318] & ~layer4_out[1319];
    assign layer5_out[6293] = layer4_out[7104];
    assign layer5_out[6294] = layer4_out[3689];
    assign layer5_out[6295] = layer4_out[6410] | layer4_out[6411];
    assign layer5_out[6296] = layer4_out[5646] & layer4_out[5647];
    assign layer5_out[6297] = ~layer4_out[3212];
    assign layer5_out[6298] = ~(layer4_out[425] ^ layer4_out[426]);
    assign layer5_out[6299] = layer4_out[5699] & ~layer4_out[5698];
    assign layer5_out[6300] = ~layer4_out[2180];
    assign layer5_out[6301] = ~(layer4_out[4753] ^ layer4_out[4754]);
    assign layer5_out[6302] = ~layer4_out[1421];
    assign layer5_out[6303] = ~layer4_out[6853];
    assign layer5_out[6304] = ~(layer4_out[3891] | layer4_out[3892]);
    assign layer5_out[6305] = layer4_out[1768] ^ layer4_out[1769];
    assign layer5_out[6306] = ~layer4_out[2720];
    assign layer5_out[6307] = ~layer4_out[2285] | layer4_out[2286];
    assign layer5_out[6308] = layer4_out[1422];
    assign layer5_out[6309] = layer4_out[3795] & ~layer4_out[3796];
    assign layer5_out[6310] = ~layer4_out[6953];
    assign layer5_out[6311] = ~layer4_out[615];
    assign layer5_out[6312] = ~layer4_out[2447] | layer4_out[2446];
    assign layer5_out[6313] = ~(layer4_out[7311] & layer4_out[7312]);
    assign layer5_out[6314] = ~layer4_out[4444];
    assign layer5_out[6315] = ~(layer4_out[1497] & layer4_out[1498]);
    assign layer5_out[6316] = layer4_out[2917];
    assign layer5_out[6317] = ~layer4_out[5400];
    assign layer5_out[6318] = layer4_out[106];
    assign layer5_out[6319] = layer4_out[4351] ^ layer4_out[4352];
    assign layer5_out[6320] = ~(layer4_out[4691] ^ layer4_out[4692]);
    assign layer5_out[6321] = layer4_out[1778];
    assign layer5_out[6322] = layer4_out[6088];
    assign layer5_out[6323] = ~(layer4_out[6297] ^ layer4_out[6298]);
    assign layer5_out[6324] = layer4_out[1371] & layer4_out[1372];
    assign layer5_out[6325] = ~(layer4_out[5275] | layer4_out[5276]);
    assign layer5_out[6326] = ~layer4_out[4005];
    assign layer5_out[6327] = ~layer4_out[2595];
    assign layer5_out[6328] = layer4_out[7619];
    assign layer5_out[6329] = ~layer4_out[3113];
    assign layer5_out[6330] = ~layer4_out[5039];
    assign layer5_out[6331] = layer4_out[5321] & layer4_out[5322];
    assign layer5_out[6332] = layer4_out[2269] ^ layer4_out[2270];
    assign layer5_out[6333] = ~layer4_out[5956];
    assign layer5_out[6334] = layer4_out[5765] ^ layer4_out[5766];
    assign layer5_out[6335] = ~(layer4_out[2612] ^ layer4_out[2613]);
    assign layer5_out[6336] = ~layer4_out[1019] | layer4_out[1018];
    assign layer5_out[6337] = ~layer4_out[5441];
    assign layer5_out[6338] = layer4_out[4702] & ~layer4_out[4701];
    assign layer5_out[6339] = ~layer4_out[6285] | layer4_out[6286];
    assign layer5_out[6340] = layer4_out[7358] & ~layer4_out[7357];
    assign layer5_out[6341] = ~layer4_out[1836];
    assign layer5_out[6342] = ~(layer4_out[7472] | layer4_out[7473]);
    assign layer5_out[6343] = ~layer4_out[5622];
    assign layer5_out[6344] = layer4_out[5867];
    assign layer5_out[6345] = ~layer4_out[980];
    assign layer5_out[6346] = layer4_out[6828] & layer4_out[6829];
    assign layer5_out[6347] = layer4_out[4573];
    assign layer5_out[6348] = ~layer4_out[7030];
    assign layer5_out[6349] = ~(layer4_out[123] ^ layer4_out[124]);
    assign layer5_out[6350] = ~layer4_out[4288];
    assign layer5_out[6351] = ~layer4_out[2088];
    assign layer5_out[6352] = ~layer4_out[2899] | layer4_out[2900];
    assign layer5_out[6353] = layer4_out[3547] & ~layer4_out[3546];
    assign layer5_out[6354] = ~layer4_out[3228];
    assign layer5_out[6355] = layer4_out[5971] ^ layer4_out[5972];
    assign layer5_out[6356] = ~layer4_out[4984];
    assign layer5_out[6357] = layer4_out[3148];
    assign layer5_out[6358] = layer4_out[2043] ^ layer4_out[2044];
    assign layer5_out[6359] = ~layer4_out[7840];
    assign layer5_out[6360] = layer4_out[5365];
    assign layer5_out[6361] = layer4_out[1314];
    assign layer5_out[6362] = ~layer4_out[5428];
    assign layer5_out[6363] = layer4_out[5458] ^ layer4_out[5459];
    assign layer5_out[6364] = ~layer4_out[1992];
    assign layer5_out[6365] = ~(layer4_out[7600] & layer4_out[7601]);
    assign layer5_out[6366] = ~(layer4_out[4208] | layer4_out[4209]);
    assign layer5_out[6367] = ~layer4_out[5916];
    assign layer5_out[6368] = layer4_out[4838] & ~layer4_out[4837];
    assign layer5_out[6369] = ~layer4_out[4248];
    assign layer5_out[6370] = layer4_out[791] & ~layer4_out[792];
    assign layer5_out[6371] = layer4_out[7138] ^ layer4_out[7139];
    assign layer5_out[6372] = layer4_out[2234] | layer4_out[2235];
    assign layer5_out[6373] = ~(layer4_out[139] ^ layer4_out[140]);
    assign layer5_out[6374] = ~layer4_out[603] | layer4_out[602];
    assign layer5_out[6375] = ~layer4_out[1114];
    assign layer5_out[6376] = ~layer4_out[2872];
    assign layer5_out[6377] = ~layer4_out[5614];
    assign layer5_out[6378] = layer4_out[687] ^ layer4_out[688];
    assign layer5_out[6379] = layer4_out[779];
    assign layer5_out[6380] = ~layer4_out[6948];
    assign layer5_out[6381] = ~layer4_out[1756];
    assign layer5_out[6382] = layer4_out[7212] & ~layer4_out[7213];
    assign layer5_out[6383] = layer4_out[2531] ^ layer4_out[2532];
    assign layer5_out[6384] = layer4_out[2701] & ~layer4_out[2702];
    assign layer5_out[6385] = layer4_out[5834] ^ layer4_out[5835];
    assign layer5_out[6386] = layer4_out[5203] & ~layer4_out[5204];
    assign layer5_out[6387] = ~layer4_out[2007];
    assign layer5_out[6388] = ~(layer4_out[1122] ^ layer4_out[1123]);
    assign layer5_out[6389] = ~layer4_out[5465];
    assign layer5_out[6390] = ~(layer4_out[1236] ^ layer4_out[1237]);
    assign layer5_out[6391] = layer4_out[1737];
    assign layer5_out[6392] = layer4_out[7088];
    assign layer5_out[6393] = ~layer4_out[6931];
    assign layer5_out[6394] = ~layer4_out[7717];
    assign layer5_out[6395] = layer4_out[7394] & ~layer4_out[7393];
    assign layer5_out[6396] = layer4_out[4463] ^ layer4_out[4464];
    assign layer5_out[6397] = layer4_out[1093];
    assign layer5_out[6398] = ~layer4_out[1444];
    assign layer5_out[6399] = ~layer4_out[6012] | layer4_out[6011];
    assign layer5_out[6400] = layer4_out[22] & layer4_out[23];
    assign layer5_out[6401] = ~layer4_out[7033];
    assign layer5_out[6402] = ~layer4_out[3046];
    assign layer5_out[6403] = ~(layer4_out[2114] ^ layer4_out[2115]);
    assign layer5_out[6404] = layer4_out[7089] ^ layer4_out[7090];
    assign layer5_out[6405] = ~layer4_out[1231];
    assign layer5_out[6406] = ~layer4_out[7173];
    assign layer5_out[6407] = ~(layer4_out[1043] ^ layer4_out[1044]);
    assign layer5_out[6408] = layer4_out[1639] & layer4_out[1640];
    assign layer5_out[6409] = layer4_out[5087];
    assign layer5_out[6410] = layer4_out[2812];
    assign layer5_out[6411] = layer4_out[7940];
    assign layer5_out[6412] = layer4_out[4431] ^ layer4_out[4432];
    assign layer5_out[6413] = ~(layer4_out[6883] ^ layer4_out[6884]);
    assign layer5_out[6414] = layer4_out[4441] | layer4_out[4442];
    assign layer5_out[6415] = layer4_out[7398] ^ layer4_out[7399];
    assign layer5_out[6416] = ~(layer4_out[5051] ^ layer4_out[5052]);
    assign layer5_out[6417] = ~(layer4_out[5199] ^ layer4_out[5200]);
    assign layer5_out[6418] = ~(layer4_out[3196] | layer4_out[3197]);
    assign layer5_out[6419] = ~layer4_out[2619];
    assign layer5_out[6420] = ~(layer4_out[3115] ^ layer4_out[3116]);
    assign layer5_out[6421] = layer4_out[6392] ^ layer4_out[6393];
    assign layer5_out[6422] = ~layer4_out[3414];
    assign layer5_out[6423] = layer4_out[7479];
    assign layer5_out[6424] = ~layer4_out[3633];
    assign layer5_out[6425] = ~layer4_out[4680];
    assign layer5_out[6426] = ~(layer4_out[3681] ^ layer4_out[3682]);
    assign layer5_out[6427] = ~layer4_out[1349] | layer4_out[1350];
    assign layer5_out[6428] = ~layer4_out[1416] | layer4_out[1415];
    assign layer5_out[6429] = layer4_out[7772];
    assign layer5_out[6430] = layer4_out[1330];
    assign layer5_out[6431] = ~layer4_out[2479];
    assign layer5_out[6432] = layer4_out[3825];
    assign layer5_out[6433] = layer4_out[2837];
    assign layer5_out[6434] = layer4_out[1190] ^ layer4_out[1191];
    assign layer5_out[6435] = layer4_out[590] & ~layer4_out[589];
    assign layer5_out[6436] = layer4_out[7064] | layer4_out[7065];
    assign layer5_out[6437] = layer4_out[284] | layer4_out[285];
    assign layer5_out[6438] = layer4_out[6714];
    assign layer5_out[6439] = layer4_out[6530] & layer4_out[6531];
    assign layer5_out[6440] = ~layer4_out[7487];
    assign layer5_out[6441] = ~(layer4_out[4367] ^ layer4_out[4368]);
    assign layer5_out[6442] = ~(layer4_out[2244] & layer4_out[2245]);
    assign layer5_out[6443] = ~layer4_out[3387] | layer4_out[3386];
    assign layer5_out[6444] = layer4_out[4833] ^ layer4_out[4834];
    assign layer5_out[6445] = layer4_out[6450];
    assign layer5_out[6446] = ~layer4_out[5047];
    assign layer5_out[6447] = layer4_out[6221] & ~layer4_out[6222];
    assign layer5_out[6448] = layer4_out[4591];
    assign layer5_out[6449] = ~(layer4_out[1640] ^ layer4_out[1641]);
    assign layer5_out[6450] = layer4_out[5733] ^ layer4_out[5734];
    assign layer5_out[6451] = layer4_out[5279] ^ layer4_out[5280];
    assign layer5_out[6452] = ~(layer4_out[232] & layer4_out[233]);
    assign layer5_out[6453] = layer4_out[3283] | layer4_out[3284];
    assign layer5_out[6454] = layer4_out[4214] ^ layer4_out[4215];
    assign layer5_out[6455] = layer4_out[2545] | layer4_out[2546];
    assign layer5_out[6456] = layer4_out[3487];
    assign layer5_out[6457] = layer4_out[7359];
    assign layer5_out[6458] = layer4_out[1979] ^ layer4_out[1980];
    assign layer5_out[6459] = layer4_out[6971] ^ layer4_out[6972];
    assign layer5_out[6460] = ~layer4_out[2896];
    assign layer5_out[6461] = layer4_out[2543] ^ layer4_out[2544];
    assign layer5_out[6462] = layer4_out[5508] | layer4_out[5509];
    assign layer5_out[6463] = ~layer4_out[3509] | layer4_out[3510];
    assign layer5_out[6464] = ~layer4_out[2650];
    assign layer5_out[6465] = layer4_out[1169] ^ layer4_out[1170];
    assign layer5_out[6466] = layer4_out[2066] & ~layer4_out[2067];
    assign layer5_out[6467] = ~layer4_out[6940] | layer4_out[6941];
    assign layer5_out[6468] = ~layer4_out[3441];
    assign layer5_out[6469] = layer4_out[870];
    assign layer5_out[6470] = layer4_out[2765];
    assign layer5_out[6471] = layer4_out[4021] ^ layer4_out[4022];
    assign layer5_out[6472] = layer4_out[2173] & ~layer4_out[2174];
    assign layer5_out[6473] = ~(layer4_out[7896] ^ layer4_out[7897]);
    assign layer5_out[6474] = ~layer4_out[3200] | layer4_out[3199];
    assign layer5_out[6475] = layer4_out[5208] & ~layer4_out[5209];
    assign layer5_out[6476] = ~(layer4_out[6588] ^ layer4_out[6589]);
    assign layer5_out[6477] = ~layer4_out[7850] | layer4_out[7849];
    assign layer5_out[6478] = ~layer4_out[1296];
    assign layer5_out[6479] = ~(layer4_out[6955] ^ layer4_out[6956]);
    assign layer5_out[6480] = ~(layer4_out[1815] ^ layer4_out[1816]);
    assign layer5_out[6481] = ~layer4_out[7620];
    assign layer5_out[6482] = ~layer4_out[5223];
    assign layer5_out[6483] = ~(layer4_out[2161] ^ layer4_out[2162]);
    assign layer5_out[6484] = ~layer4_out[3254];
    assign layer5_out[6485] = ~layer4_out[3373];
    assign layer5_out[6486] = layer4_out[1358];
    assign layer5_out[6487] = ~layer4_out[7475];
    assign layer5_out[6488] = ~layer4_out[901] | layer4_out[902];
    assign layer5_out[6489] = layer4_out[2951];
    assign layer5_out[6490] = ~layer4_out[5876];
    assign layer5_out[6491] = ~(layer4_out[4217] ^ layer4_out[4218]);
    assign layer5_out[6492] = ~layer4_out[4197];
    assign layer5_out[6493] = layer4_out[2066] & ~layer4_out[2065];
    assign layer5_out[6494] = layer4_out[7983];
    assign layer5_out[6495] = ~(layer4_out[708] ^ layer4_out[709]);
    assign layer5_out[6496] = layer4_out[4458];
    assign layer5_out[6497] = ~layer4_out[1051] | layer4_out[1052];
    assign layer5_out[6498] = ~layer4_out[4451];
    assign layer5_out[6499] = ~(layer4_out[163] | layer4_out[164]);
    assign layer5_out[6500] = ~(layer4_out[7743] ^ layer4_out[7744]);
    assign layer5_out[6501] = ~(layer4_out[903] | layer4_out[904]);
    assign layer5_out[6502] = ~(layer4_out[2480] ^ layer4_out[2481]);
    assign layer5_out[6503] = ~(layer4_out[864] ^ layer4_out[865]);
    assign layer5_out[6504] = ~(layer4_out[6236] | layer4_out[6237]);
    assign layer5_out[6505] = ~layer4_out[3322] | layer4_out[3321];
    assign layer5_out[6506] = layer4_out[5226] & ~layer4_out[5227];
    assign layer5_out[6507] = ~layer4_out[4849];
    assign layer5_out[6508] = layer4_out[7965];
    assign layer5_out[6509] = ~layer4_out[3392];
    assign layer5_out[6510] = layer4_out[7542];
    assign layer5_out[6511] = ~layer4_out[2012];
    assign layer5_out[6512] = ~(layer4_out[4139] | layer4_out[4140]);
    assign layer5_out[6513] = ~(layer4_out[341] | layer4_out[342]);
    assign layer5_out[6514] = ~layer4_out[5439];
    assign layer5_out[6515] = layer4_out[6871];
    assign layer5_out[6516] = layer4_out[380] & ~layer4_out[381];
    assign layer5_out[6517] = ~layer4_out[3301];
    assign layer5_out[6518] = layer4_out[6528] & ~layer4_out[6527];
    assign layer5_out[6519] = layer4_out[1008] | layer4_out[1009];
    assign layer5_out[6520] = ~layer4_out[2139];
    assign layer5_out[6521] = ~layer4_out[6328] | layer4_out[6329];
    assign layer5_out[6522] = layer4_out[5273];
    assign layer5_out[6523] = layer4_out[97];
    assign layer5_out[6524] = ~(layer4_out[684] ^ layer4_out[685]);
    assign layer5_out[6525] = layer4_out[2724] & layer4_out[2725];
    assign layer5_out[6526] = ~layer4_out[5252] | layer4_out[5251];
    assign layer5_out[6527] = ~(layer4_out[970] ^ layer4_out[971]);
    assign layer5_out[6528] = layer4_out[5033];
    assign layer5_out[6529] = ~(layer4_out[7877] ^ layer4_out[7878]);
    assign layer5_out[6530] = ~(layer4_out[4244] ^ layer4_out[4245]);
    assign layer5_out[6531] = layer4_out[1495] ^ layer4_out[1496];
    assign layer5_out[6532] = ~layer4_out[4284] | layer4_out[4285];
    assign layer5_out[6533] = layer4_out[3766] | layer4_out[3767];
    assign layer5_out[6534] = ~layer4_out[391];
    assign layer5_out[6535] = layer4_out[7782] | layer4_out[7783];
    assign layer5_out[6536] = ~layer4_out[6181];
    assign layer5_out[6537] = ~(layer4_out[1795] ^ layer4_out[1796]);
    assign layer5_out[6538] = ~layer4_out[6502];
    assign layer5_out[6539] = ~layer4_out[4857];
    assign layer5_out[6540] = layer4_out[3166];
    assign layer5_out[6541] = layer4_out[2742] & ~layer4_out[2741];
    assign layer5_out[6542] = layer4_out[138] & ~layer4_out[137];
    assign layer5_out[6543] = layer4_out[4364];
    assign layer5_out[6544] = layer4_out[3879] & layer4_out[3880];
    assign layer5_out[6545] = layer4_out[4190] | layer4_out[4191];
    assign layer5_out[6546] = ~layer4_out[6070];
    assign layer5_out[6547] = layer4_out[5328];
    assign layer5_out[6548] = layer4_out[6574];
    assign layer5_out[6549] = ~layer4_out[4958] | layer4_out[4959];
    assign layer5_out[6550] = ~layer4_out[660];
    assign layer5_out[6551] = ~layer4_out[5206];
    assign layer5_out[6552] = ~layer4_out[901];
    assign layer5_out[6553] = ~layer4_out[100];
    assign layer5_out[6554] = ~layer4_out[1663] | layer4_out[1664];
    assign layer5_out[6555] = layer4_out[7554];
    assign layer5_out[6556] = layer4_out[7744];
    assign layer5_out[6557] = layer4_out[2963];
    assign layer5_out[6558] = ~layer4_out[730];
    assign layer5_out[6559] = layer4_out[594];
    assign layer5_out[6560] = layer4_out[2179];
    assign layer5_out[6561] = layer4_out[6825] ^ layer4_out[6826];
    assign layer5_out[6562] = layer4_out[6076] ^ layer4_out[6077];
    assign layer5_out[6563] = layer4_out[2789];
    assign layer5_out[6564] = ~layer4_out[2587];
    assign layer5_out[6565] = layer4_out[772] ^ layer4_out[773];
    assign layer5_out[6566] = layer4_out[6799];
    assign layer5_out[6567] = ~layer4_out[2547] | layer4_out[2548];
    assign layer5_out[6568] = ~(layer4_out[5323] & layer4_out[5324]);
    assign layer5_out[6569] = layer4_out[2186];
    assign layer5_out[6570] = layer4_out[6871];
    assign layer5_out[6571] = ~layer4_out[2954];
    assign layer5_out[6572] = ~(layer4_out[3814] & layer4_out[3815]);
    assign layer5_out[6573] = ~(layer4_out[273] & layer4_out[274]);
    assign layer5_out[6574] = layer4_out[4267] & layer4_out[4268];
    assign layer5_out[6575] = ~(layer4_out[5651] ^ layer4_out[5652]);
    assign layer5_out[6576] = ~(layer4_out[4661] | layer4_out[4662]);
    assign layer5_out[6577] = layer4_out[5259];
    assign layer5_out[6578] = ~layer4_out[2064];
    assign layer5_out[6579] = layer4_out[4078] ^ layer4_out[4079];
    assign layer5_out[6580] = layer4_out[6136];
    assign layer5_out[6581] = ~(layer4_out[1910] ^ layer4_out[1911]);
    assign layer5_out[6582] = ~layer4_out[5499];
    assign layer5_out[6583] = ~layer4_out[1915] | layer4_out[1916];
    assign layer5_out[6584] = ~layer4_out[7993];
    assign layer5_out[6585] = layer4_out[1855] & layer4_out[1856];
    assign layer5_out[6586] = ~layer4_out[2683] | layer4_out[2684];
    assign layer5_out[6587] = layer4_out[6035];
    assign layer5_out[6588] = ~layer4_out[1793];
    assign layer5_out[6589] = ~layer4_out[4649];
    assign layer5_out[6590] = layer4_out[6722] & ~layer4_out[6723];
    assign layer5_out[6591] = layer4_out[6382];
    assign layer5_out[6592] = layer4_out[3922] & ~layer4_out[3923];
    assign layer5_out[6593] = layer4_out[4071];
    assign layer5_out[6594] = layer4_out[1882] ^ layer4_out[1883];
    assign layer5_out[6595] = ~(layer4_out[471] ^ layer4_out[472]);
    assign layer5_out[6596] = layer4_out[5806];
    assign layer5_out[6597] = layer4_out[1161] ^ layer4_out[1162];
    assign layer5_out[6598] = ~layer4_out[6156];
    assign layer5_out[6599] = layer4_out[5744];
    assign layer5_out[6600] = ~layer4_out[7529] | layer4_out[7530];
    assign layer5_out[6601] = layer4_out[284];
    assign layer5_out[6602] = layer4_out[733];
    assign layer5_out[6603] = ~layer4_out[1667];
    assign layer5_out[6604] = ~layer4_out[3344] | layer4_out[3343];
    assign layer5_out[6605] = ~layer4_out[2817] | layer4_out[2818];
    assign layer5_out[6606] = layer4_out[5289];
    assign layer5_out[6607] = layer4_out[4700];
    assign layer5_out[6608] = ~(layer4_out[1919] | layer4_out[1920]);
    assign layer5_out[6609] = layer4_out[3207];
    assign layer5_out[6610] = ~(layer4_out[4937] ^ layer4_out[4938]);
    assign layer5_out[6611] = layer4_out[2578] ^ layer4_out[2579];
    assign layer5_out[6612] = ~layer4_out[2893] | layer4_out[2894];
    assign layer5_out[6613] = ~layer4_out[5051] | layer4_out[5050];
    assign layer5_out[6614] = layer4_out[1854];
    assign layer5_out[6615] = ~(layer4_out[6846] ^ layer4_out[6847]);
    assign layer5_out[6616] = ~(layer4_out[797] & layer4_out[798]);
    assign layer5_out[6617] = layer4_out[6514];
    assign layer5_out[6618] = ~layer4_out[6094];
    assign layer5_out[6619] = ~layer4_out[5118];
    assign layer5_out[6620] = layer4_out[3777];
    assign layer5_out[6621] = ~layer4_out[191];
    assign layer5_out[6622] = ~layer4_out[4177];
    assign layer5_out[6623] = layer4_out[2137];
    assign layer5_out[6624] = layer4_out[1205];
    assign layer5_out[6625] = layer4_out[4946] | layer4_out[4947];
    assign layer5_out[6626] = layer4_out[6253];
    assign layer5_out[6627] = ~(layer4_out[7533] | layer4_out[7534]);
    assign layer5_out[6628] = layer4_out[5658];
    assign layer5_out[6629] = layer4_out[911] & ~layer4_out[910];
    assign layer5_out[6630] = ~(layer4_out[7112] ^ layer4_out[7113]);
    assign layer5_out[6631] = ~(layer4_out[3915] ^ layer4_out[3916]);
    assign layer5_out[6632] = layer4_out[1387];
    assign layer5_out[6633] = layer4_out[236] ^ layer4_out[237];
    assign layer5_out[6634] = layer4_out[1053];
    assign layer5_out[6635] = ~(layer4_out[2327] ^ layer4_out[2328]);
    assign layer5_out[6636] = ~layer4_out[6349] | layer4_out[6350];
    assign layer5_out[6637] = ~(layer4_out[7832] ^ layer4_out[7833]);
    assign layer5_out[6638] = layer4_out[7750] ^ layer4_out[7751];
    assign layer5_out[6639] = layer4_out[2410] ^ layer4_out[2411];
    assign layer5_out[6640] = layer4_out[4878] & layer4_out[4879];
    assign layer5_out[6641] = layer4_out[3580];
    assign layer5_out[6642] = layer4_out[5093] ^ layer4_out[5094];
    assign layer5_out[6643] = layer4_out[2022];
    assign layer5_out[6644] = ~(layer4_out[3053] ^ layer4_out[3054]);
    assign layer5_out[6645] = layer4_out[408];
    assign layer5_out[6646] = layer4_out[4449];
    assign layer5_out[6647] = layer4_out[1600] ^ layer4_out[1601];
    assign layer5_out[6648] = ~layer4_out[187] | layer4_out[186];
    assign layer5_out[6649] = ~layer4_out[5060];
    assign layer5_out[6650] = layer4_out[2102];
    assign layer5_out[6651] = ~layer4_out[6923];
    assign layer5_out[6652] = ~(layer4_out[2713] | layer4_out[2714]);
    assign layer5_out[6653] = layer4_out[4473];
    assign layer5_out[6654] = layer4_out[1325];
    assign layer5_out[6655] = ~(layer4_out[998] ^ layer4_out[999]);
    assign layer5_out[6656] = ~layer4_out[726];
    assign layer5_out[6657] = layer4_out[991] ^ layer4_out[992];
    assign layer5_out[6658] = layer4_out[1404];
    assign layer5_out[6659] = layer4_out[6863];
    assign layer5_out[6660] = layer4_out[2172];
    assign layer5_out[6661] = layer4_out[2051] & ~layer4_out[2050];
    assign layer5_out[6662] = layer4_out[1189];
    assign layer5_out[6663] = layer4_out[7752] & layer4_out[7753];
    assign layer5_out[6664] = layer4_out[5108] ^ layer4_out[5109];
    assign layer5_out[6665] = layer4_out[5631] ^ layer4_out[5632];
    assign layer5_out[6666] = ~(layer4_out[5663] | layer4_out[5664]);
    assign layer5_out[6667] = ~(layer4_out[3432] & layer4_out[3433]);
    assign layer5_out[6668] = ~(layer4_out[3967] ^ layer4_out[3968]);
    assign layer5_out[6669] = layer4_out[2375];
    assign layer5_out[6670] = layer4_out[3402] & layer4_out[3403];
    assign layer5_out[6671] = ~layer4_out[4885] | layer4_out[4886];
    assign layer5_out[6672] = ~(layer4_out[1301] ^ layer4_out[1302]);
    assign layer5_out[6673] = layer4_out[565] & layer4_out[566];
    assign layer5_out[6674] = layer4_out[5273];
    assign layer5_out[6675] = ~(layer4_out[1321] ^ layer4_out[1322]);
    assign layer5_out[6676] = layer4_out[2500] & layer4_out[2501];
    assign layer5_out[6677] = layer4_out[3284] ^ layer4_out[3285];
    assign layer5_out[6678] = ~layer4_out[1440];
    assign layer5_out[6679] = ~(layer4_out[6559] | layer4_out[6560]);
    assign layer5_out[6680] = ~layer4_out[1010] | layer4_out[1009];
    assign layer5_out[6681] = ~layer4_out[4762] | layer4_out[4761];
    assign layer5_out[6682] = ~(layer4_out[7588] ^ layer4_out[7589]);
    assign layer5_out[6683] = layer4_out[1455] & ~layer4_out[1454];
    assign layer5_out[6684] = layer4_out[485] & layer4_out[486];
    assign layer5_out[6685] = layer4_out[803] & ~layer4_out[802];
    assign layer5_out[6686] = layer4_out[7297];
    assign layer5_out[6687] = ~layer4_out[2547] | layer4_out[2546];
    assign layer5_out[6688] = ~(layer4_out[3927] ^ layer4_out[3928]);
    assign layer5_out[6689] = layer4_out[5281] ^ layer4_out[5282];
    assign layer5_out[6690] = ~layer4_out[662];
    assign layer5_out[6691] = ~layer4_out[1178] | layer4_out[1179];
    assign layer5_out[6692] = ~(layer4_out[6617] ^ layer4_out[6618]);
    assign layer5_out[6693] = ~layer4_out[2849] | layer4_out[2848];
    assign layer5_out[6694] = ~layer4_out[7742] | layer4_out[7741];
    assign layer5_out[6695] = ~layer4_out[440];
    assign layer5_out[6696] = ~layer4_out[1518];
    assign layer5_out[6697] = layer4_out[6664];
    assign layer5_out[6698] = layer4_out[7];
    assign layer5_out[6699] = ~(layer4_out[1563] ^ layer4_out[1564]);
    assign layer5_out[6700] = layer4_out[4737] ^ layer4_out[4738];
    assign layer5_out[6701] = ~layer4_out[5692] | layer4_out[5693];
    assign layer5_out[6702] = ~layer4_out[2527];
    assign layer5_out[6703] = layer4_out[7790];
    assign layer5_out[6704] = ~(layer4_out[7241] & layer4_out[7242]);
    assign layer5_out[6705] = ~layer4_out[456];
    assign layer5_out[6706] = ~layer4_out[2349];
    assign layer5_out[6707] = layer4_out[49] ^ layer4_out[50];
    assign layer5_out[6708] = ~(layer4_out[6054] & layer4_out[6055]);
    assign layer5_out[6709] = layer4_out[1434];
    assign layer5_out[6710] = ~layer4_out[10];
    assign layer5_out[6711] = layer4_out[4135];
    assign layer5_out[6712] = layer4_out[6756];
    assign layer5_out[6713] = layer4_out[3556];
    assign layer5_out[6714] = ~(layer4_out[2267] & layer4_out[2268]);
    assign layer5_out[6715] = ~layer4_out[1575];
    assign layer5_out[6716] = layer4_out[5176] ^ layer4_out[5177];
    assign layer5_out[6717] = layer4_out[7772];
    assign layer5_out[6718] = ~layer4_out[3603];
    assign layer5_out[6719] = layer4_out[5854];
    assign layer5_out[6720] = layer4_out[1636] & layer4_out[1637];
    assign layer5_out[6721] = ~(layer4_out[6000] ^ layer4_out[6001]);
    assign layer5_out[6722] = layer4_out[2028];
    assign layer5_out[6723] = layer4_out[271];
    assign layer5_out[6724] = layer4_out[2613] ^ layer4_out[2614];
    assign layer5_out[6725] = ~layer4_out[3196] | layer4_out[3195];
    assign layer5_out[6726] = ~layer4_out[861];
    assign layer5_out[6727] = layer4_out[7674] ^ layer4_out[7675];
    assign layer5_out[6728] = ~(layer4_out[1658] ^ layer4_out[1659]);
    assign layer5_out[6729] = layer4_out[5737] & ~layer4_out[5738];
    assign layer5_out[6730] = ~(layer4_out[297] | layer4_out[298]);
    assign layer5_out[6731] = ~(layer4_out[664] & layer4_out[665]);
    assign layer5_out[6732] = layer4_out[5470] & ~layer4_out[5469];
    assign layer5_out[6733] = ~(layer4_out[6116] | layer4_out[6117]);
    assign layer5_out[6734] = ~(layer4_out[1601] ^ layer4_out[1602]);
    assign layer5_out[6735] = ~layer4_out[5515];
    assign layer5_out[6736] = layer4_out[4203];
    assign layer5_out[6737] = layer4_out[786];
    assign layer5_out[6738] = layer4_out[7270];
    assign layer5_out[6739] = layer4_out[770];
    assign layer5_out[6740] = ~layer4_out[6913] | layer4_out[6914];
    assign layer5_out[6741] = layer4_out[1775] ^ layer4_out[1776];
    assign layer5_out[6742] = layer4_out[5898] & ~layer4_out[5899];
    assign layer5_out[6743] = layer4_out[4342] ^ layer4_out[4343];
    assign layer5_out[6744] = ~layer4_out[4305] | layer4_out[4304];
    assign layer5_out[6745] = layer4_out[6725];
    assign layer5_out[6746] = layer4_out[4166] & layer4_out[4167];
    assign layer5_out[6747] = layer4_out[1922] ^ layer4_out[1923];
    assign layer5_out[6748] = ~layer4_out[2784] | layer4_out[2783];
    assign layer5_out[6749] = ~(layer4_out[5040] ^ layer4_out[5041]);
    assign layer5_out[6750] = layer4_out[6954] ^ layer4_out[6955];
    assign layer5_out[6751] = layer4_out[7615] & ~layer4_out[7614];
    assign layer5_out[6752] = layer4_out[7389];
    assign layer5_out[6753] = ~layer4_out[6696];
    assign layer5_out[6754] = layer4_out[6821] ^ layer4_out[6822];
    assign layer5_out[6755] = ~(layer4_out[1778] | layer4_out[1779]);
    assign layer5_out[6756] = layer4_out[347];
    assign layer5_out[6757] = layer4_out[7082];
    assign layer5_out[6758] = ~layer4_out[6005];
    assign layer5_out[6759] = ~layer4_out[1850] | layer4_out[1849];
    assign layer5_out[6760] = layer4_out[3259];
    assign layer5_out[6761] = layer4_out[7169] & layer4_out[7170];
    assign layer5_out[6762] = ~layer4_out[788] | layer4_out[787];
    assign layer5_out[6763] = layer4_out[1942] ^ layer4_out[1943];
    assign layer5_out[6764] = layer4_out[6931];
    assign layer5_out[6765] = layer4_out[3890];
    assign layer5_out[6766] = ~layer4_out[4964];
    assign layer5_out[6767] = ~layer4_out[7876] | layer4_out[7877];
    assign layer5_out[6768] = ~(layer4_out[4509] ^ layer4_out[4510]);
    assign layer5_out[6769] = layer4_out[3481] & ~layer4_out[3482];
    assign layer5_out[6770] = layer4_out[2501] | layer4_out[2502];
    assign layer5_out[6771] = layer4_out[4523] & layer4_out[4524];
    assign layer5_out[6772] = layer4_out[4439];
    assign layer5_out[6773] = ~layer4_out[7298];
    assign layer5_out[6774] = layer4_out[2128] | layer4_out[2129];
    assign layer5_out[6775] = ~(layer4_out[2238] | layer4_out[2239]);
    assign layer5_out[6776] = layer4_out[6702] ^ layer4_out[6703];
    assign layer5_out[6777] = ~(layer4_out[7201] & layer4_out[7202]);
    assign layer5_out[6778] = layer4_out[2163];
    assign layer5_out[6779] = layer4_out[4184] & ~layer4_out[4185];
    assign layer5_out[6780] = layer4_out[5029];
    assign layer5_out[6781] = ~layer4_out[4397] | layer4_out[4398];
    assign layer5_out[6782] = ~(layer4_out[340] & layer4_out[341]);
    assign layer5_out[6783] = layer4_out[194] & layer4_out[195];
    assign layer5_out[6784] = layer4_out[4518] & ~layer4_out[4517];
    assign layer5_out[6785] = ~(layer4_out[6389] & layer4_out[6390]);
    assign layer5_out[6786] = ~layer4_out[1231];
    assign layer5_out[6787] = ~(layer4_out[2650] | layer4_out[2651]);
    assign layer5_out[6788] = layer4_out[4298];
    assign layer5_out[6789] = ~(layer4_out[591] ^ layer4_out[592]);
    assign layer5_out[6790] = layer4_out[4604];
    assign layer5_out[6791] = layer4_out[5173] & layer4_out[5174];
    assign layer5_out[6792] = ~(layer4_out[6585] & layer4_out[6586]);
    assign layer5_out[6793] = ~layer4_out[857];
    assign layer5_out[6794] = layer4_out[4888];
    assign layer5_out[6795] = layer4_out[6892];
    assign layer5_out[6796] = ~layer4_out[7911];
    assign layer5_out[6797] = layer4_out[5201];
    assign layer5_out[6798] = ~layer4_out[2336];
    assign layer5_out[6799] = ~(layer4_out[7684] ^ layer4_out[7685]);
    assign layer5_out[6800] = layer4_out[6265] | layer4_out[6266];
    assign layer5_out[6801] = layer4_out[2560] & ~layer4_out[2561];
    assign layer5_out[6802] = layer4_out[1019];
    assign layer5_out[6803] = layer4_out[1946];
    assign layer5_out[6804] = layer4_out[6887] ^ layer4_out[6888];
    assign layer5_out[6805] = ~layer4_out[4185] | layer4_out[4186];
    assign layer5_out[6806] = ~(layer4_out[5707] | layer4_out[5708]);
    assign layer5_out[6807] = layer4_out[3063] ^ layer4_out[3064];
    assign layer5_out[6808] = layer4_out[1707];
    assign layer5_out[6809] = ~(layer4_out[4335] ^ layer4_out[4336]);
    assign layer5_out[6810] = layer4_out[2688];
    assign layer5_out[6811] = layer4_out[5785];
    assign layer5_out[6812] = ~layer4_out[2130] | layer4_out[2129];
    assign layer5_out[6813] = ~(layer4_out[5358] ^ layer4_out[5359]);
    assign layer5_out[6814] = ~(layer4_out[79] ^ layer4_out[80]);
    assign layer5_out[6815] = layer4_out[4171];
    assign layer5_out[6816] = ~(layer4_out[5333] ^ layer4_out[5334]);
    assign layer5_out[6817] = layer4_out[379] | layer4_out[380];
    assign layer5_out[6818] = ~(layer4_out[3761] ^ layer4_out[3762]);
    assign layer5_out[6819] = layer4_out[1398];
    assign layer5_out[6820] = ~(layer4_out[6342] ^ layer4_out[6343]);
    assign layer5_out[6821] = ~layer4_out[7786] | layer4_out[7787];
    assign layer5_out[6822] = ~(layer4_out[2157] | layer4_out[2158]);
    assign layer5_out[6823] = ~layer4_out[1688];
    assign layer5_out[6824] = ~layer4_out[5134];
    assign layer5_out[6825] = ~layer4_out[644];
    assign layer5_out[6826] = ~layer4_out[1375] | layer4_out[1374];
    assign layer5_out[6827] = layer4_out[126];
    assign layer5_out[6828] = ~layer4_out[7465] | layer4_out[7466];
    assign layer5_out[6829] = ~layer4_out[18] | layer4_out[17];
    assign layer5_out[6830] = ~(layer4_out[7274] ^ layer4_out[7275]);
    assign layer5_out[6831] = layer4_out[4934];
    assign layer5_out[6832] = layer4_out[6689];
    assign layer5_out[6833] = layer4_out[3896] ^ layer4_out[3897];
    assign layer5_out[6834] = layer4_out[6557] ^ layer4_out[6558];
    assign layer5_out[6835] = layer4_out[7612] | layer4_out[7613];
    assign layer5_out[6836] = layer4_out[2107];
    assign layer5_out[6837] = ~(layer4_out[774] | layer4_out[775]);
    assign layer5_out[6838] = ~layer4_out[825] | layer4_out[824];
    assign layer5_out[6839] = layer4_out[23] & layer4_out[24];
    assign layer5_out[6840] = ~layer4_out[5099] | layer4_out[5100];
    assign layer5_out[6841] = ~(layer4_out[6242] ^ layer4_out[6243]);
    assign layer5_out[6842] = layer4_out[5987] ^ layer4_out[5988];
    assign layer5_out[6843] = layer4_out[1291];
    assign layer5_out[6844] = ~(layer4_out[2019] ^ layer4_out[2020]);
    assign layer5_out[6845] = ~(layer4_out[5761] ^ layer4_out[5762]);
    assign layer5_out[6846] = layer4_out[4527] ^ layer4_out[4528];
    assign layer5_out[6847] = ~layer4_out[5451];
    assign layer5_out[6848] = ~(layer4_out[5365] | layer4_out[5366]);
    assign layer5_out[6849] = ~(layer4_out[1732] ^ layer4_out[1733]);
    assign layer5_out[6850] = ~(layer4_out[783] | layer4_out[784]);
    assign layer5_out[6851] = layer4_out[2213] | layer4_out[2214];
    assign layer5_out[6852] = layer4_out[4582];
    assign layer5_out[6853] = ~layer4_out[1247];
    assign layer5_out[6854] = ~(layer4_out[7162] | layer4_out[7163]);
    assign layer5_out[6855] = ~(layer4_out[7003] ^ layer4_out[7004]);
    assign layer5_out[6856] = ~(layer4_out[997] ^ layer4_out[998]);
    assign layer5_out[6857] = ~(layer4_out[2013] ^ layer4_out[2014]);
    assign layer5_out[6858] = ~layer4_out[7935] | layer4_out[7936];
    assign layer5_out[6859] = layer4_out[4114] | layer4_out[4115];
    assign layer5_out[6860] = layer4_out[6731] ^ layer4_out[6732];
    assign layer5_out[6861] = ~(layer4_out[3073] ^ layer4_out[3074]);
    assign layer5_out[6862] = layer4_out[3628] & ~layer4_out[3629];
    assign layer5_out[6863] = ~layer4_out[7265];
    assign layer5_out[6864] = layer4_out[1441] & ~layer4_out[1440];
    assign layer5_out[6865] = layer4_out[5849] ^ layer4_out[5850];
    assign layer5_out[6866] = ~layer4_out[3188];
    assign layer5_out[6867] = layer4_out[7756] & ~layer4_out[7755];
    assign layer5_out[6868] = layer4_out[1377] ^ layer4_out[1378];
    assign layer5_out[6869] = ~(layer4_out[3184] | layer4_out[3185]);
    assign layer5_out[6870] = ~(layer4_out[4908] ^ layer4_out[4909]);
    assign layer5_out[6871] = ~(layer4_out[5706] ^ layer4_out[5707]);
    assign layer5_out[6872] = ~layer4_out[866];
    assign layer5_out[6873] = ~(layer4_out[7978] ^ layer4_out[7979]);
    assign layer5_out[6874] = layer4_out[5086];
    assign layer5_out[6875] = ~(layer4_out[1763] ^ layer4_out[1764]);
    assign layer5_out[6876] = layer4_out[6084] & ~layer4_out[6083];
    assign layer5_out[6877] = layer4_out[6229] ^ layer4_out[6230];
    assign layer5_out[6878] = ~(layer4_out[5768] ^ layer4_out[5769]);
    assign layer5_out[6879] = layer4_out[3596] | layer4_out[3597];
    assign layer5_out[6880] = layer4_out[6494];
    assign layer5_out[6881] = layer4_out[4303] & layer4_out[4304];
    assign layer5_out[6882] = ~(layer4_out[5512] ^ layer4_out[5513]);
    assign layer5_out[6883] = layer4_out[7693];
    assign layer5_out[6884] = ~layer4_out[2346] | layer4_out[2345];
    assign layer5_out[6885] = layer4_out[3578];
    assign layer5_out[6886] = ~layer4_out[7876];
    assign layer5_out[6887] = ~(layer4_out[2494] | layer4_out[2495]);
    assign layer5_out[6888] = layer4_out[5429] ^ layer4_out[5430];
    assign layer5_out[6889] = layer4_out[5589] & ~layer4_out[5590];
    assign layer5_out[6890] = layer4_out[7784];
    assign layer5_out[6891] = ~(layer4_out[56] ^ layer4_out[57]);
    assign layer5_out[6892] = layer4_out[4859] | layer4_out[4860];
    assign layer5_out[6893] = ~layer4_out[6916];
    assign layer5_out[6894] = layer4_out[2991];
    assign layer5_out[6895] = ~(layer4_out[4206] ^ layer4_out[4207]);
    assign layer5_out[6896] = layer4_out[7449] | layer4_out[7450];
    assign layer5_out[6897] = ~(layer4_out[3990] ^ layer4_out[3991]);
    assign layer5_out[6898] = layer4_out[3324] ^ layer4_out[3325];
    assign layer5_out[6899] = layer4_out[2414] & ~layer4_out[2413];
    assign layer5_out[6900] = layer4_out[7344] ^ layer4_out[7345];
    assign layer5_out[6901] = layer4_out[4044];
    assign layer5_out[6902] = layer4_out[1582] ^ layer4_out[1583];
    assign layer5_out[6903] = ~layer4_out[4411] | layer4_out[4412];
    assign layer5_out[6904] = layer4_out[3358] | layer4_out[3359];
    assign layer5_out[6905] = layer4_out[4221];
    assign layer5_out[6906] = ~(layer4_out[1964] ^ layer4_out[1965]);
    assign layer5_out[6907] = ~layer4_out[3559] | layer4_out[3560];
    assign layer5_out[6908] = layer4_out[6233] & ~layer4_out[6234];
    assign layer5_out[6909] = ~layer4_out[3383];
    assign layer5_out[6910] = layer4_out[2562] ^ layer4_out[2563];
    assign layer5_out[6911] = ~layer4_out[7203];
    assign layer5_out[6912] = layer4_out[1556] ^ layer4_out[1557];
    assign layer5_out[6913] = layer4_out[2083];
    assign layer5_out[6914] = layer4_out[6126] ^ layer4_out[6127];
    assign layer5_out[6915] = ~layer4_out[299];
    assign layer5_out[6916] = ~layer4_out[4248];
    assign layer5_out[6917] = ~(layer4_out[7438] ^ layer4_out[7439]);
    assign layer5_out[6918] = layer4_out[1751];
    assign layer5_out[6919] = ~(layer4_out[757] & layer4_out[758]);
    assign layer5_out[6920] = layer4_out[6395] & layer4_out[6396];
    assign layer5_out[6921] = layer4_out[6187] ^ layer4_out[6188];
    assign layer5_out[6922] = ~layer4_out[4804] | layer4_out[4805];
    assign layer5_out[6923] = ~(layer4_out[3263] & layer4_out[3264]);
    assign layer5_out[6924] = layer4_out[5863];
    assign layer5_out[6925] = layer4_out[7461];
    assign layer5_out[6926] = ~layer4_out[1236];
    assign layer5_out[6927] = layer4_out[69] ^ layer4_out[70];
    assign layer5_out[6928] = layer4_out[6493];
    assign layer5_out[6929] = layer4_out[795] & ~layer4_out[794];
    assign layer5_out[6930] = ~layer4_out[6384];
    assign layer5_out[6931] = layer4_out[4570];
    assign layer5_out[6932] = ~layer4_out[4956] | layer4_out[4957];
    assign layer5_out[6933] = layer4_out[5589];
    assign layer5_out[6934] = ~layer4_out[3688];
    assign layer5_out[6935] = layer4_out[4846] & ~layer4_out[4845];
    assign layer5_out[6936] = layer4_out[4101] ^ layer4_out[4102];
    assign layer5_out[6937] = layer4_out[710] ^ layer4_out[711];
    assign layer5_out[6938] = layer4_out[1274] & ~layer4_out[1273];
    assign layer5_out[6939] = ~(layer4_out[3249] ^ layer4_out[3250]);
    assign layer5_out[6940] = ~layer4_out[7097];
    assign layer5_out[6941] = layer4_out[6738] ^ layer4_out[6739];
    assign layer5_out[6942] = ~layer4_out[6857] | layer4_out[6858];
    assign layer5_out[6943] = layer4_out[5336] | layer4_out[5337];
    assign layer5_out[6944] = layer4_out[394];
    assign layer5_out[6945] = layer4_out[4773] ^ layer4_out[4774];
    assign layer5_out[6946] = layer4_out[3192] | layer4_out[3193];
    assign layer5_out[6947] = ~layer4_out[239];
    assign layer5_out[6948] = ~layer4_out[223] | layer4_out[224];
    assign layer5_out[6949] = ~layer4_out[4849];
    assign layer5_out[6950] = ~layer4_out[3783];
    assign layer5_out[6951] = layer4_out[4428] ^ layer4_out[4429];
    assign layer5_out[6952] = ~layer4_out[2865];
    assign layer5_out[6953] = ~layer4_out[3701] | layer4_out[3702];
    assign layer5_out[6954] = ~layer4_out[3263];
    assign layer5_out[6955] = ~(layer4_out[7106] & layer4_out[7107]);
    assign layer5_out[6956] = ~layer4_out[2655] | layer4_out[2654];
    assign layer5_out[6957] = ~(layer4_out[2710] & layer4_out[2711]);
    assign layer5_out[6958] = layer4_out[4052] ^ layer4_out[4053];
    assign layer5_out[6959] = ~(layer4_out[455] & layer4_out[456]);
    assign layer5_out[6960] = layer4_out[6347];
    assign layer5_out[6961] = ~layer4_out[1457];
    assign layer5_out[6962] = ~(layer4_out[2920] ^ layer4_out[2921]);
    assign layer5_out[6963] = layer4_out[3170] | layer4_out[3171];
    assign layer5_out[6964] = ~(layer4_out[5752] | layer4_out[5753]);
    assign layer5_out[6965] = ~(layer4_out[353] ^ layer4_out[354]);
    assign layer5_out[6966] = ~layer4_out[2604];
    assign layer5_out[6967] = ~layer4_out[6269];
    assign layer5_out[6968] = layer4_out[2694] | layer4_out[2695];
    assign layer5_out[6969] = layer4_out[1797] & ~layer4_out[1796];
    assign layer5_out[6970] = ~layer4_out[758];
    assign layer5_out[6971] = layer4_out[3077];
    assign layer5_out[6972] = layer4_out[3895] ^ layer4_out[3896];
    assign layer5_out[6973] = ~layer4_out[1002] | layer4_out[1001];
    assign layer5_out[6974] = ~(layer4_out[443] ^ layer4_out[444]);
    assign layer5_out[6975] = ~layer4_out[2439];
    assign layer5_out[6976] = layer4_out[6719] ^ layer4_out[6720];
    assign layer5_out[6977] = layer4_out[4126];
    assign layer5_out[6978] = ~(layer4_out[6774] | layer4_out[6775]);
    assign layer5_out[6979] = layer4_out[607];
    assign layer5_out[6980] = layer4_out[3471] ^ layer4_out[3472];
    assign layer5_out[6981] = layer4_out[3754];
    assign layer5_out[6982] = layer4_out[5174];
    assign layer5_out[6983] = layer4_out[1387];
    assign layer5_out[6984] = ~layer4_out[2676];
    assign layer5_out[6985] = layer4_out[837] ^ layer4_out[838];
    assign layer5_out[6986] = layer4_out[984] & ~layer4_out[983];
    assign layer5_out[6987] = ~(layer4_out[5284] ^ layer4_out[5285]);
    assign layer5_out[6988] = layer4_out[4086];
    assign layer5_out[6989] = layer4_out[5233] | layer4_out[5234];
    assign layer5_out[6990] = ~layer4_out[6709];
    assign layer5_out[6991] = ~layer4_out[4615];
    assign layer5_out[6992] = layer4_out[1646] ^ layer4_out[1647];
    assign layer5_out[6993] = ~(layer4_out[695] ^ layer4_out[696]);
    assign layer5_out[6994] = ~layer4_out[5168];
    assign layer5_out[6995] = ~(layer4_out[3923] ^ layer4_out[3924]);
    assign layer5_out[6996] = ~layer4_out[2756];
    assign layer5_out[6997] = layer4_out[2253] & ~layer4_out[2252];
    assign layer5_out[6998] = layer4_out[2206];
    assign layer5_out[6999] = ~layer4_out[212] | layer4_out[213];
    assign layer5_out[7000] = ~(layer4_out[982] | layer4_out[983]);
    assign layer5_out[7001] = ~(layer4_out[3422] & layer4_out[3423]);
    assign layer5_out[7002] = ~layer4_out[5098];
    assign layer5_out[7003] = ~layer4_out[832];
    assign layer5_out[7004] = layer4_out[6638] | layer4_out[6639];
    assign layer5_out[7005] = ~(layer4_out[4453] ^ layer4_out[4454]);
    assign layer5_out[7006] = ~layer4_out[5235];
    assign layer5_out[7007] = layer4_out[3513];
    assign layer5_out[7008] = ~layer4_out[5397];
    assign layer5_out[7009] = ~(layer4_out[5672] ^ layer4_out[5673]);
    assign layer5_out[7010] = layer4_out[7340] & ~layer4_out[7341];
    assign layer5_out[7011] = layer4_out[6990];
    assign layer5_out[7012] = layer4_out[7221] & layer4_out[7222];
    assign layer5_out[7013] = ~layer4_out[6415];
    assign layer5_out[7014] = ~layer4_out[4908] | layer4_out[4907];
    assign layer5_out[7015] = layer4_out[7884] & ~layer4_out[7883];
    assign layer5_out[7016] = layer4_out[7893];
    assign layer5_out[7017] = ~(layer4_out[2334] ^ layer4_out[2335]);
    assign layer5_out[7018] = ~(layer4_out[4787] ^ layer4_out[4788]);
    assign layer5_out[7019] = layer4_out[5972] ^ layer4_out[5973];
    assign layer5_out[7020] = layer4_out[1552];
    assign layer5_out[7021] = ~layer4_out[5347];
    assign layer5_out[7022] = ~layer4_out[6485];
    assign layer5_out[7023] = layer4_out[1592];
    assign layer5_out[7024] = layer4_out[2615];
    assign layer5_out[7025] = layer4_out[5693] ^ layer4_out[5694];
    assign layer5_out[7026] = ~(layer4_out[5795] & layer4_out[5796]);
    assign layer5_out[7027] = layer4_out[1197] & layer4_out[1198];
    assign layer5_out[7028] = layer4_out[7558];
    assign layer5_out[7029] = ~layer4_out[1367];
    assign layer5_out[7030] = ~(layer4_out[4165] ^ layer4_out[4166]);
    assign layer5_out[7031] = ~(layer4_out[4742] | layer4_out[4743]);
    assign layer5_out[7032] = layer4_out[4969] ^ layer4_out[4970];
    assign layer5_out[7033] = layer4_out[4644];
    assign layer5_out[7034] = ~(layer4_out[7276] ^ layer4_out[7277]);
    assign layer5_out[7035] = ~layer4_out[5666];
    assign layer5_out[7036] = layer4_out[1255];
    assign layer5_out[7037] = layer4_out[5901];
    assign layer5_out[7038] = layer4_out[5188];
    assign layer5_out[7039] = ~layer4_out[7956];
    assign layer5_out[7040] = layer4_out[7297] & ~layer4_out[7298];
    assign layer5_out[7041] = ~(layer4_out[2593] ^ layer4_out[2594]);
    assign layer5_out[7042] = layer4_out[4581];
    assign layer5_out[7043] = ~layer4_out[6394];
    assign layer5_out[7044] = ~layer4_out[4211];
    assign layer5_out[7045] = ~layer4_out[5405];
    assign layer5_out[7046] = ~layer4_out[5049];
    assign layer5_out[7047] = ~layer4_out[1111];
    assign layer5_out[7048] = layer4_out[1666] & ~layer4_out[1667];
    assign layer5_out[7049] = ~layer4_out[4211];
    assign layer5_out[7050] = layer4_out[6965] & ~layer4_out[6966];
    assign layer5_out[7051] = layer4_out[6386] & layer4_out[6387];
    assign layer5_out[7052] = ~(layer4_out[4977] ^ layer4_out[4978]);
    assign layer5_out[7053] = layer4_out[7766];
    assign layer5_out[7054] = ~(layer4_out[2224] ^ layer4_out[2225]);
    assign layer5_out[7055] = layer4_out[2998] & ~layer4_out[2997];
    assign layer5_out[7056] = layer4_out[5863];
    assign layer5_out[7057] = layer4_out[258];
    assign layer5_out[7058] = ~layer4_out[2619];
    assign layer5_out[7059] = ~(layer4_out[7778] ^ layer4_out[7779]);
    assign layer5_out[7060] = layer4_out[4712] ^ layer4_out[4713];
    assign layer5_out[7061] = layer4_out[1108] ^ layer4_out[1109];
    assign layer5_out[7062] = layer4_out[4959];
    assign layer5_out[7063] = layer4_out[7131] & ~layer4_out[7130];
    assign layer5_out[7064] = ~layer4_out[6484];
    assign layer5_out[7065] = layer4_out[6734];
    assign layer5_out[7066] = layer4_out[6964];
    assign layer5_out[7067] = ~(layer4_out[72] ^ layer4_out[73]);
    assign layer5_out[7068] = layer4_out[5824] & ~layer4_out[5823];
    assign layer5_out[7069] = ~(layer4_out[6377] ^ layer4_out[6378]);
    assign layer5_out[7070] = ~(layer4_out[2346] & layer4_out[2347]);
    assign layer5_out[7071] = ~layer4_out[7164];
    assign layer5_out[7072] = ~layer4_out[1091];
    assign layer5_out[7073] = layer4_out[255] ^ layer4_out[256];
    assign layer5_out[7074] = layer4_out[1532] ^ layer4_out[1533];
    assign layer5_out[7075] = ~(layer4_out[6635] & layer4_out[6636]);
    assign layer5_out[7076] = layer4_out[1157] & ~layer4_out[1158];
    assign layer5_out[7077] = ~(layer4_out[204] ^ layer4_out[205]);
    assign layer5_out[7078] = ~(layer4_out[3022] ^ layer4_out[3023]);
    assign layer5_out[7079] = layer4_out[4116];
    assign layer5_out[7080] = layer4_out[5874];
    assign layer5_out[7081] = ~layer4_out[63];
    assign layer5_out[7082] = ~layer4_out[2373];
    assign layer5_out[7083] = layer4_out[5614];
    assign layer5_out[7084] = ~(layer4_out[1394] | layer4_out[1395]);
    assign layer5_out[7085] = layer4_out[6836] ^ layer4_out[6837];
    assign layer5_out[7086] = layer4_out[2782];
    assign layer5_out[7087] = ~layer4_out[2308];
    assign layer5_out[7088] = ~layer4_out[6896] | layer4_out[6897];
    assign layer5_out[7089] = ~(layer4_out[3558] ^ layer4_out[3559]);
    assign layer5_out[7090] = layer4_out[4755] & layer4_out[4756];
    assign layer5_out[7091] = ~layer4_out[3621];
    assign layer5_out[7092] = layer4_out[6125];
    assign layer5_out[7093] = layer4_out[3695] ^ layer4_out[3696];
    assign layer5_out[7094] = layer4_out[2854] & ~layer4_out[2853];
    assign layer5_out[7095] = ~(layer4_out[6539] ^ layer4_out[6540]);
    assign layer5_out[7096] = layer4_out[5416];
    assign layer5_out[7097] = layer4_out[3606];
    assign layer5_out[7098] = ~layer4_out[2639];
    assign layer5_out[7099] = layer4_out[6566];
    assign layer5_out[7100] = layer4_out[7913] ^ layer4_out[7914];
    assign layer5_out[7101] = ~(layer4_out[5654] ^ layer4_out[5655]);
    assign layer5_out[7102] = ~layer4_out[63];
    assign layer5_out[7103] = layer4_out[4901] & ~layer4_out[4900];
    assign layer5_out[7104] = layer4_out[4602];
    assign layer5_out[7105] = layer4_out[7687] & layer4_out[7688];
    assign layer5_out[7106] = layer4_out[149];
    assign layer5_out[7107] = layer4_out[3737];
    assign layer5_out[7108] = ~layer4_out[6301];
    assign layer5_out[7109] = ~layer4_out[7451];
    assign layer5_out[7110] = layer4_out[7237];
    assign layer5_out[7111] = layer4_out[1255];
    assign layer5_out[7112] = ~layer4_out[7505];
    assign layer5_out[7113] = layer4_out[7342];
    assign layer5_out[7114] = layer4_out[3467];
    assign layer5_out[7115] = ~(layer4_out[1400] ^ layer4_out[1401]);
    assign layer5_out[7116] = layer4_out[6685] & ~layer4_out[6686];
    assign layer5_out[7117] = ~(layer4_out[2944] ^ layer4_out[2945]);
    assign layer5_out[7118] = ~(layer4_out[4462] ^ layer4_out[4463]);
    assign layer5_out[7119] = ~(layer4_out[7894] | layer4_out[7895]);
    assign layer5_out[7120] = ~(layer4_out[4522] ^ layer4_out[4523]);
    assign layer5_out[7121] = layer4_out[1989] & ~layer4_out[1988];
    assign layer5_out[7122] = layer4_out[6399];
    assign layer5_out[7123] = layer4_out[1774];
    assign layer5_out[7124] = ~(layer4_out[3653] ^ layer4_out[3654]);
    assign layer5_out[7125] = ~layer4_out[3079];
    assign layer5_out[7126] = ~(layer4_out[649] ^ layer4_out[650]);
    assign layer5_out[7127] = layer4_out[1041] ^ layer4_out[1042];
    assign layer5_out[7128] = ~layer4_out[1367];
    assign layer5_out[7129] = ~layer4_out[2287];
    assign layer5_out[7130] = ~layer4_out[1265];
    assign layer5_out[7131] = layer4_out[244];
    assign layer5_out[7132] = ~layer4_out[6110];
    assign layer5_out[7133] = layer4_out[729] & ~layer4_out[730];
    assign layer5_out[7134] = layer4_out[1896];
    assign layer5_out[7135] = layer4_out[7286];
    assign layer5_out[7136] = ~(layer4_out[5395] | layer4_out[5396]);
    assign layer5_out[7137] = ~(layer4_out[3309] ^ layer4_out[3310]);
    assign layer5_out[7138] = layer4_out[7556];
    assign layer5_out[7139] = ~layer4_out[3296];
    assign layer5_out[7140] = layer4_out[3788] & ~layer4_out[3789];
    assign layer5_out[7141] = layer4_out[136] & ~layer4_out[135];
    assign layer5_out[7142] = ~layer4_out[5921];
    assign layer5_out[7143] = layer4_out[675] & ~layer4_out[674];
    assign layer5_out[7144] = ~layer4_out[6929];
    assign layer5_out[7145] = layer4_out[5703] | layer4_out[5704];
    assign layer5_out[7146] = ~layer4_out[6461];
    assign layer5_out[7147] = ~layer4_out[158];
    assign layer5_out[7148] = ~layer4_out[2653] | layer4_out[2654];
    assign layer5_out[7149] = ~(layer4_out[7858] ^ layer4_out[7859]);
    assign layer5_out[7150] = layer4_out[7904] & layer4_out[7905];
    assign layer5_out[7151] = layer4_out[3041] ^ layer4_out[3042];
    assign layer5_out[7152] = layer4_out[1274] & ~layer4_out[1275];
    assign layer5_out[7153] = ~(layer4_out[4922] ^ layer4_out[4923]);
    assign layer5_out[7154] = ~(layer4_out[2325] | layer4_out[2326]);
    assign layer5_out[7155] = layer4_out[6154] ^ layer4_out[6155];
    assign layer5_out[7156] = ~(layer4_out[5941] & layer4_out[5942]);
    assign layer5_out[7157] = ~(layer4_out[7616] ^ layer4_out[7617]);
    assign layer5_out[7158] = layer4_out[3216] ^ layer4_out[3217];
    assign layer5_out[7159] = ~(layer4_out[1679] | layer4_out[1680]);
    assign layer5_out[7160] = layer4_out[2022];
    assign layer5_out[7161] = layer4_out[5494];
    assign layer5_out[7162] = layer4_out[5961];
    assign layer5_out[7163] = ~layer4_out[932];
    assign layer5_out[7164] = ~(layer4_out[4648] ^ layer4_out[4649]);
    assign layer5_out[7165] = ~(layer4_out[874] ^ layer4_out[875]);
    assign layer5_out[7166] = layer4_out[7879] ^ layer4_out[7880];
    assign layer5_out[7167] = layer4_out[5967] & layer4_out[5968];
    assign layer5_out[7168] = layer4_out[2236];
    assign layer5_out[7169] = ~layer4_out[2331];
    assign layer5_out[7170] = ~layer4_out[5288];
    assign layer5_out[7171] = layer4_out[7848] ^ layer4_out[7849];
    assign layer5_out[7172] = ~layer4_out[7328] | layer4_out[7329];
    assign layer5_out[7173] = ~(layer4_out[3592] | layer4_out[3593]);
    assign layer5_out[7174] = ~(layer4_out[1461] ^ layer4_out[1462]);
    assign layer5_out[7175] = ~(layer4_out[4328] & layer4_out[4329]);
    assign layer5_out[7176] = layer4_out[6455] ^ layer4_out[6456];
    assign layer5_out[7177] = layer4_out[2329];
    assign layer5_out[7178] = layer4_out[3174] & layer4_out[3175];
    assign layer5_out[7179] = layer4_out[6664];
    assign layer5_out[7180] = layer4_out[3022];
    assign layer5_out[7181] = ~(layer4_out[2898] ^ layer4_out[2899]);
    assign layer5_out[7182] = layer4_out[1445];
    assign layer5_out[7183] = ~(layer4_out[6171] ^ layer4_out[6172]);
    assign layer5_out[7184] = ~(layer4_out[4882] ^ layer4_out[4883]);
    assign layer5_out[7185] = layer4_out[3424];
    assign layer5_out[7186] = ~layer4_out[994];
    assign layer5_out[7187] = layer4_out[1488];
    assign layer5_out[7188] = layer4_out[2952];
    assign layer5_out[7189] = ~layer4_out[1670] | layer4_out[1671];
    assign layer5_out[7190] = layer4_out[7286];
    assign layer5_out[7191] = ~layer4_out[4321] | layer4_out[4322];
    assign layer5_out[7192] = ~layer4_out[5002] | layer4_out[5001];
    assign layer5_out[7193] = ~(layer4_out[5593] ^ layer4_out[5594]);
    assign layer5_out[7194] = ~layer4_out[1860];
    assign layer5_out[7195] = ~layer4_out[7446];
    assign layer5_out[7196] = ~(layer4_out[7310] ^ layer4_out[7311]);
    assign layer5_out[7197] = ~(layer4_out[6691] ^ layer4_out[6692]);
    assign layer5_out[7198] = ~(layer4_out[6144] ^ layer4_out[6145]);
    assign layer5_out[7199] = ~(layer4_out[2644] ^ layer4_out[2645]);
    assign layer5_out[7200] = layer4_out[497] & ~layer4_out[498];
    assign layer5_out[7201] = ~layer4_out[4256];
    assign layer5_out[7202] = ~(layer4_out[7440] & layer4_out[7441]);
    assign layer5_out[7203] = layer4_out[7252];
    assign layer5_out[7204] = ~(layer4_out[5501] | layer4_out[5502]);
    assign layer5_out[7205] = ~(layer4_out[2662] ^ layer4_out[2663]);
    assign layer5_out[7206] = layer4_out[5566] | layer4_out[5567];
    assign layer5_out[7207] = ~layer4_out[1552];
    assign layer5_out[7208] = layer4_out[6986] ^ layer4_out[6987];
    assign layer5_out[7209] = layer4_out[1639];
    assign layer5_out[7210] = ~(layer4_out[7233] ^ layer4_out[7234]);
    assign layer5_out[7211] = ~layer4_out[5871];
    assign layer5_out[7212] = ~(layer4_out[809] | layer4_out[810]);
    assign layer5_out[7213] = layer4_out[4092] ^ layer4_out[4093];
    assign layer5_out[7214] = ~layer4_out[5329];
    assign layer5_out[7215] = ~(layer4_out[2351] & layer4_out[2352]);
    assign layer5_out[7216] = layer4_out[5856] & ~layer4_out[5857];
    assign layer5_out[7217] = ~layer4_out[7966];
    assign layer5_out[7218] = ~(layer4_out[4465] ^ layer4_out[4466]);
    assign layer5_out[7219] = ~(layer4_out[1523] & layer4_out[1524]);
    assign layer5_out[7220] = ~layer4_out[6757] | layer4_out[6758];
    assign layer5_out[7221] = ~(layer4_out[7503] ^ layer4_out[7504]);
    assign layer5_out[7222] = ~layer4_out[3370];
    assign layer5_out[7223] = ~(layer4_out[3841] ^ layer4_out[3842]);
    assign layer5_out[7224] = ~layer4_out[3797] | layer4_out[3798];
    assign layer5_out[7225] = layer4_out[1125];
    assign layer5_out[7226] = layer4_out[1318] & ~layer4_out[1317];
    assign layer5_out[7227] = ~(layer4_out[2922] ^ layer4_out[2923]);
    assign layer5_out[7228] = ~layer4_out[7712];
    assign layer5_out[7229] = ~(layer4_out[5726] | layer4_out[5727]);
    assign layer5_out[7230] = ~layer4_out[1078];
    assign layer5_out[7231] = layer4_out[7895] ^ layer4_out[7896];
    assign layer5_out[7232] = ~(layer4_out[314] & layer4_out[315]);
    assign layer5_out[7233] = layer4_out[318];
    assign layer5_out[7234] = layer4_out[6014];
    assign layer5_out[7235] = layer4_out[3218] & ~layer4_out[3219];
    assign layer5_out[7236] = ~layer4_out[7006];
    assign layer5_out[7237] = ~layer4_out[1366];
    assign layer5_out[7238] = layer4_out[4758];
    assign layer5_out[7239] = ~layer4_out[2846];
    assign layer5_out[7240] = layer4_out[402];
    assign layer5_out[7241] = ~(layer4_out[5193] | layer4_out[5194]);
    assign layer5_out[7242] = layer4_out[596] & ~layer4_out[595];
    assign layer5_out[7243] = ~layer4_out[2442];
    assign layer5_out[7244] = layer4_out[1849] & ~layer4_out[1848];
    assign layer5_out[7245] = ~layer4_out[2942];
    assign layer5_out[7246] = layer4_out[3746];
    assign layer5_out[7247] = layer4_out[162] & ~layer4_out[163];
    assign layer5_out[7248] = ~layer4_out[4745];
    assign layer5_out[7249] = layer4_out[4398];
    assign layer5_out[7250] = layer4_out[4912];
    assign layer5_out[7251] = ~layer4_out[7];
    assign layer5_out[7252] = ~layer4_out[7763] | layer4_out[7764];
    assign layer5_out[7253] = ~(layer4_out[4794] | layer4_out[4795]);
    assign layer5_out[7254] = layer4_out[7820];
    assign layer5_out[7255] = layer4_out[7234] | layer4_out[7235];
    assign layer5_out[7256] = layer4_out[1023] & layer4_out[1024];
    assign layer5_out[7257] = ~(layer4_out[2646] & layer4_out[2647]);
    assign layer5_out[7258] = ~(layer4_out[1782] & layer4_out[1783]);
    assign layer5_out[7259] = layer4_out[2419] & ~layer4_out[2418];
    assign layer5_out[7260] = layer4_out[6048] & ~layer4_out[6047];
    assign layer5_out[7261] = layer4_out[2292] | layer4_out[2293];
    assign layer5_out[7262] = ~layer4_out[3900];
    assign layer5_out[7263] = layer4_out[937] & ~layer4_out[936];
    assign layer5_out[7264] = layer4_out[3773] & ~layer4_out[3774];
    assign layer5_out[7265] = ~(layer4_out[4261] ^ layer4_out[4262]);
    assign layer5_out[7266] = layer4_out[1902];
    assign layer5_out[7267] = ~layer4_out[7997] | layer4_out[7998];
    assign layer5_out[7268] = layer4_out[2556] & layer4_out[2557];
    assign layer5_out[7269] = ~(layer4_out[7610] | layer4_out[7611]);
    assign layer5_out[7270] = layer4_out[1685] | layer4_out[1686];
    assign layer5_out[7271] = ~layer4_out[4586];
    assign layer5_out[7272] = ~(layer4_out[4454] | layer4_out[4455]);
    assign layer5_out[7273] = layer4_out[6065] | layer4_out[6066];
    assign layer5_out[7274] = ~(layer4_out[3006] ^ layer4_out[3007]);
    assign layer5_out[7275] = ~layer4_out[752];
    assign layer5_out[7276] = ~layer4_out[4903];
    assign layer5_out[7277] = layer4_out[7144] & ~layer4_out[7145];
    assign layer5_out[7278] = layer4_out[7813] ^ layer4_out[7814];
    assign layer5_out[7279] = layer4_out[3746] & ~layer4_out[3745];
    assign layer5_out[7280] = ~(layer4_out[7453] | layer4_out[7454]);
    assign layer5_out[7281] = ~layer4_out[10];
    assign layer5_out[7282] = ~(layer4_out[4928] ^ layer4_out[4929]);
    assign layer5_out[7283] = ~layer4_out[3542];
    assign layer5_out[7284] = ~layer4_out[6046];
    assign layer5_out[7285] = layer4_out[1592] & ~layer4_out[1591];
    assign layer5_out[7286] = ~(layer4_out[4048] ^ layer4_out[4049]);
    assign layer5_out[7287] = ~(layer4_out[6283] | layer4_out[6284]);
    assign layer5_out[7288] = ~(layer4_out[4182] ^ layer4_out[4183]);
    assign layer5_out[7289] = layer4_out[2134];
    assign layer5_out[7290] = layer4_out[61] & ~layer4_out[60];
    assign layer5_out[7291] = layer4_out[2479];
    assign layer5_out[7292] = ~(layer4_out[7898] ^ layer4_out[7899]);
    assign layer5_out[7293] = ~(layer4_out[3295] ^ layer4_out[3296]);
    assign layer5_out[7294] = layer4_out[7959] ^ layer4_out[7960];
    assign layer5_out[7295] = layer4_out[6714] & layer4_out[6715];
    assign layer5_out[7296] = ~layer4_out[2075];
    assign layer5_out[7297] = ~layer4_out[317] | layer4_out[316];
    assign layer5_out[7298] = layer4_out[5311];
    assign layer5_out[7299] = ~layer4_out[1527];
    assign layer5_out[7300] = ~layer4_out[2412];
    assign layer5_out[7301] = layer4_out[6743] ^ layer4_out[6744];
    assign layer5_out[7302] = layer4_out[7305] & layer4_out[7306];
    assign layer5_out[7303] = layer4_out[709] & layer4_out[710];
    assign layer5_out[7304] = ~layer4_out[3752];
    assign layer5_out[7305] = ~(layer4_out[4334] | layer4_out[4335]);
    assign layer5_out[7306] = ~layer4_out[7258];
    assign layer5_out[7307] = ~layer4_out[2823] | layer4_out[2822];
    assign layer5_out[7308] = ~layer4_out[6938];
    assign layer5_out[7309] = ~layer4_out[5248] | layer4_out[5249];
    assign layer5_out[7310] = layer4_out[4061] & ~layer4_out[4062];
    assign layer5_out[7311] = ~layer4_out[7256];
    assign layer5_out[7312] = layer4_out[5869] ^ layer4_out[5870];
    assign layer5_out[7313] = layer4_out[4673];
    assign layer5_out[7314] = ~(layer4_out[2648] | layer4_out[2649]);
    assign layer5_out[7315] = ~layer4_out[1981];
    assign layer5_out[7316] = ~(layer4_out[7523] ^ layer4_out[7524]);
    assign layer5_out[7317] = layer4_out[6358];
    assign layer5_out[7318] = layer4_out[3331] ^ layer4_out[3332];
    assign layer5_out[7319] = ~(layer4_out[5601] ^ layer4_out[5602]);
    assign layer5_out[7320] = ~(layer4_out[5169] & layer4_out[5170]);
    assign layer5_out[7321] = ~(layer4_out[7733] ^ layer4_out[7734]);
    assign layer5_out[7322] = ~layer4_out[7043];
    assign layer5_out[7323] = layer4_out[6920] ^ layer4_out[6921];
    assign layer5_out[7324] = layer4_out[5107] ^ layer4_out[5108];
    assign layer5_out[7325] = layer4_out[7961] ^ layer4_out[7962];
    assign layer5_out[7326] = layer4_out[7900];
    assign layer5_out[7327] = layer4_out[3912];
    assign layer5_out[7328] = layer4_out[1739] & ~layer4_out[1738];
    assign layer5_out[7329] = ~(layer4_out[7518] | layer4_out[7519]);
    assign layer5_out[7330] = layer4_out[3778] | layer4_out[3779];
    assign layer5_out[7331] = layer4_out[6518] ^ layer4_out[6519];
    assign layer5_out[7332] = ~layer4_out[3240] | layer4_out[3239];
    assign layer5_out[7333] = layer4_out[5278] & ~layer4_out[5277];
    assign layer5_out[7334] = layer4_out[2017] & ~layer4_out[2016];
    assign layer5_out[7335] = ~layer4_out[7512];
    assign layer5_out[7336] = ~layer4_out[3317] | layer4_out[3318];
    assign layer5_out[7337] = layer4_out[4034] & layer4_out[4035];
    assign layer5_out[7338] = layer4_out[4172] & ~layer4_out[4171];
    assign layer5_out[7339] = layer4_out[5997];
    assign layer5_out[7340] = layer4_out[4388];
    assign layer5_out[7341] = ~layer4_out[50];
    assign layer5_out[7342] = layer4_out[7374] & layer4_out[7375];
    assign layer5_out[7343] = ~(layer4_out[691] ^ layer4_out[692]);
    assign layer5_out[7344] = ~layer4_out[626];
    assign layer5_out[7345] = layer4_out[2705];
    assign layer5_out[7346] = ~(layer4_out[203] ^ layer4_out[204]);
    assign layer5_out[7347] = ~layer4_out[2889];
    assign layer5_out[7348] = layer4_out[5885] & ~layer4_out[5886];
    assign layer5_out[7349] = ~layer4_out[6674];
    assign layer5_out[7350] = layer4_out[4581] ^ layer4_out[4582];
    assign layer5_out[7351] = ~layer4_out[4663] | layer4_out[4662];
    assign layer5_out[7352] = ~layer4_out[6164];
    assign layer5_out[7353] = ~layer4_out[6087];
    assign layer5_out[7354] = ~(layer4_out[2887] | layer4_out[2888]);
    assign layer5_out[7355] = layer4_out[2188] ^ layer4_out[2189];
    assign layer5_out[7356] = layer4_out[5579] & ~layer4_out[5578];
    assign layer5_out[7357] = layer4_out[3128];
    assign layer5_out[7358] = layer4_out[2482] ^ layer4_out[2483];
    assign layer5_out[7359] = layer4_out[890] & layer4_out[891];
    assign layer5_out[7360] = layer4_out[5376];
    assign layer5_out[7361] = ~(layer4_out[1802] ^ layer4_out[1803]);
    assign layer5_out[7362] = ~(layer4_out[3869] ^ layer4_out[3870]);
    assign layer5_out[7363] = ~layer4_out[7454];
    assign layer5_out[7364] = layer4_out[6747] ^ layer4_out[6748];
    assign layer5_out[7365] = ~(layer4_out[7030] ^ layer4_out[7031]);
    assign layer5_out[7366] = ~(layer4_out[3187] ^ layer4_out[3188]);
    assign layer5_out[7367] = ~(layer4_out[6808] ^ layer4_out[6809]);
    assign layer5_out[7368] = layer4_out[1300] & layer4_out[1301];
    assign layer5_out[7369] = layer4_out[6036] ^ layer4_out[6037];
    assign layer5_out[7370] = layer4_out[4054] ^ layer4_out[4055];
    assign layer5_out[7371] = ~layer4_out[2755];
    assign layer5_out[7372] = layer4_out[5366];
    assign layer5_out[7373] = layer4_out[1209] ^ layer4_out[1210];
    assign layer5_out[7374] = ~layer4_out[3025];
    assign layer5_out[7375] = ~layer4_out[3011];
    assign layer5_out[7376] = layer4_out[1650] & ~layer4_out[1649];
    assign layer5_out[7377] = ~(layer4_out[6692] ^ layer4_out[6693]);
    assign layer5_out[7378] = ~layer4_out[1022];
    assign layer5_out[7379] = layer4_out[466] & ~layer4_out[465];
    assign layer5_out[7380] = layer4_out[822] | layer4_out[823];
    assign layer5_out[7381] = layer4_out[7984] ^ layer4_out[7985];
    assign layer5_out[7382] = ~(layer4_out[5384] ^ layer4_out[5385]);
    assign layer5_out[7383] = layer4_out[3650] | layer4_out[3651];
    assign layer5_out[7384] = ~layer4_out[3100];
    assign layer5_out[7385] = layer4_out[5511];
    assign layer5_out[7386] = layer4_out[5309];
    assign layer5_out[7387] = layer4_out[4125] & ~layer4_out[4124];
    assign layer5_out[7388] = layer4_out[2242] ^ layer4_out[2243];
    assign layer5_out[7389] = ~layer4_out[5267];
    assign layer5_out[7390] = layer4_out[1757] ^ layer4_out[1758];
    assign layer5_out[7391] = ~(layer4_out[4886] ^ layer4_out[4887]);
    assign layer5_out[7392] = layer4_out[2203];
    assign layer5_out[7393] = layer4_out[4554];
    assign layer5_out[7394] = ~(layer4_out[656] | layer4_out[657]);
    assign layer5_out[7395] = ~layer4_out[7697];
    assign layer5_out[7396] = ~(layer4_out[3451] ^ layer4_out[3452]);
    assign layer5_out[7397] = layer4_out[2283] ^ layer4_out[2284];
    assign layer5_out[7398] = ~layer4_out[6940];
    assign layer5_out[7399] = layer4_out[4967];
    assign layer5_out[7400] = ~(layer4_out[3449] ^ layer4_out[3450]);
    assign layer5_out[7401] = ~(layer4_out[7996] & layer4_out[7997]);
    assign layer5_out[7402] = ~(layer4_out[4422] | layer4_out[4423]);
    assign layer5_out[7403] = layer4_out[1088] & layer4_out[1089];
    assign layer5_out[7404] = ~layer4_out[6513];
    assign layer5_out[7405] = ~(layer4_out[7995] & layer4_out[7996]);
    assign layer5_out[7406] = ~layer4_out[5455];
    assign layer5_out[7407] = ~(layer4_out[4484] & layer4_out[4485]);
    assign layer5_out[7408] = layer4_out[4408] & layer4_out[4409];
    assign layer5_out[7409] = layer4_out[4739] & ~layer4_out[4740];
    assign layer5_out[7410] = layer4_out[6603] ^ layer4_out[6604];
    assign layer5_out[7411] = ~(layer4_out[3527] ^ layer4_out[3528]);
    assign layer5_out[7412] = ~layer4_out[6044];
    assign layer5_out[7413] = ~(layer4_out[4710] | layer4_out[4711]);
    assign layer5_out[7414] = ~layer4_out[3357];
    assign layer5_out[7415] = ~layer4_out[7926];
    assign layer5_out[7416] = layer4_out[7629];
    assign layer5_out[7417] = layer4_out[945] ^ layer4_out[946];
    assign layer5_out[7418] = layer4_out[5197];
    assign layer5_out[7419] = layer4_out[1436] & layer4_out[1437];
    assign layer5_out[7420] = layer4_out[1608] ^ layer4_out[1609];
    assign layer5_out[7421] = layer4_out[6978] & ~layer4_out[6979];
    assign layer5_out[7422] = ~(layer4_out[3909] ^ layer4_out[3910]);
    assign layer5_out[7423] = ~layer4_out[7294];
    assign layer5_out[7424] = ~layer4_out[5329];
    assign layer5_out[7425] = layer4_out[7869] ^ layer4_out[7870];
    assign layer5_out[7426] = layer4_out[3873] ^ layer4_out[3874];
    assign layer5_out[7427] = layer4_out[3135] & ~layer4_out[3134];
    assign layer5_out[7428] = layer4_out[1531] | layer4_out[1532];
    assign layer5_out[7429] = layer4_out[5343];
    assign layer5_out[7430] = ~(layer4_out[1229] ^ layer4_out[1230]);
    assign layer5_out[7431] = ~(layer4_out[4370] ^ layer4_out[4371]);
    assign layer5_out[7432] = ~layer4_out[363];
    assign layer5_out[7433] = layer4_out[3437];
    assign layer5_out[7434] = ~(layer4_out[1519] ^ layer4_out[1520]);
    assign layer5_out[7435] = ~(layer4_out[4687] ^ layer4_out[4688]);
    assign layer5_out[7436] = layer4_out[1881];
    assign layer5_out[7437] = ~(layer4_out[7170] & layer4_out[7171]);
    assign layer5_out[7438] = layer4_out[6260] & layer4_out[6261];
    assign layer5_out[7439] = layer4_out[3597] | layer4_out[3598];
    assign layer5_out[7440] = layer4_out[5984] | layer4_out[5985];
    assign layer5_out[7441] = layer4_out[557];
    assign layer5_out[7442] = layer4_out[2809];
    assign layer5_out[7443] = layer4_out[2393] ^ layer4_out[2394];
    assign layer5_out[7444] = layer4_out[2854] & ~layer4_out[2855];
    assign layer5_out[7445] = layer4_out[2928];
    assign layer5_out[7446] = ~layer4_out[5524];
    assign layer5_out[7447] = layer4_out[2588];
    assign layer5_out[7448] = ~layer4_out[3629];
    assign layer5_out[7449] = layer4_out[7785] ^ layer4_out[7786];
    assign layer5_out[7450] = layer4_out[2264] ^ layer4_out[2265];
    assign layer5_out[7451] = layer4_out[3337] ^ layer4_out[3338];
    assign layer5_out[7452] = layer4_out[1606];
    assign layer5_out[7453] = ~(layer4_out[4697] | layer4_out[4698]);
    assign layer5_out[7454] = ~(layer4_out[1907] ^ layer4_out[1908]);
    assign layer5_out[7455] = ~layer4_out[6839];
    assign layer5_out[7456] = ~(layer4_out[4915] ^ layer4_out[4916]);
    assign layer5_out[7457] = ~layer4_out[3476];
    assign layer5_out[7458] = ~layer4_out[1981];
    assign layer5_out[7459] = ~layer4_out[1391];
    assign layer5_out[7460] = layer4_out[618] ^ layer4_out[619];
    assign layer5_out[7461] = layer4_out[3847];
    assign layer5_out[7462] = layer4_out[3004];
    assign layer5_out[7463] = layer4_out[7018] & layer4_out[7019];
    assign layer5_out[7464] = layer4_out[1294];
    assign layer5_out[7465] = layer4_out[7779] ^ layer4_out[7780];
    assign layer5_out[7466] = layer4_out[3456] & ~layer4_out[3457];
    assign layer5_out[7467] = ~layer4_out[2068];
    assign layer5_out[7468] = ~layer4_out[1407];
    assign layer5_out[7469] = layer4_out[3353];
    assign layer5_out[7470] = ~layer4_out[210];
    assign layer5_out[7471] = layer4_out[254] ^ layer4_out[255];
    assign layer5_out[7472] = ~(layer4_out[2641] ^ layer4_out[2642]);
    assign layer5_out[7473] = ~layer4_out[1026];
    assign layer5_out[7474] = layer4_out[2872];
    assign layer5_out[7475] = layer4_out[7456];
    assign layer5_out[7476] = layer4_out[1060] ^ layer4_out[1061];
    assign layer5_out[7477] = layer4_out[1515];
    assign layer5_out[7478] = layer4_out[7317] & layer4_out[7318];
    assign layer5_out[7479] = layer4_out[150] & ~layer4_out[149];
    assign layer5_out[7480] = layer4_out[4474] & ~layer4_out[4475];
    assign layer5_out[7481] = ~(layer4_out[1469] ^ layer4_out[1470]);
    assign layer5_out[7482] = layer4_out[7531];
    assign layer5_out[7483] = layer4_out[3104];
    assign layer5_out[7484] = ~(layer4_out[4876] ^ layer4_out[4877]);
    assign layer5_out[7485] = layer4_out[1473];
    assign layer5_out[7486] = layer4_out[4780];
    assign layer5_out[7487] = layer4_out[2465];
    assign layer5_out[7488] = ~layer4_out[3529] | layer4_out[3530];
    assign layer5_out[7489] = layer4_out[6012];
    assign layer5_out[7490] = layer4_out[215];
    assign layer5_out[7491] = ~(layer4_out[3513] | layer4_out[3514]);
    assign layer5_out[7492] = ~layer4_out[7801];
    assign layer5_out[7493] = ~layer4_out[5896];
    assign layer5_out[7494] = layer4_out[36] ^ layer4_out[37];
    assign layer5_out[7495] = layer4_out[7128] & layer4_out[7129];
    assign layer5_out[7496] = layer4_out[2487] & ~layer4_out[2488];
    assign layer5_out[7497] = layer4_out[1585];
    assign layer5_out[7498] = layer4_out[2008] & ~layer4_out[2009];
    assign layer5_out[7499] = ~layer4_out[6777];
    assign layer5_out[7500] = ~(layer4_out[676] | layer4_out[677]);
    assign layer5_out[7501] = layer4_out[2778] & ~layer4_out[2777];
    assign layer5_out[7502] = layer4_out[1067];
    assign layer5_out[7503] = ~(layer4_out[582] ^ layer4_out[583]);
    assign layer5_out[7504] = layer4_out[7468];
    assign layer5_out[7505] = layer4_out[7908];
    assign layer5_out[7506] = ~layer4_out[6344] | layer4_out[6345];
    assign layer5_out[7507] = layer4_out[348];
    assign layer5_out[7508] = layer4_out[303] & ~layer4_out[302];
    assign layer5_out[7509] = layer4_out[1268];
    assign layer5_out[7510] = layer4_out[2333] ^ layer4_out[2334];
    assign layer5_out[7511] = ~layer4_out[2752];
    assign layer5_out[7512] = ~layer4_out[6876];
    assign layer5_out[7513] = layer4_out[7255];
    assign layer5_out[7514] = ~layer4_out[2460];
    assign layer5_out[7515] = ~layer4_out[1173];
    assign layer5_out[7516] = ~(layer4_out[854] & layer4_out[855]);
    assign layer5_out[7517] = layer4_out[2383] ^ layer4_out[2384];
    assign layer5_out[7518] = layer4_out[5732] | layer4_out[5733];
    assign layer5_out[7519] = ~layer4_out[6334];
    assign layer5_out[7520] = ~layer4_out[2448];
    assign layer5_out[7521] = ~layer4_out[2274];
    assign layer5_out[7522] = ~(layer4_out[7500] & layer4_out[7501]);
    assign layer5_out[7523] = ~layer4_out[5259];
    assign layer5_out[7524] = layer4_out[88] & layer4_out[89];
    assign layer5_out[7525] = ~layer4_out[6408];
    assign layer5_out[7526] = layer4_out[7433] & ~layer4_out[7434];
    assign layer5_out[7527] = layer4_out[7210];
    assign layer5_out[7528] = ~layer4_out[6697];
    assign layer5_out[7529] = ~layer4_out[3632];
    assign layer5_out[7530] = ~(layer4_out[1702] ^ layer4_out[1703]);
    assign layer5_out[7531] = layer4_out[7521];
    assign layer5_out[7532] = ~layer4_out[5851];
    assign layer5_out[7533] = ~layer4_out[6262];
    assign layer5_out[7534] = layer4_out[5388] ^ layer4_out[5389];
    assign layer5_out[7535] = layer4_out[894] ^ layer4_out[895];
    assign layer5_out[7536] = layer4_out[5798];
    assign layer5_out[7537] = layer4_out[3697] & ~layer4_out[3696];
    assign layer5_out[7538] = ~(layer4_out[2681] ^ layer4_out[2682]);
    assign layer5_out[7539] = layer4_out[999] ^ layer4_out[1000];
    assign layer5_out[7540] = layer4_out[3297];
    assign layer5_out[7541] = layer4_out[6281] ^ layer4_out[6282];
    assign layer5_out[7542] = layer4_out[475];
    assign layer5_out[7543] = layer4_out[3704];
    assign layer5_out[7544] = layer4_out[5585] & ~layer4_out[5584];
    assign layer5_out[7545] = ~layer4_out[5969];
    assign layer5_out[7546] = layer4_out[3012];
    assign layer5_out[7547] = ~layer4_out[995];
    assign layer5_out[7548] = ~layer4_out[2985];
    assign layer5_out[7549] = layer4_out[5708] | layer4_out[5709];
    assign layer5_out[7550] = layer4_out[3526];
    assign layer5_out[7551] = ~layer4_out[7522] | layer4_out[7523];
    assign layer5_out[7552] = ~(layer4_out[5802] | layer4_out[5803]);
    assign layer5_out[7553] = layer4_out[6562];
    assign layer5_out[7554] = layer4_out[4039] & ~layer4_out[4040];
    assign layer5_out[7555] = ~(layer4_out[3029] ^ layer4_out[3030]);
    assign layer5_out[7556] = ~layer4_out[4158];
    assign layer5_out[7557] = ~layer4_out[462];
    assign layer5_out[7558] = layer4_out[2474] & layer4_out[2475];
    assign layer5_out[7559] = layer4_out[5420];
    assign layer5_out[7560] = layer4_out[4730];
    assign layer5_out[7561] = layer4_out[4343] & ~layer4_out[4344];
    assign layer5_out[7562] = ~(layer4_out[768] ^ layer4_out[769]);
    assign layer5_out[7563] = layer4_out[5700];
    assign layer5_out[7564] = layer4_out[3490] ^ layer4_out[3491];
    assign layer5_out[7565] = layer4_out[5003] & ~layer4_out[5004];
    assign layer5_out[7566] = ~(layer4_out[6804] ^ layer4_out[6805]);
    assign layer5_out[7567] = layer4_out[2025] & ~layer4_out[2024];
    assign layer5_out[7568] = ~(layer4_out[6829] | layer4_out[6830]);
    assign layer5_out[7569] = ~layer4_out[3812];
    assign layer5_out[7570] = layer4_out[1750] ^ layer4_out[1751];
    assign layer5_out[7571] = layer4_out[2968] ^ layer4_out[2969];
    assign layer5_out[7572] = layer4_out[3728];
    assign layer5_out[7573] = layer4_out[6277] | layer4_out[6278];
    assign layer5_out[7574] = layer4_out[2903];
    assign layer5_out[7575] = ~(layer4_out[1698] ^ layer4_out[1699]);
    assign layer5_out[7576] = layer4_out[3458] & ~layer4_out[3457];
    assign layer5_out[7577] = layer4_out[2900] | layer4_out[2901];
    assign layer5_out[7578] = ~(layer4_out[540] | layer4_out[541]);
    assign layer5_out[7579] = layer4_out[593] ^ layer4_out[594];
    assign layer5_out[7580] = ~(layer4_out[2851] ^ layer4_out[2852]);
    assign layer5_out[7581] = ~layer4_out[6209] | layer4_out[6210];
    assign layer5_out[7582] = ~layer4_out[5435];
    assign layer5_out[7583] = ~layer4_out[3500];
    assign layer5_out[7584] = layer4_out[5376];
    assign layer5_out[7585] = ~layer4_out[5691];
    assign layer5_out[7586] = ~(layer4_out[4163] ^ layer4_out[4164]);
    assign layer5_out[7587] = layer4_out[6733] ^ layer4_out[6734];
    assign layer5_out[7588] = layer4_out[5648] & ~layer4_out[5649];
    assign layer5_out[7589] = ~layer4_out[4843];
    assign layer5_out[7590] = ~layer4_out[3960];
    assign layer5_out[7591] = layer4_out[2586];
    assign layer5_out[7592] = layer4_out[478];
    assign layer5_out[7593] = layer4_out[1761] | layer4_out[1762];
    assign layer5_out[7594] = layer4_out[948];
    assign layer5_out[7595] = layer4_out[7261] | layer4_out[7262];
    assign layer5_out[7596] = ~layer4_out[2643];
    assign layer5_out[7597] = layer4_out[5420];
    assign layer5_out[7598] = ~layer4_out[5541];
    assign layer5_out[7599] = ~(layer4_out[7704] ^ layer4_out[7705]);
    assign layer5_out[7600] = layer4_out[5100] | layer4_out[5101];
    assign layer5_out[7601] = layer4_out[2353];
    assign layer5_out[7602] = layer4_out[6495] ^ layer4_out[6496];
    assign layer5_out[7603] = layer4_out[4320] & layer4_out[4321];
    assign layer5_out[7604] = layer4_out[2578];
    assign layer5_out[7605] = ~(layer4_out[6796] ^ layer4_out[6797]);
    assign layer5_out[7606] = layer4_out[4867] & ~layer4_out[4868];
    assign layer5_out[7607] = ~(layer4_out[6900] ^ layer4_out[6901]);
    assign layer5_out[7608] = ~(layer4_out[3826] ^ layer4_out[3827]);
    assign layer5_out[7609] = layer4_out[6542] & ~layer4_out[6541];
    assign layer5_out[7610] = layer4_out[7371] & ~layer4_out[7370];
    assign layer5_out[7611] = ~layer4_out[7736];
    assign layer5_out[7612] = layer4_out[4619] ^ layer4_out[4620];
    assign layer5_out[7613] = layer4_out[4146] & layer4_out[4147];
    assign layer5_out[7614] = layer4_out[3783];
    assign layer5_out[7615] = layer4_out[4639];
    assign layer5_out[7616] = ~(layer4_out[6628] ^ layer4_out[6629]);
    assign layer5_out[7617] = layer4_out[3704] & ~layer4_out[3703];
    assign layer5_out[7618] = layer4_out[5103];
    assign layer5_out[7619] = layer4_out[6193] & ~layer4_out[6192];
    assign layer5_out[7620] = layer4_out[6274] | layer4_out[6275];
    assign layer5_out[7621] = ~(layer4_out[2909] ^ layer4_out[2910]);
    assign layer5_out[7622] = ~layer4_out[3908] | layer4_out[3909];
    assign layer5_out[7623] = layer4_out[4082] & ~layer4_out[4083];
    assign layer5_out[7624] = ~layer4_out[6314];
    assign layer5_out[7625] = layer4_out[689] ^ layer4_out[690];
    assign layer5_out[7626] = ~(layer4_out[2918] ^ layer4_out[2919]);
    assign layer5_out[7627] = layer4_out[345] ^ layer4_out[346];
    assign layer5_out[7628] = ~(layer4_out[3647] | layer4_out[3648]);
    assign layer5_out[7629] = ~(layer4_out[6893] ^ layer4_out[6894]);
    assign layer5_out[7630] = layer4_out[6977] & layer4_out[6978];
    assign layer5_out[7631] = ~(layer4_out[1241] & layer4_out[1242]);
    assign layer5_out[7632] = ~layer4_out[855];
    assign layer5_out[7633] = ~layer4_out[5780];
    assign layer5_out[7634] = layer4_out[700] & ~layer4_out[699];
    assign layer5_out[7635] = layer4_out[240];
    assign layer5_out[7636] = ~layer4_out[5958];
    assign layer5_out[7637] = layer4_out[6686] | layer4_out[6687];
    assign layer5_out[7638] = ~layer4_out[5833];
    assign layer5_out[7639] = ~layer4_out[7084];
    assign layer5_out[7640] = ~(layer4_out[1904] | layer4_out[1905]);
    assign layer5_out[7641] = layer4_out[643];
    assign layer5_out[7642] = layer4_out[336] ^ layer4_out[337];
    assign layer5_out[7643] = ~layer4_out[5010];
    assign layer5_out[7644] = ~layer4_out[5891];
    assign layer5_out[7645] = layer4_out[912] ^ layer4_out[913];
    assign layer5_out[7646] = ~layer4_out[3061];
    assign layer5_out[7647] = ~(layer4_out[820] | layer4_out[821]);
    assign layer5_out[7648] = ~layer4_out[719];
    assign layer5_out[7649] = layer4_out[1695];
    assign layer5_out[7650] = ~(layer4_out[6397] ^ layer4_out[6398]);
    assign layer5_out[7651] = layer4_out[3867];
    assign layer5_out[7652] = ~(layer4_out[2730] ^ layer4_out[2731]);
    assign layer5_out[7653] = layer4_out[5400];
    assign layer5_out[7654] = layer4_out[5464] ^ layer4_out[5465];
    assign layer5_out[7655] = layer4_out[6000];
    assign layer5_out[7656] = ~layer4_out[2716];
    assign layer5_out[7657] = layer4_out[3116] | layer4_out[3117];
    assign layer5_out[7658] = ~(layer4_out[1470] ^ layer4_out[1471]);
    assign layer5_out[7659] = layer4_out[2203];
    assign layer5_out[7660] = ~layer4_out[4854] | layer4_out[4855];
    assign layer5_out[7661] = ~(layer4_out[7292] ^ layer4_out[7293]);
    assign layer5_out[7662] = layer4_out[6645];
    assign layer5_out[7663] = layer4_out[4003] ^ layer4_out[4004];
    assign layer5_out[7664] = layer4_out[3012] & ~layer4_out[3011];
    assign layer5_out[7665] = ~(layer4_out[5096] | layer4_out[5097]);
    assign layer5_out[7666] = layer4_out[220] ^ layer4_out[221];
    assign layer5_out[7667] = layer4_out[6065];
    assign layer5_out[7668] = ~layer4_out[1918] | layer4_out[1919];
    assign layer5_out[7669] = layer4_out[3353];
    assign layer5_out[7670] = ~layer4_out[943];
    assign layer5_out[7671] = ~(layer4_out[383] | layer4_out[384]);
    assign layer5_out[7672] = layer4_out[5280] ^ layer4_out[5281];
    assign layer5_out[7673] = ~(layer4_out[7573] ^ layer4_out[7574]);
    assign layer5_out[7674] = layer4_out[1709] ^ layer4_out[1710];
    assign layer5_out[7675] = ~layer4_out[1277];
    assign layer5_out[7676] = ~(layer4_out[7889] ^ layer4_out[7890]);
    assign layer5_out[7677] = ~(layer4_out[7378] ^ layer4_out[7379]);
    assign layer5_out[7678] = layer4_out[7493];
    assign layer5_out[7679] = ~layer4_out[4045] | layer4_out[4046];
    assign layer5_out[7680] = layer4_out[6835] & layer4_out[6836];
    assign layer5_out[7681] = layer4_out[1007];
    assign layer5_out[7682] = ~(layer4_out[3669] ^ layer4_out[3670]);
    assign layer5_out[7683] = ~(layer4_out[11] ^ layer4_out[12]);
    assign layer5_out[7684] = ~(layer4_out[2042] & layer4_out[2043]);
    assign layer5_out[7685] = layer4_out[3843] ^ layer4_out[3844];
    assign layer5_out[7686] = ~layer4_out[2949];
    assign layer5_out[7687] = ~(layer4_out[6102] | layer4_out[6103]);
    assign layer5_out[7688] = layer4_out[2308];
    assign layer5_out[7689] = layer4_out[1963];
    assign layer5_out[7690] = ~(layer4_out[2769] | layer4_out[2770]);
    assign layer5_out[7691] = layer4_out[5286];
    assign layer5_out[7692] = layer4_out[1515];
    assign layer5_out[7693] = layer4_out[5767] & layer4_out[5768];
    assign layer5_out[7694] = layer4_out[5141] & layer4_out[5142];
    assign layer5_out[7695] = ~(layer4_out[7412] & layer4_out[7413]);
    assign layer5_out[7696] = layer4_out[7326] | layer4_out[7327];
    assign layer5_out[7697] = ~layer4_out[1020];
    assign layer5_out[7698] = layer4_out[2856] ^ layer4_out[2857];
    assign layer5_out[7699] = layer4_out[926] ^ layer4_out[927];
    assign layer5_out[7700] = ~layer4_out[1867];
    assign layer5_out[7701] = ~(layer4_out[1166] & layer4_out[1167]);
    assign layer5_out[7702] = ~layer4_out[7153];
    assign layer5_out[7703] = layer4_out[7018] & ~layer4_out[7017];
    assign layer5_out[7704] = layer4_out[2449] ^ layer4_out[2450];
    assign layer5_out[7705] = ~layer4_out[4070];
    assign layer5_out[7706] = layer4_out[683] & layer4_out[684];
    assign layer5_out[7707] = ~layer4_out[1383];
    assign layer5_out[7708] = ~(layer4_out[7694] ^ layer4_out[7695]);
    assign layer5_out[7709] = ~(layer4_out[7596] & layer4_out[7597]);
    assign layer5_out[7710] = ~layer4_out[3838];
    assign layer5_out[7711] = ~(layer4_out[5053] | layer4_out[5054]);
    assign layer5_out[7712] = ~layer4_out[2261] | layer4_out[2262];
    assign layer5_out[7713] = ~layer4_out[3712] | layer4_out[3713];
    assign layer5_out[7714] = layer4_out[1361];
    assign layer5_out[7715] = layer4_out[920] & layer4_out[921];
    assign layer5_out[7716] = layer4_out[6569];
    assign layer5_out[7717] = ~(layer4_out[7232] ^ layer4_out[7233]);
    assign layer5_out[7718] = layer4_out[4645];
    assign layer5_out[7719] = ~(layer4_out[7011] ^ layer4_out[7012]);
    assign layer5_out[7720] = layer4_out[7447] | layer4_out[7448];
    assign layer5_out[7721] = ~layer4_out[6273];
    assign layer5_out[7722] = ~layer4_out[7133];
    assign layer5_out[7723] = layer4_out[7982] & ~layer4_out[7981];
    assign layer5_out[7724] = ~(layer4_out[1179] | layer4_out[1180]);
    assign layer5_out[7725] = ~layer4_out[7769];
    assign layer5_out[7726] = ~layer4_out[3089];
    assign layer5_out[7727] = ~layer4_out[3174] | layer4_out[3173];
    assign layer5_out[7728] = ~layer4_out[2180] | layer4_out[2179];
    assign layer5_out[7729] = layer4_out[3437] | layer4_out[3438];
    assign layer5_out[7730] = layer4_out[985] & layer4_out[986];
    assign layer5_out[7731] = layer4_out[1493] & layer4_out[1494];
    assign layer5_out[7732] = layer4_out[7149] | layer4_out[7150];
    assign layer5_out[7733] = layer4_out[7012] & layer4_out[7013];
    assign layer5_out[7734] = layer4_out[5037];
    assign layer5_out[7735] = layer4_out[5218];
    assign layer5_out[7736] = layer4_out[2011] ^ layer4_out[2012];
    assign layer5_out[7737] = ~layer4_out[905];
    assign layer5_out[7738] = ~(layer4_out[4118] | layer4_out[4119]);
    assign layer5_out[7739] = layer4_out[6321];
    assign layer5_out[7740] = ~(layer4_out[4186] | layer4_out[4187]);
    assign layer5_out[7741] = ~layer4_out[3149];
    assign layer5_out[7742] = layer4_out[4738] & layer4_out[4739];
    assign layer5_out[7743] = layer4_out[1410] ^ layer4_out[1411];
    assign layer5_out[7744] = ~(layer4_out[7196] | layer4_out[7197]);
    assign layer5_out[7745] = ~layer4_out[4437];
    assign layer5_out[7746] = ~(layer4_out[7033] | layer4_out[7034]);
    assign layer5_out[7747] = layer4_out[7218] & layer4_out[7219];
    assign layer5_out[7748] = ~layer4_out[3089];
    assign layer5_out[7749] = ~(layer4_out[6446] ^ layer4_out[6447]);
    assign layer5_out[7750] = layer4_out[1538] & ~layer4_out[1539];
    assign layer5_out[7751] = layer4_out[994];
    assign layer5_out[7752] = layer4_out[5626];
    assign layer5_out[7753] = ~layer4_out[2361];
    assign layer5_out[7754] = ~layer4_out[5787] | layer4_out[5788];
    assign layer5_out[7755] = layer4_out[221];
    assign layer5_out[7756] = ~(layer4_out[7043] & layer4_out[7044]);
    assign layer5_out[7757] = ~(layer4_out[6325] ^ layer4_out[6326]);
    assign layer5_out[7758] = ~layer4_out[3177];
    assign layer5_out[7759] = ~(layer4_out[5620] ^ layer4_out[5621]);
    assign layer5_out[7760] = layer4_out[339];
    assign layer5_out[7761] = ~(layer4_out[2785] ^ layer4_out[2786]);
    assign layer5_out[7762] = ~(layer4_out[1808] ^ layer4_out[1809]);
    assign layer5_out[7763] = layer4_out[5507] & layer4_out[5508];
    assign layer5_out[7764] = ~(layer4_out[2855] & layer4_out[2856]);
    assign layer5_out[7765] = layer4_out[2591] & layer4_out[2592];
    assign layer5_out[7766] = ~layer4_out[210];
    assign layer5_out[7767] = layer4_out[6247] ^ layer4_out[6248];
    assign layer5_out[7768] = ~layer4_out[7040] | layer4_out[7041];
    assign layer5_out[7769] = layer4_out[3495] & layer4_out[3496];
    assign layer5_out[7770] = layer4_out[4098] ^ layer4_out[4099];
    assign layer5_out[7771] = layer4_out[2664] & ~layer4_out[2665];
    assign layer5_out[7772] = ~layer4_out[2185];
    assign layer5_out[7773] = layer4_out[4487] & ~layer4_out[4488];
    assign layer5_out[7774] = layer4_out[3246] & ~layer4_out[3245];
    assign layer5_out[7775] = ~(layer4_out[4809] | layer4_out[4810]);
    assign layer5_out[7776] = ~layer4_out[6344] | layer4_out[6343];
    assign layer5_out[7777] = ~layer4_out[1337] | layer4_out[1336];
    assign layer5_out[7778] = layer4_out[1881];
    assign layer5_out[7779] = layer4_out[1774];
    assign layer5_out[7780] = layer4_out[6690] & ~layer4_out[6691];
    assign layer5_out[7781] = ~(layer4_out[2354] ^ layer4_out[2355]);
    assign layer5_out[7782] = ~layer4_out[3179];
    assign layer5_out[7783] = ~layer4_out[5943] | layer4_out[5944];
    assign layer5_out[7784] = layer4_out[2390];
    assign layer5_out[7785] = layer4_out[4532] & ~layer4_out[4533];
    assign layer5_out[7786] = layer4_out[2263] & layer4_out[2264];
    assign layer5_out[7787] = layer4_out[545];
    assign layer5_out[7788] = ~(layer4_out[5599] ^ layer4_out[5600]);
    assign layer5_out[7789] = layer4_out[4497] ^ layer4_out[4498];
    assign layer5_out[7790] = layer4_out[5931];
    assign layer5_out[7791] = layer4_out[3983] ^ layer4_out[3984];
    assign layer5_out[7792] = layer4_out[2575] & layer4_out[2576];
    assign layer5_out[7793] = layer4_out[893];
    assign layer5_out[7794] = ~(layer4_out[3231] ^ layer4_out[3232]);
    assign layer5_out[7795] = layer4_out[5702];
    assign layer5_out[7796] = layer4_out[5902];
    assign layer5_out[7797] = ~layer4_out[5806];
    assign layer5_out[7798] = layer4_out[661];
    assign layer5_out[7799] = ~layer4_out[853];
    assign layer5_out[7800] = ~layer4_out[3242] | layer4_out[3243];
    assign layer5_out[7801] = ~layer4_out[5383];
    assign layer5_out[7802] = layer4_out[2174];
    assign layer5_out[7803] = layer4_out[1941];
    assign layer5_out[7804] = ~(layer4_out[7925] | layer4_out[7926]);
    assign layer5_out[7805] = layer4_out[3570];
    assign layer5_out[7806] = ~layer4_out[3982];
    assign layer5_out[7807] = ~layer4_out[6889];
    assign layer5_out[7808] = ~layer4_out[7615] | layer4_out[7616];
    assign layer5_out[7809] = layer4_out[180];
    assign layer5_out[7810] = layer4_out[3719];
    assign layer5_out[7811] = ~layer4_out[671];
    assign layer5_out[7812] = ~layer4_out[3712];
    assign layer5_out[7813] = ~layer4_out[4482] | layer4_out[4481];
    assign layer5_out[7814] = ~layer4_out[7499];
    assign layer5_out[7815] = layer4_out[3794];
    assign layer5_out[7816] = layer4_out[7649];
    assign layer5_out[7817] = layer4_out[7979] & layer4_out[7980];
    assign layer5_out[7818] = ~layer4_out[3383];
    assign layer5_out[7819] = ~layer4_out[4957];
    assign layer5_out[7820] = layer4_out[5205];
    assign layer5_out[7821] = ~layer4_out[1138];
    assign layer5_out[7822] = layer4_out[1448];
    assign layer5_out[7823] = layer4_out[5211];
    assign layer5_out[7824] = ~(layer4_out[4293] ^ layer4_out[4294]);
    assign layer5_out[7825] = layer4_out[775] & layer4_out[776];
    assign layer5_out[7826] = layer4_out[6533];
    assign layer5_out[7827] = layer4_out[5441];
    assign layer5_out[7828] = ~(layer4_out[5379] & layer4_out[5380]);
    assign layer5_out[7829] = ~layer4_out[6483];
    assign layer5_out[7830] = layer4_out[5045];
    assign layer5_out[7831] = layer4_out[7367] ^ layer4_out[7368];
    assign layer5_out[7832] = layer4_out[1479] & ~layer4_out[1478];
    assign layer5_out[7833] = ~(layer4_out[6646] | layer4_out[6647]);
    assign layer5_out[7834] = ~layer4_out[4096];
    assign layer5_out[7835] = layer4_out[5765];
    assign layer5_out[7836] = layer4_out[707];
    assign layer5_out[7837] = layer4_out[4939];
    assign layer5_out[7838] = ~(layer4_out[7067] ^ layer4_out[7068]);
    assign layer5_out[7839] = ~layer4_out[1859];
    assign layer5_out[7840] = layer4_out[5879] ^ layer4_out[5880];
    assign layer5_out[7841] = layer4_out[7687] & ~layer4_out[7686];
    assign layer5_out[7842] = ~(layer4_out[4289] | layer4_out[4290]);
    assign layer5_out[7843] = ~layer4_out[2749];
    assign layer5_out[7844] = layer4_out[6433] ^ layer4_out[6434];
    assign layer5_out[7845] = ~layer4_out[7258];
    assign layer5_out[7846] = layer4_out[5370] & ~layer4_out[5369];
    assign layer5_out[7847] = ~layer4_out[6990];
    assign layer5_out[7848] = ~layer4_out[6197];
    assign layer5_out[7849] = layer4_out[6554];
    assign layer5_out[7850] = ~(layer4_out[987] | layer4_out[988]);
    assign layer5_out[7851] = ~layer4_out[766];
    assign layer5_out[7852] = ~layer4_out[3596];
    assign layer5_out[7853] = layer4_out[5948] ^ layer4_out[5949];
    assign layer5_out[7854] = ~layer4_out[1588] | layer4_out[1589];
    assign layer5_out[7855] = ~(layer4_out[166] ^ layer4_out[167]);
    assign layer5_out[7856] = layer4_out[2838] ^ layer4_out[2839];
    assign layer5_out[7857] = ~layer4_out[5976] | layer4_out[5977];
    assign layer5_out[7858] = layer4_out[1263] & ~layer4_out[1264];
    assign layer5_out[7859] = layer4_out[4428] & ~layer4_out[4427];
    assign layer5_out[7860] = layer4_out[5713];
    assign layer5_out[7861] = layer4_out[6827];
    assign layer5_out[7862] = ~(layer4_out[7383] ^ layer4_out[7384]);
    assign layer5_out[7863] = ~(layer4_out[252] ^ layer4_out[253]);
    assign layer5_out[7864] = layer4_out[5936];
    assign layer5_out[7865] = layer4_out[3260] & layer4_out[3261];
    assign layer5_out[7866] = layer4_out[2240] & ~layer4_out[2241];
    assign layer5_out[7867] = layer4_out[1199] ^ layer4_out[1200];
    assign layer5_out[7868] = ~layer4_out[3994];
    assign layer5_out[7869] = ~layer4_out[6959] | layer4_out[6958];
    assign layer5_out[7870] = layer4_out[2003];
    assign layer5_out[7871] = layer4_out[720] & ~layer4_out[721];
    assign layer5_out[7872] = layer4_out[6556];
    assign layer5_out[7873] = layer4_out[1306] ^ layer4_out[1307];
    assign layer5_out[7874] = layer4_out[5912] ^ layer4_out[5913];
    assign layer5_out[7875] = layer4_out[1071];
    assign layer5_out[7876] = ~layer4_out[2674];
    assign layer5_out[7877] = ~(layer4_out[5910] ^ layer4_out[5911]);
    assign layer5_out[7878] = ~layer4_out[191];
    assign layer5_out[7879] = layer4_out[1268];
    assign layer5_out[7880] = layer4_out[2465] & layer4_out[2466];
    assign layer5_out[7881] = ~layer4_out[1484];
    assign layer5_out[7882] = layer4_out[5249] & layer4_out[5250];
    assign layer5_out[7883] = ~layer4_out[6183] | layer4_out[6182];
    assign layer5_out[7884] = ~(layer4_out[3472] ^ layer4_out[3473]);
    assign layer5_out[7885] = layer4_out[1963] & layer4_out[1964];
    assign layer5_out[7886] = ~layer4_out[2674];
    assign layer5_out[7887] = ~layer4_out[671];
    assign layer5_out[7888] = ~(layer4_out[5850] & layer4_out[5851]);
    assign layer5_out[7889] = ~(layer4_out[3055] ^ layer4_out[3056]);
    assign layer5_out[7890] = ~(layer4_out[7597] & layer4_out[7598]);
    assign layer5_out[7891] = ~layer4_out[5894] | layer4_out[5895];
    assign layer5_out[7892] = layer4_out[5604];
    assign layer5_out[7893] = layer4_out[2890] & ~layer4_out[2891];
    assign layer5_out[7894] = ~(layer4_out[5052] | layer4_out[5053]);
    assign layer5_out[7895] = layer4_out[4013] ^ layer4_out[4014];
    assign layer5_out[7896] = layer4_out[115];
    assign layer5_out[7897] = layer4_out[4937] & ~layer4_out[4936];
    assign layer5_out[7898] = layer4_out[6510] & ~layer4_out[6509];
    assign layer5_out[7899] = ~layer4_out[5394] | layer4_out[5395];
    assign layer5_out[7900] = layer4_out[7660];
    assign layer5_out[7901] = ~(layer4_out[5537] ^ layer4_out[5538]);
    assign layer5_out[7902] = ~layer4_out[6422];
    assign layer5_out[7903] = layer4_out[2001];
    assign layer5_out[7904] = layer4_out[3865];
    assign layer5_out[7905] = layer4_out[5256] ^ layer4_out[5257];
    assign layer5_out[7906] = ~(layer4_out[7846] ^ layer4_out[7847]);
    assign layer5_out[7907] = layer4_out[4806];
    assign layer5_out[7908] = layer4_out[5618];
    assign layer5_out[7909] = layer4_out[513] & ~layer4_out[512];
    assign layer5_out[7910] = ~layer4_out[4249];
    assign layer5_out[7911] = ~layer4_out[848] | layer4_out[849];
    assign layer5_out[7912] = ~layer4_out[6217];
    assign layer5_out[7913] = ~layer4_out[2846];
    assign layer5_out[7914] = layer4_out[2192] & ~layer4_out[2191];
    assign layer5_out[7915] = ~layer4_out[4790] | layer4_out[4791];
    assign layer5_out[7916] = layer4_out[6478] & layer4_out[6479];
    assign layer5_out[7917] = layer4_out[4232];
    assign layer5_out[7918] = ~(layer4_out[7056] | layer4_out[7057]);
    assign layer5_out[7919] = layer4_out[5550];
    assign layer5_out[7920] = layer4_out[2493] ^ layer4_out[2494];
    assign layer5_out[7921] = layer4_out[4394] ^ layer4_out[4395];
    assign layer5_out[7922] = layer4_out[416];
    assign layer5_out[7923] = ~(layer4_out[1177] ^ layer4_out[1178]);
    assign layer5_out[7924] = layer4_out[3837] & ~layer4_out[3836];
    assign layer5_out[7925] = ~(layer4_out[5216] ^ layer4_out[5217]);
    assign layer5_out[7926] = layer4_out[2192] & layer4_out[2193];
    assign layer5_out[7927] = layer4_out[5685];
    assign layer5_out[7928] = ~layer4_out[5821];
    assign layer5_out[7929] = ~layer4_out[7279];
    assign layer5_out[7930] = layer4_out[5373];
    assign layer5_out[7931] = layer4_out[5913] & ~layer4_out[5914];
    assign layer5_out[7932] = layer4_out[3182];
    assign layer5_out[7933] = layer4_out[2368] & layer4_out[2369];
    assign layer5_out[7934] = ~layer4_out[7903];
    assign layer5_out[7935] = ~(layer4_out[7179] ^ layer4_out[7180]);
    assign layer5_out[7936] = ~layer4_out[4346] | layer4_out[4347];
    assign layer5_out[7937] = ~(layer4_out[3051] ^ layer4_out[3052]);
    assign layer5_out[7938] = layer4_out[1562];
    assign layer5_out[7939] = layer4_out[6612] | layer4_out[6613];
    assign layer5_out[7940] = layer4_out[5736] & layer4_out[5737];
    assign layer5_out[7941] = ~layer4_out[6632];
    assign layer5_out[7942] = ~layer4_out[4888];
    assign layer5_out[7943] = layer4_out[4797];
    assign layer5_out[7944] = layer4_out[7943] & ~layer4_out[7942];
    assign layer5_out[7945] = ~layer4_out[4237];
    assign layer5_out[7946] = layer4_out[7726] & layer4_out[7727];
    assign layer5_out[7947] = ~(layer4_out[5759] ^ layer4_out[5760]);
    assign layer5_out[7948] = layer4_out[2711] ^ layer4_out[2712];
    assign layer5_out[7949] = layer4_out[388] & ~layer4_out[389];
    assign layer5_out[7950] = ~layer4_out[3535];
    assign layer5_out[7951] = ~layer4_out[4016];
    assign layer5_out[7952] = layer4_out[3432];
    assign layer5_out[7953] = ~layer4_out[6803] | layer4_out[6804];
    assign layer5_out[7954] = ~(layer4_out[4807] ^ layer4_out[4808]);
    assign layer5_out[7955] = ~(layer4_out[5125] & layer4_out[5126]);
    assign layer5_out[7956] = layer4_out[2559];
    assign layer5_out[7957] = layer4_out[7149];
    assign layer5_out[7958] = layer4_out[6310];
    assign layer5_out[7959] = ~layer4_out[3362] | layer4_out[3361];
    assign layer5_out[7960] = layer4_out[4079] ^ layer4_out[4080];
    assign layer5_out[7961] = layer4_out[7305];
    assign layer5_out[7962] = ~layer4_out[3130];
    assign layer5_out[7963] = layer4_out[7515] & ~layer4_out[7516];
    assign layer5_out[7964] = layer4_out[2388] ^ layer4_out[2389];
    assign layer5_out[7965] = ~layer4_out[2182];
    assign layer5_out[7966] = ~(layer4_out[6194] ^ layer4_out[6195]);
    assign layer5_out[7967] = layer4_out[3539] | layer4_out[3540];
    assign layer5_out[7968] = layer4_out[6697] ^ layer4_out[6698];
    assign layer5_out[7969] = ~(layer4_out[2216] ^ layer4_out[2217]);
    assign layer5_out[7970] = ~layer4_out[3575];
    assign layer5_out[7971] = ~(layer4_out[5224] ^ layer4_out[5225]);
    assign layer5_out[7972] = ~layer4_out[7990];
    assign layer5_out[7973] = layer4_out[5467] ^ layer4_out[5468];
    assign layer5_out[7974] = layer4_out[5136] & ~layer4_out[5135];
    assign layer5_out[7975] = layer4_out[3128];
    assign layer5_out[7976] = ~(layer4_out[385] ^ layer4_out[386]);
    assign layer5_out[7977] = layer4_out[4817] | layer4_out[4818];
    assign layer5_out[7978] = layer4_out[4914] ^ layer4_out[4915];
    assign layer5_out[7979] = layer4_out[4571] | layer4_out[4572];
    assign layer5_out[7980] = layer4_out[948];
    assign layer5_out[7981] = layer4_out[7353];
    assign layer5_out[7982] = layer4_out[6439] & ~layer4_out[6438];
    assign layer5_out[7983] = ~(layer4_out[2073] | layer4_out[2074]);
    assign layer5_out[7984] = ~layer4_out[754];
    assign layer5_out[7985] = ~(layer4_out[4418] | layer4_out[4419]);
    assign layer5_out[7986] = ~layer4_out[2819];
    assign layer5_out[7987] = ~layer4_out[7912];
    assign layer5_out[7988] = layer4_out[7204] ^ layer4_out[7205];
    assign layer5_out[7989] = ~(layer4_out[3232] ^ layer4_out[3233]);
    assign layer5_out[7990] = ~layer4_out[6043] | layer4_out[6042];
    assign layer5_out[7991] = ~layer4_out[4654];
    assign layer5_out[7992] = layer4_out[3584] ^ layer4_out[3585];
    assign layer5_out[7993] = layer4_out[2957] ^ layer4_out[2958];
    assign layer5_out[7994] = layer4_out[3963];
    assign layer5_out[7995] = ~(layer4_out[4192] ^ layer4_out[4193]);
    assign layer5_out[7996] = ~layer4_out[1391];
    assign layer5_out[7997] = ~(layer4_out[1388] ^ layer4_out[1389]);
    assign layer5_out[7998] = layer4_out[7729];
    assign layer5_out[7999] = layer4_out[3811] & ~layer4_out[3812];
      wire [7999:0] last_layer_output;
      assign last_layer_output = layer5_out;
      wire [9:0] result [9:0];

      assign result[0] = last_layer_output[0] + last_layer_output[1] + last_layer_output[2] + last_layer_output[3] + last_layer_output[4] + last_layer_output[5] + last_layer_output[6] + last_layer_output[7] + last_layer_output[8] + last_layer_output[9] + last_layer_output[10] + last_layer_output[11] + last_layer_output[12] + last_layer_output[13] + last_layer_output[14] + last_layer_output[15] + last_layer_output[16] + last_layer_output[17] + last_layer_output[18] + last_layer_output[19] + last_layer_output[20] + last_layer_output[21] + last_layer_output[22] + last_layer_output[23] + last_layer_output[24] + last_layer_output[25] + last_layer_output[26] + last_layer_output[27] + last_layer_output[28] + last_layer_output[29] + last_layer_output[30] + last_layer_output[31] + last_layer_output[32] + last_layer_output[33] + last_layer_output[34] + last_layer_output[35] + last_layer_output[36] + last_layer_output[37] + last_layer_output[38] + last_layer_output[39] + last_layer_output[40] + last_layer_output[41] + last_layer_output[42] + last_layer_output[43] + last_layer_output[44] + last_layer_output[45] + last_layer_output[46] + last_layer_output[47] + last_layer_output[48] + last_layer_output[49] + last_layer_output[50] + last_layer_output[51] + last_layer_output[52] + last_layer_output[53] + last_layer_output[54] + last_layer_output[55] + last_layer_output[56] + last_layer_output[57] + last_layer_output[58] + last_layer_output[59] + last_layer_output[60] + last_layer_output[61] + last_layer_output[62] + last_layer_output[63] + last_layer_output[64] + last_layer_output[65] + last_layer_output[66] + last_layer_output[67] + last_layer_output[68] + last_layer_output[69] + last_layer_output[70] + last_layer_output[71] + last_layer_output[72] + last_layer_output[73] + last_layer_output[74] + last_layer_output[75] + last_layer_output[76] + last_layer_output[77] + last_layer_output[78] + last_layer_output[79] + last_layer_output[80] + last_layer_output[81] + last_layer_output[82] + last_layer_output[83] + last_layer_output[84] + last_layer_output[85] + last_layer_output[86] + last_layer_output[87] + last_layer_output[88] + last_layer_output[89] + last_layer_output[90] + last_layer_output[91] + last_layer_output[92] + last_layer_output[93] + last_layer_output[94] + last_layer_output[95] + last_layer_output[96] + last_layer_output[97] + last_layer_output[98] + last_layer_output[99] + last_layer_output[100] + last_layer_output[101] + last_layer_output[102] + last_layer_output[103] + last_layer_output[104] + last_layer_output[105] + last_layer_output[106] + last_layer_output[107] + last_layer_output[108] + last_layer_output[109] + last_layer_output[110] + last_layer_output[111] + last_layer_output[112] + last_layer_output[113] + last_layer_output[114] + last_layer_output[115] + last_layer_output[116] + last_layer_output[117] + last_layer_output[118] + last_layer_output[119] + last_layer_output[120] + last_layer_output[121] + last_layer_output[122] + last_layer_output[123] + last_layer_output[124] + last_layer_output[125] + last_layer_output[126] + last_layer_output[127] + last_layer_output[128] + last_layer_output[129] + last_layer_output[130] + last_layer_output[131] + last_layer_output[132] + last_layer_output[133] + last_layer_output[134] + last_layer_output[135] + last_layer_output[136] + last_layer_output[137] + last_layer_output[138] + last_layer_output[139] + last_layer_output[140] + last_layer_output[141] + last_layer_output[142] + last_layer_output[143] + last_layer_output[144] + last_layer_output[145] + last_layer_output[146] + last_layer_output[147] + last_layer_output[148] + last_layer_output[149] + last_layer_output[150] + last_layer_output[151] + last_layer_output[152] + last_layer_output[153] + last_layer_output[154] + last_layer_output[155] + last_layer_output[156] + last_layer_output[157] + last_layer_output[158] + last_layer_output[159] + last_layer_output[160] + last_layer_output[161] + last_layer_output[162] + last_layer_output[163] + last_layer_output[164] + last_layer_output[165] + last_layer_output[166] + last_layer_output[167] + last_layer_output[168] + last_layer_output[169] + last_layer_output[170] + last_layer_output[171] + last_layer_output[172] + last_layer_output[173] + last_layer_output[174] + last_layer_output[175] + last_layer_output[176] + last_layer_output[177] + last_layer_output[178] + last_layer_output[179] + last_layer_output[180] + last_layer_output[181] + last_layer_output[182] + last_layer_output[183] + last_layer_output[184] + last_layer_output[185] + last_layer_output[186] + last_layer_output[187] + last_layer_output[188] + last_layer_output[189] + last_layer_output[190] + last_layer_output[191] + last_layer_output[192] + last_layer_output[193] + last_layer_output[194] + last_layer_output[195] + last_layer_output[196] + last_layer_output[197] + last_layer_output[198] + last_layer_output[199] + last_layer_output[200] + last_layer_output[201] + last_layer_output[202] + last_layer_output[203] + last_layer_output[204] + last_layer_output[205] + last_layer_output[206] + last_layer_output[207] + last_layer_output[208] + last_layer_output[209] + last_layer_output[210] + last_layer_output[211] + last_layer_output[212] + last_layer_output[213] + last_layer_output[214] + last_layer_output[215] + last_layer_output[216] + last_layer_output[217] + last_layer_output[218] + last_layer_output[219] + last_layer_output[220] + last_layer_output[221] + last_layer_output[222] + last_layer_output[223] + last_layer_output[224] + last_layer_output[225] + last_layer_output[226] + last_layer_output[227] + last_layer_output[228] + last_layer_output[229] + last_layer_output[230] + last_layer_output[231] + last_layer_output[232] + last_layer_output[233] + last_layer_output[234] + last_layer_output[235] + last_layer_output[236] + last_layer_output[237] + last_layer_output[238] + last_layer_output[239] + last_layer_output[240] + last_layer_output[241] + last_layer_output[242] + last_layer_output[243] + last_layer_output[244] + last_layer_output[245] + last_layer_output[246] + last_layer_output[247] + last_layer_output[248] + last_layer_output[249] + last_layer_output[250] + last_layer_output[251] + last_layer_output[252] + last_layer_output[253] + last_layer_output[254] + last_layer_output[255] + last_layer_output[256] + last_layer_output[257] + last_layer_output[258] + last_layer_output[259] + last_layer_output[260] + last_layer_output[261] + last_layer_output[262] + last_layer_output[263] + last_layer_output[264] + last_layer_output[265] + last_layer_output[266] + last_layer_output[267] + last_layer_output[268] + last_layer_output[269] + last_layer_output[270] + last_layer_output[271] + last_layer_output[272] + last_layer_output[273] + last_layer_output[274] + last_layer_output[275] + last_layer_output[276] + last_layer_output[277] + last_layer_output[278] + last_layer_output[279] + last_layer_output[280] + last_layer_output[281] + last_layer_output[282] + last_layer_output[283] + last_layer_output[284] + last_layer_output[285] + last_layer_output[286] + last_layer_output[287] + last_layer_output[288] + last_layer_output[289] + last_layer_output[290] + last_layer_output[291] + last_layer_output[292] + last_layer_output[293] + last_layer_output[294] + last_layer_output[295] + last_layer_output[296] + last_layer_output[297] + last_layer_output[298] + last_layer_output[299] + last_layer_output[300] + last_layer_output[301] + last_layer_output[302] + last_layer_output[303] + last_layer_output[304] + last_layer_output[305] + last_layer_output[306] + last_layer_output[307] + last_layer_output[308] + last_layer_output[309] + last_layer_output[310] + last_layer_output[311] + last_layer_output[312] + last_layer_output[313] + last_layer_output[314] + last_layer_output[315] + last_layer_output[316] + last_layer_output[317] + last_layer_output[318] + last_layer_output[319] + last_layer_output[320] + last_layer_output[321] + last_layer_output[322] + last_layer_output[323] + last_layer_output[324] + last_layer_output[325] + last_layer_output[326] + last_layer_output[327] + last_layer_output[328] + last_layer_output[329] + last_layer_output[330] + last_layer_output[331] + last_layer_output[332] + last_layer_output[333] + last_layer_output[334] + last_layer_output[335] + last_layer_output[336] + last_layer_output[337] + last_layer_output[338] + last_layer_output[339] + last_layer_output[340] + last_layer_output[341] + last_layer_output[342] + last_layer_output[343] + last_layer_output[344] + last_layer_output[345] + last_layer_output[346] + last_layer_output[347] + last_layer_output[348] + last_layer_output[349] + last_layer_output[350] + last_layer_output[351] + last_layer_output[352] + last_layer_output[353] + last_layer_output[354] + last_layer_output[355] + last_layer_output[356] + last_layer_output[357] + last_layer_output[358] + last_layer_output[359] + last_layer_output[360] + last_layer_output[361] + last_layer_output[362] + last_layer_output[363] + last_layer_output[364] + last_layer_output[365] + last_layer_output[366] + last_layer_output[367] + last_layer_output[368] + last_layer_output[369] + last_layer_output[370] + last_layer_output[371] + last_layer_output[372] + last_layer_output[373] + last_layer_output[374] + last_layer_output[375] + last_layer_output[376] + last_layer_output[377] + last_layer_output[378] + last_layer_output[379] + last_layer_output[380] + last_layer_output[381] + last_layer_output[382] + last_layer_output[383] + last_layer_output[384] + last_layer_output[385] + last_layer_output[386] + last_layer_output[387] + last_layer_output[388] + last_layer_output[389] + last_layer_output[390] + last_layer_output[391] + last_layer_output[392] + last_layer_output[393] + last_layer_output[394] + last_layer_output[395] + last_layer_output[396] + last_layer_output[397] + last_layer_output[398] + last_layer_output[399] + last_layer_output[400] + last_layer_output[401] + last_layer_output[402] + last_layer_output[403] + last_layer_output[404] + last_layer_output[405] + last_layer_output[406] + last_layer_output[407] + last_layer_output[408] + last_layer_output[409] + last_layer_output[410] + last_layer_output[411] + last_layer_output[412] + last_layer_output[413] + last_layer_output[414] + last_layer_output[415] + last_layer_output[416] + last_layer_output[417] + last_layer_output[418] + last_layer_output[419] + last_layer_output[420] + last_layer_output[421] + last_layer_output[422] + last_layer_output[423] + last_layer_output[424] + last_layer_output[425] + last_layer_output[426] + last_layer_output[427] + last_layer_output[428] + last_layer_output[429] + last_layer_output[430] + last_layer_output[431] + last_layer_output[432] + last_layer_output[433] + last_layer_output[434] + last_layer_output[435] + last_layer_output[436] + last_layer_output[437] + last_layer_output[438] + last_layer_output[439] + last_layer_output[440] + last_layer_output[441] + last_layer_output[442] + last_layer_output[443] + last_layer_output[444] + last_layer_output[445] + last_layer_output[446] + last_layer_output[447] + last_layer_output[448] + last_layer_output[449] + last_layer_output[450] + last_layer_output[451] + last_layer_output[452] + last_layer_output[453] + last_layer_output[454] + last_layer_output[455] + last_layer_output[456] + last_layer_output[457] + last_layer_output[458] + last_layer_output[459] + last_layer_output[460] + last_layer_output[461] + last_layer_output[462] + last_layer_output[463] + last_layer_output[464] + last_layer_output[465] + last_layer_output[466] + last_layer_output[467] + last_layer_output[468] + last_layer_output[469] + last_layer_output[470] + last_layer_output[471] + last_layer_output[472] + last_layer_output[473] + last_layer_output[474] + last_layer_output[475] + last_layer_output[476] + last_layer_output[477] + last_layer_output[478] + last_layer_output[479] + last_layer_output[480] + last_layer_output[481] + last_layer_output[482] + last_layer_output[483] + last_layer_output[484] + last_layer_output[485] + last_layer_output[486] + last_layer_output[487] + last_layer_output[488] + last_layer_output[489] + last_layer_output[490] + last_layer_output[491] + last_layer_output[492] + last_layer_output[493] + last_layer_output[494] + last_layer_output[495] + last_layer_output[496] + last_layer_output[497] + last_layer_output[498] + last_layer_output[499] + last_layer_output[500] + last_layer_output[501] + last_layer_output[502] + last_layer_output[503] + last_layer_output[504] + last_layer_output[505] + last_layer_output[506] + last_layer_output[507] + last_layer_output[508] + last_layer_output[509] + last_layer_output[510] + last_layer_output[511] + last_layer_output[512] + last_layer_output[513] + last_layer_output[514] + last_layer_output[515] + last_layer_output[516] + last_layer_output[517] + last_layer_output[518] + last_layer_output[519] + last_layer_output[520] + last_layer_output[521] + last_layer_output[522] + last_layer_output[523] + last_layer_output[524] + last_layer_output[525] + last_layer_output[526] + last_layer_output[527] + last_layer_output[528] + last_layer_output[529] + last_layer_output[530] + last_layer_output[531] + last_layer_output[532] + last_layer_output[533] + last_layer_output[534] + last_layer_output[535] + last_layer_output[536] + last_layer_output[537] + last_layer_output[538] + last_layer_output[539] + last_layer_output[540] + last_layer_output[541] + last_layer_output[542] + last_layer_output[543] + last_layer_output[544] + last_layer_output[545] + last_layer_output[546] + last_layer_output[547] + last_layer_output[548] + last_layer_output[549] + last_layer_output[550] + last_layer_output[551] + last_layer_output[552] + last_layer_output[553] + last_layer_output[554] + last_layer_output[555] + last_layer_output[556] + last_layer_output[557] + last_layer_output[558] + last_layer_output[559] + last_layer_output[560] + last_layer_output[561] + last_layer_output[562] + last_layer_output[563] + last_layer_output[564] + last_layer_output[565] + last_layer_output[566] + last_layer_output[567] + last_layer_output[568] + last_layer_output[569] + last_layer_output[570] + last_layer_output[571] + last_layer_output[572] + last_layer_output[573] + last_layer_output[574] + last_layer_output[575] + last_layer_output[576] + last_layer_output[577] + last_layer_output[578] + last_layer_output[579] + last_layer_output[580] + last_layer_output[581] + last_layer_output[582] + last_layer_output[583] + last_layer_output[584] + last_layer_output[585] + last_layer_output[586] + last_layer_output[587] + last_layer_output[588] + last_layer_output[589] + last_layer_output[590] + last_layer_output[591] + last_layer_output[592] + last_layer_output[593] + last_layer_output[594] + last_layer_output[595] + last_layer_output[596] + last_layer_output[597] + last_layer_output[598] + last_layer_output[599] + last_layer_output[600] + last_layer_output[601] + last_layer_output[602] + last_layer_output[603] + last_layer_output[604] + last_layer_output[605] + last_layer_output[606] + last_layer_output[607] + last_layer_output[608] + last_layer_output[609] + last_layer_output[610] + last_layer_output[611] + last_layer_output[612] + last_layer_output[613] + last_layer_output[614] + last_layer_output[615] + last_layer_output[616] + last_layer_output[617] + last_layer_output[618] + last_layer_output[619] + last_layer_output[620] + last_layer_output[621] + last_layer_output[622] + last_layer_output[623] + last_layer_output[624] + last_layer_output[625] + last_layer_output[626] + last_layer_output[627] + last_layer_output[628] + last_layer_output[629] + last_layer_output[630] + last_layer_output[631] + last_layer_output[632] + last_layer_output[633] + last_layer_output[634] + last_layer_output[635] + last_layer_output[636] + last_layer_output[637] + last_layer_output[638] + last_layer_output[639] + last_layer_output[640] + last_layer_output[641] + last_layer_output[642] + last_layer_output[643] + last_layer_output[644] + last_layer_output[645] + last_layer_output[646] + last_layer_output[647] + last_layer_output[648] + last_layer_output[649] + last_layer_output[650] + last_layer_output[651] + last_layer_output[652] + last_layer_output[653] + last_layer_output[654] + last_layer_output[655] + last_layer_output[656] + last_layer_output[657] + last_layer_output[658] + last_layer_output[659] + last_layer_output[660] + last_layer_output[661] + last_layer_output[662] + last_layer_output[663] + last_layer_output[664] + last_layer_output[665] + last_layer_output[666] + last_layer_output[667] + last_layer_output[668] + last_layer_output[669] + last_layer_output[670] + last_layer_output[671] + last_layer_output[672] + last_layer_output[673] + last_layer_output[674] + last_layer_output[675] + last_layer_output[676] + last_layer_output[677] + last_layer_output[678] + last_layer_output[679] + last_layer_output[680] + last_layer_output[681] + last_layer_output[682] + last_layer_output[683] + last_layer_output[684] + last_layer_output[685] + last_layer_output[686] + last_layer_output[687] + last_layer_output[688] + last_layer_output[689] + last_layer_output[690] + last_layer_output[691] + last_layer_output[692] + last_layer_output[693] + last_layer_output[694] + last_layer_output[695] + last_layer_output[696] + last_layer_output[697] + last_layer_output[698] + last_layer_output[699] + last_layer_output[700] + last_layer_output[701] + last_layer_output[702] + last_layer_output[703] + last_layer_output[704] + last_layer_output[705] + last_layer_output[706] + last_layer_output[707] + last_layer_output[708] + last_layer_output[709] + last_layer_output[710] + last_layer_output[711] + last_layer_output[712] + last_layer_output[713] + last_layer_output[714] + last_layer_output[715] + last_layer_output[716] + last_layer_output[717] + last_layer_output[718] + last_layer_output[719] + last_layer_output[720] + last_layer_output[721] + last_layer_output[722] + last_layer_output[723] + last_layer_output[724] + last_layer_output[725] + last_layer_output[726] + last_layer_output[727] + last_layer_output[728] + last_layer_output[729] + last_layer_output[730] + last_layer_output[731] + last_layer_output[732] + last_layer_output[733] + last_layer_output[734] + last_layer_output[735] + last_layer_output[736] + last_layer_output[737] + last_layer_output[738] + last_layer_output[739] + last_layer_output[740] + last_layer_output[741] + last_layer_output[742] + last_layer_output[743] + last_layer_output[744] + last_layer_output[745] + last_layer_output[746] + last_layer_output[747] + last_layer_output[748] + last_layer_output[749] + last_layer_output[750] + last_layer_output[751] + last_layer_output[752] + last_layer_output[753] + last_layer_output[754] + last_layer_output[755] + last_layer_output[756] + last_layer_output[757] + last_layer_output[758] + last_layer_output[759] + last_layer_output[760] + last_layer_output[761] + last_layer_output[762] + last_layer_output[763] + last_layer_output[764] + last_layer_output[765] + last_layer_output[766] + last_layer_output[767] + last_layer_output[768] + last_layer_output[769] + last_layer_output[770] + last_layer_output[771] + last_layer_output[772] + last_layer_output[773] + last_layer_output[774] + last_layer_output[775] + last_layer_output[776] + last_layer_output[777] + last_layer_output[778] + last_layer_output[779] + last_layer_output[780] + last_layer_output[781] + last_layer_output[782] + last_layer_output[783] + last_layer_output[784] + last_layer_output[785] + last_layer_output[786] + last_layer_output[787] + last_layer_output[788] + last_layer_output[789] + last_layer_output[790] + last_layer_output[791] + last_layer_output[792] + last_layer_output[793] + last_layer_output[794] + last_layer_output[795] + last_layer_output[796] + last_layer_output[797] + last_layer_output[798] + last_layer_output[799];
      assign result[1] = last_layer_output[800] + last_layer_output[801] + last_layer_output[802] + last_layer_output[803] + last_layer_output[804] + last_layer_output[805] + last_layer_output[806] + last_layer_output[807] + last_layer_output[808] + last_layer_output[809] + last_layer_output[810] + last_layer_output[811] + last_layer_output[812] + last_layer_output[813] + last_layer_output[814] + last_layer_output[815] + last_layer_output[816] + last_layer_output[817] + last_layer_output[818] + last_layer_output[819] + last_layer_output[820] + last_layer_output[821] + last_layer_output[822] + last_layer_output[823] + last_layer_output[824] + last_layer_output[825] + last_layer_output[826] + last_layer_output[827] + last_layer_output[828] + last_layer_output[829] + last_layer_output[830] + last_layer_output[831] + last_layer_output[832] + last_layer_output[833] + last_layer_output[834] + last_layer_output[835] + last_layer_output[836] + last_layer_output[837] + last_layer_output[838] + last_layer_output[839] + last_layer_output[840] + last_layer_output[841] + last_layer_output[842] + last_layer_output[843] + last_layer_output[844] + last_layer_output[845] + last_layer_output[846] + last_layer_output[847] + last_layer_output[848] + last_layer_output[849] + last_layer_output[850] + last_layer_output[851] + last_layer_output[852] + last_layer_output[853] + last_layer_output[854] + last_layer_output[855] + last_layer_output[856] + last_layer_output[857] + last_layer_output[858] + last_layer_output[859] + last_layer_output[860] + last_layer_output[861] + last_layer_output[862] + last_layer_output[863] + last_layer_output[864] + last_layer_output[865] + last_layer_output[866] + last_layer_output[867] + last_layer_output[868] + last_layer_output[869] + last_layer_output[870] + last_layer_output[871] + last_layer_output[872] + last_layer_output[873] + last_layer_output[874] + last_layer_output[875] + last_layer_output[876] + last_layer_output[877] + last_layer_output[878] + last_layer_output[879] + last_layer_output[880] + last_layer_output[881] + last_layer_output[882] + last_layer_output[883] + last_layer_output[884] + last_layer_output[885] + last_layer_output[886] + last_layer_output[887] + last_layer_output[888] + last_layer_output[889] + last_layer_output[890] + last_layer_output[891] + last_layer_output[892] + last_layer_output[893] + last_layer_output[894] + last_layer_output[895] + last_layer_output[896] + last_layer_output[897] + last_layer_output[898] + last_layer_output[899] + last_layer_output[900] + last_layer_output[901] + last_layer_output[902] + last_layer_output[903] + last_layer_output[904] + last_layer_output[905] + last_layer_output[906] + last_layer_output[907] + last_layer_output[908] + last_layer_output[909] + last_layer_output[910] + last_layer_output[911] + last_layer_output[912] + last_layer_output[913] + last_layer_output[914] + last_layer_output[915] + last_layer_output[916] + last_layer_output[917] + last_layer_output[918] + last_layer_output[919] + last_layer_output[920] + last_layer_output[921] + last_layer_output[922] + last_layer_output[923] + last_layer_output[924] + last_layer_output[925] + last_layer_output[926] + last_layer_output[927] + last_layer_output[928] + last_layer_output[929] + last_layer_output[930] + last_layer_output[931] + last_layer_output[932] + last_layer_output[933] + last_layer_output[934] + last_layer_output[935] + last_layer_output[936] + last_layer_output[937] + last_layer_output[938] + last_layer_output[939] + last_layer_output[940] + last_layer_output[941] + last_layer_output[942] + last_layer_output[943] + last_layer_output[944] + last_layer_output[945] + last_layer_output[946] + last_layer_output[947] + last_layer_output[948] + last_layer_output[949] + last_layer_output[950] + last_layer_output[951] + last_layer_output[952] + last_layer_output[953] + last_layer_output[954] + last_layer_output[955] + last_layer_output[956] + last_layer_output[957] + last_layer_output[958] + last_layer_output[959] + last_layer_output[960] + last_layer_output[961] + last_layer_output[962] + last_layer_output[963] + last_layer_output[964] + last_layer_output[965] + last_layer_output[966] + last_layer_output[967] + last_layer_output[968] + last_layer_output[969] + last_layer_output[970] + last_layer_output[971] + last_layer_output[972] + last_layer_output[973] + last_layer_output[974] + last_layer_output[975] + last_layer_output[976] + last_layer_output[977] + last_layer_output[978] + last_layer_output[979] + last_layer_output[980] + last_layer_output[981] + last_layer_output[982] + last_layer_output[983] + last_layer_output[984] + last_layer_output[985] + last_layer_output[986] + last_layer_output[987] + last_layer_output[988] + last_layer_output[989] + last_layer_output[990] + last_layer_output[991] + last_layer_output[992] + last_layer_output[993] + last_layer_output[994] + last_layer_output[995] + last_layer_output[996] + last_layer_output[997] + last_layer_output[998] + last_layer_output[999] + last_layer_output[1000] + last_layer_output[1001] + last_layer_output[1002] + last_layer_output[1003] + last_layer_output[1004] + last_layer_output[1005] + last_layer_output[1006] + last_layer_output[1007] + last_layer_output[1008] + last_layer_output[1009] + last_layer_output[1010] + last_layer_output[1011] + last_layer_output[1012] + last_layer_output[1013] + last_layer_output[1014] + last_layer_output[1015] + last_layer_output[1016] + last_layer_output[1017] + last_layer_output[1018] + last_layer_output[1019] + last_layer_output[1020] + last_layer_output[1021] + last_layer_output[1022] + last_layer_output[1023] + last_layer_output[1024] + last_layer_output[1025] + last_layer_output[1026] + last_layer_output[1027] + last_layer_output[1028] + last_layer_output[1029] + last_layer_output[1030] + last_layer_output[1031] + last_layer_output[1032] + last_layer_output[1033] + last_layer_output[1034] + last_layer_output[1035] + last_layer_output[1036] + last_layer_output[1037] + last_layer_output[1038] + last_layer_output[1039] + last_layer_output[1040] + last_layer_output[1041] + last_layer_output[1042] + last_layer_output[1043] + last_layer_output[1044] + last_layer_output[1045] + last_layer_output[1046] + last_layer_output[1047] + last_layer_output[1048] + last_layer_output[1049] + last_layer_output[1050] + last_layer_output[1051] + last_layer_output[1052] + last_layer_output[1053] + last_layer_output[1054] + last_layer_output[1055] + last_layer_output[1056] + last_layer_output[1057] + last_layer_output[1058] + last_layer_output[1059] + last_layer_output[1060] + last_layer_output[1061] + last_layer_output[1062] + last_layer_output[1063] + last_layer_output[1064] + last_layer_output[1065] + last_layer_output[1066] + last_layer_output[1067] + last_layer_output[1068] + last_layer_output[1069] + last_layer_output[1070] + last_layer_output[1071] + last_layer_output[1072] + last_layer_output[1073] + last_layer_output[1074] + last_layer_output[1075] + last_layer_output[1076] + last_layer_output[1077] + last_layer_output[1078] + last_layer_output[1079] + last_layer_output[1080] + last_layer_output[1081] + last_layer_output[1082] + last_layer_output[1083] + last_layer_output[1084] + last_layer_output[1085] + last_layer_output[1086] + last_layer_output[1087] + last_layer_output[1088] + last_layer_output[1089] + last_layer_output[1090] + last_layer_output[1091] + last_layer_output[1092] + last_layer_output[1093] + last_layer_output[1094] + last_layer_output[1095] + last_layer_output[1096] + last_layer_output[1097] + last_layer_output[1098] + last_layer_output[1099] + last_layer_output[1100] + last_layer_output[1101] + last_layer_output[1102] + last_layer_output[1103] + last_layer_output[1104] + last_layer_output[1105] + last_layer_output[1106] + last_layer_output[1107] + last_layer_output[1108] + last_layer_output[1109] + last_layer_output[1110] + last_layer_output[1111] + last_layer_output[1112] + last_layer_output[1113] + last_layer_output[1114] + last_layer_output[1115] + last_layer_output[1116] + last_layer_output[1117] + last_layer_output[1118] + last_layer_output[1119] + last_layer_output[1120] + last_layer_output[1121] + last_layer_output[1122] + last_layer_output[1123] + last_layer_output[1124] + last_layer_output[1125] + last_layer_output[1126] + last_layer_output[1127] + last_layer_output[1128] + last_layer_output[1129] + last_layer_output[1130] + last_layer_output[1131] + last_layer_output[1132] + last_layer_output[1133] + last_layer_output[1134] + last_layer_output[1135] + last_layer_output[1136] + last_layer_output[1137] + last_layer_output[1138] + last_layer_output[1139] + last_layer_output[1140] + last_layer_output[1141] + last_layer_output[1142] + last_layer_output[1143] + last_layer_output[1144] + last_layer_output[1145] + last_layer_output[1146] + last_layer_output[1147] + last_layer_output[1148] + last_layer_output[1149] + last_layer_output[1150] + last_layer_output[1151] + last_layer_output[1152] + last_layer_output[1153] + last_layer_output[1154] + last_layer_output[1155] + last_layer_output[1156] + last_layer_output[1157] + last_layer_output[1158] + last_layer_output[1159] + last_layer_output[1160] + last_layer_output[1161] + last_layer_output[1162] + last_layer_output[1163] + last_layer_output[1164] + last_layer_output[1165] + last_layer_output[1166] + last_layer_output[1167] + last_layer_output[1168] + last_layer_output[1169] + last_layer_output[1170] + last_layer_output[1171] + last_layer_output[1172] + last_layer_output[1173] + last_layer_output[1174] + last_layer_output[1175] + last_layer_output[1176] + last_layer_output[1177] + last_layer_output[1178] + last_layer_output[1179] + last_layer_output[1180] + last_layer_output[1181] + last_layer_output[1182] + last_layer_output[1183] + last_layer_output[1184] + last_layer_output[1185] + last_layer_output[1186] + last_layer_output[1187] + last_layer_output[1188] + last_layer_output[1189] + last_layer_output[1190] + last_layer_output[1191] + last_layer_output[1192] + last_layer_output[1193] + last_layer_output[1194] + last_layer_output[1195] + last_layer_output[1196] + last_layer_output[1197] + last_layer_output[1198] + last_layer_output[1199] + last_layer_output[1200] + last_layer_output[1201] + last_layer_output[1202] + last_layer_output[1203] + last_layer_output[1204] + last_layer_output[1205] + last_layer_output[1206] + last_layer_output[1207] + last_layer_output[1208] + last_layer_output[1209] + last_layer_output[1210] + last_layer_output[1211] + last_layer_output[1212] + last_layer_output[1213] + last_layer_output[1214] + last_layer_output[1215] + last_layer_output[1216] + last_layer_output[1217] + last_layer_output[1218] + last_layer_output[1219] + last_layer_output[1220] + last_layer_output[1221] + last_layer_output[1222] + last_layer_output[1223] + last_layer_output[1224] + last_layer_output[1225] + last_layer_output[1226] + last_layer_output[1227] + last_layer_output[1228] + last_layer_output[1229] + last_layer_output[1230] + last_layer_output[1231] + last_layer_output[1232] + last_layer_output[1233] + last_layer_output[1234] + last_layer_output[1235] + last_layer_output[1236] + last_layer_output[1237] + last_layer_output[1238] + last_layer_output[1239] + last_layer_output[1240] + last_layer_output[1241] + last_layer_output[1242] + last_layer_output[1243] + last_layer_output[1244] + last_layer_output[1245] + last_layer_output[1246] + last_layer_output[1247] + last_layer_output[1248] + last_layer_output[1249] + last_layer_output[1250] + last_layer_output[1251] + last_layer_output[1252] + last_layer_output[1253] + last_layer_output[1254] + last_layer_output[1255] + last_layer_output[1256] + last_layer_output[1257] + last_layer_output[1258] + last_layer_output[1259] + last_layer_output[1260] + last_layer_output[1261] + last_layer_output[1262] + last_layer_output[1263] + last_layer_output[1264] + last_layer_output[1265] + last_layer_output[1266] + last_layer_output[1267] + last_layer_output[1268] + last_layer_output[1269] + last_layer_output[1270] + last_layer_output[1271] + last_layer_output[1272] + last_layer_output[1273] + last_layer_output[1274] + last_layer_output[1275] + last_layer_output[1276] + last_layer_output[1277] + last_layer_output[1278] + last_layer_output[1279] + last_layer_output[1280] + last_layer_output[1281] + last_layer_output[1282] + last_layer_output[1283] + last_layer_output[1284] + last_layer_output[1285] + last_layer_output[1286] + last_layer_output[1287] + last_layer_output[1288] + last_layer_output[1289] + last_layer_output[1290] + last_layer_output[1291] + last_layer_output[1292] + last_layer_output[1293] + last_layer_output[1294] + last_layer_output[1295] + last_layer_output[1296] + last_layer_output[1297] + last_layer_output[1298] + last_layer_output[1299] + last_layer_output[1300] + last_layer_output[1301] + last_layer_output[1302] + last_layer_output[1303] + last_layer_output[1304] + last_layer_output[1305] + last_layer_output[1306] + last_layer_output[1307] + last_layer_output[1308] + last_layer_output[1309] + last_layer_output[1310] + last_layer_output[1311] + last_layer_output[1312] + last_layer_output[1313] + last_layer_output[1314] + last_layer_output[1315] + last_layer_output[1316] + last_layer_output[1317] + last_layer_output[1318] + last_layer_output[1319] + last_layer_output[1320] + last_layer_output[1321] + last_layer_output[1322] + last_layer_output[1323] + last_layer_output[1324] + last_layer_output[1325] + last_layer_output[1326] + last_layer_output[1327] + last_layer_output[1328] + last_layer_output[1329] + last_layer_output[1330] + last_layer_output[1331] + last_layer_output[1332] + last_layer_output[1333] + last_layer_output[1334] + last_layer_output[1335] + last_layer_output[1336] + last_layer_output[1337] + last_layer_output[1338] + last_layer_output[1339] + last_layer_output[1340] + last_layer_output[1341] + last_layer_output[1342] + last_layer_output[1343] + last_layer_output[1344] + last_layer_output[1345] + last_layer_output[1346] + last_layer_output[1347] + last_layer_output[1348] + last_layer_output[1349] + last_layer_output[1350] + last_layer_output[1351] + last_layer_output[1352] + last_layer_output[1353] + last_layer_output[1354] + last_layer_output[1355] + last_layer_output[1356] + last_layer_output[1357] + last_layer_output[1358] + last_layer_output[1359] + last_layer_output[1360] + last_layer_output[1361] + last_layer_output[1362] + last_layer_output[1363] + last_layer_output[1364] + last_layer_output[1365] + last_layer_output[1366] + last_layer_output[1367] + last_layer_output[1368] + last_layer_output[1369] + last_layer_output[1370] + last_layer_output[1371] + last_layer_output[1372] + last_layer_output[1373] + last_layer_output[1374] + last_layer_output[1375] + last_layer_output[1376] + last_layer_output[1377] + last_layer_output[1378] + last_layer_output[1379] + last_layer_output[1380] + last_layer_output[1381] + last_layer_output[1382] + last_layer_output[1383] + last_layer_output[1384] + last_layer_output[1385] + last_layer_output[1386] + last_layer_output[1387] + last_layer_output[1388] + last_layer_output[1389] + last_layer_output[1390] + last_layer_output[1391] + last_layer_output[1392] + last_layer_output[1393] + last_layer_output[1394] + last_layer_output[1395] + last_layer_output[1396] + last_layer_output[1397] + last_layer_output[1398] + last_layer_output[1399] + last_layer_output[1400] + last_layer_output[1401] + last_layer_output[1402] + last_layer_output[1403] + last_layer_output[1404] + last_layer_output[1405] + last_layer_output[1406] + last_layer_output[1407] + last_layer_output[1408] + last_layer_output[1409] + last_layer_output[1410] + last_layer_output[1411] + last_layer_output[1412] + last_layer_output[1413] + last_layer_output[1414] + last_layer_output[1415] + last_layer_output[1416] + last_layer_output[1417] + last_layer_output[1418] + last_layer_output[1419] + last_layer_output[1420] + last_layer_output[1421] + last_layer_output[1422] + last_layer_output[1423] + last_layer_output[1424] + last_layer_output[1425] + last_layer_output[1426] + last_layer_output[1427] + last_layer_output[1428] + last_layer_output[1429] + last_layer_output[1430] + last_layer_output[1431] + last_layer_output[1432] + last_layer_output[1433] + last_layer_output[1434] + last_layer_output[1435] + last_layer_output[1436] + last_layer_output[1437] + last_layer_output[1438] + last_layer_output[1439] + last_layer_output[1440] + last_layer_output[1441] + last_layer_output[1442] + last_layer_output[1443] + last_layer_output[1444] + last_layer_output[1445] + last_layer_output[1446] + last_layer_output[1447] + last_layer_output[1448] + last_layer_output[1449] + last_layer_output[1450] + last_layer_output[1451] + last_layer_output[1452] + last_layer_output[1453] + last_layer_output[1454] + last_layer_output[1455] + last_layer_output[1456] + last_layer_output[1457] + last_layer_output[1458] + last_layer_output[1459] + last_layer_output[1460] + last_layer_output[1461] + last_layer_output[1462] + last_layer_output[1463] + last_layer_output[1464] + last_layer_output[1465] + last_layer_output[1466] + last_layer_output[1467] + last_layer_output[1468] + last_layer_output[1469] + last_layer_output[1470] + last_layer_output[1471] + last_layer_output[1472] + last_layer_output[1473] + last_layer_output[1474] + last_layer_output[1475] + last_layer_output[1476] + last_layer_output[1477] + last_layer_output[1478] + last_layer_output[1479] + last_layer_output[1480] + last_layer_output[1481] + last_layer_output[1482] + last_layer_output[1483] + last_layer_output[1484] + last_layer_output[1485] + last_layer_output[1486] + last_layer_output[1487] + last_layer_output[1488] + last_layer_output[1489] + last_layer_output[1490] + last_layer_output[1491] + last_layer_output[1492] + last_layer_output[1493] + last_layer_output[1494] + last_layer_output[1495] + last_layer_output[1496] + last_layer_output[1497] + last_layer_output[1498] + last_layer_output[1499] + last_layer_output[1500] + last_layer_output[1501] + last_layer_output[1502] + last_layer_output[1503] + last_layer_output[1504] + last_layer_output[1505] + last_layer_output[1506] + last_layer_output[1507] + last_layer_output[1508] + last_layer_output[1509] + last_layer_output[1510] + last_layer_output[1511] + last_layer_output[1512] + last_layer_output[1513] + last_layer_output[1514] + last_layer_output[1515] + last_layer_output[1516] + last_layer_output[1517] + last_layer_output[1518] + last_layer_output[1519] + last_layer_output[1520] + last_layer_output[1521] + last_layer_output[1522] + last_layer_output[1523] + last_layer_output[1524] + last_layer_output[1525] + last_layer_output[1526] + last_layer_output[1527] + last_layer_output[1528] + last_layer_output[1529] + last_layer_output[1530] + last_layer_output[1531] + last_layer_output[1532] + last_layer_output[1533] + last_layer_output[1534] + last_layer_output[1535] + last_layer_output[1536] + last_layer_output[1537] + last_layer_output[1538] + last_layer_output[1539] + last_layer_output[1540] + last_layer_output[1541] + last_layer_output[1542] + last_layer_output[1543] + last_layer_output[1544] + last_layer_output[1545] + last_layer_output[1546] + last_layer_output[1547] + last_layer_output[1548] + last_layer_output[1549] + last_layer_output[1550] + last_layer_output[1551] + last_layer_output[1552] + last_layer_output[1553] + last_layer_output[1554] + last_layer_output[1555] + last_layer_output[1556] + last_layer_output[1557] + last_layer_output[1558] + last_layer_output[1559] + last_layer_output[1560] + last_layer_output[1561] + last_layer_output[1562] + last_layer_output[1563] + last_layer_output[1564] + last_layer_output[1565] + last_layer_output[1566] + last_layer_output[1567] + last_layer_output[1568] + last_layer_output[1569] + last_layer_output[1570] + last_layer_output[1571] + last_layer_output[1572] + last_layer_output[1573] + last_layer_output[1574] + last_layer_output[1575] + last_layer_output[1576] + last_layer_output[1577] + last_layer_output[1578] + last_layer_output[1579] + last_layer_output[1580] + last_layer_output[1581] + last_layer_output[1582] + last_layer_output[1583] + last_layer_output[1584] + last_layer_output[1585] + last_layer_output[1586] + last_layer_output[1587] + last_layer_output[1588] + last_layer_output[1589] + last_layer_output[1590] + last_layer_output[1591] + last_layer_output[1592] + last_layer_output[1593] + last_layer_output[1594] + last_layer_output[1595] + last_layer_output[1596] + last_layer_output[1597] + last_layer_output[1598] + last_layer_output[1599];
      assign result[2] = last_layer_output[1600] + last_layer_output[1601] + last_layer_output[1602] + last_layer_output[1603] + last_layer_output[1604] + last_layer_output[1605] + last_layer_output[1606] + last_layer_output[1607] + last_layer_output[1608] + last_layer_output[1609] + last_layer_output[1610] + last_layer_output[1611] + last_layer_output[1612] + last_layer_output[1613] + last_layer_output[1614] + last_layer_output[1615] + last_layer_output[1616] + last_layer_output[1617] + last_layer_output[1618] + last_layer_output[1619] + last_layer_output[1620] + last_layer_output[1621] + last_layer_output[1622] + last_layer_output[1623] + last_layer_output[1624] + last_layer_output[1625] + last_layer_output[1626] + last_layer_output[1627] + last_layer_output[1628] + last_layer_output[1629] + last_layer_output[1630] + last_layer_output[1631] + last_layer_output[1632] + last_layer_output[1633] + last_layer_output[1634] + last_layer_output[1635] + last_layer_output[1636] + last_layer_output[1637] + last_layer_output[1638] + last_layer_output[1639] + last_layer_output[1640] + last_layer_output[1641] + last_layer_output[1642] + last_layer_output[1643] + last_layer_output[1644] + last_layer_output[1645] + last_layer_output[1646] + last_layer_output[1647] + last_layer_output[1648] + last_layer_output[1649] + last_layer_output[1650] + last_layer_output[1651] + last_layer_output[1652] + last_layer_output[1653] + last_layer_output[1654] + last_layer_output[1655] + last_layer_output[1656] + last_layer_output[1657] + last_layer_output[1658] + last_layer_output[1659] + last_layer_output[1660] + last_layer_output[1661] + last_layer_output[1662] + last_layer_output[1663] + last_layer_output[1664] + last_layer_output[1665] + last_layer_output[1666] + last_layer_output[1667] + last_layer_output[1668] + last_layer_output[1669] + last_layer_output[1670] + last_layer_output[1671] + last_layer_output[1672] + last_layer_output[1673] + last_layer_output[1674] + last_layer_output[1675] + last_layer_output[1676] + last_layer_output[1677] + last_layer_output[1678] + last_layer_output[1679] + last_layer_output[1680] + last_layer_output[1681] + last_layer_output[1682] + last_layer_output[1683] + last_layer_output[1684] + last_layer_output[1685] + last_layer_output[1686] + last_layer_output[1687] + last_layer_output[1688] + last_layer_output[1689] + last_layer_output[1690] + last_layer_output[1691] + last_layer_output[1692] + last_layer_output[1693] + last_layer_output[1694] + last_layer_output[1695] + last_layer_output[1696] + last_layer_output[1697] + last_layer_output[1698] + last_layer_output[1699] + last_layer_output[1700] + last_layer_output[1701] + last_layer_output[1702] + last_layer_output[1703] + last_layer_output[1704] + last_layer_output[1705] + last_layer_output[1706] + last_layer_output[1707] + last_layer_output[1708] + last_layer_output[1709] + last_layer_output[1710] + last_layer_output[1711] + last_layer_output[1712] + last_layer_output[1713] + last_layer_output[1714] + last_layer_output[1715] + last_layer_output[1716] + last_layer_output[1717] + last_layer_output[1718] + last_layer_output[1719] + last_layer_output[1720] + last_layer_output[1721] + last_layer_output[1722] + last_layer_output[1723] + last_layer_output[1724] + last_layer_output[1725] + last_layer_output[1726] + last_layer_output[1727] + last_layer_output[1728] + last_layer_output[1729] + last_layer_output[1730] + last_layer_output[1731] + last_layer_output[1732] + last_layer_output[1733] + last_layer_output[1734] + last_layer_output[1735] + last_layer_output[1736] + last_layer_output[1737] + last_layer_output[1738] + last_layer_output[1739] + last_layer_output[1740] + last_layer_output[1741] + last_layer_output[1742] + last_layer_output[1743] + last_layer_output[1744] + last_layer_output[1745] + last_layer_output[1746] + last_layer_output[1747] + last_layer_output[1748] + last_layer_output[1749] + last_layer_output[1750] + last_layer_output[1751] + last_layer_output[1752] + last_layer_output[1753] + last_layer_output[1754] + last_layer_output[1755] + last_layer_output[1756] + last_layer_output[1757] + last_layer_output[1758] + last_layer_output[1759] + last_layer_output[1760] + last_layer_output[1761] + last_layer_output[1762] + last_layer_output[1763] + last_layer_output[1764] + last_layer_output[1765] + last_layer_output[1766] + last_layer_output[1767] + last_layer_output[1768] + last_layer_output[1769] + last_layer_output[1770] + last_layer_output[1771] + last_layer_output[1772] + last_layer_output[1773] + last_layer_output[1774] + last_layer_output[1775] + last_layer_output[1776] + last_layer_output[1777] + last_layer_output[1778] + last_layer_output[1779] + last_layer_output[1780] + last_layer_output[1781] + last_layer_output[1782] + last_layer_output[1783] + last_layer_output[1784] + last_layer_output[1785] + last_layer_output[1786] + last_layer_output[1787] + last_layer_output[1788] + last_layer_output[1789] + last_layer_output[1790] + last_layer_output[1791] + last_layer_output[1792] + last_layer_output[1793] + last_layer_output[1794] + last_layer_output[1795] + last_layer_output[1796] + last_layer_output[1797] + last_layer_output[1798] + last_layer_output[1799] + last_layer_output[1800] + last_layer_output[1801] + last_layer_output[1802] + last_layer_output[1803] + last_layer_output[1804] + last_layer_output[1805] + last_layer_output[1806] + last_layer_output[1807] + last_layer_output[1808] + last_layer_output[1809] + last_layer_output[1810] + last_layer_output[1811] + last_layer_output[1812] + last_layer_output[1813] + last_layer_output[1814] + last_layer_output[1815] + last_layer_output[1816] + last_layer_output[1817] + last_layer_output[1818] + last_layer_output[1819] + last_layer_output[1820] + last_layer_output[1821] + last_layer_output[1822] + last_layer_output[1823] + last_layer_output[1824] + last_layer_output[1825] + last_layer_output[1826] + last_layer_output[1827] + last_layer_output[1828] + last_layer_output[1829] + last_layer_output[1830] + last_layer_output[1831] + last_layer_output[1832] + last_layer_output[1833] + last_layer_output[1834] + last_layer_output[1835] + last_layer_output[1836] + last_layer_output[1837] + last_layer_output[1838] + last_layer_output[1839] + last_layer_output[1840] + last_layer_output[1841] + last_layer_output[1842] + last_layer_output[1843] + last_layer_output[1844] + last_layer_output[1845] + last_layer_output[1846] + last_layer_output[1847] + last_layer_output[1848] + last_layer_output[1849] + last_layer_output[1850] + last_layer_output[1851] + last_layer_output[1852] + last_layer_output[1853] + last_layer_output[1854] + last_layer_output[1855] + last_layer_output[1856] + last_layer_output[1857] + last_layer_output[1858] + last_layer_output[1859] + last_layer_output[1860] + last_layer_output[1861] + last_layer_output[1862] + last_layer_output[1863] + last_layer_output[1864] + last_layer_output[1865] + last_layer_output[1866] + last_layer_output[1867] + last_layer_output[1868] + last_layer_output[1869] + last_layer_output[1870] + last_layer_output[1871] + last_layer_output[1872] + last_layer_output[1873] + last_layer_output[1874] + last_layer_output[1875] + last_layer_output[1876] + last_layer_output[1877] + last_layer_output[1878] + last_layer_output[1879] + last_layer_output[1880] + last_layer_output[1881] + last_layer_output[1882] + last_layer_output[1883] + last_layer_output[1884] + last_layer_output[1885] + last_layer_output[1886] + last_layer_output[1887] + last_layer_output[1888] + last_layer_output[1889] + last_layer_output[1890] + last_layer_output[1891] + last_layer_output[1892] + last_layer_output[1893] + last_layer_output[1894] + last_layer_output[1895] + last_layer_output[1896] + last_layer_output[1897] + last_layer_output[1898] + last_layer_output[1899] + last_layer_output[1900] + last_layer_output[1901] + last_layer_output[1902] + last_layer_output[1903] + last_layer_output[1904] + last_layer_output[1905] + last_layer_output[1906] + last_layer_output[1907] + last_layer_output[1908] + last_layer_output[1909] + last_layer_output[1910] + last_layer_output[1911] + last_layer_output[1912] + last_layer_output[1913] + last_layer_output[1914] + last_layer_output[1915] + last_layer_output[1916] + last_layer_output[1917] + last_layer_output[1918] + last_layer_output[1919] + last_layer_output[1920] + last_layer_output[1921] + last_layer_output[1922] + last_layer_output[1923] + last_layer_output[1924] + last_layer_output[1925] + last_layer_output[1926] + last_layer_output[1927] + last_layer_output[1928] + last_layer_output[1929] + last_layer_output[1930] + last_layer_output[1931] + last_layer_output[1932] + last_layer_output[1933] + last_layer_output[1934] + last_layer_output[1935] + last_layer_output[1936] + last_layer_output[1937] + last_layer_output[1938] + last_layer_output[1939] + last_layer_output[1940] + last_layer_output[1941] + last_layer_output[1942] + last_layer_output[1943] + last_layer_output[1944] + last_layer_output[1945] + last_layer_output[1946] + last_layer_output[1947] + last_layer_output[1948] + last_layer_output[1949] + last_layer_output[1950] + last_layer_output[1951] + last_layer_output[1952] + last_layer_output[1953] + last_layer_output[1954] + last_layer_output[1955] + last_layer_output[1956] + last_layer_output[1957] + last_layer_output[1958] + last_layer_output[1959] + last_layer_output[1960] + last_layer_output[1961] + last_layer_output[1962] + last_layer_output[1963] + last_layer_output[1964] + last_layer_output[1965] + last_layer_output[1966] + last_layer_output[1967] + last_layer_output[1968] + last_layer_output[1969] + last_layer_output[1970] + last_layer_output[1971] + last_layer_output[1972] + last_layer_output[1973] + last_layer_output[1974] + last_layer_output[1975] + last_layer_output[1976] + last_layer_output[1977] + last_layer_output[1978] + last_layer_output[1979] + last_layer_output[1980] + last_layer_output[1981] + last_layer_output[1982] + last_layer_output[1983] + last_layer_output[1984] + last_layer_output[1985] + last_layer_output[1986] + last_layer_output[1987] + last_layer_output[1988] + last_layer_output[1989] + last_layer_output[1990] + last_layer_output[1991] + last_layer_output[1992] + last_layer_output[1993] + last_layer_output[1994] + last_layer_output[1995] + last_layer_output[1996] + last_layer_output[1997] + last_layer_output[1998] + last_layer_output[1999] + last_layer_output[2000] + last_layer_output[2001] + last_layer_output[2002] + last_layer_output[2003] + last_layer_output[2004] + last_layer_output[2005] + last_layer_output[2006] + last_layer_output[2007] + last_layer_output[2008] + last_layer_output[2009] + last_layer_output[2010] + last_layer_output[2011] + last_layer_output[2012] + last_layer_output[2013] + last_layer_output[2014] + last_layer_output[2015] + last_layer_output[2016] + last_layer_output[2017] + last_layer_output[2018] + last_layer_output[2019] + last_layer_output[2020] + last_layer_output[2021] + last_layer_output[2022] + last_layer_output[2023] + last_layer_output[2024] + last_layer_output[2025] + last_layer_output[2026] + last_layer_output[2027] + last_layer_output[2028] + last_layer_output[2029] + last_layer_output[2030] + last_layer_output[2031] + last_layer_output[2032] + last_layer_output[2033] + last_layer_output[2034] + last_layer_output[2035] + last_layer_output[2036] + last_layer_output[2037] + last_layer_output[2038] + last_layer_output[2039] + last_layer_output[2040] + last_layer_output[2041] + last_layer_output[2042] + last_layer_output[2043] + last_layer_output[2044] + last_layer_output[2045] + last_layer_output[2046] + last_layer_output[2047] + last_layer_output[2048] + last_layer_output[2049] + last_layer_output[2050] + last_layer_output[2051] + last_layer_output[2052] + last_layer_output[2053] + last_layer_output[2054] + last_layer_output[2055] + last_layer_output[2056] + last_layer_output[2057] + last_layer_output[2058] + last_layer_output[2059] + last_layer_output[2060] + last_layer_output[2061] + last_layer_output[2062] + last_layer_output[2063] + last_layer_output[2064] + last_layer_output[2065] + last_layer_output[2066] + last_layer_output[2067] + last_layer_output[2068] + last_layer_output[2069] + last_layer_output[2070] + last_layer_output[2071] + last_layer_output[2072] + last_layer_output[2073] + last_layer_output[2074] + last_layer_output[2075] + last_layer_output[2076] + last_layer_output[2077] + last_layer_output[2078] + last_layer_output[2079] + last_layer_output[2080] + last_layer_output[2081] + last_layer_output[2082] + last_layer_output[2083] + last_layer_output[2084] + last_layer_output[2085] + last_layer_output[2086] + last_layer_output[2087] + last_layer_output[2088] + last_layer_output[2089] + last_layer_output[2090] + last_layer_output[2091] + last_layer_output[2092] + last_layer_output[2093] + last_layer_output[2094] + last_layer_output[2095] + last_layer_output[2096] + last_layer_output[2097] + last_layer_output[2098] + last_layer_output[2099] + last_layer_output[2100] + last_layer_output[2101] + last_layer_output[2102] + last_layer_output[2103] + last_layer_output[2104] + last_layer_output[2105] + last_layer_output[2106] + last_layer_output[2107] + last_layer_output[2108] + last_layer_output[2109] + last_layer_output[2110] + last_layer_output[2111] + last_layer_output[2112] + last_layer_output[2113] + last_layer_output[2114] + last_layer_output[2115] + last_layer_output[2116] + last_layer_output[2117] + last_layer_output[2118] + last_layer_output[2119] + last_layer_output[2120] + last_layer_output[2121] + last_layer_output[2122] + last_layer_output[2123] + last_layer_output[2124] + last_layer_output[2125] + last_layer_output[2126] + last_layer_output[2127] + last_layer_output[2128] + last_layer_output[2129] + last_layer_output[2130] + last_layer_output[2131] + last_layer_output[2132] + last_layer_output[2133] + last_layer_output[2134] + last_layer_output[2135] + last_layer_output[2136] + last_layer_output[2137] + last_layer_output[2138] + last_layer_output[2139] + last_layer_output[2140] + last_layer_output[2141] + last_layer_output[2142] + last_layer_output[2143] + last_layer_output[2144] + last_layer_output[2145] + last_layer_output[2146] + last_layer_output[2147] + last_layer_output[2148] + last_layer_output[2149] + last_layer_output[2150] + last_layer_output[2151] + last_layer_output[2152] + last_layer_output[2153] + last_layer_output[2154] + last_layer_output[2155] + last_layer_output[2156] + last_layer_output[2157] + last_layer_output[2158] + last_layer_output[2159] + last_layer_output[2160] + last_layer_output[2161] + last_layer_output[2162] + last_layer_output[2163] + last_layer_output[2164] + last_layer_output[2165] + last_layer_output[2166] + last_layer_output[2167] + last_layer_output[2168] + last_layer_output[2169] + last_layer_output[2170] + last_layer_output[2171] + last_layer_output[2172] + last_layer_output[2173] + last_layer_output[2174] + last_layer_output[2175] + last_layer_output[2176] + last_layer_output[2177] + last_layer_output[2178] + last_layer_output[2179] + last_layer_output[2180] + last_layer_output[2181] + last_layer_output[2182] + last_layer_output[2183] + last_layer_output[2184] + last_layer_output[2185] + last_layer_output[2186] + last_layer_output[2187] + last_layer_output[2188] + last_layer_output[2189] + last_layer_output[2190] + last_layer_output[2191] + last_layer_output[2192] + last_layer_output[2193] + last_layer_output[2194] + last_layer_output[2195] + last_layer_output[2196] + last_layer_output[2197] + last_layer_output[2198] + last_layer_output[2199] + last_layer_output[2200] + last_layer_output[2201] + last_layer_output[2202] + last_layer_output[2203] + last_layer_output[2204] + last_layer_output[2205] + last_layer_output[2206] + last_layer_output[2207] + last_layer_output[2208] + last_layer_output[2209] + last_layer_output[2210] + last_layer_output[2211] + last_layer_output[2212] + last_layer_output[2213] + last_layer_output[2214] + last_layer_output[2215] + last_layer_output[2216] + last_layer_output[2217] + last_layer_output[2218] + last_layer_output[2219] + last_layer_output[2220] + last_layer_output[2221] + last_layer_output[2222] + last_layer_output[2223] + last_layer_output[2224] + last_layer_output[2225] + last_layer_output[2226] + last_layer_output[2227] + last_layer_output[2228] + last_layer_output[2229] + last_layer_output[2230] + last_layer_output[2231] + last_layer_output[2232] + last_layer_output[2233] + last_layer_output[2234] + last_layer_output[2235] + last_layer_output[2236] + last_layer_output[2237] + last_layer_output[2238] + last_layer_output[2239] + last_layer_output[2240] + last_layer_output[2241] + last_layer_output[2242] + last_layer_output[2243] + last_layer_output[2244] + last_layer_output[2245] + last_layer_output[2246] + last_layer_output[2247] + last_layer_output[2248] + last_layer_output[2249] + last_layer_output[2250] + last_layer_output[2251] + last_layer_output[2252] + last_layer_output[2253] + last_layer_output[2254] + last_layer_output[2255] + last_layer_output[2256] + last_layer_output[2257] + last_layer_output[2258] + last_layer_output[2259] + last_layer_output[2260] + last_layer_output[2261] + last_layer_output[2262] + last_layer_output[2263] + last_layer_output[2264] + last_layer_output[2265] + last_layer_output[2266] + last_layer_output[2267] + last_layer_output[2268] + last_layer_output[2269] + last_layer_output[2270] + last_layer_output[2271] + last_layer_output[2272] + last_layer_output[2273] + last_layer_output[2274] + last_layer_output[2275] + last_layer_output[2276] + last_layer_output[2277] + last_layer_output[2278] + last_layer_output[2279] + last_layer_output[2280] + last_layer_output[2281] + last_layer_output[2282] + last_layer_output[2283] + last_layer_output[2284] + last_layer_output[2285] + last_layer_output[2286] + last_layer_output[2287] + last_layer_output[2288] + last_layer_output[2289] + last_layer_output[2290] + last_layer_output[2291] + last_layer_output[2292] + last_layer_output[2293] + last_layer_output[2294] + last_layer_output[2295] + last_layer_output[2296] + last_layer_output[2297] + last_layer_output[2298] + last_layer_output[2299] + last_layer_output[2300] + last_layer_output[2301] + last_layer_output[2302] + last_layer_output[2303] + last_layer_output[2304] + last_layer_output[2305] + last_layer_output[2306] + last_layer_output[2307] + last_layer_output[2308] + last_layer_output[2309] + last_layer_output[2310] + last_layer_output[2311] + last_layer_output[2312] + last_layer_output[2313] + last_layer_output[2314] + last_layer_output[2315] + last_layer_output[2316] + last_layer_output[2317] + last_layer_output[2318] + last_layer_output[2319] + last_layer_output[2320] + last_layer_output[2321] + last_layer_output[2322] + last_layer_output[2323] + last_layer_output[2324] + last_layer_output[2325] + last_layer_output[2326] + last_layer_output[2327] + last_layer_output[2328] + last_layer_output[2329] + last_layer_output[2330] + last_layer_output[2331] + last_layer_output[2332] + last_layer_output[2333] + last_layer_output[2334] + last_layer_output[2335] + last_layer_output[2336] + last_layer_output[2337] + last_layer_output[2338] + last_layer_output[2339] + last_layer_output[2340] + last_layer_output[2341] + last_layer_output[2342] + last_layer_output[2343] + last_layer_output[2344] + last_layer_output[2345] + last_layer_output[2346] + last_layer_output[2347] + last_layer_output[2348] + last_layer_output[2349] + last_layer_output[2350] + last_layer_output[2351] + last_layer_output[2352] + last_layer_output[2353] + last_layer_output[2354] + last_layer_output[2355] + last_layer_output[2356] + last_layer_output[2357] + last_layer_output[2358] + last_layer_output[2359] + last_layer_output[2360] + last_layer_output[2361] + last_layer_output[2362] + last_layer_output[2363] + last_layer_output[2364] + last_layer_output[2365] + last_layer_output[2366] + last_layer_output[2367] + last_layer_output[2368] + last_layer_output[2369] + last_layer_output[2370] + last_layer_output[2371] + last_layer_output[2372] + last_layer_output[2373] + last_layer_output[2374] + last_layer_output[2375] + last_layer_output[2376] + last_layer_output[2377] + last_layer_output[2378] + last_layer_output[2379] + last_layer_output[2380] + last_layer_output[2381] + last_layer_output[2382] + last_layer_output[2383] + last_layer_output[2384] + last_layer_output[2385] + last_layer_output[2386] + last_layer_output[2387] + last_layer_output[2388] + last_layer_output[2389] + last_layer_output[2390] + last_layer_output[2391] + last_layer_output[2392] + last_layer_output[2393] + last_layer_output[2394] + last_layer_output[2395] + last_layer_output[2396] + last_layer_output[2397] + last_layer_output[2398] + last_layer_output[2399];
      assign result[3] = last_layer_output[2400] + last_layer_output[2401] + last_layer_output[2402] + last_layer_output[2403] + last_layer_output[2404] + last_layer_output[2405] + last_layer_output[2406] + last_layer_output[2407] + last_layer_output[2408] + last_layer_output[2409] + last_layer_output[2410] + last_layer_output[2411] + last_layer_output[2412] + last_layer_output[2413] + last_layer_output[2414] + last_layer_output[2415] + last_layer_output[2416] + last_layer_output[2417] + last_layer_output[2418] + last_layer_output[2419] + last_layer_output[2420] + last_layer_output[2421] + last_layer_output[2422] + last_layer_output[2423] + last_layer_output[2424] + last_layer_output[2425] + last_layer_output[2426] + last_layer_output[2427] + last_layer_output[2428] + last_layer_output[2429] + last_layer_output[2430] + last_layer_output[2431] + last_layer_output[2432] + last_layer_output[2433] + last_layer_output[2434] + last_layer_output[2435] + last_layer_output[2436] + last_layer_output[2437] + last_layer_output[2438] + last_layer_output[2439] + last_layer_output[2440] + last_layer_output[2441] + last_layer_output[2442] + last_layer_output[2443] + last_layer_output[2444] + last_layer_output[2445] + last_layer_output[2446] + last_layer_output[2447] + last_layer_output[2448] + last_layer_output[2449] + last_layer_output[2450] + last_layer_output[2451] + last_layer_output[2452] + last_layer_output[2453] + last_layer_output[2454] + last_layer_output[2455] + last_layer_output[2456] + last_layer_output[2457] + last_layer_output[2458] + last_layer_output[2459] + last_layer_output[2460] + last_layer_output[2461] + last_layer_output[2462] + last_layer_output[2463] + last_layer_output[2464] + last_layer_output[2465] + last_layer_output[2466] + last_layer_output[2467] + last_layer_output[2468] + last_layer_output[2469] + last_layer_output[2470] + last_layer_output[2471] + last_layer_output[2472] + last_layer_output[2473] + last_layer_output[2474] + last_layer_output[2475] + last_layer_output[2476] + last_layer_output[2477] + last_layer_output[2478] + last_layer_output[2479] + last_layer_output[2480] + last_layer_output[2481] + last_layer_output[2482] + last_layer_output[2483] + last_layer_output[2484] + last_layer_output[2485] + last_layer_output[2486] + last_layer_output[2487] + last_layer_output[2488] + last_layer_output[2489] + last_layer_output[2490] + last_layer_output[2491] + last_layer_output[2492] + last_layer_output[2493] + last_layer_output[2494] + last_layer_output[2495] + last_layer_output[2496] + last_layer_output[2497] + last_layer_output[2498] + last_layer_output[2499] + last_layer_output[2500] + last_layer_output[2501] + last_layer_output[2502] + last_layer_output[2503] + last_layer_output[2504] + last_layer_output[2505] + last_layer_output[2506] + last_layer_output[2507] + last_layer_output[2508] + last_layer_output[2509] + last_layer_output[2510] + last_layer_output[2511] + last_layer_output[2512] + last_layer_output[2513] + last_layer_output[2514] + last_layer_output[2515] + last_layer_output[2516] + last_layer_output[2517] + last_layer_output[2518] + last_layer_output[2519] + last_layer_output[2520] + last_layer_output[2521] + last_layer_output[2522] + last_layer_output[2523] + last_layer_output[2524] + last_layer_output[2525] + last_layer_output[2526] + last_layer_output[2527] + last_layer_output[2528] + last_layer_output[2529] + last_layer_output[2530] + last_layer_output[2531] + last_layer_output[2532] + last_layer_output[2533] + last_layer_output[2534] + last_layer_output[2535] + last_layer_output[2536] + last_layer_output[2537] + last_layer_output[2538] + last_layer_output[2539] + last_layer_output[2540] + last_layer_output[2541] + last_layer_output[2542] + last_layer_output[2543] + last_layer_output[2544] + last_layer_output[2545] + last_layer_output[2546] + last_layer_output[2547] + last_layer_output[2548] + last_layer_output[2549] + last_layer_output[2550] + last_layer_output[2551] + last_layer_output[2552] + last_layer_output[2553] + last_layer_output[2554] + last_layer_output[2555] + last_layer_output[2556] + last_layer_output[2557] + last_layer_output[2558] + last_layer_output[2559] + last_layer_output[2560] + last_layer_output[2561] + last_layer_output[2562] + last_layer_output[2563] + last_layer_output[2564] + last_layer_output[2565] + last_layer_output[2566] + last_layer_output[2567] + last_layer_output[2568] + last_layer_output[2569] + last_layer_output[2570] + last_layer_output[2571] + last_layer_output[2572] + last_layer_output[2573] + last_layer_output[2574] + last_layer_output[2575] + last_layer_output[2576] + last_layer_output[2577] + last_layer_output[2578] + last_layer_output[2579] + last_layer_output[2580] + last_layer_output[2581] + last_layer_output[2582] + last_layer_output[2583] + last_layer_output[2584] + last_layer_output[2585] + last_layer_output[2586] + last_layer_output[2587] + last_layer_output[2588] + last_layer_output[2589] + last_layer_output[2590] + last_layer_output[2591] + last_layer_output[2592] + last_layer_output[2593] + last_layer_output[2594] + last_layer_output[2595] + last_layer_output[2596] + last_layer_output[2597] + last_layer_output[2598] + last_layer_output[2599] + last_layer_output[2600] + last_layer_output[2601] + last_layer_output[2602] + last_layer_output[2603] + last_layer_output[2604] + last_layer_output[2605] + last_layer_output[2606] + last_layer_output[2607] + last_layer_output[2608] + last_layer_output[2609] + last_layer_output[2610] + last_layer_output[2611] + last_layer_output[2612] + last_layer_output[2613] + last_layer_output[2614] + last_layer_output[2615] + last_layer_output[2616] + last_layer_output[2617] + last_layer_output[2618] + last_layer_output[2619] + last_layer_output[2620] + last_layer_output[2621] + last_layer_output[2622] + last_layer_output[2623] + last_layer_output[2624] + last_layer_output[2625] + last_layer_output[2626] + last_layer_output[2627] + last_layer_output[2628] + last_layer_output[2629] + last_layer_output[2630] + last_layer_output[2631] + last_layer_output[2632] + last_layer_output[2633] + last_layer_output[2634] + last_layer_output[2635] + last_layer_output[2636] + last_layer_output[2637] + last_layer_output[2638] + last_layer_output[2639] + last_layer_output[2640] + last_layer_output[2641] + last_layer_output[2642] + last_layer_output[2643] + last_layer_output[2644] + last_layer_output[2645] + last_layer_output[2646] + last_layer_output[2647] + last_layer_output[2648] + last_layer_output[2649] + last_layer_output[2650] + last_layer_output[2651] + last_layer_output[2652] + last_layer_output[2653] + last_layer_output[2654] + last_layer_output[2655] + last_layer_output[2656] + last_layer_output[2657] + last_layer_output[2658] + last_layer_output[2659] + last_layer_output[2660] + last_layer_output[2661] + last_layer_output[2662] + last_layer_output[2663] + last_layer_output[2664] + last_layer_output[2665] + last_layer_output[2666] + last_layer_output[2667] + last_layer_output[2668] + last_layer_output[2669] + last_layer_output[2670] + last_layer_output[2671] + last_layer_output[2672] + last_layer_output[2673] + last_layer_output[2674] + last_layer_output[2675] + last_layer_output[2676] + last_layer_output[2677] + last_layer_output[2678] + last_layer_output[2679] + last_layer_output[2680] + last_layer_output[2681] + last_layer_output[2682] + last_layer_output[2683] + last_layer_output[2684] + last_layer_output[2685] + last_layer_output[2686] + last_layer_output[2687] + last_layer_output[2688] + last_layer_output[2689] + last_layer_output[2690] + last_layer_output[2691] + last_layer_output[2692] + last_layer_output[2693] + last_layer_output[2694] + last_layer_output[2695] + last_layer_output[2696] + last_layer_output[2697] + last_layer_output[2698] + last_layer_output[2699] + last_layer_output[2700] + last_layer_output[2701] + last_layer_output[2702] + last_layer_output[2703] + last_layer_output[2704] + last_layer_output[2705] + last_layer_output[2706] + last_layer_output[2707] + last_layer_output[2708] + last_layer_output[2709] + last_layer_output[2710] + last_layer_output[2711] + last_layer_output[2712] + last_layer_output[2713] + last_layer_output[2714] + last_layer_output[2715] + last_layer_output[2716] + last_layer_output[2717] + last_layer_output[2718] + last_layer_output[2719] + last_layer_output[2720] + last_layer_output[2721] + last_layer_output[2722] + last_layer_output[2723] + last_layer_output[2724] + last_layer_output[2725] + last_layer_output[2726] + last_layer_output[2727] + last_layer_output[2728] + last_layer_output[2729] + last_layer_output[2730] + last_layer_output[2731] + last_layer_output[2732] + last_layer_output[2733] + last_layer_output[2734] + last_layer_output[2735] + last_layer_output[2736] + last_layer_output[2737] + last_layer_output[2738] + last_layer_output[2739] + last_layer_output[2740] + last_layer_output[2741] + last_layer_output[2742] + last_layer_output[2743] + last_layer_output[2744] + last_layer_output[2745] + last_layer_output[2746] + last_layer_output[2747] + last_layer_output[2748] + last_layer_output[2749] + last_layer_output[2750] + last_layer_output[2751] + last_layer_output[2752] + last_layer_output[2753] + last_layer_output[2754] + last_layer_output[2755] + last_layer_output[2756] + last_layer_output[2757] + last_layer_output[2758] + last_layer_output[2759] + last_layer_output[2760] + last_layer_output[2761] + last_layer_output[2762] + last_layer_output[2763] + last_layer_output[2764] + last_layer_output[2765] + last_layer_output[2766] + last_layer_output[2767] + last_layer_output[2768] + last_layer_output[2769] + last_layer_output[2770] + last_layer_output[2771] + last_layer_output[2772] + last_layer_output[2773] + last_layer_output[2774] + last_layer_output[2775] + last_layer_output[2776] + last_layer_output[2777] + last_layer_output[2778] + last_layer_output[2779] + last_layer_output[2780] + last_layer_output[2781] + last_layer_output[2782] + last_layer_output[2783] + last_layer_output[2784] + last_layer_output[2785] + last_layer_output[2786] + last_layer_output[2787] + last_layer_output[2788] + last_layer_output[2789] + last_layer_output[2790] + last_layer_output[2791] + last_layer_output[2792] + last_layer_output[2793] + last_layer_output[2794] + last_layer_output[2795] + last_layer_output[2796] + last_layer_output[2797] + last_layer_output[2798] + last_layer_output[2799] + last_layer_output[2800] + last_layer_output[2801] + last_layer_output[2802] + last_layer_output[2803] + last_layer_output[2804] + last_layer_output[2805] + last_layer_output[2806] + last_layer_output[2807] + last_layer_output[2808] + last_layer_output[2809] + last_layer_output[2810] + last_layer_output[2811] + last_layer_output[2812] + last_layer_output[2813] + last_layer_output[2814] + last_layer_output[2815] + last_layer_output[2816] + last_layer_output[2817] + last_layer_output[2818] + last_layer_output[2819] + last_layer_output[2820] + last_layer_output[2821] + last_layer_output[2822] + last_layer_output[2823] + last_layer_output[2824] + last_layer_output[2825] + last_layer_output[2826] + last_layer_output[2827] + last_layer_output[2828] + last_layer_output[2829] + last_layer_output[2830] + last_layer_output[2831] + last_layer_output[2832] + last_layer_output[2833] + last_layer_output[2834] + last_layer_output[2835] + last_layer_output[2836] + last_layer_output[2837] + last_layer_output[2838] + last_layer_output[2839] + last_layer_output[2840] + last_layer_output[2841] + last_layer_output[2842] + last_layer_output[2843] + last_layer_output[2844] + last_layer_output[2845] + last_layer_output[2846] + last_layer_output[2847] + last_layer_output[2848] + last_layer_output[2849] + last_layer_output[2850] + last_layer_output[2851] + last_layer_output[2852] + last_layer_output[2853] + last_layer_output[2854] + last_layer_output[2855] + last_layer_output[2856] + last_layer_output[2857] + last_layer_output[2858] + last_layer_output[2859] + last_layer_output[2860] + last_layer_output[2861] + last_layer_output[2862] + last_layer_output[2863] + last_layer_output[2864] + last_layer_output[2865] + last_layer_output[2866] + last_layer_output[2867] + last_layer_output[2868] + last_layer_output[2869] + last_layer_output[2870] + last_layer_output[2871] + last_layer_output[2872] + last_layer_output[2873] + last_layer_output[2874] + last_layer_output[2875] + last_layer_output[2876] + last_layer_output[2877] + last_layer_output[2878] + last_layer_output[2879] + last_layer_output[2880] + last_layer_output[2881] + last_layer_output[2882] + last_layer_output[2883] + last_layer_output[2884] + last_layer_output[2885] + last_layer_output[2886] + last_layer_output[2887] + last_layer_output[2888] + last_layer_output[2889] + last_layer_output[2890] + last_layer_output[2891] + last_layer_output[2892] + last_layer_output[2893] + last_layer_output[2894] + last_layer_output[2895] + last_layer_output[2896] + last_layer_output[2897] + last_layer_output[2898] + last_layer_output[2899] + last_layer_output[2900] + last_layer_output[2901] + last_layer_output[2902] + last_layer_output[2903] + last_layer_output[2904] + last_layer_output[2905] + last_layer_output[2906] + last_layer_output[2907] + last_layer_output[2908] + last_layer_output[2909] + last_layer_output[2910] + last_layer_output[2911] + last_layer_output[2912] + last_layer_output[2913] + last_layer_output[2914] + last_layer_output[2915] + last_layer_output[2916] + last_layer_output[2917] + last_layer_output[2918] + last_layer_output[2919] + last_layer_output[2920] + last_layer_output[2921] + last_layer_output[2922] + last_layer_output[2923] + last_layer_output[2924] + last_layer_output[2925] + last_layer_output[2926] + last_layer_output[2927] + last_layer_output[2928] + last_layer_output[2929] + last_layer_output[2930] + last_layer_output[2931] + last_layer_output[2932] + last_layer_output[2933] + last_layer_output[2934] + last_layer_output[2935] + last_layer_output[2936] + last_layer_output[2937] + last_layer_output[2938] + last_layer_output[2939] + last_layer_output[2940] + last_layer_output[2941] + last_layer_output[2942] + last_layer_output[2943] + last_layer_output[2944] + last_layer_output[2945] + last_layer_output[2946] + last_layer_output[2947] + last_layer_output[2948] + last_layer_output[2949] + last_layer_output[2950] + last_layer_output[2951] + last_layer_output[2952] + last_layer_output[2953] + last_layer_output[2954] + last_layer_output[2955] + last_layer_output[2956] + last_layer_output[2957] + last_layer_output[2958] + last_layer_output[2959] + last_layer_output[2960] + last_layer_output[2961] + last_layer_output[2962] + last_layer_output[2963] + last_layer_output[2964] + last_layer_output[2965] + last_layer_output[2966] + last_layer_output[2967] + last_layer_output[2968] + last_layer_output[2969] + last_layer_output[2970] + last_layer_output[2971] + last_layer_output[2972] + last_layer_output[2973] + last_layer_output[2974] + last_layer_output[2975] + last_layer_output[2976] + last_layer_output[2977] + last_layer_output[2978] + last_layer_output[2979] + last_layer_output[2980] + last_layer_output[2981] + last_layer_output[2982] + last_layer_output[2983] + last_layer_output[2984] + last_layer_output[2985] + last_layer_output[2986] + last_layer_output[2987] + last_layer_output[2988] + last_layer_output[2989] + last_layer_output[2990] + last_layer_output[2991] + last_layer_output[2992] + last_layer_output[2993] + last_layer_output[2994] + last_layer_output[2995] + last_layer_output[2996] + last_layer_output[2997] + last_layer_output[2998] + last_layer_output[2999] + last_layer_output[3000] + last_layer_output[3001] + last_layer_output[3002] + last_layer_output[3003] + last_layer_output[3004] + last_layer_output[3005] + last_layer_output[3006] + last_layer_output[3007] + last_layer_output[3008] + last_layer_output[3009] + last_layer_output[3010] + last_layer_output[3011] + last_layer_output[3012] + last_layer_output[3013] + last_layer_output[3014] + last_layer_output[3015] + last_layer_output[3016] + last_layer_output[3017] + last_layer_output[3018] + last_layer_output[3019] + last_layer_output[3020] + last_layer_output[3021] + last_layer_output[3022] + last_layer_output[3023] + last_layer_output[3024] + last_layer_output[3025] + last_layer_output[3026] + last_layer_output[3027] + last_layer_output[3028] + last_layer_output[3029] + last_layer_output[3030] + last_layer_output[3031] + last_layer_output[3032] + last_layer_output[3033] + last_layer_output[3034] + last_layer_output[3035] + last_layer_output[3036] + last_layer_output[3037] + last_layer_output[3038] + last_layer_output[3039] + last_layer_output[3040] + last_layer_output[3041] + last_layer_output[3042] + last_layer_output[3043] + last_layer_output[3044] + last_layer_output[3045] + last_layer_output[3046] + last_layer_output[3047] + last_layer_output[3048] + last_layer_output[3049] + last_layer_output[3050] + last_layer_output[3051] + last_layer_output[3052] + last_layer_output[3053] + last_layer_output[3054] + last_layer_output[3055] + last_layer_output[3056] + last_layer_output[3057] + last_layer_output[3058] + last_layer_output[3059] + last_layer_output[3060] + last_layer_output[3061] + last_layer_output[3062] + last_layer_output[3063] + last_layer_output[3064] + last_layer_output[3065] + last_layer_output[3066] + last_layer_output[3067] + last_layer_output[3068] + last_layer_output[3069] + last_layer_output[3070] + last_layer_output[3071] + last_layer_output[3072] + last_layer_output[3073] + last_layer_output[3074] + last_layer_output[3075] + last_layer_output[3076] + last_layer_output[3077] + last_layer_output[3078] + last_layer_output[3079] + last_layer_output[3080] + last_layer_output[3081] + last_layer_output[3082] + last_layer_output[3083] + last_layer_output[3084] + last_layer_output[3085] + last_layer_output[3086] + last_layer_output[3087] + last_layer_output[3088] + last_layer_output[3089] + last_layer_output[3090] + last_layer_output[3091] + last_layer_output[3092] + last_layer_output[3093] + last_layer_output[3094] + last_layer_output[3095] + last_layer_output[3096] + last_layer_output[3097] + last_layer_output[3098] + last_layer_output[3099] + last_layer_output[3100] + last_layer_output[3101] + last_layer_output[3102] + last_layer_output[3103] + last_layer_output[3104] + last_layer_output[3105] + last_layer_output[3106] + last_layer_output[3107] + last_layer_output[3108] + last_layer_output[3109] + last_layer_output[3110] + last_layer_output[3111] + last_layer_output[3112] + last_layer_output[3113] + last_layer_output[3114] + last_layer_output[3115] + last_layer_output[3116] + last_layer_output[3117] + last_layer_output[3118] + last_layer_output[3119] + last_layer_output[3120] + last_layer_output[3121] + last_layer_output[3122] + last_layer_output[3123] + last_layer_output[3124] + last_layer_output[3125] + last_layer_output[3126] + last_layer_output[3127] + last_layer_output[3128] + last_layer_output[3129] + last_layer_output[3130] + last_layer_output[3131] + last_layer_output[3132] + last_layer_output[3133] + last_layer_output[3134] + last_layer_output[3135] + last_layer_output[3136] + last_layer_output[3137] + last_layer_output[3138] + last_layer_output[3139] + last_layer_output[3140] + last_layer_output[3141] + last_layer_output[3142] + last_layer_output[3143] + last_layer_output[3144] + last_layer_output[3145] + last_layer_output[3146] + last_layer_output[3147] + last_layer_output[3148] + last_layer_output[3149] + last_layer_output[3150] + last_layer_output[3151] + last_layer_output[3152] + last_layer_output[3153] + last_layer_output[3154] + last_layer_output[3155] + last_layer_output[3156] + last_layer_output[3157] + last_layer_output[3158] + last_layer_output[3159] + last_layer_output[3160] + last_layer_output[3161] + last_layer_output[3162] + last_layer_output[3163] + last_layer_output[3164] + last_layer_output[3165] + last_layer_output[3166] + last_layer_output[3167] + last_layer_output[3168] + last_layer_output[3169] + last_layer_output[3170] + last_layer_output[3171] + last_layer_output[3172] + last_layer_output[3173] + last_layer_output[3174] + last_layer_output[3175] + last_layer_output[3176] + last_layer_output[3177] + last_layer_output[3178] + last_layer_output[3179] + last_layer_output[3180] + last_layer_output[3181] + last_layer_output[3182] + last_layer_output[3183] + last_layer_output[3184] + last_layer_output[3185] + last_layer_output[3186] + last_layer_output[3187] + last_layer_output[3188] + last_layer_output[3189] + last_layer_output[3190] + last_layer_output[3191] + last_layer_output[3192] + last_layer_output[3193] + last_layer_output[3194] + last_layer_output[3195] + last_layer_output[3196] + last_layer_output[3197] + last_layer_output[3198] + last_layer_output[3199];
      assign result[4] = last_layer_output[3200] + last_layer_output[3201] + last_layer_output[3202] + last_layer_output[3203] + last_layer_output[3204] + last_layer_output[3205] + last_layer_output[3206] + last_layer_output[3207] + last_layer_output[3208] + last_layer_output[3209] + last_layer_output[3210] + last_layer_output[3211] + last_layer_output[3212] + last_layer_output[3213] + last_layer_output[3214] + last_layer_output[3215] + last_layer_output[3216] + last_layer_output[3217] + last_layer_output[3218] + last_layer_output[3219] + last_layer_output[3220] + last_layer_output[3221] + last_layer_output[3222] + last_layer_output[3223] + last_layer_output[3224] + last_layer_output[3225] + last_layer_output[3226] + last_layer_output[3227] + last_layer_output[3228] + last_layer_output[3229] + last_layer_output[3230] + last_layer_output[3231] + last_layer_output[3232] + last_layer_output[3233] + last_layer_output[3234] + last_layer_output[3235] + last_layer_output[3236] + last_layer_output[3237] + last_layer_output[3238] + last_layer_output[3239] + last_layer_output[3240] + last_layer_output[3241] + last_layer_output[3242] + last_layer_output[3243] + last_layer_output[3244] + last_layer_output[3245] + last_layer_output[3246] + last_layer_output[3247] + last_layer_output[3248] + last_layer_output[3249] + last_layer_output[3250] + last_layer_output[3251] + last_layer_output[3252] + last_layer_output[3253] + last_layer_output[3254] + last_layer_output[3255] + last_layer_output[3256] + last_layer_output[3257] + last_layer_output[3258] + last_layer_output[3259] + last_layer_output[3260] + last_layer_output[3261] + last_layer_output[3262] + last_layer_output[3263] + last_layer_output[3264] + last_layer_output[3265] + last_layer_output[3266] + last_layer_output[3267] + last_layer_output[3268] + last_layer_output[3269] + last_layer_output[3270] + last_layer_output[3271] + last_layer_output[3272] + last_layer_output[3273] + last_layer_output[3274] + last_layer_output[3275] + last_layer_output[3276] + last_layer_output[3277] + last_layer_output[3278] + last_layer_output[3279] + last_layer_output[3280] + last_layer_output[3281] + last_layer_output[3282] + last_layer_output[3283] + last_layer_output[3284] + last_layer_output[3285] + last_layer_output[3286] + last_layer_output[3287] + last_layer_output[3288] + last_layer_output[3289] + last_layer_output[3290] + last_layer_output[3291] + last_layer_output[3292] + last_layer_output[3293] + last_layer_output[3294] + last_layer_output[3295] + last_layer_output[3296] + last_layer_output[3297] + last_layer_output[3298] + last_layer_output[3299] + last_layer_output[3300] + last_layer_output[3301] + last_layer_output[3302] + last_layer_output[3303] + last_layer_output[3304] + last_layer_output[3305] + last_layer_output[3306] + last_layer_output[3307] + last_layer_output[3308] + last_layer_output[3309] + last_layer_output[3310] + last_layer_output[3311] + last_layer_output[3312] + last_layer_output[3313] + last_layer_output[3314] + last_layer_output[3315] + last_layer_output[3316] + last_layer_output[3317] + last_layer_output[3318] + last_layer_output[3319] + last_layer_output[3320] + last_layer_output[3321] + last_layer_output[3322] + last_layer_output[3323] + last_layer_output[3324] + last_layer_output[3325] + last_layer_output[3326] + last_layer_output[3327] + last_layer_output[3328] + last_layer_output[3329] + last_layer_output[3330] + last_layer_output[3331] + last_layer_output[3332] + last_layer_output[3333] + last_layer_output[3334] + last_layer_output[3335] + last_layer_output[3336] + last_layer_output[3337] + last_layer_output[3338] + last_layer_output[3339] + last_layer_output[3340] + last_layer_output[3341] + last_layer_output[3342] + last_layer_output[3343] + last_layer_output[3344] + last_layer_output[3345] + last_layer_output[3346] + last_layer_output[3347] + last_layer_output[3348] + last_layer_output[3349] + last_layer_output[3350] + last_layer_output[3351] + last_layer_output[3352] + last_layer_output[3353] + last_layer_output[3354] + last_layer_output[3355] + last_layer_output[3356] + last_layer_output[3357] + last_layer_output[3358] + last_layer_output[3359] + last_layer_output[3360] + last_layer_output[3361] + last_layer_output[3362] + last_layer_output[3363] + last_layer_output[3364] + last_layer_output[3365] + last_layer_output[3366] + last_layer_output[3367] + last_layer_output[3368] + last_layer_output[3369] + last_layer_output[3370] + last_layer_output[3371] + last_layer_output[3372] + last_layer_output[3373] + last_layer_output[3374] + last_layer_output[3375] + last_layer_output[3376] + last_layer_output[3377] + last_layer_output[3378] + last_layer_output[3379] + last_layer_output[3380] + last_layer_output[3381] + last_layer_output[3382] + last_layer_output[3383] + last_layer_output[3384] + last_layer_output[3385] + last_layer_output[3386] + last_layer_output[3387] + last_layer_output[3388] + last_layer_output[3389] + last_layer_output[3390] + last_layer_output[3391] + last_layer_output[3392] + last_layer_output[3393] + last_layer_output[3394] + last_layer_output[3395] + last_layer_output[3396] + last_layer_output[3397] + last_layer_output[3398] + last_layer_output[3399] + last_layer_output[3400] + last_layer_output[3401] + last_layer_output[3402] + last_layer_output[3403] + last_layer_output[3404] + last_layer_output[3405] + last_layer_output[3406] + last_layer_output[3407] + last_layer_output[3408] + last_layer_output[3409] + last_layer_output[3410] + last_layer_output[3411] + last_layer_output[3412] + last_layer_output[3413] + last_layer_output[3414] + last_layer_output[3415] + last_layer_output[3416] + last_layer_output[3417] + last_layer_output[3418] + last_layer_output[3419] + last_layer_output[3420] + last_layer_output[3421] + last_layer_output[3422] + last_layer_output[3423] + last_layer_output[3424] + last_layer_output[3425] + last_layer_output[3426] + last_layer_output[3427] + last_layer_output[3428] + last_layer_output[3429] + last_layer_output[3430] + last_layer_output[3431] + last_layer_output[3432] + last_layer_output[3433] + last_layer_output[3434] + last_layer_output[3435] + last_layer_output[3436] + last_layer_output[3437] + last_layer_output[3438] + last_layer_output[3439] + last_layer_output[3440] + last_layer_output[3441] + last_layer_output[3442] + last_layer_output[3443] + last_layer_output[3444] + last_layer_output[3445] + last_layer_output[3446] + last_layer_output[3447] + last_layer_output[3448] + last_layer_output[3449] + last_layer_output[3450] + last_layer_output[3451] + last_layer_output[3452] + last_layer_output[3453] + last_layer_output[3454] + last_layer_output[3455] + last_layer_output[3456] + last_layer_output[3457] + last_layer_output[3458] + last_layer_output[3459] + last_layer_output[3460] + last_layer_output[3461] + last_layer_output[3462] + last_layer_output[3463] + last_layer_output[3464] + last_layer_output[3465] + last_layer_output[3466] + last_layer_output[3467] + last_layer_output[3468] + last_layer_output[3469] + last_layer_output[3470] + last_layer_output[3471] + last_layer_output[3472] + last_layer_output[3473] + last_layer_output[3474] + last_layer_output[3475] + last_layer_output[3476] + last_layer_output[3477] + last_layer_output[3478] + last_layer_output[3479] + last_layer_output[3480] + last_layer_output[3481] + last_layer_output[3482] + last_layer_output[3483] + last_layer_output[3484] + last_layer_output[3485] + last_layer_output[3486] + last_layer_output[3487] + last_layer_output[3488] + last_layer_output[3489] + last_layer_output[3490] + last_layer_output[3491] + last_layer_output[3492] + last_layer_output[3493] + last_layer_output[3494] + last_layer_output[3495] + last_layer_output[3496] + last_layer_output[3497] + last_layer_output[3498] + last_layer_output[3499] + last_layer_output[3500] + last_layer_output[3501] + last_layer_output[3502] + last_layer_output[3503] + last_layer_output[3504] + last_layer_output[3505] + last_layer_output[3506] + last_layer_output[3507] + last_layer_output[3508] + last_layer_output[3509] + last_layer_output[3510] + last_layer_output[3511] + last_layer_output[3512] + last_layer_output[3513] + last_layer_output[3514] + last_layer_output[3515] + last_layer_output[3516] + last_layer_output[3517] + last_layer_output[3518] + last_layer_output[3519] + last_layer_output[3520] + last_layer_output[3521] + last_layer_output[3522] + last_layer_output[3523] + last_layer_output[3524] + last_layer_output[3525] + last_layer_output[3526] + last_layer_output[3527] + last_layer_output[3528] + last_layer_output[3529] + last_layer_output[3530] + last_layer_output[3531] + last_layer_output[3532] + last_layer_output[3533] + last_layer_output[3534] + last_layer_output[3535] + last_layer_output[3536] + last_layer_output[3537] + last_layer_output[3538] + last_layer_output[3539] + last_layer_output[3540] + last_layer_output[3541] + last_layer_output[3542] + last_layer_output[3543] + last_layer_output[3544] + last_layer_output[3545] + last_layer_output[3546] + last_layer_output[3547] + last_layer_output[3548] + last_layer_output[3549] + last_layer_output[3550] + last_layer_output[3551] + last_layer_output[3552] + last_layer_output[3553] + last_layer_output[3554] + last_layer_output[3555] + last_layer_output[3556] + last_layer_output[3557] + last_layer_output[3558] + last_layer_output[3559] + last_layer_output[3560] + last_layer_output[3561] + last_layer_output[3562] + last_layer_output[3563] + last_layer_output[3564] + last_layer_output[3565] + last_layer_output[3566] + last_layer_output[3567] + last_layer_output[3568] + last_layer_output[3569] + last_layer_output[3570] + last_layer_output[3571] + last_layer_output[3572] + last_layer_output[3573] + last_layer_output[3574] + last_layer_output[3575] + last_layer_output[3576] + last_layer_output[3577] + last_layer_output[3578] + last_layer_output[3579] + last_layer_output[3580] + last_layer_output[3581] + last_layer_output[3582] + last_layer_output[3583] + last_layer_output[3584] + last_layer_output[3585] + last_layer_output[3586] + last_layer_output[3587] + last_layer_output[3588] + last_layer_output[3589] + last_layer_output[3590] + last_layer_output[3591] + last_layer_output[3592] + last_layer_output[3593] + last_layer_output[3594] + last_layer_output[3595] + last_layer_output[3596] + last_layer_output[3597] + last_layer_output[3598] + last_layer_output[3599] + last_layer_output[3600] + last_layer_output[3601] + last_layer_output[3602] + last_layer_output[3603] + last_layer_output[3604] + last_layer_output[3605] + last_layer_output[3606] + last_layer_output[3607] + last_layer_output[3608] + last_layer_output[3609] + last_layer_output[3610] + last_layer_output[3611] + last_layer_output[3612] + last_layer_output[3613] + last_layer_output[3614] + last_layer_output[3615] + last_layer_output[3616] + last_layer_output[3617] + last_layer_output[3618] + last_layer_output[3619] + last_layer_output[3620] + last_layer_output[3621] + last_layer_output[3622] + last_layer_output[3623] + last_layer_output[3624] + last_layer_output[3625] + last_layer_output[3626] + last_layer_output[3627] + last_layer_output[3628] + last_layer_output[3629] + last_layer_output[3630] + last_layer_output[3631] + last_layer_output[3632] + last_layer_output[3633] + last_layer_output[3634] + last_layer_output[3635] + last_layer_output[3636] + last_layer_output[3637] + last_layer_output[3638] + last_layer_output[3639] + last_layer_output[3640] + last_layer_output[3641] + last_layer_output[3642] + last_layer_output[3643] + last_layer_output[3644] + last_layer_output[3645] + last_layer_output[3646] + last_layer_output[3647] + last_layer_output[3648] + last_layer_output[3649] + last_layer_output[3650] + last_layer_output[3651] + last_layer_output[3652] + last_layer_output[3653] + last_layer_output[3654] + last_layer_output[3655] + last_layer_output[3656] + last_layer_output[3657] + last_layer_output[3658] + last_layer_output[3659] + last_layer_output[3660] + last_layer_output[3661] + last_layer_output[3662] + last_layer_output[3663] + last_layer_output[3664] + last_layer_output[3665] + last_layer_output[3666] + last_layer_output[3667] + last_layer_output[3668] + last_layer_output[3669] + last_layer_output[3670] + last_layer_output[3671] + last_layer_output[3672] + last_layer_output[3673] + last_layer_output[3674] + last_layer_output[3675] + last_layer_output[3676] + last_layer_output[3677] + last_layer_output[3678] + last_layer_output[3679] + last_layer_output[3680] + last_layer_output[3681] + last_layer_output[3682] + last_layer_output[3683] + last_layer_output[3684] + last_layer_output[3685] + last_layer_output[3686] + last_layer_output[3687] + last_layer_output[3688] + last_layer_output[3689] + last_layer_output[3690] + last_layer_output[3691] + last_layer_output[3692] + last_layer_output[3693] + last_layer_output[3694] + last_layer_output[3695] + last_layer_output[3696] + last_layer_output[3697] + last_layer_output[3698] + last_layer_output[3699] + last_layer_output[3700] + last_layer_output[3701] + last_layer_output[3702] + last_layer_output[3703] + last_layer_output[3704] + last_layer_output[3705] + last_layer_output[3706] + last_layer_output[3707] + last_layer_output[3708] + last_layer_output[3709] + last_layer_output[3710] + last_layer_output[3711] + last_layer_output[3712] + last_layer_output[3713] + last_layer_output[3714] + last_layer_output[3715] + last_layer_output[3716] + last_layer_output[3717] + last_layer_output[3718] + last_layer_output[3719] + last_layer_output[3720] + last_layer_output[3721] + last_layer_output[3722] + last_layer_output[3723] + last_layer_output[3724] + last_layer_output[3725] + last_layer_output[3726] + last_layer_output[3727] + last_layer_output[3728] + last_layer_output[3729] + last_layer_output[3730] + last_layer_output[3731] + last_layer_output[3732] + last_layer_output[3733] + last_layer_output[3734] + last_layer_output[3735] + last_layer_output[3736] + last_layer_output[3737] + last_layer_output[3738] + last_layer_output[3739] + last_layer_output[3740] + last_layer_output[3741] + last_layer_output[3742] + last_layer_output[3743] + last_layer_output[3744] + last_layer_output[3745] + last_layer_output[3746] + last_layer_output[3747] + last_layer_output[3748] + last_layer_output[3749] + last_layer_output[3750] + last_layer_output[3751] + last_layer_output[3752] + last_layer_output[3753] + last_layer_output[3754] + last_layer_output[3755] + last_layer_output[3756] + last_layer_output[3757] + last_layer_output[3758] + last_layer_output[3759] + last_layer_output[3760] + last_layer_output[3761] + last_layer_output[3762] + last_layer_output[3763] + last_layer_output[3764] + last_layer_output[3765] + last_layer_output[3766] + last_layer_output[3767] + last_layer_output[3768] + last_layer_output[3769] + last_layer_output[3770] + last_layer_output[3771] + last_layer_output[3772] + last_layer_output[3773] + last_layer_output[3774] + last_layer_output[3775] + last_layer_output[3776] + last_layer_output[3777] + last_layer_output[3778] + last_layer_output[3779] + last_layer_output[3780] + last_layer_output[3781] + last_layer_output[3782] + last_layer_output[3783] + last_layer_output[3784] + last_layer_output[3785] + last_layer_output[3786] + last_layer_output[3787] + last_layer_output[3788] + last_layer_output[3789] + last_layer_output[3790] + last_layer_output[3791] + last_layer_output[3792] + last_layer_output[3793] + last_layer_output[3794] + last_layer_output[3795] + last_layer_output[3796] + last_layer_output[3797] + last_layer_output[3798] + last_layer_output[3799] + last_layer_output[3800] + last_layer_output[3801] + last_layer_output[3802] + last_layer_output[3803] + last_layer_output[3804] + last_layer_output[3805] + last_layer_output[3806] + last_layer_output[3807] + last_layer_output[3808] + last_layer_output[3809] + last_layer_output[3810] + last_layer_output[3811] + last_layer_output[3812] + last_layer_output[3813] + last_layer_output[3814] + last_layer_output[3815] + last_layer_output[3816] + last_layer_output[3817] + last_layer_output[3818] + last_layer_output[3819] + last_layer_output[3820] + last_layer_output[3821] + last_layer_output[3822] + last_layer_output[3823] + last_layer_output[3824] + last_layer_output[3825] + last_layer_output[3826] + last_layer_output[3827] + last_layer_output[3828] + last_layer_output[3829] + last_layer_output[3830] + last_layer_output[3831] + last_layer_output[3832] + last_layer_output[3833] + last_layer_output[3834] + last_layer_output[3835] + last_layer_output[3836] + last_layer_output[3837] + last_layer_output[3838] + last_layer_output[3839] + last_layer_output[3840] + last_layer_output[3841] + last_layer_output[3842] + last_layer_output[3843] + last_layer_output[3844] + last_layer_output[3845] + last_layer_output[3846] + last_layer_output[3847] + last_layer_output[3848] + last_layer_output[3849] + last_layer_output[3850] + last_layer_output[3851] + last_layer_output[3852] + last_layer_output[3853] + last_layer_output[3854] + last_layer_output[3855] + last_layer_output[3856] + last_layer_output[3857] + last_layer_output[3858] + last_layer_output[3859] + last_layer_output[3860] + last_layer_output[3861] + last_layer_output[3862] + last_layer_output[3863] + last_layer_output[3864] + last_layer_output[3865] + last_layer_output[3866] + last_layer_output[3867] + last_layer_output[3868] + last_layer_output[3869] + last_layer_output[3870] + last_layer_output[3871] + last_layer_output[3872] + last_layer_output[3873] + last_layer_output[3874] + last_layer_output[3875] + last_layer_output[3876] + last_layer_output[3877] + last_layer_output[3878] + last_layer_output[3879] + last_layer_output[3880] + last_layer_output[3881] + last_layer_output[3882] + last_layer_output[3883] + last_layer_output[3884] + last_layer_output[3885] + last_layer_output[3886] + last_layer_output[3887] + last_layer_output[3888] + last_layer_output[3889] + last_layer_output[3890] + last_layer_output[3891] + last_layer_output[3892] + last_layer_output[3893] + last_layer_output[3894] + last_layer_output[3895] + last_layer_output[3896] + last_layer_output[3897] + last_layer_output[3898] + last_layer_output[3899] + last_layer_output[3900] + last_layer_output[3901] + last_layer_output[3902] + last_layer_output[3903] + last_layer_output[3904] + last_layer_output[3905] + last_layer_output[3906] + last_layer_output[3907] + last_layer_output[3908] + last_layer_output[3909] + last_layer_output[3910] + last_layer_output[3911] + last_layer_output[3912] + last_layer_output[3913] + last_layer_output[3914] + last_layer_output[3915] + last_layer_output[3916] + last_layer_output[3917] + last_layer_output[3918] + last_layer_output[3919] + last_layer_output[3920] + last_layer_output[3921] + last_layer_output[3922] + last_layer_output[3923] + last_layer_output[3924] + last_layer_output[3925] + last_layer_output[3926] + last_layer_output[3927] + last_layer_output[3928] + last_layer_output[3929] + last_layer_output[3930] + last_layer_output[3931] + last_layer_output[3932] + last_layer_output[3933] + last_layer_output[3934] + last_layer_output[3935] + last_layer_output[3936] + last_layer_output[3937] + last_layer_output[3938] + last_layer_output[3939] + last_layer_output[3940] + last_layer_output[3941] + last_layer_output[3942] + last_layer_output[3943] + last_layer_output[3944] + last_layer_output[3945] + last_layer_output[3946] + last_layer_output[3947] + last_layer_output[3948] + last_layer_output[3949] + last_layer_output[3950] + last_layer_output[3951] + last_layer_output[3952] + last_layer_output[3953] + last_layer_output[3954] + last_layer_output[3955] + last_layer_output[3956] + last_layer_output[3957] + last_layer_output[3958] + last_layer_output[3959] + last_layer_output[3960] + last_layer_output[3961] + last_layer_output[3962] + last_layer_output[3963] + last_layer_output[3964] + last_layer_output[3965] + last_layer_output[3966] + last_layer_output[3967] + last_layer_output[3968] + last_layer_output[3969] + last_layer_output[3970] + last_layer_output[3971] + last_layer_output[3972] + last_layer_output[3973] + last_layer_output[3974] + last_layer_output[3975] + last_layer_output[3976] + last_layer_output[3977] + last_layer_output[3978] + last_layer_output[3979] + last_layer_output[3980] + last_layer_output[3981] + last_layer_output[3982] + last_layer_output[3983] + last_layer_output[3984] + last_layer_output[3985] + last_layer_output[3986] + last_layer_output[3987] + last_layer_output[3988] + last_layer_output[3989] + last_layer_output[3990] + last_layer_output[3991] + last_layer_output[3992] + last_layer_output[3993] + last_layer_output[3994] + last_layer_output[3995] + last_layer_output[3996] + last_layer_output[3997] + last_layer_output[3998] + last_layer_output[3999];
      assign result[5] = last_layer_output[4000] + last_layer_output[4001] + last_layer_output[4002] + last_layer_output[4003] + last_layer_output[4004] + last_layer_output[4005] + last_layer_output[4006] + last_layer_output[4007] + last_layer_output[4008] + last_layer_output[4009] + last_layer_output[4010] + last_layer_output[4011] + last_layer_output[4012] + last_layer_output[4013] + last_layer_output[4014] + last_layer_output[4015] + last_layer_output[4016] + last_layer_output[4017] + last_layer_output[4018] + last_layer_output[4019] + last_layer_output[4020] + last_layer_output[4021] + last_layer_output[4022] + last_layer_output[4023] + last_layer_output[4024] + last_layer_output[4025] + last_layer_output[4026] + last_layer_output[4027] + last_layer_output[4028] + last_layer_output[4029] + last_layer_output[4030] + last_layer_output[4031] + last_layer_output[4032] + last_layer_output[4033] + last_layer_output[4034] + last_layer_output[4035] + last_layer_output[4036] + last_layer_output[4037] + last_layer_output[4038] + last_layer_output[4039] + last_layer_output[4040] + last_layer_output[4041] + last_layer_output[4042] + last_layer_output[4043] + last_layer_output[4044] + last_layer_output[4045] + last_layer_output[4046] + last_layer_output[4047] + last_layer_output[4048] + last_layer_output[4049] + last_layer_output[4050] + last_layer_output[4051] + last_layer_output[4052] + last_layer_output[4053] + last_layer_output[4054] + last_layer_output[4055] + last_layer_output[4056] + last_layer_output[4057] + last_layer_output[4058] + last_layer_output[4059] + last_layer_output[4060] + last_layer_output[4061] + last_layer_output[4062] + last_layer_output[4063] + last_layer_output[4064] + last_layer_output[4065] + last_layer_output[4066] + last_layer_output[4067] + last_layer_output[4068] + last_layer_output[4069] + last_layer_output[4070] + last_layer_output[4071] + last_layer_output[4072] + last_layer_output[4073] + last_layer_output[4074] + last_layer_output[4075] + last_layer_output[4076] + last_layer_output[4077] + last_layer_output[4078] + last_layer_output[4079] + last_layer_output[4080] + last_layer_output[4081] + last_layer_output[4082] + last_layer_output[4083] + last_layer_output[4084] + last_layer_output[4085] + last_layer_output[4086] + last_layer_output[4087] + last_layer_output[4088] + last_layer_output[4089] + last_layer_output[4090] + last_layer_output[4091] + last_layer_output[4092] + last_layer_output[4093] + last_layer_output[4094] + last_layer_output[4095] + last_layer_output[4096] + last_layer_output[4097] + last_layer_output[4098] + last_layer_output[4099] + last_layer_output[4100] + last_layer_output[4101] + last_layer_output[4102] + last_layer_output[4103] + last_layer_output[4104] + last_layer_output[4105] + last_layer_output[4106] + last_layer_output[4107] + last_layer_output[4108] + last_layer_output[4109] + last_layer_output[4110] + last_layer_output[4111] + last_layer_output[4112] + last_layer_output[4113] + last_layer_output[4114] + last_layer_output[4115] + last_layer_output[4116] + last_layer_output[4117] + last_layer_output[4118] + last_layer_output[4119] + last_layer_output[4120] + last_layer_output[4121] + last_layer_output[4122] + last_layer_output[4123] + last_layer_output[4124] + last_layer_output[4125] + last_layer_output[4126] + last_layer_output[4127] + last_layer_output[4128] + last_layer_output[4129] + last_layer_output[4130] + last_layer_output[4131] + last_layer_output[4132] + last_layer_output[4133] + last_layer_output[4134] + last_layer_output[4135] + last_layer_output[4136] + last_layer_output[4137] + last_layer_output[4138] + last_layer_output[4139] + last_layer_output[4140] + last_layer_output[4141] + last_layer_output[4142] + last_layer_output[4143] + last_layer_output[4144] + last_layer_output[4145] + last_layer_output[4146] + last_layer_output[4147] + last_layer_output[4148] + last_layer_output[4149] + last_layer_output[4150] + last_layer_output[4151] + last_layer_output[4152] + last_layer_output[4153] + last_layer_output[4154] + last_layer_output[4155] + last_layer_output[4156] + last_layer_output[4157] + last_layer_output[4158] + last_layer_output[4159] + last_layer_output[4160] + last_layer_output[4161] + last_layer_output[4162] + last_layer_output[4163] + last_layer_output[4164] + last_layer_output[4165] + last_layer_output[4166] + last_layer_output[4167] + last_layer_output[4168] + last_layer_output[4169] + last_layer_output[4170] + last_layer_output[4171] + last_layer_output[4172] + last_layer_output[4173] + last_layer_output[4174] + last_layer_output[4175] + last_layer_output[4176] + last_layer_output[4177] + last_layer_output[4178] + last_layer_output[4179] + last_layer_output[4180] + last_layer_output[4181] + last_layer_output[4182] + last_layer_output[4183] + last_layer_output[4184] + last_layer_output[4185] + last_layer_output[4186] + last_layer_output[4187] + last_layer_output[4188] + last_layer_output[4189] + last_layer_output[4190] + last_layer_output[4191] + last_layer_output[4192] + last_layer_output[4193] + last_layer_output[4194] + last_layer_output[4195] + last_layer_output[4196] + last_layer_output[4197] + last_layer_output[4198] + last_layer_output[4199] + last_layer_output[4200] + last_layer_output[4201] + last_layer_output[4202] + last_layer_output[4203] + last_layer_output[4204] + last_layer_output[4205] + last_layer_output[4206] + last_layer_output[4207] + last_layer_output[4208] + last_layer_output[4209] + last_layer_output[4210] + last_layer_output[4211] + last_layer_output[4212] + last_layer_output[4213] + last_layer_output[4214] + last_layer_output[4215] + last_layer_output[4216] + last_layer_output[4217] + last_layer_output[4218] + last_layer_output[4219] + last_layer_output[4220] + last_layer_output[4221] + last_layer_output[4222] + last_layer_output[4223] + last_layer_output[4224] + last_layer_output[4225] + last_layer_output[4226] + last_layer_output[4227] + last_layer_output[4228] + last_layer_output[4229] + last_layer_output[4230] + last_layer_output[4231] + last_layer_output[4232] + last_layer_output[4233] + last_layer_output[4234] + last_layer_output[4235] + last_layer_output[4236] + last_layer_output[4237] + last_layer_output[4238] + last_layer_output[4239] + last_layer_output[4240] + last_layer_output[4241] + last_layer_output[4242] + last_layer_output[4243] + last_layer_output[4244] + last_layer_output[4245] + last_layer_output[4246] + last_layer_output[4247] + last_layer_output[4248] + last_layer_output[4249] + last_layer_output[4250] + last_layer_output[4251] + last_layer_output[4252] + last_layer_output[4253] + last_layer_output[4254] + last_layer_output[4255] + last_layer_output[4256] + last_layer_output[4257] + last_layer_output[4258] + last_layer_output[4259] + last_layer_output[4260] + last_layer_output[4261] + last_layer_output[4262] + last_layer_output[4263] + last_layer_output[4264] + last_layer_output[4265] + last_layer_output[4266] + last_layer_output[4267] + last_layer_output[4268] + last_layer_output[4269] + last_layer_output[4270] + last_layer_output[4271] + last_layer_output[4272] + last_layer_output[4273] + last_layer_output[4274] + last_layer_output[4275] + last_layer_output[4276] + last_layer_output[4277] + last_layer_output[4278] + last_layer_output[4279] + last_layer_output[4280] + last_layer_output[4281] + last_layer_output[4282] + last_layer_output[4283] + last_layer_output[4284] + last_layer_output[4285] + last_layer_output[4286] + last_layer_output[4287] + last_layer_output[4288] + last_layer_output[4289] + last_layer_output[4290] + last_layer_output[4291] + last_layer_output[4292] + last_layer_output[4293] + last_layer_output[4294] + last_layer_output[4295] + last_layer_output[4296] + last_layer_output[4297] + last_layer_output[4298] + last_layer_output[4299] + last_layer_output[4300] + last_layer_output[4301] + last_layer_output[4302] + last_layer_output[4303] + last_layer_output[4304] + last_layer_output[4305] + last_layer_output[4306] + last_layer_output[4307] + last_layer_output[4308] + last_layer_output[4309] + last_layer_output[4310] + last_layer_output[4311] + last_layer_output[4312] + last_layer_output[4313] + last_layer_output[4314] + last_layer_output[4315] + last_layer_output[4316] + last_layer_output[4317] + last_layer_output[4318] + last_layer_output[4319] + last_layer_output[4320] + last_layer_output[4321] + last_layer_output[4322] + last_layer_output[4323] + last_layer_output[4324] + last_layer_output[4325] + last_layer_output[4326] + last_layer_output[4327] + last_layer_output[4328] + last_layer_output[4329] + last_layer_output[4330] + last_layer_output[4331] + last_layer_output[4332] + last_layer_output[4333] + last_layer_output[4334] + last_layer_output[4335] + last_layer_output[4336] + last_layer_output[4337] + last_layer_output[4338] + last_layer_output[4339] + last_layer_output[4340] + last_layer_output[4341] + last_layer_output[4342] + last_layer_output[4343] + last_layer_output[4344] + last_layer_output[4345] + last_layer_output[4346] + last_layer_output[4347] + last_layer_output[4348] + last_layer_output[4349] + last_layer_output[4350] + last_layer_output[4351] + last_layer_output[4352] + last_layer_output[4353] + last_layer_output[4354] + last_layer_output[4355] + last_layer_output[4356] + last_layer_output[4357] + last_layer_output[4358] + last_layer_output[4359] + last_layer_output[4360] + last_layer_output[4361] + last_layer_output[4362] + last_layer_output[4363] + last_layer_output[4364] + last_layer_output[4365] + last_layer_output[4366] + last_layer_output[4367] + last_layer_output[4368] + last_layer_output[4369] + last_layer_output[4370] + last_layer_output[4371] + last_layer_output[4372] + last_layer_output[4373] + last_layer_output[4374] + last_layer_output[4375] + last_layer_output[4376] + last_layer_output[4377] + last_layer_output[4378] + last_layer_output[4379] + last_layer_output[4380] + last_layer_output[4381] + last_layer_output[4382] + last_layer_output[4383] + last_layer_output[4384] + last_layer_output[4385] + last_layer_output[4386] + last_layer_output[4387] + last_layer_output[4388] + last_layer_output[4389] + last_layer_output[4390] + last_layer_output[4391] + last_layer_output[4392] + last_layer_output[4393] + last_layer_output[4394] + last_layer_output[4395] + last_layer_output[4396] + last_layer_output[4397] + last_layer_output[4398] + last_layer_output[4399] + last_layer_output[4400] + last_layer_output[4401] + last_layer_output[4402] + last_layer_output[4403] + last_layer_output[4404] + last_layer_output[4405] + last_layer_output[4406] + last_layer_output[4407] + last_layer_output[4408] + last_layer_output[4409] + last_layer_output[4410] + last_layer_output[4411] + last_layer_output[4412] + last_layer_output[4413] + last_layer_output[4414] + last_layer_output[4415] + last_layer_output[4416] + last_layer_output[4417] + last_layer_output[4418] + last_layer_output[4419] + last_layer_output[4420] + last_layer_output[4421] + last_layer_output[4422] + last_layer_output[4423] + last_layer_output[4424] + last_layer_output[4425] + last_layer_output[4426] + last_layer_output[4427] + last_layer_output[4428] + last_layer_output[4429] + last_layer_output[4430] + last_layer_output[4431] + last_layer_output[4432] + last_layer_output[4433] + last_layer_output[4434] + last_layer_output[4435] + last_layer_output[4436] + last_layer_output[4437] + last_layer_output[4438] + last_layer_output[4439] + last_layer_output[4440] + last_layer_output[4441] + last_layer_output[4442] + last_layer_output[4443] + last_layer_output[4444] + last_layer_output[4445] + last_layer_output[4446] + last_layer_output[4447] + last_layer_output[4448] + last_layer_output[4449] + last_layer_output[4450] + last_layer_output[4451] + last_layer_output[4452] + last_layer_output[4453] + last_layer_output[4454] + last_layer_output[4455] + last_layer_output[4456] + last_layer_output[4457] + last_layer_output[4458] + last_layer_output[4459] + last_layer_output[4460] + last_layer_output[4461] + last_layer_output[4462] + last_layer_output[4463] + last_layer_output[4464] + last_layer_output[4465] + last_layer_output[4466] + last_layer_output[4467] + last_layer_output[4468] + last_layer_output[4469] + last_layer_output[4470] + last_layer_output[4471] + last_layer_output[4472] + last_layer_output[4473] + last_layer_output[4474] + last_layer_output[4475] + last_layer_output[4476] + last_layer_output[4477] + last_layer_output[4478] + last_layer_output[4479] + last_layer_output[4480] + last_layer_output[4481] + last_layer_output[4482] + last_layer_output[4483] + last_layer_output[4484] + last_layer_output[4485] + last_layer_output[4486] + last_layer_output[4487] + last_layer_output[4488] + last_layer_output[4489] + last_layer_output[4490] + last_layer_output[4491] + last_layer_output[4492] + last_layer_output[4493] + last_layer_output[4494] + last_layer_output[4495] + last_layer_output[4496] + last_layer_output[4497] + last_layer_output[4498] + last_layer_output[4499] + last_layer_output[4500] + last_layer_output[4501] + last_layer_output[4502] + last_layer_output[4503] + last_layer_output[4504] + last_layer_output[4505] + last_layer_output[4506] + last_layer_output[4507] + last_layer_output[4508] + last_layer_output[4509] + last_layer_output[4510] + last_layer_output[4511] + last_layer_output[4512] + last_layer_output[4513] + last_layer_output[4514] + last_layer_output[4515] + last_layer_output[4516] + last_layer_output[4517] + last_layer_output[4518] + last_layer_output[4519] + last_layer_output[4520] + last_layer_output[4521] + last_layer_output[4522] + last_layer_output[4523] + last_layer_output[4524] + last_layer_output[4525] + last_layer_output[4526] + last_layer_output[4527] + last_layer_output[4528] + last_layer_output[4529] + last_layer_output[4530] + last_layer_output[4531] + last_layer_output[4532] + last_layer_output[4533] + last_layer_output[4534] + last_layer_output[4535] + last_layer_output[4536] + last_layer_output[4537] + last_layer_output[4538] + last_layer_output[4539] + last_layer_output[4540] + last_layer_output[4541] + last_layer_output[4542] + last_layer_output[4543] + last_layer_output[4544] + last_layer_output[4545] + last_layer_output[4546] + last_layer_output[4547] + last_layer_output[4548] + last_layer_output[4549] + last_layer_output[4550] + last_layer_output[4551] + last_layer_output[4552] + last_layer_output[4553] + last_layer_output[4554] + last_layer_output[4555] + last_layer_output[4556] + last_layer_output[4557] + last_layer_output[4558] + last_layer_output[4559] + last_layer_output[4560] + last_layer_output[4561] + last_layer_output[4562] + last_layer_output[4563] + last_layer_output[4564] + last_layer_output[4565] + last_layer_output[4566] + last_layer_output[4567] + last_layer_output[4568] + last_layer_output[4569] + last_layer_output[4570] + last_layer_output[4571] + last_layer_output[4572] + last_layer_output[4573] + last_layer_output[4574] + last_layer_output[4575] + last_layer_output[4576] + last_layer_output[4577] + last_layer_output[4578] + last_layer_output[4579] + last_layer_output[4580] + last_layer_output[4581] + last_layer_output[4582] + last_layer_output[4583] + last_layer_output[4584] + last_layer_output[4585] + last_layer_output[4586] + last_layer_output[4587] + last_layer_output[4588] + last_layer_output[4589] + last_layer_output[4590] + last_layer_output[4591] + last_layer_output[4592] + last_layer_output[4593] + last_layer_output[4594] + last_layer_output[4595] + last_layer_output[4596] + last_layer_output[4597] + last_layer_output[4598] + last_layer_output[4599] + last_layer_output[4600] + last_layer_output[4601] + last_layer_output[4602] + last_layer_output[4603] + last_layer_output[4604] + last_layer_output[4605] + last_layer_output[4606] + last_layer_output[4607] + last_layer_output[4608] + last_layer_output[4609] + last_layer_output[4610] + last_layer_output[4611] + last_layer_output[4612] + last_layer_output[4613] + last_layer_output[4614] + last_layer_output[4615] + last_layer_output[4616] + last_layer_output[4617] + last_layer_output[4618] + last_layer_output[4619] + last_layer_output[4620] + last_layer_output[4621] + last_layer_output[4622] + last_layer_output[4623] + last_layer_output[4624] + last_layer_output[4625] + last_layer_output[4626] + last_layer_output[4627] + last_layer_output[4628] + last_layer_output[4629] + last_layer_output[4630] + last_layer_output[4631] + last_layer_output[4632] + last_layer_output[4633] + last_layer_output[4634] + last_layer_output[4635] + last_layer_output[4636] + last_layer_output[4637] + last_layer_output[4638] + last_layer_output[4639] + last_layer_output[4640] + last_layer_output[4641] + last_layer_output[4642] + last_layer_output[4643] + last_layer_output[4644] + last_layer_output[4645] + last_layer_output[4646] + last_layer_output[4647] + last_layer_output[4648] + last_layer_output[4649] + last_layer_output[4650] + last_layer_output[4651] + last_layer_output[4652] + last_layer_output[4653] + last_layer_output[4654] + last_layer_output[4655] + last_layer_output[4656] + last_layer_output[4657] + last_layer_output[4658] + last_layer_output[4659] + last_layer_output[4660] + last_layer_output[4661] + last_layer_output[4662] + last_layer_output[4663] + last_layer_output[4664] + last_layer_output[4665] + last_layer_output[4666] + last_layer_output[4667] + last_layer_output[4668] + last_layer_output[4669] + last_layer_output[4670] + last_layer_output[4671] + last_layer_output[4672] + last_layer_output[4673] + last_layer_output[4674] + last_layer_output[4675] + last_layer_output[4676] + last_layer_output[4677] + last_layer_output[4678] + last_layer_output[4679] + last_layer_output[4680] + last_layer_output[4681] + last_layer_output[4682] + last_layer_output[4683] + last_layer_output[4684] + last_layer_output[4685] + last_layer_output[4686] + last_layer_output[4687] + last_layer_output[4688] + last_layer_output[4689] + last_layer_output[4690] + last_layer_output[4691] + last_layer_output[4692] + last_layer_output[4693] + last_layer_output[4694] + last_layer_output[4695] + last_layer_output[4696] + last_layer_output[4697] + last_layer_output[4698] + last_layer_output[4699] + last_layer_output[4700] + last_layer_output[4701] + last_layer_output[4702] + last_layer_output[4703] + last_layer_output[4704] + last_layer_output[4705] + last_layer_output[4706] + last_layer_output[4707] + last_layer_output[4708] + last_layer_output[4709] + last_layer_output[4710] + last_layer_output[4711] + last_layer_output[4712] + last_layer_output[4713] + last_layer_output[4714] + last_layer_output[4715] + last_layer_output[4716] + last_layer_output[4717] + last_layer_output[4718] + last_layer_output[4719] + last_layer_output[4720] + last_layer_output[4721] + last_layer_output[4722] + last_layer_output[4723] + last_layer_output[4724] + last_layer_output[4725] + last_layer_output[4726] + last_layer_output[4727] + last_layer_output[4728] + last_layer_output[4729] + last_layer_output[4730] + last_layer_output[4731] + last_layer_output[4732] + last_layer_output[4733] + last_layer_output[4734] + last_layer_output[4735] + last_layer_output[4736] + last_layer_output[4737] + last_layer_output[4738] + last_layer_output[4739] + last_layer_output[4740] + last_layer_output[4741] + last_layer_output[4742] + last_layer_output[4743] + last_layer_output[4744] + last_layer_output[4745] + last_layer_output[4746] + last_layer_output[4747] + last_layer_output[4748] + last_layer_output[4749] + last_layer_output[4750] + last_layer_output[4751] + last_layer_output[4752] + last_layer_output[4753] + last_layer_output[4754] + last_layer_output[4755] + last_layer_output[4756] + last_layer_output[4757] + last_layer_output[4758] + last_layer_output[4759] + last_layer_output[4760] + last_layer_output[4761] + last_layer_output[4762] + last_layer_output[4763] + last_layer_output[4764] + last_layer_output[4765] + last_layer_output[4766] + last_layer_output[4767] + last_layer_output[4768] + last_layer_output[4769] + last_layer_output[4770] + last_layer_output[4771] + last_layer_output[4772] + last_layer_output[4773] + last_layer_output[4774] + last_layer_output[4775] + last_layer_output[4776] + last_layer_output[4777] + last_layer_output[4778] + last_layer_output[4779] + last_layer_output[4780] + last_layer_output[4781] + last_layer_output[4782] + last_layer_output[4783] + last_layer_output[4784] + last_layer_output[4785] + last_layer_output[4786] + last_layer_output[4787] + last_layer_output[4788] + last_layer_output[4789] + last_layer_output[4790] + last_layer_output[4791] + last_layer_output[4792] + last_layer_output[4793] + last_layer_output[4794] + last_layer_output[4795] + last_layer_output[4796] + last_layer_output[4797] + last_layer_output[4798] + last_layer_output[4799];
      assign result[6] = last_layer_output[4800] + last_layer_output[4801] + last_layer_output[4802] + last_layer_output[4803] + last_layer_output[4804] + last_layer_output[4805] + last_layer_output[4806] + last_layer_output[4807] + last_layer_output[4808] + last_layer_output[4809] + last_layer_output[4810] + last_layer_output[4811] + last_layer_output[4812] + last_layer_output[4813] + last_layer_output[4814] + last_layer_output[4815] + last_layer_output[4816] + last_layer_output[4817] + last_layer_output[4818] + last_layer_output[4819] + last_layer_output[4820] + last_layer_output[4821] + last_layer_output[4822] + last_layer_output[4823] + last_layer_output[4824] + last_layer_output[4825] + last_layer_output[4826] + last_layer_output[4827] + last_layer_output[4828] + last_layer_output[4829] + last_layer_output[4830] + last_layer_output[4831] + last_layer_output[4832] + last_layer_output[4833] + last_layer_output[4834] + last_layer_output[4835] + last_layer_output[4836] + last_layer_output[4837] + last_layer_output[4838] + last_layer_output[4839] + last_layer_output[4840] + last_layer_output[4841] + last_layer_output[4842] + last_layer_output[4843] + last_layer_output[4844] + last_layer_output[4845] + last_layer_output[4846] + last_layer_output[4847] + last_layer_output[4848] + last_layer_output[4849] + last_layer_output[4850] + last_layer_output[4851] + last_layer_output[4852] + last_layer_output[4853] + last_layer_output[4854] + last_layer_output[4855] + last_layer_output[4856] + last_layer_output[4857] + last_layer_output[4858] + last_layer_output[4859] + last_layer_output[4860] + last_layer_output[4861] + last_layer_output[4862] + last_layer_output[4863] + last_layer_output[4864] + last_layer_output[4865] + last_layer_output[4866] + last_layer_output[4867] + last_layer_output[4868] + last_layer_output[4869] + last_layer_output[4870] + last_layer_output[4871] + last_layer_output[4872] + last_layer_output[4873] + last_layer_output[4874] + last_layer_output[4875] + last_layer_output[4876] + last_layer_output[4877] + last_layer_output[4878] + last_layer_output[4879] + last_layer_output[4880] + last_layer_output[4881] + last_layer_output[4882] + last_layer_output[4883] + last_layer_output[4884] + last_layer_output[4885] + last_layer_output[4886] + last_layer_output[4887] + last_layer_output[4888] + last_layer_output[4889] + last_layer_output[4890] + last_layer_output[4891] + last_layer_output[4892] + last_layer_output[4893] + last_layer_output[4894] + last_layer_output[4895] + last_layer_output[4896] + last_layer_output[4897] + last_layer_output[4898] + last_layer_output[4899] + last_layer_output[4900] + last_layer_output[4901] + last_layer_output[4902] + last_layer_output[4903] + last_layer_output[4904] + last_layer_output[4905] + last_layer_output[4906] + last_layer_output[4907] + last_layer_output[4908] + last_layer_output[4909] + last_layer_output[4910] + last_layer_output[4911] + last_layer_output[4912] + last_layer_output[4913] + last_layer_output[4914] + last_layer_output[4915] + last_layer_output[4916] + last_layer_output[4917] + last_layer_output[4918] + last_layer_output[4919] + last_layer_output[4920] + last_layer_output[4921] + last_layer_output[4922] + last_layer_output[4923] + last_layer_output[4924] + last_layer_output[4925] + last_layer_output[4926] + last_layer_output[4927] + last_layer_output[4928] + last_layer_output[4929] + last_layer_output[4930] + last_layer_output[4931] + last_layer_output[4932] + last_layer_output[4933] + last_layer_output[4934] + last_layer_output[4935] + last_layer_output[4936] + last_layer_output[4937] + last_layer_output[4938] + last_layer_output[4939] + last_layer_output[4940] + last_layer_output[4941] + last_layer_output[4942] + last_layer_output[4943] + last_layer_output[4944] + last_layer_output[4945] + last_layer_output[4946] + last_layer_output[4947] + last_layer_output[4948] + last_layer_output[4949] + last_layer_output[4950] + last_layer_output[4951] + last_layer_output[4952] + last_layer_output[4953] + last_layer_output[4954] + last_layer_output[4955] + last_layer_output[4956] + last_layer_output[4957] + last_layer_output[4958] + last_layer_output[4959] + last_layer_output[4960] + last_layer_output[4961] + last_layer_output[4962] + last_layer_output[4963] + last_layer_output[4964] + last_layer_output[4965] + last_layer_output[4966] + last_layer_output[4967] + last_layer_output[4968] + last_layer_output[4969] + last_layer_output[4970] + last_layer_output[4971] + last_layer_output[4972] + last_layer_output[4973] + last_layer_output[4974] + last_layer_output[4975] + last_layer_output[4976] + last_layer_output[4977] + last_layer_output[4978] + last_layer_output[4979] + last_layer_output[4980] + last_layer_output[4981] + last_layer_output[4982] + last_layer_output[4983] + last_layer_output[4984] + last_layer_output[4985] + last_layer_output[4986] + last_layer_output[4987] + last_layer_output[4988] + last_layer_output[4989] + last_layer_output[4990] + last_layer_output[4991] + last_layer_output[4992] + last_layer_output[4993] + last_layer_output[4994] + last_layer_output[4995] + last_layer_output[4996] + last_layer_output[4997] + last_layer_output[4998] + last_layer_output[4999] + last_layer_output[5000] + last_layer_output[5001] + last_layer_output[5002] + last_layer_output[5003] + last_layer_output[5004] + last_layer_output[5005] + last_layer_output[5006] + last_layer_output[5007] + last_layer_output[5008] + last_layer_output[5009] + last_layer_output[5010] + last_layer_output[5011] + last_layer_output[5012] + last_layer_output[5013] + last_layer_output[5014] + last_layer_output[5015] + last_layer_output[5016] + last_layer_output[5017] + last_layer_output[5018] + last_layer_output[5019] + last_layer_output[5020] + last_layer_output[5021] + last_layer_output[5022] + last_layer_output[5023] + last_layer_output[5024] + last_layer_output[5025] + last_layer_output[5026] + last_layer_output[5027] + last_layer_output[5028] + last_layer_output[5029] + last_layer_output[5030] + last_layer_output[5031] + last_layer_output[5032] + last_layer_output[5033] + last_layer_output[5034] + last_layer_output[5035] + last_layer_output[5036] + last_layer_output[5037] + last_layer_output[5038] + last_layer_output[5039] + last_layer_output[5040] + last_layer_output[5041] + last_layer_output[5042] + last_layer_output[5043] + last_layer_output[5044] + last_layer_output[5045] + last_layer_output[5046] + last_layer_output[5047] + last_layer_output[5048] + last_layer_output[5049] + last_layer_output[5050] + last_layer_output[5051] + last_layer_output[5052] + last_layer_output[5053] + last_layer_output[5054] + last_layer_output[5055] + last_layer_output[5056] + last_layer_output[5057] + last_layer_output[5058] + last_layer_output[5059] + last_layer_output[5060] + last_layer_output[5061] + last_layer_output[5062] + last_layer_output[5063] + last_layer_output[5064] + last_layer_output[5065] + last_layer_output[5066] + last_layer_output[5067] + last_layer_output[5068] + last_layer_output[5069] + last_layer_output[5070] + last_layer_output[5071] + last_layer_output[5072] + last_layer_output[5073] + last_layer_output[5074] + last_layer_output[5075] + last_layer_output[5076] + last_layer_output[5077] + last_layer_output[5078] + last_layer_output[5079] + last_layer_output[5080] + last_layer_output[5081] + last_layer_output[5082] + last_layer_output[5083] + last_layer_output[5084] + last_layer_output[5085] + last_layer_output[5086] + last_layer_output[5087] + last_layer_output[5088] + last_layer_output[5089] + last_layer_output[5090] + last_layer_output[5091] + last_layer_output[5092] + last_layer_output[5093] + last_layer_output[5094] + last_layer_output[5095] + last_layer_output[5096] + last_layer_output[5097] + last_layer_output[5098] + last_layer_output[5099] + last_layer_output[5100] + last_layer_output[5101] + last_layer_output[5102] + last_layer_output[5103] + last_layer_output[5104] + last_layer_output[5105] + last_layer_output[5106] + last_layer_output[5107] + last_layer_output[5108] + last_layer_output[5109] + last_layer_output[5110] + last_layer_output[5111] + last_layer_output[5112] + last_layer_output[5113] + last_layer_output[5114] + last_layer_output[5115] + last_layer_output[5116] + last_layer_output[5117] + last_layer_output[5118] + last_layer_output[5119] + last_layer_output[5120] + last_layer_output[5121] + last_layer_output[5122] + last_layer_output[5123] + last_layer_output[5124] + last_layer_output[5125] + last_layer_output[5126] + last_layer_output[5127] + last_layer_output[5128] + last_layer_output[5129] + last_layer_output[5130] + last_layer_output[5131] + last_layer_output[5132] + last_layer_output[5133] + last_layer_output[5134] + last_layer_output[5135] + last_layer_output[5136] + last_layer_output[5137] + last_layer_output[5138] + last_layer_output[5139] + last_layer_output[5140] + last_layer_output[5141] + last_layer_output[5142] + last_layer_output[5143] + last_layer_output[5144] + last_layer_output[5145] + last_layer_output[5146] + last_layer_output[5147] + last_layer_output[5148] + last_layer_output[5149] + last_layer_output[5150] + last_layer_output[5151] + last_layer_output[5152] + last_layer_output[5153] + last_layer_output[5154] + last_layer_output[5155] + last_layer_output[5156] + last_layer_output[5157] + last_layer_output[5158] + last_layer_output[5159] + last_layer_output[5160] + last_layer_output[5161] + last_layer_output[5162] + last_layer_output[5163] + last_layer_output[5164] + last_layer_output[5165] + last_layer_output[5166] + last_layer_output[5167] + last_layer_output[5168] + last_layer_output[5169] + last_layer_output[5170] + last_layer_output[5171] + last_layer_output[5172] + last_layer_output[5173] + last_layer_output[5174] + last_layer_output[5175] + last_layer_output[5176] + last_layer_output[5177] + last_layer_output[5178] + last_layer_output[5179] + last_layer_output[5180] + last_layer_output[5181] + last_layer_output[5182] + last_layer_output[5183] + last_layer_output[5184] + last_layer_output[5185] + last_layer_output[5186] + last_layer_output[5187] + last_layer_output[5188] + last_layer_output[5189] + last_layer_output[5190] + last_layer_output[5191] + last_layer_output[5192] + last_layer_output[5193] + last_layer_output[5194] + last_layer_output[5195] + last_layer_output[5196] + last_layer_output[5197] + last_layer_output[5198] + last_layer_output[5199] + last_layer_output[5200] + last_layer_output[5201] + last_layer_output[5202] + last_layer_output[5203] + last_layer_output[5204] + last_layer_output[5205] + last_layer_output[5206] + last_layer_output[5207] + last_layer_output[5208] + last_layer_output[5209] + last_layer_output[5210] + last_layer_output[5211] + last_layer_output[5212] + last_layer_output[5213] + last_layer_output[5214] + last_layer_output[5215] + last_layer_output[5216] + last_layer_output[5217] + last_layer_output[5218] + last_layer_output[5219] + last_layer_output[5220] + last_layer_output[5221] + last_layer_output[5222] + last_layer_output[5223] + last_layer_output[5224] + last_layer_output[5225] + last_layer_output[5226] + last_layer_output[5227] + last_layer_output[5228] + last_layer_output[5229] + last_layer_output[5230] + last_layer_output[5231] + last_layer_output[5232] + last_layer_output[5233] + last_layer_output[5234] + last_layer_output[5235] + last_layer_output[5236] + last_layer_output[5237] + last_layer_output[5238] + last_layer_output[5239] + last_layer_output[5240] + last_layer_output[5241] + last_layer_output[5242] + last_layer_output[5243] + last_layer_output[5244] + last_layer_output[5245] + last_layer_output[5246] + last_layer_output[5247] + last_layer_output[5248] + last_layer_output[5249] + last_layer_output[5250] + last_layer_output[5251] + last_layer_output[5252] + last_layer_output[5253] + last_layer_output[5254] + last_layer_output[5255] + last_layer_output[5256] + last_layer_output[5257] + last_layer_output[5258] + last_layer_output[5259] + last_layer_output[5260] + last_layer_output[5261] + last_layer_output[5262] + last_layer_output[5263] + last_layer_output[5264] + last_layer_output[5265] + last_layer_output[5266] + last_layer_output[5267] + last_layer_output[5268] + last_layer_output[5269] + last_layer_output[5270] + last_layer_output[5271] + last_layer_output[5272] + last_layer_output[5273] + last_layer_output[5274] + last_layer_output[5275] + last_layer_output[5276] + last_layer_output[5277] + last_layer_output[5278] + last_layer_output[5279] + last_layer_output[5280] + last_layer_output[5281] + last_layer_output[5282] + last_layer_output[5283] + last_layer_output[5284] + last_layer_output[5285] + last_layer_output[5286] + last_layer_output[5287] + last_layer_output[5288] + last_layer_output[5289] + last_layer_output[5290] + last_layer_output[5291] + last_layer_output[5292] + last_layer_output[5293] + last_layer_output[5294] + last_layer_output[5295] + last_layer_output[5296] + last_layer_output[5297] + last_layer_output[5298] + last_layer_output[5299] + last_layer_output[5300] + last_layer_output[5301] + last_layer_output[5302] + last_layer_output[5303] + last_layer_output[5304] + last_layer_output[5305] + last_layer_output[5306] + last_layer_output[5307] + last_layer_output[5308] + last_layer_output[5309] + last_layer_output[5310] + last_layer_output[5311] + last_layer_output[5312] + last_layer_output[5313] + last_layer_output[5314] + last_layer_output[5315] + last_layer_output[5316] + last_layer_output[5317] + last_layer_output[5318] + last_layer_output[5319] + last_layer_output[5320] + last_layer_output[5321] + last_layer_output[5322] + last_layer_output[5323] + last_layer_output[5324] + last_layer_output[5325] + last_layer_output[5326] + last_layer_output[5327] + last_layer_output[5328] + last_layer_output[5329] + last_layer_output[5330] + last_layer_output[5331] + last_layer_output[5332] + last_layer_output[5333] + last_layer_output[5334] + last_layer_output[5335] + last_layer_output[5336] + last_layer_output[5337] + last_layer_output[5338] + last_layer_output[5339] + last_layer_output[5340] + last_layer_output[5341] + last_layer_output[5342] + last_layer_output[5343] + last_layer_output[5344] + last_layer_output[5345] + last_layer_output[5346] + last_layer_output[5347] + last_layer_output[5348] + last_layer_output[5349] + last_layer_output[5350] + last_layer_output[5351] + last_layer_output[5352] + last_layer_output[5353] + last_layer_output[5354] + last_layer_output[5355] + last_layer_output[5356] + last_layer_output[5357] + last_layer_output[5358] + last_layer_output[5359] + last_layer_output[5360] + last_layer_output[5361] + last_layer_output[5362] + last_layer_output[5363] + last_layer_output[5364] + last_layer_output[5365] + last_layer_output[5366] + last_layer_output[5367] + last_layer_output[5368] + last_layer_output[5369] + last_layer_output[5370] + last_layer_output[5371] + last_layer_output[5372] + last_layer_output[5373] + last_layer_output[5374] + last_layer_output[5375] + last_layer_output[5376] + last_layer_output[5377] + last_layer_output[5378] + last_layer_output[5379] + last_layer_output[5380] + last_layer_output[5381] + last_layer_output[5382] + last_layer_output[5383] + last_layer_output[5384] + last_layer_output[5385] + last_layer_output[5386] + last_layer_output[5387] + last_layer_output[5388] + last_layer_output[5389] + last_layer_output[5390] + last_layer_output[5391] + last_layer_output[5392] + last_layer_output[5393] + last_layer_output[5394] + last_layer_output[5395] + last_layer_output[5396] + last_layer_output[5397] + last_layer_output[5398] + last_layer_output[5399] + last_layer_output[5400] + last_layer_output[5401] + last_layer_output[5402] + last_layer_output[5403] + last_layer_output[5404] + last_layer_output[5405] + last_layer_output[5406] + last_layer_output[5407] + last_layer_output[5408] + last_layer_output[5409] + last_layer_output[5410] + last_layer_output[5411] + last_layer_output[5412] + last_layer_output[5413] + last_layer_output[5414] + last_layer_output[5415] + last_layer_output[5416] + last_layer_output[5417] + last_layer_output[5418] + last_layer_output[5419] + last_layer_output[5420] + last_layer_output[5421] + last_layer_output[5422] + last_layer_output[5423] + last_layer_output[5424] + last_layer_output[5425] + last_layer_output[5426] + last_layer_output[5427] + last_layer_output[5428] + last_layer_output[5429] + last_layer_output[5430] + last_layer_output[5431] + last_layer_output[5432] + last_layer_output[5433] + last_layer_output[5434] + last_layer_output[5435] + last_layer_output[5436] + last_layer_output[5437] + last_layer_output[5438] + last_layer_output[5439] + last_layer_output[5440] + last_layer_output[5441] + last_layer_output[5442] + last_layer_output[5443] + last_layer_output[5444] + last_layer_output[5445] + last_layer_output[5446] + last_layer_output[5447] + last_layer_output[5448] + last_layer_output[5449] + last_layer_output[5450] + last_layer_output[5451] + last_layer_output[5452] + last_layer_output[5453] + last_layer_output[5454] + last_layer_output[5455] + last_layer_output[5456] + last_layer_output[5457] + last_layer_output[5458] + last_layer_output[5459] + last_layer_output[5460] + last_layer_output[5461] + last_layer_output[5462] + last_layer_output[5463] + last_layer_output[5464] + last_layer_output[5465] + last_layer_output[5466] + last_layer_output[5467] + last_layer_output[5468] + last_layer_output[5469] + last_layer_output[5470] + last_layer_output[5471] + last_layer_output[5472] + last_layer_output[5473] + last_layer_output[5474] + last_layer_output[5475] + last_layer_output[5476] + last_layer_output[5477] + last_layer_output[5478] + last_layer_output[5479] + last_layer_output[5480] + last_layer_output[5481] + last_layer_output[5482] + last_layer_output[5483] + last_layer_output[5484] + last_layer_output[5485] + last_layer_output[5486] + last_layer_output[5487] + last_layer_output[5488] + last_layer_output[5489] + last_layer_output[5490] + last_layer_output[5491] + last_layer_output[5492] + last_layer_output[5493] + last_layer_output[5494] + last_layer_output[5495] + last_layer_output[5496] + last_layer_output[5497] + last_layer_output[5498] + last_layer_output[5499] + last_layer_output[5500] + last_layer_output[5501] + last_layer_output[5502] + last_layer_output[5503] + last_layer_output[5504] + last_layer_output[5505] + last_layer_output[5506] + last_layer_output[5507] + last_layer_output[5508] + last_layer_output[5509] + last_layer_output[5510] + last_layer_output[5511] + last_layer_output[5512] + last_layer_output[5513] + last_layer_output[5514] + last_layer_output[5515] + last_layer_output[5516] + last_layer_output[5517] + last_layer_output[5518] + last_layer_output[5519] + last_layer_output[5520] + last_layer_output[5521] + last_layer_output[5522] + last_layer_output[5523] + last_layer_output[5524] + last_layer_output[5525] + last_layer_output[5526] + last_layer_output[5527] + last_layer_output[5528] + last_layer_output[5529] + last_layer_output[5530] + last_layer_output[5531] + last_layer_output[5532] + last_layer_output[5533] + last_layer_output[5534] + last_layer_output[5535] + last_layer_output[5536] + last_layer_output[5537] + last_layer_output[5538] + last_layer_output[5539] + last_layer_output[5540] + last_layer_output[5541] + last_layer_output[5542] + last_layer_output[5543] + last_layer_output[5544] + last_layer_output[5545] + last_layer_output[5546] + last_layer_output[5547] + last_layer_output[5548] + last_layer_output[5549] + last_layer_output[5550] + last_layer_output[5551] + last_layer_output[5552] + last_layer_output[5553] + last_layer_output[5554] + last_layer_output[5555] + last_layer_output[5556] + last_layer_output[5557] + last_layer_output[5558] + last_layer_output[5559] + last_layer_output[5560] + last_layer_output[5561] + last_layer_output[5562] + last_layer_output[5563] + last_layer_output[5564] + last_layer_output[5565] + last_layer_output[5566] + last_layer_output[5567] + last_layer_output[5568] + last_layer_output[5569] + last_layer_output[5570] + last_layer_output[5571] + last_layer_output[5572] + last_layer_output[5573] + last_layer_output[5574] + last_layer_output[5575] + last_layer_output[5576] + last_layer_output[5577] + last_layer_output[5578] + last_layer_output[5579] + last_layer_output[5580] + last_layer_output[5581] + last_layer_output[5582] + last_layer_output[5583] + last_layer_output[5584] + last_layer_output[5585] + last_layer_output[5586] + last_layer_output[5587] + last_layer_output[5588] + last_layer_output[5589] + last_layer_output[5590] + last_layer_output[5591] + last_layer_output[5592] + last_layer_output[5593] + last_layer_output[5594] + last_layer_output[5595] + last_layer_output[5596] + last_layer_output[5597] + last_layer_output[5598] + last_layer_output[5599];
      assign result[7] = last_layer_output[5600] + last_layer_output[5601] + last_layer_output[5602] + last_layer_output[5603] + last_layer_output[5604] + last_layer_output[5605] + last_layer_output[5606] + last_layer_output[5607] + last_layer_output[5608] + last_layer_output[5609] + last_layer_output[5610] + last_layer_output[5611] + last_layer_output[5612] + last_layer_output[5613] + last_layer_output[5614] + last_layer_output[5615] + last_layer_output[5616] + last_layer_output[5617] + last_layer_output[5618] + last_layer_output[5619] + last_layer_output[5620] + last_layer_output[5621] + last_layer_output[5622] + last_layer_output[5623] + last_layer_output[5624] + last_layer_output[5625] + last_layer_output[5626] + last_layer_output[5627] + last_layer_output[5628] + last_layer_output[5629] + last_layer_output[5630] + last_layer_output[5631] + last_layer_output[5632] + last_layer_output[5633] + last_layer_output[5634] + last_layer_output[5635] + last_layer_output[5636] + last_layer_output[5637] + last_layer_output[5638] + last_layer_output[5639] + last_layer_output[5640] + last_layer_output[5641] + last_layer_output[5642] + last_layer_output[5643] + last_layer_output[5644] + last_layer_output[5645] + last_layer_output[5646] + last_layer_output[5647] + last_layer_output[5648] + last_layer_output[5649] + last_layer_output[5650] + last_layer_output[5651] + last_layer_output[5652] + last_layer_output[5653] + last_layer_output[5654] + last_layer_output[5655] + last_layer_output[5656] + last_layer_output[5657] + last_layer_output[5658] + last_layer_output[5659] + last_layer_output[5660] + last_layer_output[5661] + last_layer_output[5662] + last_layer_output[5663] + last_layer_output[5664] + last_layer_output[5665] + last_layer_output[5666] + last_layer_output[5667] + last_layer_output[5668] + last_layer_output[5669] + last_layer_output[5670] + last_layer_output[5671] + last_layer_output[5672] + last_layer_output[5673] + last_layer_output[5674] + last_layer_output[5675] + last_layer_output[5676] + last_layer_output[5677] + last_layer_output[5678] + last_layer_output[5679] + last_layer_output[5680] + last_layer_output[5681] + last_layer_output[5682] + last_layer_output[5683] + last_layer_output[5684] + last_layer_output[5685] + last_layer_output[5686] + last_layer_output[5687] + last_layer_output[5688] + last_layer_output[5689] + last_layer_output[5690] + last_layer_output[5691] + last_layer_output[5692] + last_layer_output[5693] + last_layer_output[5694] + last_layer_output[5695] + last_layer_output[5696] + last_layer_output[5697] + last_layer_output[5698] + last_layer_output[5699] + last_layer_output[5700] + last_layer_output[5701] + last_layer_output[5702] + last_layer_output[5703] + last_layer_output[5704] + last_layer_output[5705] + last_layer_output[5706] + last_layer_output[5707] + last_layer_output[5708] + last_layer_output[5709] + last_layer_output[5710] + last_layer_output[5711] + last_layer_output[5712] + last_layer_output[5713] + last_layer_output[5714] + last_layer_output[5715] + last_layer_output[5716] + last_layer_output[5717] + last_layer_output[5718] + last_layer_output[5719] + last_layer_output[5720] + last_layer_output[5721] + last_layer_output[5722] + last_layer_output[5723] + last_layer_output[5724] + last_layer_output[5725] + last_layer_output[5726] + last_layer_output[5727] + last_layer_output[5728] + last_layer_output[5729] + last_layer_output[5730] + last_layer_output[5731] + last_layer_output[5732] + last_layer_output[5733] + last_layer_output[5734] + last_layer_output[5735] + last_layer_output[5736] + last_layer_output[5737] + last_layer_output[5738] + last_layer_output[5739] + last_layer_output[5740] + last_layer_output[5741] + last_layer_output[5742] + last_layer_output[5743] + last_layer_output[5744] + last_layer_output[5745] + last_layer_output[5746] + last_layer_output[5747] + last_layer_output[5748] + last_layer_output[5749] + last_layer_output[5750] + last_layer_output[5751] + last_layer_output[5752] + last_layer_output[5753] + last_layer_output[5754] + last_layer_output[5755] + last_layer_output[5756] + last_layer_output[5757] + last_layer_output[5758] + last_layer_output[5759] + last_layer_output[5760] + last_layer_output[5761] + last_layer_output[5762] + last_layer_output[5763] + last_layer_output[5764] + last_layer_output[5765] + last_layer_output[5766] + last_layer_output[5767] + last_layer_output[5768] + last_layer_output[5769] + last_layer_output[5770] + last_layer_output[5771] + last_layer_output[5772] + last_layer_output[5773] + last_layer_output[5774] + last_layer_output[5775] + last_layer_output[5776] + last_layer_output[5777] + last_layer_output[5778] + last_layer_output[5779] + last_layer_output[5780] + last_layer_output[5781] + last_layer_output[5782] + last_layer_output[5783] + last_layer_output[5784] + last_layer_output[5785] + last_layer_output[5786] + last_layer_output[5787] + last_layer_output[5788] + last_layer_output[5789] + last_layer_output[5790] + last_layer_output[5791] + last_layer_output[5792] + last_layer_output[5793] + last_layer_output[5794] + last_layer_output[5795] + last_layer_output[5796] + last_layer_output[5797] + last_layer_output[5798] + last_layer_output[5799] + last_layer_output[5800] + last_layer_output[5801] + last_layer_output[5802] + last_layer_output[5803] + last_layer_output[5804] + last_layer_output[5805] + last_layer_output[5806] + last_layer_output[5807] + last_layer_output[5808] + last_layer_output[5809] + last_layer_output[5810] + last_layer_output[5811] + last_layer_output[5812] + last_layer_output[5813] + last_layer_output[5814] + last_layer_output[5815] + last_layer_output[5816] + last_layer_output[5817] + last_layer_output[5818] + last_layer_output[5819] + last_layer_output[5820] + last_layer_output[5821] + last_layer_output[5822] + last_layer_output[5823] + last_layer_output[5824] + last_layer_output[5825] + last_layer_output[5826] + last_layer_output[5827] + last_layer_output[5828] + last_layer_output[5829] + last_layer_output[5830] + last_layer_output[5831] + last_layer_output[5832] + last_layer_output[5833] + last_layer_output[5834] + last_layer_output[5835] + last_layer_output[5836] + last_layer_output[5837] + last_layer_output[5838] + last_layer_output[5839] + last_layer_output[5840] + last_layer_output[5841] + last_layer_output[5842] + last_layer_output[5843] + last_layer_output[5844] + last_layer_output[5845] + last_layer_output[5846] + last_layer_output[5847] + last_layer_output[5848] + last_layer_output[5849] + last_layer_output[5850] + last_layer_output[5851] + last_layer_output[5852] + last_layer_output[5853] + last_layer_output[5854] + last_layer_output[5855] + last_layer_output[5856] + last_layer_output[5857] + last_layer_output[5858] + last_layer_output[5859] + last_layer_output[5860] + last_layer_output[5861] + last_layer_output[5862] + last_layer_output[5863] + last_layer_output[5864] + last_layer_output[5865] + last_layer_output[5866] + last_layer_output[5867] + last_layer_output[5868] + last_layer_output[5869] + last_layer_output[5870] + last_layer_output[5871] + last_layer_output[5872] + last_layer_output[5873] + last_layer_output[5874] + last_layer_output[5875] + last_layer_output[5876] + last_layer_output[5877] + last_layer_output[5878] + last_layer_output[5879] + last_layer_output[5880] + last_layer_output[5881] + last_layer_output[5882] + last_layer_output[5883] + last_layer_output[5884] + last_layer_output[5885] + last_layer_output[5886] + last_layer_output[5887] + last_layer_output[5888] + last_layer_output[5889] + last_layer_output[5890] + last_layer_output[5891] + last_layer_output[5892] + last_layer_output[5893] + last_layer_output[5894] + last_layer_output[5895] + last_layer_output[5896] + last_layer_output[5897] + last_layer_output[5898] + last_layer_output[5899] + last_layer_output[5900] + last_layer_output[5901] + last_layer_output[5902] + last_layer_output[5903] + last_layer_output[5904] + last_layer_output[5905] + last_layer_output[5906] + last_layer_output[5907] + last_layer_output[5908] + last_layer_output[5909] + last_layer_output[5910] + last_layer_output[5911] + last_layer_output[5912] + last_layer_output[5913] + last_layer_output[5914] + last_layer_output[5915] + last_layer_output[5916] + last_layer_output[5917] + last_layer_output[5918] + last_layer_output[5919] + last_layer_output[5920] + last_layer_output[5921] + last_layer_output[5922] + last_layer_output[5923] + last_layer_output[5924] + last_layer_output[5925] + last_layer_output[5926] + last_layer_output[5927] + last_layer_output[5928] + last_layer_output[5929] + last_layer_output[5930] + last_layer_output[5931] + last_layer_output[5932] + last_layer_output[5933] + last_layer_output[5934] + last_layer_output[5935] + last_layer_output[5936] + last_layer_output[5937] + last_layer_output[5938] + last_layer_output[5939] + last_layer_output[5940] + last_layer_output[5941] + last_layer_output[5942] + last_layer_output[5943] + last_layer_output[5944] + last_layer_output[5945] + last_layer_output[5946] + last_layer_output[5947] + last_layer_output[5948] + last_layer_output[5949] + last_layer_output[5950] + last_layer_output[5951] + last_layer_output[5952] + last_layer_output[5953] + last_layer_output[5954] + last_layer_output[5955] + last_layer_output[5956] + last_layer_output[5957] + last_layer_output[5958] + last_layer_output[5959] + last_layer_output[5960] + last_layer_output[5961] + last_layer_output[5962] + last_layer_output[5963] + last_layer_output[5964] + last_layer_output[5965] + last_layer_output[5966] + last_layer_output[5967] + last_layer_output[5968] + last_layer_output[5969] + last_layer_output[5970] + last_layer_output[5971] + last_layer_output[5972] + last_layer_output[5973] + last_layer_output[5974] + last_layer_output[5975] + last_layer_output[5976] + last_layer_output[5977] + last_layer_output[5978] + last_layer_output[5979] + last_layer_output[5980] + last_layer_output[5981] + last_layer_output[5982] + last_layer_output[5983] + last_layer_output[5984] + last_layer_output[5985] + last_layer_output[5986] + last_layer_output[5987] + last_layer_output[5988] + last_layer_output[5989] + last_layer_output[5990] + last_layer_output[5991] + last_layer_output[5992] + last_layer_output[5993] + last_layer_output[5994] + last_layer_output[5995] + last_layer_output[5996] + last_layer_output[5997] + last_layer_output[5998] + last_layer_output[5999] + last_layer_output[6000] + last_layer_output[6001] + last_layer_output[6002] + last_layer_output[6003] + last_layer_output[6004] + last_layer_output[6005] + last_layer_output[6006] + last_layer_output[6007] + last_layer_output[6008] + last_layer_output[6009] + last_layer_output[6010] + last_layer_output[6011] + last_layer_output[6012] + last_layer_output[6013] + last_layer_output[6014] + last_layer_output[6015] + last_layer_output[6016] + last_layer_output[6017] + last_layer_output[6018] + last_layer_output[6019] + last_layer_output[6020] + last_layer_output[6021] + last_layer_output[6022] + last_layer_output[6023] + last_layer_output[6024] + last_layer_output[6025] + last_layer_output[6026] + last_layer_output[6027] + last_layer_output[6028] + last_layer_output[6029] + last_layer_output[6030] + last_layer_output[6031] + last_layer_output[6032] + last_layer_output[6033] + last_layer_output[6034] + last_layer_output[6035] + last_layer_output[6036] + last_layer_output[6037] + last_layer_output[6038] + last_layer_output[6039] + last_layer_output[6040] + last_layer_output[6041] + last_layer_output[6042] + last_layer_output[6043] + last_layer_output[6044] + last_layer_output[6045] + last_layer_output[6046] + last_layer_output[6047] + last_layer_output[6048] + last_layer_output[6049] + last_layer_output[6050] + last_layer_output[6051] + last_layer_output[6052] + last_layer_output[6053] + last_layer_output[6054] + last_layer_output[6055] + last_layer_output[6056] + last_layer_output[6057] + last_layer_output[6058] + last_layer_output[6059] + last_layer_output[6060] + last_layer_output[6061] + last_layer_output[6062] + last_layer_output[6063] + last_layer_output[6064] + last_layer_output[6065] + last_layer_output[6066] + last_layer_output[6067] + last_layer_output[6068] + last_layer_output[6069] + last_layer_output[6070] + last_layer_output[6071] + last_layer_output[6072] + last_layer_output[6073] + last_layer_output[6074] + last_layer_output[6075] + last_layer_output[6076] + last_layer_output[6077] + last_layer_output[6078] + last_layer_output[6079] + last_layer_output[6080] + last_layer_output[6081] + last_layer_output[6082] + last_layer_output[6083] + last_layer_output[6084] + last_layer_output[6085] + last_layer_output[6086] + last_layer_output[6087] + last_layer_output[6088] + last_layer_output[6089] + last_layer_output[6090] + last_layer_output[6091] + last_layer_output[6092] + last_layer_output[6093] + last_layer_output[6094] + last_layer_output[6095] + last_layer_output[6096] + last_layer_output[6097] + last_layer_output[6098] + last_layer_output[6099] + last_layer_output[6100] + last_layer_output[6101] + last_layer_output[6102] + last_layer_output[6103] + last_layer_output[6104] + last_layer_output[6105] + last_layer_output[6106] + last_layer_output[6107] + last_layer_output[6108] + last_layer_output[6109] + last_layer_output[6110] + last_layer_output[6111] + last_layer_output[6112] + last_layer_output[6113] + last_layer_output[6114] + last_layer_output[6115] + last_layer_output[6116] + last_layer_output[6117] + last_layer_output[6118] + last_layer_output[6119] + last_layer_output[6120] + last_layer_output[6121] + last_layer_output[6122] + last_layer_output[6123] + last_layer_output[6124] + last_layer_output[6125] + last_layer_output[6126] + last_layer_output[6127] + last_layer_output[6128] + last_layer_output[6129] + last_layer_output[6130] + last_layer_output[6131] + last_layer_output[6132] + last_layer_output[6133] + last_layer_output[6134] + last_layer_output[6135] + last_layer_output[6136] + last_layer_output[6137] + last_layer_output[6138] + last_layer_output[6139] + last_layer_output[6140] + last_layer_output[6141] + last_layer_output[6142] + last_layer_output[6143] + last_layer_output[6144] + last_layer_output[6145] + last_layer_output[6146] + last_layer_output[6147] + last_layer_output[6148] + last_layer_output[6149] + last_layer_output[6150] + last_layer_output[6151] + last_layer_output[6152] + last_layer_output[6153] + last_layer_output[6154] + last_layer_output[6155] + last_layer_output[6156] + last_layer_output[6157] + last_layer_output[6158] + last_layer_output[6159] + last_layer_output[6160] + last_layer_output[6161] + last_layer_output[6162] + last_layer_output[6163] + last_layer_output[6164] + last_layer_output[6165] + last_layer_output[6166] + last_layer_output[6167] + last_layer_output[6168] + last_layer_output[6169] + last_layer_output[6170] + last_layer_output[6171] + last_layer_output[6172] + last_layer_output[6173] + last_layer_output[6174] + last_layer_output[6175] + last_layer_output[6176] + last_layer_output[6177] + last_layer_output[6178] + last_layer_output[6179] + last_layer_output[6180] + last_layer_output[6181] + last_layer_output[6182] + last_layer_output[6183] + last_layer_output[6184] + last_layer_output[6185] + last_layer_output[6186] + last_layer_output[6187] + last_layer_output[6188] + last_layer_output[6189] + last_layer_output[6190] + last_layer_output[6191] + last_layer_output[6192] + last_layer_output[6193] + last_layer_output[6194] + last_layer_output[6195] + last_layer_output[6196] + last_layer_output[6197] + last_layer_output[6198] + last_layer_output[6199] + last_layer_output[6200] + last_layer_output[6201] + last_layer_output[6202] + last_layer_output[6203] + last_layer_output[6204] + last_layer_output[6205] + last_layer_output[6206] + last_layer_output[6207] + last_layer_output[6208] + last_layer_output[6209] + last_layer_output[6210] + last_layer_output[6211] + last_layer_output[6212] + last_layer_output[6213] + last_layer_output[6214] + last_layer_output[6215] + last_layer_output[6216] + last_layer_output[6217] + last_layer_output[6218] + last_layer_output[6219] + last_layer_output[6220] + last_layer_output[6221] + last_layer_output[6222] + last_layer_output[6223] + last_layer_output[6224] + last_layer_output[6225] + last_layer_output[6226] + last_layer_output[6227] + last_layer_output[6228] + last_layer_output[6229] + last_layer_output[6230] + last_layer_output[6231] + last_layer_output[6232] + last_layer_output[6233] + last_layer_output[6234] + last_layer_output[6235] + last_layer_output[6236] + last_layer_output[6237] + last_layer_output[6238] + last_layer_output[6239] + last_layer_output[6240] + last_layer_output[6241] + last_layer_output[6242] + last_layer_output[6243] + last_layer_output[6244] + last_layer_output[6245] + last_layer_output[6246] + last_layer_output[6247] + last_layer_output[6248] + last_layer_output[6249] + last_layer_output[6250] + last_layer_output[6251] + last_layer_output[6252] + last_layer_output[6253] + last_layer_output[6254] + last_layer_output[6255] + last_layer_output[6256] + last_layer_output[6257] + last_layer_output[6258] + last_layer_output[6259] + last_layer_output[6260] + last_layer_output[6261] + last_layer_output[6262] + last_layer_output[6263] + last_layer_output[6264] + last_layer_output[6265] + last_layer_output[6266] + last_layer_output[6267] + last_layer_output[6268] + last_layer_output[6269] + last_layer_output[6270] + last_layer_output[6271] + last_layer_output[6272] + last_layer_output[6273] + last_layer_output[6274] + last_layer_output[6275] + last_layer_output[6276] + last_layer_output[6277] + last_layer_output[6278] + last_layer_output[6279] + last_layer_output[6280] + last_layer_output[6281] + last_layer_output[6282] + last_layer_output[6283] + last_layer_output[6284] + last_layer_output[6285] + last_layer_output[6286] + last_layer_output[6287] + last_layer_output[6288] + last_layer_output[6289] + last_layer_output[6290] + last_layer_output[6291] + last_layer_output[6292] + last_layer_output[6293] + last_layer_output[6294] + last_layer_output[6295] + last_layer_output[6296] + last_layer_output[6297] + last_layer_output[6298] + last_layer_output[6299] + last_layer_output[6300] + last_layer_output[6301] + last_layer_output[6302] + last_layer_output[6303] + last_layer_output[6304] + last_layer_output[6305] + last_layer_output[6306] + last_layer_output[6307] + last_layer_output[6308] + last_layer_output[6309] + last_layer_output[6310] + last_layer_output[6311] + last_layer_output[6312] + last_layer_output[6313] + last_layer_output[6314] + last_layer_output[6315] + last_layer_output[6316] + last_layer_output[6317] + last_layer_output[6318] + last_layer_output[6319] + last_layer_output[6320] + last_layer_output[6321] + last_layer_output[6322] + last_layer_output[6323] + last_layer_output[6324] + last_layer_output[6325] + last_layer_output[6326] + last_layer_output[6327] + last_layer_output[6328] + last_layer_output[6329] + last_layer_output[6330] + last_layer_output[6331] + last_layer_output[6332] + last_layer_output[6333] + last_layer_output[6334] + last_layer_output[6335] + last_layer_output[6336] + last_layer_output[6337] + last_layer_output[6338] + last_layer_output[6339] + last_layer_output[6340] + last_layer_output[6341] + last_layer_output[6342] + last_layer_output[6343] + last_layer_output[6344] + last_layer_output[6345] + last_layer_output[6346] + last_layer_output[6347] + last_layer_output[6348] + last_layer_output[6349] + last_layer_output[6350] + last_layer_output[6351] + last_layer_output[6352] + last_layer_output[6353] + last_layer_output[6354] + last_layer_output[6355] + last_layer_output[6356] + last_layer_output[6357] + last_layer_output[6358] + last_layer_output[6359] + last_layer_output[6360] + last_layer_output[6361] + last_layer_output[6362] + last_layer_output[6363] + last_layer_output[6364] + last_layer_output[6365] + last_layer_output[6366] + last_layer_output[6367] + last_layer_output[6368] + last_layer_output[6369] + last_layer_output[6370] + last_layer_output[6371] + last_layer_output[6372] + last_layer_output[6373] + last_layer_output[6374] + last_layer_output[6375] + last_layer_output[6376] + last_layer_output[6377] + last_layer_output[6378] + last_layer_output[6379] + last_layer_output[6380] + last_layer_output[6381] + last_layer_output[6382] + last_layer_output[6383] + last_layer_output[6384] + last_layer_output[6385] + last_layer_output[6386] + last_layer_output[6387] + last_layer_output[6388] + last_layer_output[6389] + last_layer_output[6390] + last_layer_output[6391] + last_layer_output[6392] + last_layer_output[6393] + last_layer_output[6394] + last_layer_output[6395] + last_layer_output[6396] + last_layer_output[6397] + last_layer_output[6398] + last_layer_output[6399];
      assign result[8] = last_layer_output[6400] + last_layer_output[6401] + last_layer_output[6402] + last_layer_output[6403] + last_layer_output[6404] + last_layer_output[6405] + last_layer_output[6406] + last_layer_output[6407] + last_layer_output[6408] + last_layer_output[6409] + last_layer_output[6410] + last_layer_output[6411] + last_layer_output[6412] + last_layer_output[6413] + last_layer_output[6414] + last_layer_output[6415] + last_layer_output[6416] + last_layer_output[6417] + last_layer_output[6418] + last_layer_output[6419] + last_layer_output[6420] + last_layer_output[6421] + last_layer_output[6422] + last_layer_output[6423] + last_layer_output[6424] + last_layer_output[6425] + last_layer_output[6426] + last_layer_output[6427] + last_layer_output[6428] + last_layer_output[6429] + last_layer_output[6430] + last_layer_output[6431] + last_layer_output[6432] + last_layer_output[6433] + last_layer_output[6434] + last_layer_output[6435] + last_layer_output[6436] + last_layer_output[6437] + last_layer_output[6438] + last_layer_output[6439] + last_layer_output[6440] + last_layer_output[6441] + last_layer_output[6442] + last_layer_output[6443] + last_layer_output[6444] + last_layer_output[6445] + last_layer_output[6446] + last_layer_output[6447] + last_layer_output[6448] + last_layer_output[6449] + last_layer_output[6450] + last_layer_output[6451] + last_layer_output[6452] + last_layer_output[6453] + last_layer_output[6454] + last_layer_output[6455] + last_layer_output[6456] + last_layer_output[6457] + last_layer_output[6458] + last_layer_output[6459] + last_layer_output[6460] + last_layer_output[6461] + last_layer_output[6462] + last_layer_output[6463] + last_layer_output[6464] + last_layer_output[6465] + last_layer_output[6466] + last_layer_output[6467] + last_layer_output[6468] + last_layer_output[6469] + last_layer_output[6470] + last_layer_output[6471] + last_layer_output[6472] + last_layer_output[6473] + last_layer_output[6474] + last_layer_output[6475] + last_layer_output[6476] + last_layer_output[6477] + last_layer_output[6478] + last_layer_output[6479] + last_layer_output[6480] + last_layer_output[6481] + last_layer_output[6482] + last_layer_output[6483] + last_layer_output[6484] + last_layer_output[6485] + last_layer_output[6486] + last_layer_output[6487] + last_layer_output[6488] + last_layer_output[6489] + last_layer_output[6490] + last_layer_output[6491] + last_layer_output[6492] + last_layer_output[6493] + last_layer_output[6494] + last_layer_output[6495] + last_layer_output[6496] + last_layer_output[6497] + last_layer_output[6498] + last_layer_output[6499] + last_layer_output[6500] + last_layer_output[6501] + last_layer_output[6502] + last_layer_output[6503] + last_layer_output[6504] + last_layer_output[6505] + last_layer_output[6506] + last_layer_output[6507] + last_layer_output[6508] + last_layer_output[6509] + last_layer_output[6510] + last_layer_output[6511] + last_layer_output[6512] + last_layer_output[6513] + last_layer_output[6514] + last_layer_output[6515] + last_layer_output[6516] + last_layer_output[6517] + last_layer_output[6518] + last_layer_output[6519] + last_layer_output[6520] + last_layer_output[6521] + last_layer_output[6522] + last_layer_output[6523] + last_layer_output[6524] + last_layer_output[6525] + last_layer_output[6526] + last_layer_output[6527] + last_layer_output[6528] + last_layer_output[6529] + last_layer_output[6530] + last_layer_output[6531] + last_layer_output[6532] + last_layer_output[6533] + last_layer_output[6534] + last_layer_output[6535] + last_layer_output[6536] + last_layer_output[6537] + last_layer_output[6538] + last_layer_output[6539] + last_layer_output[6540] + last_layer_output[6541] + last_layer_output[6542] + last_layer_output[6543] + last_layer_output[6544] + last_layer_output[6545] + last_layer_output[6546] + last_layer_output[6547] + last_layer_output[6548] + last_layer_output[6549] + last_layer_output[6550] + last_layer_output[6551] + last_layer_output[6552] + last_layer_output[6553] + last_layer_output[6554] + last_layer_output[6555] + last_layer_output[6556] + last_layer_output[6557] + last_layer_output[6558] + last_layer_output[6559] + last_layer_output[6560] + last_layer_output[6561] + last_layer_output[6562] + last_layer_output[6563] + last_layer_output[6564] + last_layer_output[6565] + last_layer_output[6566] + last_layer_output[6567] + last_layer_output[6568] + last_layer_output[6569] + last_layer_output[6570] + last_layer_output[6571] + last_layer_output[6572] + last_layer_output[6573] + last_layer_output[6574] + last_layer_output[6575] + last_layer_output[6576] + last_layer_output[6577] + last_layer_output[6578] + last_layer_output[6579] + last_layer_output[6580] + last_layer_output[6581] + last_layer_output[6582] + last_layer_output[6583] + last_layer_output[6584] + last_layer_output[6585] + last_layer_output[6586] + last_layer_output[6587] + last_layer_output[6588] + last_layer_output[6589] + last_layer_output[6590] + last_layer_output[6591] + last_layer_output[6592] + last_layer_output[6593] + last_layer_output[6594] + last_layer_output[6595] + last_layer_output[6596] + last_layer_output[6597] + last_layer_output[6598] + last_layer_output[6599] + last_layer_output[6600] + last_layer_output[6601] + last_layer_output[6602] + last_layer_output[6603] + last_layer_output[6604] + last_layer_output[6605] + last_layer_output[6606] + last_layer_output[6607] + last_layer_output[6608] + last_layer_output[6609] + last_layer_output[6610] + last_layer_output[6611] + last_layer_output[6612] + last_layer_output[6613] + last_layer_output[6614] + last_layer_output[6615] + last_layer_output[6616] + last_layer_output[6617] + last_layer_output[6618] + last_layer_output[6619] + last_layer_output[6620] + last_layer_output[6621] + last_layer_output[6622] + last_layer_output[6623] + last_layer_output[6624] + last_layer_output[6625] + last_layer_output[6626] + last_layer_output[6627] + last_layer_output[6628] + last_layer_output[6629] + last_layer_output[6630] + last_layer_output[6631] + last_layer_output[6632] + last_layer_output[6633] + last_layer_output[6634] + last_layer_output[6635] + last_layer_output[6636] + last_layer_output[6637] + last_layer_output[6638] + last_layer_output[6639] + last_layer_output[6640] + last_layer_output[6641] + last_layer_output[6642] + last_layer_output[6643] + last_layer_output[6644] + last_layer_output[6645] + last_layer_output[6646] + last_layer_output[6647] + last_layer_output[6648] + last_layer_output[6649] + last_layer_output[6650] + last_layer_output[6651] + last_layer_output[6652] + last_layer_output[6653] + last_layer_output[6654] + last_layer_output[6655] + last_layer_output[6656] + last_layer_output[6657] + last_layer_output[6658] + last_layer_output[6659] + last_layer_output[6660] + last_layer_output[6661] + last_layer_output[6662] + last_layer_output[6663] + last_layer_output[6664] + last_layer_output[6665] + last_layer_output[6666] + last_layer_output[6667] + last_layer_output[6668] + last_layer_output[6669] + last_layer_output[6670] + last_layer_output[6671] + last_layer_output[6672] + last_layer_output[6673] + last_layer_output[6674] + last_layer_output[6675] + last_layer_output[6676] + last_layer_output[6677] + last_layer_output[6678] + last_layer_output[6679] + last_layer_output[6680] + last_layer_output[6681] + last_layer_output[6682] + last_layer_output[6683] + last_layer_output[6684] + last_layer_output[6685] + last_layer_output[6686] + last_layer_output[6687] + last_layer_output[6688] + last_layer_output[6689] + last_layer_output[6690] + last_layer_output[6691] + last_layer_output[6692] + last_layer_output[6693] + last_layer_output[6694] + last_layer_output[6695] + last_layer_output[6696] + last_layer_output[6697] + last_layer_output[6698] + last_layer_output[6699] + last_layer_output[6700] + last_layer_output[6701] + last_layer_output[6702] + last_layer_output[6703] + last_layer_output[6704] + last_layer_output[6705] + last_layer_output[6706] + last_layer_output[6707] + last_layer_output[6708] + last_layer_output[6709] + last_layer_output[6710] + last_layer_output[6711] + last_layer_output[6712] + last_layer_output[6713] + last_layer_output[6714] + last_layer_output[6715] + last_layer_output[6716] + last_layer_output[6717] + last_layer_output[6718] + last_layer_output[6719] + last_layer_output[6720] + last_layer_output[6721] + last_layer_output[6722] + last_layer_output[6723] + last_layer_output[6724] + last_layer_output[6725] + last_layer_output[6726] + last_layer_output[6727] + last_layer_output[6728] + last_layer_output[6729] + last_layer_output[6730] + last_layer_output[6731] + last_layer_output[6732] + last_layer_output[6733] + last_layer_output[6734] + last_layer_output[6735] + last_layer_output[6736] + last_layer_output[6737] + last_layer_output[6738] + last_layer_output[6739] + last_layer_output[6740] + last_layer_output[6741] + last_layer_output[6742] + last_layer_output[6743] + last_layer_output[6744] + last_layer_output[6745] + last_layer_output[6746] + last_layer_output[6747] + last_layer_output[6748] + last_layer_output[6749] + last_layer_output[6750] + last_layer_output[6751] + last_layer_output[6752] + last_layer_output[6753] + last_layer_output[6754] + last_layer_output[6755] + last_layer_output[6756] + last_layer_output[6757] + last_layer_output[6758] + last_layer_output[6759] + last_layer_output[6760] + last_layer_output[6761] + last_layer_output[6762] + last_layer_output[6763] + last_layer_output[6764] + last_layer_output[6765] + last_layer_output[6766] + last_layer_output[6767] + last_layer_output[6768] + last_layer_output[6769] + last_layer_output[6770] + last_layer_output[6771] + last_layer_output[6772] + last_layer_output[6773] + last_layer_output[6774] + last_layer_output[6775] + last_layer_output[6776] + last_layer_output[6777] + last_layer_output[6778] + last_layer_output[6779] + last_layer_output[6780] + last_layer_output[6781] + last_layer_output[6782] + last_layer_output[6783] + last_layer_output[6784] + last_layer_output[6785] + last_layer_output[6786] + last_layer_output[6787] + last_layer_output[6788] + last_layer_output[6789] + last_layer_output[6790] + last_layer_output[6791] + last_layer_output[6792] + last_layer_output[6793] + last_layer_output[6794] + last_layer_output[6795] + last_layer_output[6796] + last_layer_output[6797] + last_layer_output[6798] + last_layer_output[6799] + last_layer_output[6800] + last_layer_output[6801] + last_layer_output[6802] + last_layer_output[6803] + last_layer_output[6804] + last_layer_output[6805] + last_layer_output[6806] + last_layer_output[6807] + last_layer_output[6808] + last_layer_output[6809] + last_layer_output[6810] + last_layer_output[6811] + last_layer_output[6812] + last_layer_output[6813] + last_layer_output[6814] + last_layer_output[6815] + last_layer_output[6816] + last_layer_output[6817] + last_layer_output[6818] + last_layer_output[6819] + last_layer_output[6820] + last_layer_output[6821] + last_layer_output[6822] + last_layer_output[6823] + last_layer_output[6824] + last_layer_output[6825] + last_layer_output[6826] + last_layer_output[6827] + last_layer_output[6828] + last_layer_output[6829] + last_layer_output[6830] + last_layer_output[6831] + last_layer_output[6832] + last_layer_output[6833] + last_layer_output[6834] + last_layer_output[6835] + last_layer_output[6836] + last_layer_output[6837] + last_layer_output[6838] + last_layer_output[6839] + last_layer_output[6840] + last_layer_output[6841] + last_layer_output[6842] + last_layer_output[6843] + last_layer_output[6844] + last_layer_output[6845] + last_layer_output[6846] + last_layer_output[6847] + last_layer_output[6848] + last_layer_output[6849] + last_layer_output[6850] + last_layer_output[6851] + last_layer_output[6852] + last_layer_output[6853] + last_layer_output[6854] + last_layer_output[6855] + last_layer_output[6856] + last_layer_output[6857] + last_layer_output[6858] + last_layer_output[6859] + last_layer_output[6860] + last_layer_output[6861] + last_layer_output[6862] + last_layer_output[6863] + last_layer_output[6864] + last_layer_output[6865] + last_layer_output[6866] + last_layer_output[6867] + last_layer_output[6868] + last_layer_output[6869] + last_layer_output[6870] + last_layer_output[6871] + last_layer_output[6872] + last_layer_output[6873] + last_layer_output[6874] + last_layer_output[6875] + last_layer_output[6876] + last_layer_output[6877] + last_layer_output[6878] + last_layer_output[6879] + last_layer_output[6880] + last_layer_output[6881] + last_layer_output[6882] + last_layer_output[6883] + last_layer_output[6884] + last_layer_output[6885] + last_layer_output[6886] + last_layer_output[6887] + last_layer_output[6888] + last_layer_output[6889] + last_layer_output[6890] + last_layer_output[6891] + last_layer_output[6892] + last_layer_output[6893] + last_layer_output[6894] + last_layer_output[6895] + last_layer_output[6896] + last_layer_output[6897] + last_layer_output[6898] + last_layer_output[6899] + last_layer_output[6900] + last_layer_output[6901] + last_layer_output[6902] + last_layer_output[6903] + last_layer_output[6904] + last_layer_output[6905] + last_layer_output[6906] + last_layer_output[6907] + last_layer_output[6908] + last_layer_output[6909] + last_layer_output[6910] + last_layer_output[6911] + last_layer_output[6912] + last_layer_output[6913] + last_layer_output[6914] + last_layer_output[6915] + last_layer_output[6916] + last_layer_output[6917] + last_layer_output[6918] + last_layer_output[6919] + last_layer_output[6920] + last_layer_output[6921] + last_layer_output[6922] + last_layer_output[6923] + last_layer_output[6924] + last_layer_output[6925] + last_layer_output[6926] + last_layer_output[6927] + last_layer_output[6928] + last_layer_output[6929] + last_layer_output[6930] + last_layer_output[6931] + last_layer_output[6932] + last_layer_output[6933] + last_layer_output[6934] + last_layer_output[6935] + last_layer_output[6936] + last_layer_output[6937] + last_layer_output[6938] + last_layer_output[6939] + last_layer_output[6940] + last_layer_output[6941] + last_layer_output[6942] + last_layer_output[6943] + last_layer_output[6944] + last_layer_output[6945] + last_layer_output[6946] + last_layer_output[6947] + last_layer_output[6948] + last_layer_output[6949] + last_layer_output[6950] + last_layer_output[6951] + last_layer_output[6952] + last_layer_output[6953] + last_layer_output[6954] + last_layer_output[6955] + last_layer_output[6956] + last_layer_output[6957] + last_layer_output[6958] + last_layer_output[6959] + last_layer_output[6960] + last_layer_output[6961] + last_layer_output[6962] + last_layer_output[6963] + last_layer_output[6964] + last_layer_output[6965] + last_layer_output[6966] + last_layer_output[6967] + last_layer_output[6968] + last_layer_output[6969] + last_layer_output[6970] + last_layer_output[6971] + last_layer_output[6972] + last_layer_output[6973] + last_layer_output[6974] + last_layer_output[6975] + last_layer_output[6976] + last_layer_output[6977] + last_layer_output[6978] + last_layer_output[6979] + last_layer_output[6980] + last_layer_output[6981] + last_layer_output[6982] + last_layer_output[6983] + last_layer_output[6984] + last_layer_output[6985] + last_layer_output[6986] + last_layer_output[6987] + last_layer_output[6988] + last_layer_output[6989] + last_layer_output[6990] + last_layer_output[6991] + last_layer_output[6992] + last_layer_output[6993] + last_layer_output[6994] + last_layer_output[6995] + last_layer_output[6996] + last_layer_output[6997] + last_layer_output[6998] + last_layer_output[6999] + last_layer_output[7000] + last_layer_output[7001] + last_layer_output[7002] + last_layer_output[7003] + last_layer_output[7004] + last_layer_output[7005] + last_layer_output[7006] + last_layer_output[7007] + last_layer_output[7008] + last_layer_output[7009] + last_layer_output[7010] + last_layer_output[7011] + last_layer_output[7012] + last_layer_output[7013] + last_layer_output[7014] + last_layer_output[7015] + last_layer_output[7016] + last_layer_output[7017] + last_layer_output[7018] + last_layer_output[7019] + last_layer_output[7020] + last_layer_output[7021] + last_layer_output[7022] + last_layer_output[7023] + last_layer_output[7024] + last_layer_output[7025] + last_layer_output[7026] + last_layer_output[7027] + last_layer_output[7028] + last_layer_output[7029] + last_layer_output[7030] + last_layer_output[7031] + last_layer_output[7032] + last_layer_output[7033] + last_layer_output[7034] + last_layer_output[7035] + last_layer_output[7036] + last_layer_output[7037] + last_layer_output[7038] + last_layer_output[7039] + last_layer_output[7040] + last_layer_output[7041] + last_layer_output[7042] + last_layer_output[7043] + last_layer_output[7044] + last_layer_output[7045] + last_layer_output[7046] + last_layer_output[7047] + last_layer_output[7048] + last_layer_output[7049] + last_layer_output[7050] + last_layer_output[7051] + last_layer_output[7052] + last_layer_output[7053] + last_layer_output[7054] + last_layer_output[7055] + last_layer_output[7056] + last_layer_output[7057] + last_layer_output[7058] + last_layer_output[7059] + last_layer_output[7060] + last_layer_output[7061] + last_layer_output[7062] + last_layer_output[7063] + last_layer_output[7064] + last_layer_output[7065] + last_layer_output[7066] + last_layer_output[7067] + last_layer_output[7068] + last_layer_output[7069] + last_layer_output[7070] + last_layer_output[7071] + last_layer_output[7072] + last_layer_output[7073] + last_layer_output[7074] + last_layer_output[7075] + last_layer_output[7076] + last_layer_output[7077] + last_layer_output[7078] + last_layer_output[7079] + last_layer_output[7080] + last_layer_output[7081] + last_layer_output[7082] + last_layer_output[7083] + last_layer_output[7084] + last_layer_output[7085] + last_layer_output[7086] + last_layer_output[7087] + last_layer_output[7088] + last_layer_output[7089] + last_layer_output[7090] + last_layer_output[7091] + last_layer_output[7092] + last_layer_output[7093] + last_layer_output[7094] + last_layer_output[7095] + last_layer_output[7096] + last_layer_output[7097] + last_layer_output[7098] + last_layer_output[7099] + last_layer_output[7100] + last_layer_output[7101] + last_layer_output[7102] + last_layer_output[7103] + last_layer_output[7104] + last_layer_output[7105] + last_layer_output[7106] + last_layer_output[7107] + last_layer_output[7108] + last_layer_output[7109] + last_layer_output[7110] + last_layer_output[7111] + last_layer_output[7112] + last_layer_output[7113] + last_layer_output[7114] + last_layer_output[7115] + last_layer_output[7116] + last_layer_output[7117] + last_layer_output[7118] + last_layer_output[7119] + last_layer_output[7120] + last_layer_output[7121] + last_layer_output[7122] + last_layer_output[7123] + last_layer_output[7124] + last_layer_output[7125] + last_layer_output[7126] + last_layer_output[7127] + last_layer_output[7128] + last_layer_output[7129] + last_layer_output[7130] + last_layer_output[7131] + last_layer_output[7132] + last_layer_output[7133] + last_layer_output[7134] + last_layer_output[7135] + last_layer_output[7136] + last_layer_output[7137] + last_layer_output[7138] + last_layer_output[7139] + last_layer_output[7140] + last_layer_output[7141] + last_layer_output[7142] + last_layer_output[7143] + last_layer_output[7144] + last_layer_output[7145] + last_layer_output[7146] + last_layer_output[7147] + last_layer_output[7148] + last_layer_output[7149] + last_layer_output[7150] + last_layer_output[7151] + last_layer_output[7152] + last_layer_output[7153] + last_layer_output[7154] + last_layer_output[7155] + last_layer_output[7156] + last_layer_output[7157] + last_layer_output[7158] + last_layer_output[7159] + last_layer_output[7160] + last_layer_output[7161] + last_layer_output[7162] + last_layer_output[7163] + last_layer_output[7164] + last_layer_output[7165] + last_layer_output[7166] + last_layer_output[7167] + last_layer_output[7168] + last_layer_output[7169] + last_layer_output[7170] + last_layer_output[7171] + last_layer_output[7172] + last_layer_output[7173] + last_layer_output[7174] + last_layer_output[7175] + last_layer_output[7176] + last_layer_output[7177] + last_layer_output[7178] + last_layer_output[7179] + last_layer_output[7180] + last_layer_output[7181] + last_layer_output[7182] + last_layer_output[7183] + last_layer_output[7184] + last_layer_output[7185] + last_layer_output[7186] + last_layer_output[7187] + last_layer_output[7188] + last_layer_output[7189] + last_layer_output[7190] + last_layer_output[7191] + last_layer_output[7192] + last_layer_output[7193] + last_layer_output[7194] + last_layer_output[7195] + last_layer_output[7196] + last_layer_output[7197] + last_layer_output[7198] + last_layer_output[7199];
      assign result[9] = last_layer_output[7200] + last_layer_output[7201] + last_layer_output[7202] + last_layer_output[7203] + last_layer_output[7204] + last_layer_output[7205] + last_layer_output[7206] + last_layer_output[7207] + last_layer_output[7208] + last_layer_output[7209] + last_layer_output[7210] + last_layer_output[7211] + last_layer_output[7212] + last_layer_output[7213] + last_layer_output[7214] + last_layer_output[7215] + last_layer_output[7216] + last_layer_output[7217] + last_layer_output[7218] + last_layer_output[7219] + last_layer_output[7220] + last_layer_output[7221] + last_layer_output[7222] + last_layer_output[7223] + last_layer_output[7224] + last_layer_output[7225] + last_layer_output[7226] + last_layer_output[7227] + last_layer_output[7228] + last_layer_output[7229] + last_layer_output[7230] + last_layer_output[7231] + last_layer_output[7232] + last_layer_output[7233] + last_layer_output[7234] + last_layer_output[7235] + last_layer_output[7236] + last_layer_output[7237] + last_layer_output[7238] + last_layer_output[7239] + last_layer_output[7240] + last_layer_output[7241] + last_layer_output[7242] + last_layer_output[7243] + last_layer_output[7244] + last_layer_output[7245] + last_layer_output[7246] + last_layer_output[7247] + last_layer_output[7248] + last_layer_output[7249] + last_layer_output[7250] + last_layer_output[7251] + last_layer_output[7252] + last_layer_output[7253] + last_layer_output[7254] + last_layer_output[7255] + last_layer_output[7256] + last_layer_output[7257] + last_layer_output[7258] + last_layer_output[7259] + last_layer_output[7260] + last_layer_output[7261] + last_layer_output[7262] + last_layer_output[7263] + last_layer_output[7264] + last_layer_output[7265] + last_layer_output[7266] + last_layer_output[7267] + last_layer_output[7268] + last_layer_output[7269] + last_layer_output[7270] + last_layer_output[7271] + last_layer_output[7272] + last_layer_output[7273] + last_layer_output[7274] + last_layer_output[7275] + last_layer_output[7276] + last_layer_output[7277] + last_layer_output[7278] + last_layer_output[7279] + last_layer_output[7280] + last_layer_output[7281] + last_layer_output[7282] + last_layer_output[7283] + last_layer_output[7284] + last_layer_output[7285] + last_layer_output[7286] + last_layer_output[7287] + last_layer_output[7288] + last_layer_output[7289] + last_layer_output[7290] + last_layer_output[7291] + last_layer_output[7292] + last_layer_output[7293] + last_layer_output[7294] + last_layer_output[7295] + last_layer_output[7296] + last_layer_output[7297] + last_layer_output[7298] + last_layer_output[7299] + last_layer_output[7300] + last_layer_output[7301] + last_layer_output[7302] + last_layer_output[7303] + last_layer_output[7304] + last_layer_output[7305] + last_layer_output[7306] + last_layer_output[7307] + last_layer_output[7308] + last_layer_output[7309] + last_layer_output[7310] + last_layer_output[7311] + last_layer_output[7312] + last_layer_output[7313] + last_layer_output[7314] + last_layer_output[7315] + last_layer_output[7316] + last_layer_output[7317] + last_layer_output[7318] + last_layer_output[7319] + last_layer_output[7320] + last_layer_output[7321] + last_layer_output[7322] + last_layer_output[7323] + last_layer_output[7324] + last_layer_output[7325] + last_layer_output[7326] + last_layer_output[7327] + last_layer_output[7328] + last_layer_output[7329] + last_layer_output[7330] + last_layer_output[7331] + last_layer_output[7332] + last_layer_output[7333] + last_layer_output[7334] + last_layer_output[7335] + last_layer_output[7336] + last_layer_output[7337] + last_layer_output[7338] + last_layer_output[7339] + last_layer_output[7340] + last_layer_output[7341] + last_layer_output[7342] + last_layer_output[7343] + last_layer_output[7344] + last_layer_output[7345] + last_layer_output[7346] + last_layer_output[7347] + last_layer_output[7348] + last_layer_output[7349] + last_layer_output[7350] + last_layer_output[7351] + last_layer_output[7352] + last_layer_output[7353] + last_layer_output[7354] + last_layer_output[7355] + last_layer_output[7356] + last_layer_output[7357] + last_layer_output[7358] + last_layer_output[7359] + last_layer_output[7360] + last_layer_output[7361] + last_layer_output[7362] + last_layer_output[7363] + last_layer_output[7364] + last_layer_output[7365] + last_layer_output[7366] + last_layer_output[7367] + last_layer_output[7368] + last_layer_output[7369] + last_layer_output[7370] + last_layer_output[7371] + last_layer_output[7372] + last_layer_output[7373] + last_layer_output[7374] + last_layer_output[7375] + last_layer_output[7376] + last_layer_output[7377] + last_layer_output[7378] + last_layer_output[7379] + last_layer_output[7380] + last_layer_output[7381] + last_layer_output[7382] + last_layer_output[7383] + last_layer_output[7384] + last_layer_output[7385] + last_layer_output[7386] + last_layer_output[7387] + last_layer_output[7388] + last_layer_output[7389] + last_layer_output[7390] + last_layer_output[7391] + last_layer_output[7392] + last_layer_output[7393] + last_layer_output[7394] + last_layer_output[7395] + last_layer_output[7396] + last_layer_output[7397] + last_layer_output[7398] + last_layer_output[7399] + last_layer_output[7400] + last_layer_output[7401] + last_layer_output[7402] + last_layer_output[7403] + last_layer_output[7404] + last_layer_output[7405] + last_layer_output[7406] + last_layer_output[7407] + last_layer_output[7408] + last_layer_output[7409] + last_layer_output[7410] + last_layer_output[7411] + last_layer_output[7412] + last_layer_output[7413] + last_layer_output[7414] + last_layer_output[7415] + last_layer_output[7416] + last_layer_output[7417] + last_layer_output[7418] + last_layer_output[7419] + last_layer_output[7420] + last_layer_output[7421] + last_layer_output[7422] + last_layer_output[7423] + last_layer_output[7424] + last_layer_output[7425] + last_layer_output[7426] + last_layer_output[7427] + last_layer_output[7428] + last_layer_output[7429] + last_layer_output[7430] + last_layer_output[7431] + last_layer_output[7432] + last_layer_output[7433] + last_layer_output[7434] + last_layer_output[7435] + last_layer_output[7436] + last_layer_output[7437] + last_layer_output[7438] + last_layer_output[7439] + last_layer_output[7440] + last_layer_output[7441] + last_layer_output[7442] + last_layer_output[7443] + last_layer_output[7444] + last_layer_output[7445] + last_layer_output[7446] + last_layer_output[7447] + last_layer_output[7448] + last_layer_output[7449] + last_layer_output[7450] + last_layer_output[7451] + last_layer_output[7452] + last_layer_output[7453] + last_layer_output[7454] + last_layer_output[7455] + last_layer_output[7456] + last_layer_output[7457] + last_layer_output[7458] + last_layer_output[7459] + last_layer_output[7460] + last_layer_output[7461] + last_layer_output[7462] + last_layer_output[7463] + last_layer_output[7464] + last_layer_output[7465] + last_layer_output[7466] + last_layer_output[7467] + last_layer_output[7468] + last_layer_output[7469] + last_layer_output[7470] + last_layer_output[7471] + last_layer_output[7472] + last_layer_output[7473] + last_layer_output[7474] + last_layer_output[7475] + last_layer_output[7476] + last_layer_output[7477] + last_layer_output[7478] + last_layer_output[7479] + last_layer_output[7480] + last_layer_output[7481] + last_layer_output[7482] + last_layer_output[7483] + last_layer_output[7484] + last_layer_output[7485] + last_layer_output[7486] + last_layer_output[7487] + last_layer_output[7488] + last_layer_output[7489] + last_layer_output[7490] + last_layer_output[7491] + last_layer_output[7492] + last_layer_output[7493] + last_layer_output[7494] + last_layer_output[7495] + last_layer_output[7496] + last_layer_output[7497] + last_layer_output[7498] + last_layer_output[7499] + last_layer_output[7500] + last_layer_output[7501] + last_layer_output[7502] + last_layer_output[7503] + last_layer_output[7504] + last_layer_output[7505] + last_layer_output[7506] + last_layer_output[7507] + last_layer_output[7508] + last_layer_output[7509] + last_layer_output[7510] + last_layer_output[7511] + last_layer_output[7512] + last_layer_output[7513] + last_layer_output[7514] + last_layer_output[7515] + last_layer_output[7516] + last_layer_output[7517] + last_layer_output[7518] + last_layer_output[7519] + last_layer_output[7520] + last_layer_output[7521] + last_layer_output[7522] + last_layer_output[7523] + last_layer_output[7524] + last_layer_output[7525] + last_layer_output[7526] + last_layer_output[7527] + last_layer_output[7528] + last_layer_output[7529] + last_layer_output[7530] + last_layer_output[7531] + last_layer_output[7532] + last_layer_output[7533] + last_layer_output[7534] + last_layer_output[7535] + last_layer_output[7536] + last_layer_output[7537] + last_layer_output[7538] + last_layer_output[7539] + last_layer_output[7540] + last_layer_output[7541] + last_layer_output[7542] + last_layer_output[7543] + last_layer_output[7544] + last_layer_output[7545] + last_layer_output[7546] + last_layer_output[7547] + last_layer_output[7548] + last_layer_output[7549] + last_layer_output[7550] + last_layer_output[7551] + last_layer_output[7552] + last_layer_output[7553] + last_layer_output[7554] + last_layer_output[7555] + last_layer_output[7556] + last_layer_output[7557] + last_layer_output[7558] + last_layer_output[7559] + last_layer_output[7560] + last_layer_output[7561] + last_layer_output[7562] + last_layer_output[7563] + last_layer_output[7564] + last_layer_output[7565] + last_layer_output[7566] + last_layer_output[7567] + last_layer_output[7568] + last_layer_output[7569] + last_layer_output[7570] + last_layer_output[7571] + last_layer_output[7572] + last_layer_output[7573] + last_layer_output[7574] + last_layer_output[7575] + last_layer_output[7576] + last_layer_output[7577] + last_layer_output[7578] + last_layer_output[7579] + last_layer_output[7580] + last_layer_output[7581] + last_layer_output[7582] + last_layer_output[7583] + last_layer_output[7584] + last_layer_output[7585] + last_layer_output[7586] + last_layer_output[7587] + last_layer_output[7588] + last_layer_output[7589] + last_layer_output[7590] + last_layer_output[7591] + last_layer_output[7592] + last_layer_output[7593] + last_layer_output[7594] + last_layer_output[7595] + last_layer_output[7596] + last_layer_output[7597] + last_layer_output[7598] + last_layer_output[7599] + last_layer_output[7600] + last_layer_output[7601] + last_layer_output[7602] + last_layer_output[7603] + last_layer_output[7604] + last_layer_output[7605] + last_layer_output[7606] + last_layer_output[7607] + last_layer_output[7608] + last_layer_output[7609] + last_layer_output[7610] + last_layer_output[7611] + last_layer_output[7612] + last_layer_output[7613] + last_layer_output[7614] + last_layer_output[7615] + last_layer_output[7616] + last_layer_output[7617] + last_layer_output[7618] + last_layer_output[7619] + last_layer_output[7620] + last_layer_output[7621] + last_layer_output[7622] + last_layer_output[7623] + last_layer_output[7624] + last_layer_output[7625] + last_layer_output[7626] + last_layer_output[7627] + last_layer_output[7628] + last_layer_output[7629] + last_layer_output[7630] + last_layer_output[7631] + last_layer_output[7632] + last_layer_output[7633] + last_layer_output[7634] + last_layer_output[7635] + last_layer_output[7636] + last_layer_output[7637] + last_layer_output[7638] + last_layer_output[7639] + last_layer_output[7640] + last_layer_output[7641] + last_layer_output[7642] + last_layer_output[7643] + last_layer_output[7644] + last_layer_output[7645] + last_layer_output[7646] + last_layer_output[7647] + last_layer_output[7648] + last_layer_output[7649] + last_layer_output[7650] + last_layer_output[7651] + last_layer_output[7652] + last_layer_output[7653] + last_layer_output[7654] + last_layer_output[7655] + last_layer_output[7656] + last_layer_output[7657] + last_layer_output[7658] + last_layer_output[7659] + last_layer_output[7660] + last_layer_output[7661] + last_layer_output[7662] + last_layer_output[7663] + last_layer_output[7664] + last_layer_output[7665] + last_layer_output[7666] + last_layer_output[7667] + last_layer_output[7668] + last_layer_output[7669] + last_layer_output[7670] + last_layer_output[7671] + last_layer_output[7672] + last_layer_output[7673] + last_layer_output[7674] + last_layer_output[7675] + last_layer_output[7676] + last_layer_output[7677] + last_layer_output[7678] + last_layer_output[7679] + last_layer_output[7680] + last_layer_output[7681] + last_layer_output[7682] + last_layer_output[7683] + last_layer_output[7684] + last_layer_output[7685] + last_layer_output[7686] + last_layer_output[7687] + last_layer_output[7688] + last_layer_output[7689] + last_layer_output[7690] + last_layer_output[7691] + last_layer_output[7692] + last_layer_output[7693] + last_layer_output[7694] + last_layer_output[7695] + last_layer_output[7696] + last_layer_output[7697] + last_layer_output[7698] + last_layer_output[7699] + last_layer_output[7700] + last_layer_output[7701] + last_layer_output[7702] + last_layer_output[7703] + last_layer_output[7704] + last_layer_output[7705] + last_layer_output[7706] + last_layer_output[7707] + last_layer_output[7708] + last_layer_output[7709] + last_layer_output[7710] + last_layer_output[7711] + last_layer_output[7712] + last_layer_output[7713] + last_layer_output[7714] + last_layer_output[7715] + last_layer_output[7716] + last_layer_output[7717] + last_layer_output[7718] + last_layer_output[7719] + last_layer_output[7720] + last_layer_output[7721] + last_layer_output[7722] + last_layer_output[7723] + last_layer_output[7724] + last_layer_output[7725] + last_layer_output[7726] + last_layer_output[7727] + last_layer_output[7728] + last_layer_output[7729] + last_layer_output[7730] + last_layer_output[7731] + last_layer_output[7732] + last_layer_output[7733] + last_layer_output[7734] + last_layer_output[7735] + last_layer_output[7736] + last_layer_output[7737] + last_layer_output[7738] + last_layer_output[7739] + last_layer_output[7740] + last_layer_output[7741] + last_layer_output[7742] + last_layer_output[7743] + last_layer_output[7744] + last_layer_output[7745] + last_layer_output[7746] + last_layer_output[7747] + last_layer_output[7748] + last_layer_output[7749] + last_layer_output[7750] + last_layer_output[7751] + last_layer_output[7752] + last_layer_output[7753] + last_layer_output[7754] + last_layer_output[7755] + last_layer_output[7756] + last_layer_output[7757] + last_layer_output[7758] + last_layer_output[7759] + last_layer_output[7760] + last_layer_output[7761] + last_layer_output[7762] + last_layer_output[7763] + last_layer_output[7764] + last_layer_output[7765] + last_layer_output[7766] + last_layer_output[7767] + last_layer_output[7768] + last_layer_output[7769] + last_layer_output[7770] + last_layer_output[7771] + last_layer_output[7772] + last_layer_output[7773] + last_layer_output[7774] + last_layer_output[7775] + last_layer_output[7776] + last_layer_output[7777] + last_layer_output[7778] + last_layer_output[7779] + last_layer_output[7780] + last_layer_output[7781] + last_layer_output[7782] + last_layer_output[7783] + last_layer_output[7784] + last_layer_output[7785] + last_layer_output[7786] + last_layer_output[7787] + last_layer_output[7788] + last_layer_output[7789] + last_layer_output[7790] + last_layer_output[7791] + last_layer_output[7792] + last_layer_output[7793] + last_layer_output[7794] + last_layer_output[7795] + last_layer_output[7796] + last_layer_output[7797] + last_layer_output[7798] + last_layer_output[7799] + last_layer_output[7800] + last_layer_output[7801] + last_layer_output[7802] + last_layer_output[7803] + last_layer_output[7804] + last_layer_output[7805] + last_layer_output[7806] + last_layer_output[7807] + last_layer_output[7808] + last_layer_output[7809] + last_layer_output[7810] + last_layer_output[7811] + last_layer_output[7812] + last_layer_output[7813] + last_layer_output[7814] + last_layer_output[7815] + last_layer_output[7816] + last_layer_output[7817] + last_layer_output[7818] + last_layer_output[7819] + last_layer_output[7820] + last_layer_output[7821] + last_layer_output[7822] + last_layer_output[7823] + last_layer_output[7824] + last_layer_output[7825] + last_layer_output[7826] + last_layer_output[7827] + last_layer_output[7828] + last_layer_output[7829] + last_layer_output[7830] + last_layer_output[7831] + last_layer_output[7832] + last_layer_output[7833] + last_layer_output[7834] + last_layer_output[7835] + last_layer_output[7836] + last_layer_output[7837] + last_layer_output[7838] + last_layer_output[7839] + last_layer_output[7840] + last_layer_output[7841] + last_layer_output[7842] + last_layer_output[7843] + last_layer_output[7844] + last_layer_output[7845] + last_layer_output[7846] + last_layer_output[7847] + last_layer_output[7848] + last_layer_output[7849] + last_layer_output[7850] + last_layer_output[7851] + last_layer_output[7852] + last_layer_output[7853] + last_layer_output[7854] + last_layer_output[7855] + last_layer_output[7856] + last_layer_output[7857] + last_layer_output[7858] + last_layer_output[7859] + last_layer_output[7860] + last_layer_output[7861] + last_layer_output[7862] + last_layer_output[7863] + last_layer_output[7864] + last_layer_output[7865] + last_layer_output[7866] + last_layer_output[7867] + last_layer_output[7868] + last_layer_output[7869] + last_layer_output[7870] + last_layer_output[7871] + last_layer_output[7872] + last_layer_output[7873] + last_layer_output[7874] + last_layer_output[7875] + last_layer_output[7876] + last_layer_output[7877] + last_layer_output[7878] + last_layer_output[7879] + last_layer_output[7880] + last_layer_output[7881] + last_layer_output[7882] + last_layer_output[7883] + last_layer_output[7884] + last_layer_output[7885] + last_layer_output[7886] + last_layer_output[7887] + last_layer_output[7888] + last_layer_output[7889] + last_layer_output[7890] + last_layer_output[7891] + last_layer_output[7892] + last_layer_output[7893] + last_layer_output[7894] + last_layer_output[7895] + last_layer_output[7896] + last_layer_output[7897] + last_layer_output[7898] + last_layer_output[7899] + last_layer_output[7900] + last_layer_output[7901] + last_layer_output[7902] + last_layer_output[7903] + last_layer_output[7904] + last_layer_output[7905] + last_layer_output[7906] + last_layer_output[7907] + last_layer_output[7908] + last_layer_output[7909] + last_layer_output[7910] + last_layer_output[7911] + last_layer_output[7912] + last_layer_output[7913] + last_layer_output[7914] + last_layer_output[7915] + last_layer_output[7916] + last_layer_output[7917] + last_layer_output[7918] + last_layer_output[7919] + last_layer_output[7920] + last_layer_output[7921] + last_layer_output[7922] + last_layer_output[7923] + last_layer_output[7924] + last_layer_output[7925] + last_layer_output[7926] + last_layer_output[7927] + last_layer_output[7928] + last_layer_output[7929] + last_layer_output[7930] + last_layer_output[7931] + last_layer_output[7932] + last_layer_output[7933] + last_layer_output[7934] + last_layer_output[7935] + last_layer_output[7936] + last_layer_output[7937] + last_layer_output[7938] + last_layer_output[7939] + last_layer_output[7940] + last_layer_output[7941] + last_layer_output[7942] + last_layer_output[7943] + last_layer_output[7944] + last_layer_output[7945] + last_layer_output[7946] + last_layer_output[7947] + last_layer_output[7948] + last_layer_output[7949] + last_layer_output[7950] + last_layer_output[7951] + last_layer_output[7952] + last_layer_output[7953] + last_layer_output[7954] + last_layer_output[7955] + last_layer_output[7956] + last_layer_output[7957] + last_layer_output[7958] + last_layer_output[7959] + last_layer_output[7960] + last_layer_output[7961] + last_layer_output[7962] + last_layer_output[7963] + last_layer_output[7964] + last_layer_output[7965] + last_layer_output[7966] + last_layer_output[7967] + last_layer_output[7968] + last_layer_output[7969] + last_layer_output[7970] + last_layer_output[7971] + last_layer_output[7972] + last_layer_output[7973] + last_layer_output[7974] + last_layer_output[7975] + last_layer_output[7976] + last_layer_output[7977] + last_layer_output[7978] + last_layer_output[7979] + last_layer_output[7980] + last_layer_output[7981] + last_layer_output[7982] + last_layer_output[7983] + last_layer_output[7984] + last_layer_output[7985] + last_layer_output[7986] + last_layer_output[7987] + last_layer_output[7988] + last_layer_output[7989] + last_layer_output[7990] + last_layer_output[7991] + last_layer_output[7992] + last_layer_output[7993] + last_layer_output[7994] + last_layer_output[7995] + last_layer_output[7996] + last_layer_output[7997] + last_layer_output[7998] + last_layer_output[7999];
      assign y[99:90]=result[0];
      assign y[89:80]=result[1];
      assign y[79:70]=result[2];
      assign y[69:60]=result[3];
      assign y[59:50]=result[4];
      assign y[49:40]=result[5];
      assign y[39:30]=result[6];
      assign y[29:20]=result[7];
      assign y[19:10]=result[8];
      assign y[9:0]=result[9];
endmodule
