module logic_network (    input wire [399:0] x,
    output wire [49:0] y
);
      wire [199:0] layer0_out;
      wire [199:0] layer1_out;
      wire [199:0] layer2_out;
      wire [199:0] layer3_out;
    assign layer0_out[0] = ~x[306];
    assign layer0_out[1] = ~(x[164] | x[165]);
    assign layer0_out[2] = ~(x[150] | x[151]);
    assign layer0_out[3] = x[46] | x[47];
    assign layer0_out[4] = x[291] & ~x[290];
    assign layer0_out[5] = ~x[311] | x[310];
    assign layer0_out[6] = ~x[80] | x[81];
    assign layer0_out[7] = ~(x[176] | x[177]);
    assign layer0_out[8] = 1'b0;
    assign layer0_out[9] = x[142] | x[143];
    assign layer0_out[10] = x[274] | x[275];
    assign layer0_out[11] = 1'b1;
    assign layer0_out[12] = ~x[93];
    assign layer0_out[13] = 1'b1;
    assign layer0_out[14] = 1'b1;
    assign layer0_out[15] = ~x[84];
    assign layer0_out[16] = x[82] ^ x[83];
    assign layer0_out[17] = x[266] | x[267];
    assign layer0_out[18] = 1'b1;
    assign layer0_out[19] = ~(x[184] | x[185]);
    assign layer0_out[20] = 1'b0;
    assign layer0_out[21] = x[129];
    assign layer0_out[22] = 1'b1;
    assign layer0_out[23] = x[190];
    assign layer0_out[24] = 1'b0;
    assign layer0_out[25] = 1'b1;
    assign layer0_out[26] = x[216] | x[217];
    assign layer0_out[27] = ~(x[300] | x[301]);
    assign layer0_out[28] = ~(x[188] | x[189]);
    assign layer0_out[29] = x[364] | x[365];
    assign layer0_out[30] = 1'b1;
    assign layer0_out[31] = ~(x[250] | x[251]);
    assign layer0_out[32] = x[76] | x[77];
    assign layer0_out[33] = x[194] & x[195];
    assign layer0_out[34] = 1'b1;
    assign layer0_out[35] = x[104] | x[105];
    assign layer0_out[36] = ~(x[248] | x[249]);
    assign layer0_out[37] = 1'b0;
    assign layer0_out[38] = x[236] | x[237];
    assign layer0_out[39] = ~(x[238] | x[239]);
    assign layer0_out[40] = x[15];
    assign layer0_out[41] = ~x[6] | x[7];
    assign layer0_out[42] = x[346];
    assign layer0_out[43] = x[172];
    assign layer0_out[44] = x[140] & ~x[141];
    assign layer0_out[45] = x[271];
    assign layer0_out[46] = 1'b0;
    assign layer0_out[47] = 1'b0;
    assign layer0_out[48] = x[348];
    assign layer0_out[49] = 1'b0;
    assign layer0_out[50] = x[278] | x[279];
    assign layer0_out[51] = x[74] | x[75];
    assign layer0_out[52] = x[334] | x[335];
    assign layer0_out[53] = x[262] | x[263];
    assign layer0_out[54] = ~(x[386] | x[387]);
    assign layer0_out[55] = ~(x[90] | x[91]);
    assign layer0_out[56] = ~x[317] | x[316];
    assign layer0_out[57] = x[181];
    assign layer0_out[58] = 1'b0;
    assign layer0_out[59] = ~(x[394] | x[395]);
    assign layer0_out[60] = ~x[41] | x[40];
    assign layer0_out[61] = x[242] | x[243];
    assign layer0_out[62] = x[158] | x[159];
    assign layer0_out[63] = x[3] & ~x[2];
    assign layer0_out[64] = x[44] | x[45];
    assign layer0_out[65] = x[264] | x[265];
    assign layer0_out[66] = x[370] & x[371];
    assign layer0_out[67] = x[350] | x[351];
    assign layer0_out[68] = 1'b1;
    assign layer0_out[69] = x[166] | x[167];
    assign layer0_out[70] = x[204] | x[205];
    assign layer0_out[71] = ~x[138];
    assign layer0_out[72] = ~x[110];
    assign layer0_out[73] = 1'b0;
    assign layer0_out[74] = ~(x[30] | x[31]);
    assign layer0_out[75] = ~x[168];
    assign layer0_out[76] = ~x[235];
    assign layer0_out[77] = ~(x[246] | x[247]);
    assign layer0_out[78] = 1'b0;
    assign layer0_out[79] = ~(x[284] | x[285]);
    assign layer0_out[80] = ~(x[124] | x[125]);
    assign layer0_out[81] = x[201];
    assign layer0_out[82] = x[118] ^ x[119];
    assign layer0_out[83] = ~x[29];
    assign layer0_out[84] = x[207];
    assign layer0_out[85] = 1'b0;
    assign layer0_out[86] = ~(x[202] | x[203]);
    assign layer0_out[87] = ~x[148];
    assign layer0_out[88] = ~x[113];
    assign layer0_out[89] = ~(x[152] | x[153]);
    assign layer0_out[90] = ~x[9] | x[8];
    assign layer0_out[91] = x[34] & x[35];
    assign layer0_out[92] = 1'b1;
    assign layer0_out[93] = 1'b1;
    assign layer0_out[94] = ~(x[170] | x[171]);
    assign layer0_out[95] = x[240] | x[241];
    assign layer0_out[96] = ~x[100] | x[101];
    assign layer0_out[97] = 1'b0;
    assign layer0_out[98] = ~(x[20] ^ x[21]);
    assign layer0_out[99] = x[126];
    assign layer0_out[100] = x[372] | x[373];
    assign layer0_out[101] = ~(x[106] | x[107]);
    assign layer0_out[102] = 1'b0;
    assign layer0_out[103] = ~(x[302] | x[303]);
    assign layer0_out[104] = ~(x[382] & x[383]);
    assign layer0_out[105] = ~(x[282] | x[283]);
    assign layer0_out[106] = ~x[221];
    assign layer0_out[107] = ~x[27];
    assign layer0_out[108] = x[280] | x[281];
    assign layer0_out[109] = x[322] | x[323];
    assign layer0_out[110] = 1'b1;
    assign layer0_out[111] = x[342] | x[343];
    assign layer0_out[112] = 1'b1;
    assign layer0_out[113] = x[344] | x[345];
    assign layer0_out[114] = 1'b0;
    assign layer0_out[115] = ~(x[218] | x[219]);
    assign layer0_out[116] = x[198] | x[199];
    assign layer0_out[117] = ~(x[222] | x[223]);
    assign layer0_out[118] = ~x[333];
    assign layer0_out[119] = x[276] | x[277];
    assign layer0_out[120] = x[48];
    assign layer0_out[121] = 1'b1;
    assign layer0_out[122] = x[286] | x[287];
    assign layer0_out[123] = x[53];
    assign layer0_out[124] = ~(x[54] | x[55]);
    assign layer0_out[125] = x[186] | x[187];
    assign layer0_out[126] = ~(x[174] | x[175]);
    assign layer0_out[127] = x[340] | x[341];
    assign layer0_out[128] = ~x[390];
    assign layer0_out[129] = x[388] | x[389];
    assign layer0_out[130] = ~(x[42] & x[43]);
    assign layer0_out[131] = x[154] | x[155];
    assign layer0_out[132] = ~(x[356] | x[357]);
    assign layer0_out[133] = ~(x[298] | x[299]);
    assign layer0_out[134] = ~(x[320] | x[321]);
    assign layer0_out[135] = x[366] | x[367];
    assign layer0_out[136] = ~(x[244] | x[245]);
    assign layer0_out[137] = ~x[209];
    assign layer0_out[138] = 1'b1;
    assign layer0_out[139] = x[324] | x[325];
    assign layer0_out[140] = x[147];
    assign layer0_out[141] = ~(x[0] ^ x[1]);
    assign layer0_out[142] = ~x[61];
    assign layer0_out[143] = ~x[259] | x[258];
    assign layer0_out[144] = x[224] | x[225];
    assign layer0_out[145] = x[36] | x[37];
    assign layer0_out[146] = ~(x[380] | x[381]);
    assign layer0_out[147] = 1'b1;
    assign layer0_out[148] = ~(x[136] | x[137]);
    assign layer0_out[149] = x[294] | x[295];
    assign layer0_out[150] = 1'b1;
    assign layer0_out[151] = ~(x[256] | x[257]);
    assign layer0_out[152] = x[318] | x[319];
    assign layer0_out[153] = 1'b1;
    assign layer0_out[154] = 1'b1;
    assign layer0_out[155] = x[162] | x[163];
    assign layer0_out[156] = ~(x[22] ^ x[23]);
    assign layer0_out[157] = x[98] & ~x[99];
    assign layer0_out[158] = x[308] | x[309];
    assign layer0_out[159] = ~(x[96] | x[97]);
    assign layer0_out[160] = ~(x[254] | x[255]);
    assign layer0_out[161] = x[229];
    assign layer0_out[162] = x[12] | x[13];
    assign layer0_out[163] = 1'b0;
    assign layer0_out[164] = ~(x[24] | x[25]);
    assign layer0_out[165] = ~(x[66] | x[67]);
    assign layer0_out[166] = ~(x[296] | x[297]);
    assign layer0_out[167] = x[196] | x[197];
    assign layer0_out[168] = ~(x[358] & x[359]);
    assign layer0_out[169] = x[134] | x[135];
    assign layer0_out[170] = x[95];
    assign layer0_out[171] = x[313];
    assign layer0_out[172] = ~(x[132] | x[133]);
    assign layer0_out[173] = x[114] | x[115];
    assign layer0_out[174] = ~x[17] | x[16];
    assign layer0_out[175] = x[272];
    assign layer0_out[176] = x[233];
    assign layer0_out[177] = ~(x[384] | x[385]);
    assign layer0_out[178] = x[56] | x[57];
    assign layer0_out[179] = x[116] | x[117];
    assign layer0_out[180] = ~x[59];
    assign layer0_out[181] = 1'b0;
    assign layer0_out[182] = ~(x[288] | x[289]);
    assign layer0_out[183] = x[32] & x[33];
    assign layer0_out[184] = x[304];
    assign layer0_out[185] = ~(x[38] | x[39]);
    assign layer0_out[186] = 1'b1;
    assign layer0_out[187] = ~x[399] | x[398];
    assign layer0_out[188] = x[378] | x[379];
    assign layer0_out[189] = 1'b0;
    assign layer0_out[190] = x[130] | x[131];
    assign layer0_out[191] = ~x[102];
    assign layer0_out[192] = x[214] | x[215];
    assign layer0_out[193] = x[336] | x[337];
    assign layer0_out[194] = 1'b0;
    assign layer0_out[195] = x[355];
    assign layer0_out[196] = ~x[231];
    assign layer0_out[197] = x[368] & x[369];
    assign layer0_out[198] = x[78] | x[79];
    assign layer0_out[199] = x[226];
    assign layer1_out[0] = layer0_out[188];
    assign layer1_out[1] = ~layer0_out[61];
    assign layer1_out[2] = layer0_out[4] & ~layer0_out[5];
    assign layer1_out[3] = layer0_out[15] & ~layer0_out[16];
    assign layer1_out[4] = 1'b0;
    assign layer1_out[5] = layer0_out[166];
    assign layer1_out[6] = layer0_out[139];
    assign layer1_out[7] = ~(layer0_out[52] | layer0_out[53]);
    assign layer1_out[8] = ~layer0_out[116] | layer0_out[117];
    assign layer1_out[9] = layer0_out[111];
    assign layer1_out[10] = ~layer0_out[174] | layer0_out[173];
    assign layer1_out[11] = 1'b0;
    assign layer1_out[12] = ~layer0_out[45];
    assign layer1_out[13] = ~layer0_out[135];
    assign layer1_out[14] = ~layer0_out[131];
    assign layer1_out[15] = layer0_out[155];
    assign layer1_out[16] = ~(layer0_out[89] | layer0_out[90]);
    assign layer1_out[17] = layer0_out[185];
    assign layer1_out[18] = ~(layer0_out[47] | layer0_out[48]);
    assign layer1_out[19] = ~(layer0_out[141] ^ layer0_out[142]);
    assign layer1_out[20] = ~(layer0_out[79] & layer0_out[80]);
    assign layer1_out[21] = layer0_out[94];
    assign layer1_out[22] = layer0_out[67];
    assign layer1_out[23] = ~layer0_out[135] | layer0_out[136];
    assign layer1_out[24] = 1'b1;
    assign layer1_out[25] = ~layer0_out[113];
    assign layer1_out[26] = 1'b1;
    assign layer1_out[27] = ~layer0_out[86];
    assign layer1_out[28] = ~layer0_out[7];
    assign layer1_out[29] = ~(layer0_out[69] | layer0_out[70]);
    assign layer1_out[30] = ~layer0_out[146];
    assign layer1_out[31] = layer0_out[95];
    assign layer1_out[32] = layer0_out[152];
    assign layer1_out[33] = ~layer0_out[91];
    assign layer1_out[34] = layer0_out[106] & ~layer0_out[107];
    assign layer1_out[35] = layer0_out[182];
    assign layer1_out[36] = layer0_out[19];
    assign layer1_out[37] = ~(layer0_out[49] & layer0_out[50]);
    assign layer1_out[38] = ~layer0_out[164] | layer0_out[165];
    assign layer1_out[39] = layer0_out[13] | layer0_out[14];
    assign layer1_out[40] = ~layer0_out[77];
    assign layer1_out[41] = layer0_out[102] | layer0_out[103];
    assign layer1_out[42] = layer0_out[142];
    assign layer1_out[43] = 1'b1;
    assign layer1_out[44] = 1'b0;
    assign layer1_out[45] = 1'b1;
    assign layer1_out[46] = layer0_out[17];
    assign layer1_out[47] = ~layer0_out[101];
    assign layer1_out[48] = ~layer0_out[133] | layer0_out[134];
    assign layer1_out[49] = layer0_out[51] & ~layer0_out[50];
    assign layer1_out[50] = layer0_out[148] & layer0_out[149];
    assign layer1_out[51] = ~layer0_out[66];
    assign layer1_out[52] = ~(layer0_out[190] | layer0_out[191]);
    assign layer1_out[53] = layer0_out[0];
    assign layer1_out[54] = ~layer0_out[122];
    assign layer1_out[55] = ~layer0_out[151];
    assign layer1_out[56] = layer0_out[191] & ~layer0_out[192];
    assign layer1_out[57] = ~layer0_out[79];
    assign layer1_out[58] = layer0_out[160];
    assign layer1_out[59] = layer0_out[132] & layer0_out[133];
    assign layer1_out[60] = layer0_out[55] ^ layer0_out[56];
    assign layer1_out[61] = ~(layer0_out[73] ^ layer0_out[74]);
    assign layer1_out[62] = layer0_out[185];
    assign layer1_out[63] = ~layer0_out[123];
    assign layer1_out[64] = 1'b0;
    assign layer1_out[65] = layer0_out[41] & ~layer0_out[42];
    assign layer1_out[66] = ~(layer0_out[37] & layer0_out[38]);
    assign layer1_out[67] = layer0_out[19];
    assign layer1_out[68] = layer0_out[172];
    assign layer1_out[69] = layer0_out[44] & layer0_out[45];
    assign layer1_out[70] = ~(layer0_out[0] & layer0_out[2]);
    assign layer1_out[71] = layer0_out[17] & layer0_out[18];
    assign layer1_out[72] = ~layer0_out[126] | layer0_out[127];
    assign layer1_out[73] = layer0_out[35];
    assign layer1_out[74] = layer0_out[36] | layer0_out[37];
    assign layer1_out[75] = ~layer0_out[65];
    assign layer1_out[76] = layer0_out[83] & ~layer0_out[82];
    assign layer1_out[77] = layer0_out[193];
    assign layer1_out[78] = 1'b1;
    assign layer1_out[79] = layer0_out[129] & layer0_out[130];
    assign layer1_out[80] = layer0_out[109];
    assign layer1_out[81] = ~layer0_out[163] | layer0_out[164];
    assign layer1_out[82] = layer0_out[166] & ~layer0_out[167];
    assign layer1_out[83] = layer0_out[48] & ~layer0_out[49];
    assign layer1_out[84] = ~layer0_out[130] | layer0_out[131];
    assign layer1_out[85] = layer0_out[186] | layer0_out[187];
    assign layer1_out[86] = layer0_out[27] & ~layer0_out[26];
    assign layer1_out[87] = ~layer0_out[5] | layer0_out[6];
    assign layer1_out[88] = layer0_out[62];
    assign layer1_out[89] = layer0_out[117] & ~layer0_out[118];
    assign layer1_out[90] = ~layer0_out[29];
    assign layer1_out[91] = ~(layer0_out[169] | layer0_out[170]);
    assign layer1_out[92] = ~layer0_out[27] | layer0_out[28];
    assign layer1_out[93] = layer0_out[107] & ~layer0_out[108];
    assign layer1_out[94] = ~layer0_out[21];
    assign layer1_out[95] = layer0_out[125];
    assign layer1_out[96] = layer0_out[9];
    assign layer1_out[97] = layer0_out[151] & ~layer0_out[152];
    assign layer1_out[98] = ~(layer0_out[179] | layer0_out[180]);
    assign layer1_out[99] = layer0_out[32];
    assign layer1_out[100] = layer0_out[64] & ~layer0_out[65];
    assign layer1_out[101] = layer0_out[137];
    assign layer1_out[102] = 1'b0;
    assign layer1_out[103] = layer0_out[10];
    assign layer1_out[104] = layer0_out[170] | layer0_out[171];
    assign layer1_out[105] = layer0_out[178] | layer0_out[179];
    assign layer1_out[106] = layer0_out[28] & ~layer0_out[29];
    assign layer1_out[107] = layer0_out[81];
    assign layer1_out[108] = layer0_out[193];
    assign layer1_out[109] = ~layer0_out[8] | layer0_out[9];
    assign layer1_out[110] = layer0_out[85];
    assign layer1_out[111] = layer0_out[149] & layer0_out[150];
    assign layer1_out[112] = ~layer0_out[92];
    assign layer1_out[113] = layer0_out[129];
    assign layer1_out[114] = layer0_out[182];
    assign layer1_out[115] = ~layer0_out[120];
    assign layer1_out[116] = ~layer0_out[43] | layer0_out[44];
    assign layer1_out[117] = layer0_out[162];
    assign layer1_out[118] = layer0_out[22] & ~layer0_out[23];
    assign layer1_out[119] = layer0_out[69];
    assign layer1_out[120] = ~(layer0_out[140] & layer0_out[141]);
    assign layer1_out[121] = layer0_out[71] & ~layer0_out[70];
    assign layer1_out[122] = layer0_out[197];
    assign layer1_out[123] = layer0_out[195];
    assign layer1_out[124] = layer0_out[61] | layer0_out[62];
    assign layer1_out[125] = ~layer0_out[58];
    assign layer1_out[126] = layer0_out[12];
    assign layer1_out[127] = ~layer0_out[72];
    assign layer1_out[128] = layer0_out[104] & layer0_out[105];
    assign layer1_out[129] = ~layer0_out[54] | layer0_out[53];
    assign layer1_out[130] = layer0_out[155];
    assign layer1_out[131] = layer0_out[91] & ~layer0_out[92];
    assign layer1_out[132] = ~layer0_out[78];
    assign layer1_out[133] = ~layer0_out[120] | layer0_out[119];
    assign layer1_out[134] = ~(layer0_out[153] | layer0_out[154]);
    assign layer1_out[135] = layer0_out[54] & layer0_out[55];
    assign layer1_out[136] = layer0_out[196];
    assign layer1_out[137] = layer0_out[59];
    assign layer1_out[138] = ~(layer0_out[72] | layer0_out[73]);
    assign layer1_out[139] = ~layer0_out[138] | layer0_out[139];
    assign layer1_out[140] = ~layer0_out[181] | layer0_out[180];
    assign layer1_out[141] = 1'b0;
    assign layer1_out[142] = ~(layer0_out[198] | layer0_out[199]);
    assign layer1_out[143] = ~layer0_out[3];
    assign layer1_out[144] = ~(layer0_out[35] | layer0_out[36]);
    assign layer1_out[145] = ~(layer0_out[105] & layer0_out[106]);
    assign layer1_out[146] = 1'b0;
    assign layer1_out[147] = layer0_out[6] & layer0_out[7];
    assign layer1_out[148] = ~(layer0_out[127] & layer0_out[128]);
    assign layer1_out[149] = ~(layer0_out[75] & layer0_out[76]);
    assign layer1_out[150] = layer0_out[58];
    assign layer1_out[151] = ~(layer0_out[158] & layer0_out[159]);
    assign layer1_out[152] = layer0_out[43];
    assign layer1_out[153] = layer0_out[51] & ~layer0_out[52];
    assign layer1_out[154] = layer0_out[167] & layer0_out[168];
    assign layer1_out[155] = layer0_out[23];
    assign layer1_out[156] = layer0_out[74] | layer0_out[75];
    assign layer1_out[157] = layer0_out[172];
    assign layer1_out[158] = ~layer0_out[144];
    assign layer1_out[159] = ~layer0_out[24] | layer0_out[25];
    assign layer1_out[160] = layer0_out[63] | layer0_out[64];
    assign layer1_out[161] = layer0_out[125] | layer0_out[126];
    assign layer1_out[162] = layer0_out[113];
    assign layer1_out[163] = layer0_out[12] | layer0_out[13];
    assign layer1_out[164] = layer0_out[100] & ~layer0_out[99];
    assign layer1_out[165] = layer0_out[147];
    assign layer1_out[166] = 1'b1;
    assign layer1_out[167] = layer0_out[158];
    assign layer1_out[168] = layer0_out[30];
    assign layer1_out[169] = ~layer0_out[177] | layer0_out[178];
    assign layer1_out[170] = layer0_out[168] & ~layer0_out[169];
    assign layer1_out[171] = ~layer0_out[159] | layer0_out[160];
    assign layer1_out[172] = layer0_out[144] & ~layer0_out[145];
    assign layer1_out[173] = 1'b0;
    assign layer1_out[174] = layer0_out[175];
    assign layer1_out[175] = ~(layer0_out[176] | layer0_out[177]);
    assign layer1_out[176] = layer0_out[146] & ~layer0_out[145];
    assign layer1_out[177] = ~layer0_out[88];
    assign layer1_out[178] = layer0_out[138] & ~layer0_out[137];
    assign layer1_out[179] = layer0_out[88] & layer0_out[89];
    assign layer1_out[180] = layer0_out[93] | layer0_out[94];
    assign layer1_out[181] = 1'b1;
    assign layer1_out[182] = layer0_out[184];
    assign layer1_out[183] = ~layer0_out[124] | layer0_out[123];
    assign layer1_out[184] = ~(layer0_out[196] | layer0_out[197]);
    assign layer1_out[185] = layer0_out[80] & ~layer0_out[81];
    assign layer1_out[186] = layer0_out[39] & ~layer0_out[38];
    assign layer1_out[187] = ~layer0_out[2] | layer0_out[1];
    assign layer1_out[188] = ~layer0_out[84] | layer0_out[83];
    assign layer1_out[189] = ~layer0_out[118] | layer0_out[119];
    assign layer1_out[190] = ~(layer0_out[39] & layer0_out[40]);
    assign layer1_out[191] = layer0_out[109] & layer0_out[110];
    assign layer1_out[192] = ~layer0_out[31];
    assign layer1_out[193] = ~layer0_out[115] | layer0_out[116];
    assign layer1_out[194] = ~layer0_out[87];
    assign layer1_out[195] = 1'b0;
    assign layer1_out[196] = ~layer0_out[111];
    assign layer1_out[197] = layer0_out[103] & layer0_out[104];
    assign layer1_out[198] = layer0_out[2];
    assign layer1_out[199] = 1'b1;
    assign layer2_out[0] = ~layer1_out[15];
    assign layer2_out[1] = ~layer1_out[113];
    assign layer2_out[2] = layer1_out[27];
    assign layer2_out[3] = layer1_out[25];
    assign layer2_out[4] = layer1_out[198];
    assign layer2_out[5] = ~layer1_out[198];
    assign layer2_out[6] = layer1_out[83];
    assign layer2_out[7] = ~layer1_out[120] | layer1_out[119];
    assign layer2_out[8] = layer1_out[194] & ~layer1_out[193];
    assign layer2_out[9] = layer1_out[14];
    assign layer2_out[10] = layer1_out[46];
    assign layer2_out[11] = layer1_out[167];
    assign layer2_out[12] = ~layer1_out[100];
    assign layer2_out[13] = layer1_out[17] | layer1_out[18];
    assign layer2_out[14] = layer1_out[188] & ~layer1_out[187];
    assign layer2_out[15] = 1'b1;
    assign layer2_out[16] = layer1_out[155] & ~layer1_out[154];
    assign layer2_out[17] = layer1_out[51];
    assign layer2_out[18] = layer1_out[79] | layer1_out[80];
    assign layer2_out[19] = layer1_out[96];
    assign layer2_out[20] = ~(layer1_out[108] ^ layer1_out[109]);
    assign layer2_out[21] = layer1_out[121];
    assign layer2_out[22] = layer1_out[91];
    assign layer2_out[23] = ~layer1_out[114];
    assign layer2_out[24] = layer1_out[182];
    assign layer2_out[25] = ~layer1_out[44] | layer1_out[45];
    assign layer2_out[26] = ~layer1_out[119];
    assign layer2_out[27] = ~(layer1_out[180] | layer1_out[181]);
    assign layer2_out[28] = ~layer1_out[153];
    assign layer2_out[29] = ~layer1_out[103];
    assign layer2_out[30] = ~layer1_out[41] | layer1_out[40];
    assign layer2_out[31] = ~(layer1_out[196] & layer1_out[197]);
    assign layer2_out[32] = layer1_out[186];
    assign layer2_out[33] = ~layer1_out[89];
    assign layer2_out[34] = layer1_out[126];
    assign layer2_out[35] = layer1_out[3] ^ layer1_out[4];
    assign layer2_out[36] = layer1_out[97];
    assign layer2_out[37] = ~layer1_out[20];
    assign layer2_out[38] = layer1_out[50];
    assign layer2_out[39] = layer1_out[141];
    assign layer2_out[40] = layer1_out[58];
    assign layer2_out[41] = ~(layer1_out[10] ^ layer1_out[11]);
    assign layer2_out[42] = layer1_out[12] | layer1_out[13];
    assign layer2_out[43] = ~layer1_out[109];
    assign layer2_out[44] = ~layer1_out[167];
    assign layer2_out[45] = layer1_out[156];
    assign layer2_out[46] = ~layer1_out[128];
    assign layer2_out[47] = layer1_out[7] & layer1_out[8];
    assign layer2_out[48] = layer1_out[29];
    assign layer2_out[49] = layer1_out[90] & ~layer1_out[89];
    assign layer2_out[50] = ~(layer1_out[173] & layer1_out[174]);
    assign layer2_out[51] = layer1_out[135];
    assign layer2_out[52] = 1'b0;
    assign layer2_out[53] = layer1_out[118];
    assign layer2_out[54] = layer1_out[57];
    assign layer2_out[55] = layer1_out[116];
    assign layer2_out[56] = layer1_out[121];
    assign layer2_out[57] = layer1_out[128];
    assign layer2_out[58] = layer1_out[72] | layer1_out[73];
    assign layer2_out[59] = ~layer1_out[46];
    assign layer2_out[60] = ~layer1_out[194];
    assign layer2_out[61] = ~(layer1_out[104] | layer1_out[105]);
    assign layer2_out[62] = layer1_out[151] & layer1_out[152];
    assign layer2_out[63] = ~layer1_out[6];
    assign layer2_out[64] = ~(layer1_out[150] & layer1_out[151]);
    assign layer2_out[65] = ~layer1_out[67];
    assign layer2_out[66] = layer1_out[92];
    assign layer2_out[67] = layer1_out[196];
    assign layer2_out[68] = layer1_out[154];
    assign layer2_out[69] = layer1_out[51] & ~layer1_out[50];
    assign layer2_out[70] = ~layer1_out[175];
    assign layer2_out[71] = ~layer1_out[174];
    assign layer2_out[72] = layer1_out[136] & ~layer1_out[135];
    assign layer2_out[73] = layer1_out[111];
    assign layer2_out[74] = ~layer1_out[53];
    assign layer2_out[75] = ~layer1_out[100] | layer1_out[99];
    assign layer2_out[76] = layer1_out[62];
    assign layer2_out[77] = layer1_out[64] & layer1_out[65];
    assign layer2_out[78] = layer1_out[144] & ~layer1_out[145];
    assign layer2_out[79] = layer1_out[186] & ~layer1_out[187];
    assign layer2_out[80] = layer1_out[38];
    assign layer2_out[81] = layer1_out[94] & layer1_out[95];
    assign layer2_out[82] = layer1_out[114] | layer1_out[115];
    assign layer2_out[83] = ~layer1_out[171] | layer1_out[172];
    assign layer2_out[84] = layer1_out[26] | layer1_out[27];
    assign layer2_out[85] = layer1_out[170];
    assign layer2_out[86] = ~layer1_out[111];
    assign layer2_out[87] = ~layer1_out[164];
    assign layer2_out[88] = ~(layer1_out[48] & layer1_out[49]);
    assign layer2_out[89] = layer1_out[144];
    assign layer2_out[90] = layer1_out[136] & layer1_out[137];
    assign layer2_out[91] = layer1_out[59] & layer1_out[60];
    assign layer2_out[92] = ~layer1_out[93];
    assign layer2_out[93] = ~(layer1_out[123] | layer1_out[124]);
    assign layer2_out[94] = ~layer1_out[67];
    assign layer2_out[95] = layer1_out[184] & ~layer1_out[185];
    assign layer2_out[96] = layer1_out[15] & ~layer1_out[16];
    assign layer2_out[97] = ~layer1_out[188] | layer1_out[189];
    assign layer2_out[98] = layer1_out[176] | layer1_out[177];
    assign layer2_out[99] = ~layer1_out[157];
    assign layer2_out[100] = ~layer1_out[183];
    assign layer2_out[101] = ~(layer1_out[34] | layer1_out[35]);
    assign layer2_out[102] = layer1_out[79];
    assign layer2_out[103] = layer1_out[54];
    assign layer2_out[104] = layer1_out[57];
    assign layer2_out[105] = layer1_out[88];
    assign layer2_out[106] = ~layer1_out[162];
    assign layer2_out[107] = layer1_out[98] ^ layer1_out[99];
    assign layer2_out[108] = ~layer1_out[193];
    assign layer2_out[109] = ~(layer1_out[41] & layer1_out[42]);
    assign layer2_out[110] = layer1_out[23];
    assign layer2_out[111] = layer1_out[162];
    assign layer2_out[112] = layer1_out[137];
    assign layer2_out[113] = layer1_out[179];
    assign layer2_out[114] = ~(layer1_out[158] ^ layer1_out[159]);
    assign layer2_out[115] = ~(layer1_out[190] & layer1_out[191]);
    assign layer2_out[116] = layer1_out[108] & ~layer1_out[107];
    assign layer2_out[117] = layer1_out[33] & layer1_out[34];
    assign layer2_out[118] = layer1_out[64];
    assign layer2_out[119] = ~layer1_out[65];
    assign layer2_out[120] = ~(layer1_out[18] & layer1_out[19]);
    assign layer2_out[121] = ~layer1_out[81] | layer1_out[80];
    assign layer2_out[122] = ~(layer1_out[141] & layer1_out[142]);
    assign layer2_out[123] = layer1_out[28];
    assign layer2_out[124] = ~(layer1_out[95] | layer1_out[96]);
    assign layer2_out[125] = layer1_out[139] ^ layer1_out[140];
    assign layer2_out[126] = 1'b1;
    assign layer2_out[127] = ~layer1_out[25];
    assign layer2_out[128] = 1'b0;
    assign layer2_out[129] = layer1_out[133] | layer1_out[134];
    assign layer2_out[130] = ~layer1_out[48] | layer1_out[47];
    assign layer2_out[131] = ~layer1_out[129] | layer1_out[130];
    assign layer2_out[132] = ~layer1_out[166] | layer1_out[165];
    assign layer2_out[133] = ~(layer1_out[55] | layer1_out[56]);
    assign layer2_out[134] = ~layer1_out[156];
    assign layer2_out[135] = ~layer1_out[169];
    assign layer2_out[136] = layer1_out[42] & ~layer1_out[43];
    assign layer2_out[137] = layer1_out[148] & layer1_out[149];
    assign layer2_out[138] = layer1_out[81] ^ layer1_out[82];
    assign layer2_out[139] = ~(layer1_out[147] ^ layer1_out[148]);
    assign layer2_out[140] = ~layer1_out[22] | layer1_out[21];
    assign layer2_out[141] = layer1_out[86];
    assign layer2_out[142] = ~(layer1_out[32] ^ layer1_out[33]);
    assign layer2_out[143] = ~(layer1_out[101] ^ layer1_out[102]);
    assign layer2_out[144] = ~layer1_out[178];
    assign layer2_out[145] = ~(layer1_out[142] & layer1_out[143]);
    assign layer2_out[146] = ~layer1_out[8] | layer1_out[9];
    assign layer2_out[147] = ~layer1_out[17];
    assign layer2_out[148] = layer1_out[37] & layer1_out[38];
    assign layer2_out[149] = layer1_out[76];
    assign layer2_out[150] = ~(layer1_out[70] | layer1_out[71]);
    assign layer2_out[151] = ~layer1_out[132] | layer1_out[133];
    assign layer2_out[152] = layer1_out[75];
    assign layer2_out[153] = ~layer1_out[106] | layer1_out[107];
    assign layer2_out[154] = layer1_out[105] | layer1_out[106];
    assign layer2_out[155] = layer1_out[83];
    assign layer2_out[156] = layer1_out[86];
    assign layer2_out[157] = layer1_out[61] & ~layer1_out[60];
    assign layer2_out[158] = layer1_out[11] ^ layer1_out[12];
    assign layer2_out[159] = ~layer1_out[44] | layer1_out[43];
    assign layer2_out[160] = layer1_out[70];
    assign layer2_out[161] = layer1_out[36];
    assign layer2_out[162] = ~layer1_out[0] | layer1_out[1];
    assign layer2_out[163] = layer1_out[74];
    assign layer2_out[164] = layer1_out[139];
    assign layer2_out[165] = layer1_out[7];
    assign layer2_out[166] = layer1_out[130];
    assign layer2_out[167] = ~layer1_out[93];
    assign layer2_out[168] = layer1_out[2];
    assign layer2_out[169] = layer1_out[177];
    assign layer2_out[170] = ~layer1_out[170];
    assign layer2_out[171] = ~(layer1_out[146] & layer1_out[147]);
    assign layer2_out[172] = layer1_out[10] & ~layer1_out[9];
    assign layer2_out[173] = ~layer1_out[116];
    assign layer2_out[174] = layer1_out[172] | layer1_out[173];
    assign layer2_out[175] = layer1_out[161] & ~layer1_out[160];
    assign layer2_out[176] = ~layer1_out[68];
    assign layer2_out[177] = ~layer1_out[72];
    assign layer2_out[178] = ~layer1_out[40];
    assign layer2_out[179] = layer1_out[145];
    assign layer2_out[180] = layer1_out[31] & ~layer1_out[32];
    assign layer2_out[181] = layer1_out[5];
    assign layer2_out[182] = layer1_out[124];
    assign layer2_out[183] = layer1_out[30];
    assign layer2_out[184] = layer1_out[123];
    assign layer2_out[185] = ~layer1_out[192] | layer1_out[191];
    assign layer2_out[186] = layer1_out[84] ^ layer1_out[85];
    assign layer2_out[187] = ~layer1_out[76];
    assign layer2_out[188] = ~layer1_out[20];
    assign layer2_out[189] = layer1_out[3];
    assign layer2_out[190] = layer1_out[36];
    assign layer2_out[191] = layer1_out[1] & ~layer1_out[2];
    assign layer2_out[192] = ~layer1_out[159] | layer1_out[160];
    assign layer2_out[193] = layer1_out[54] & layer1_out[55];
    assign layer2_out[194] = ~layer1_out[149] | layer1_out[150];
    assign layer2_out[195] = layer1_out[125];
    assign layer2_out[196] = ~layer1_out[23];
    assign layer2_out[197] = ~layer1_out[103];
    assign layer2_out[198] = layer1_out[61];
    assign layer2_out[199] = layer1_out[131] & ~layer1_out[132];
    assign layer3_out[0] = ~layer2_out[181] | layer2_out[180];
    assign layer3_out[1] = layer2_out[65];
    assign layer3_out[2] = layer2_out[31] & ~layer2_out[32];
    assign layer3_out[3] = layer2_out[121];
    assign layer3_out[4] = layer2_out[90] & ~layer2_out[89];
    assign layer3_out[5] = ~(layer2_out[122] ^ layer2_out[123]);
    assign layer3_out[6] = layer2_out[14];
    assign layer3_out[7] = layer2_out[144] & ~layer2_out[143];
    assign layer3_out[8] = layer2_out[68];
    assign layer3_out[9] = ~layer2_out[156];
    assign layer3_out[10] = layer2_out[111];
    assign layer3_out[11] = ~layer2_out[99];
    assign layer3_out[12] = ~layer2_out[86];
    assign layer3_out[13] = layer2_out[182];
    assign layer3_out[14] = ~layer2_out[106];
    assign layer3_out[15] = layer2_out[146];
    assign layer3_out[16] = layer2_out[127];
    assign layer3_out[17] = ~layer2_out[21];
    assign layer3_out[18] = layer2_out[164] & ~layer2_out[165];
    assign layer3_out[19] = ~(layer2_out[114] & layer2_out[115]);
    assign layer3_out[20] = layer2_out[91];
    assign layer3_out[21] = layer2_out[177];
    assign layer3_out[22] = layer2_out[78];
    assign layer3_out[23] = layer2_out[98] & ~layer2_out[97];
    assign layer3_out[24] = layer2_out[22] & layer2_out[23];
    assign layer3_out[25] = layer2_out[48];
    assign layer3_out[26] = layer2_out[143];
    assign layer3_out[27] = layer2_out[47] & layer2_out[48];
    assign layer3_out[28] = layer2_out[125];
    assign layer3_out[29] = layer2_out[194];
    assign layer3_out[30] = layer2_out[61];
    assign layer3_out[31] = layer2_out[23] & ~layer2_out[24];
    assign layer3_out[32] = layer2_out[188];
    assign layer3_out[33] = layer2_out[41] & layer2_out[42];
    assign layer3_out[34] = ~layer2_out[92];
    assign layer3_out[35] = layer2_out[21] & layer2_out[22];
    assign layer3_out[36] = layer2_out[160] & layer2_out[161];
    assign layer3_out[37] = ~layer2_out[145];
    assign layer3_out[38] = layer2_out[101];
    assign layer3_out[39] = ~layer2_out[58];
    assign layer3_out[40] = layer2_out[55] & layer2_out[56];
    assign layer3_out[41] = layer2_out[184];
    assign layer3_out[42] = layer2_out[124] & ~layer2_out[125];
    assign layer3_out[43] = ~layer2_out[158];
    assign layer3_out[44] = ~(layer2_out[102] | layer2_out[103]);
    assign layer3_out[45] = ~layer2_out[33];
    assign layer3_out[46] = layer2_out[116];
    assign layer3_out[47] = layer2_out[53];
    assign layer3_out[48] = layer2_out[66] & ~layer2_out[65];
    assign layer3_out[49] = layer2_out[117];
    assign layer3_out[50] = layer2_out[133];
    assign layer3_out[51] = ~layer2_out[137];
    assign layer3_out[52] = layer2_out[41];
    assign layer3_out[53] = ~layer2_out[175];
    assign layer3_out[54] = layer2_out[66] & ~layer2_out[67];
    assign layer3_out[55] = ~layer2_out[115] | layer2_out[116];
    assign layer3_out[56] = layer2_out[119];
    assign layer3_out[57] = ~layer2_out[178];
    assign layer3_out[58] = ~layer2_out[154];
    assign layer3_out[59] = ~(layer2_out[2] | layer2_out[3]);
    assign layer3_out[60] = layer2_out[193];
    assign layer3_out[61] = layer2_out[62];
    assign layer3_out[62] = layer2_out[0] & ~layer2_out[2];
    assign layer3_out[63] = layer2_out[50] ^ layer2_out[51];
    assign layer3_out[64] = layer2_out[71];
    assign layer3_out[65] = ~(layer2_out[10] | layer2_out[11]);
    assign layer3_out[66] = ~(layer2_out[12] & layer2_out[13]);
    assign layer3_out[67] = ~layer2_out[14];
    assign layer3_out[68] = layer2_out[167] & ~layer2_out[166];
    assign layer3_out[69] = layer2_out[193];
    assign layer3_out[70] = layer2_out[73] & ~layer2_out[74];
    assign layer3_out[71] = ~layer2_out[69];
    assign layer3_out[72] = ~layer2_out[87];
    assign layer3_out[73] = ~(layer2_out[29] | layer2_out[30]);
    assign layer3_out[74] = layer2_out[5];
    assign layer3_out[75] = layer2_out[114] & ~layer2_out[113];
    assign layer3_out[76] = ~layer2_out[140];
    assign layer3_out[77] = layer2_out[37];
    assign layer3_out[78] = layer2_out[120];
    assign layer3_out[79] = layer2_out[185];
    assign layer3_out[80] = ~layer2_out[190];
    assign layer3_out[81] = ~layer2_out[18];
    assign layer3_out[82] = layer2_out[63];
    assign layer3_out[83] = ~(layer2_out[198] ^ layer2_out[199]);
    assign layer3_out[84] = layer2_out[95] | layer2_out[96];
    assign layer3_out[85] = layer2_out[17] & ~layer2_out[18];
    assign layer3_out[86] = layer2_out[44];
    assign layer3_out[87] = layer2_out[36] & ~layer2_out[35];
    assign layer3_out[88] = layer2_out[57] & ~layer2_out[56];
    assign layer3_out[89] = ~layer2_out[0];
    assign layer3_out[90] = layer2_out[169];
    assign layer3_out[91] = layer2_out[51];
    assign layer3_out[92] = layer2_out[171] & layer2_out[172];
    assign layer3_out[93] = ~layer2_out[198];
    assign layer3_out[94] = ~layer2_out[155];
    assign layer3_out[95] = layer2_out[126] & ~layer2_out[127];
    assign layer3_out[96] = ~(layer2_out[49] ^ layer2_out[50]);
    assign layer3_out[97] = ~layer2_out[167];
    assign layer3_out[98] = layer2_out[81];
    assign layer3_out[99] = ~layer2_out[158];
    assign layer3_out[100] = ~(layer2_out[75] & layer2_out[76]);
    assign layer3_out[101] = ~layer2_out[170];
    assign layer3_out[102] = layer2_out[147];
    assign layer3_out[103] = layer2_out[185] & ~layer2_out[184];
    assign layer3_out[104] = ~layer2_out[141] | layer2_out[142];
    assign layer3_out[105] = layer2_out[103] & ~layer2_out[104];
    assign layer3_out[106] = layer2_out[32];
    assign layer3_out[107] = layer2_out[59] & ~layer2_out[60];
    assign layer3_out[108] = layer2_out[191] & ~layer2_out[190];
    assign layer3_out[109] = ~layer2_out[99];
    assign layer3_out[110] = layer2_out[72];
    assign layer3_out[111] = layer2_out[94];
    assign layer3_out[112] = layer2_out[163] & layer2_out[164];
    assign layer3_out[113] = layer2_out[36] & ~layer2_out[37];
    assign layer3_out[114] = layer2_out[130];
    assign layer3_out[115] = ~layer2_out[76];
    assign layer3_out[116] = layer2_out[96];
    assign layer3_out[117] = ~(layer2_out[105] | layer2_out[106]);
    assign layer3_out[118] = layer2_out[79];
    assign layer3_out[119] = layer2_out[9] & ~layer2_out[10];
    assign layer3_out[120] = layer2_out[100];
    assign layer3_out[121] = layer2_out[38];
    assign layer3_out[122] = ~layer2_out[1];
    assign layer3_out[123] = ~layer2_out[110];
    assign layer3_out[124] = ~layer2_out[192];
    assign layer3_out[125] = ~(layer2_out[169] | layer2_out[170]);
    assign layer3_out[126] = layer2_out[83] & layer2_out[84];
    assign layer3_out[127] = layer2_out[85];
    assign layer3_out[128] = layer2_out[129];
    assign layer3_out[129] = layer2_out[179] ^ layer2_out[180];
    assign layer3_out[130] = ~layer2_out[5];
    assign layer3_out[131] = layer2_out[113];
    assign layer3_out[132] = layer2_out[6];
    assign layer3_out[133] = ~layer2_out[42];
    assign layer3_out[134] = ~layer2_out[40];
    assign layer3_out[135] = layer2_out[174] & ~layer2_out[173];
    assign layer3_out[136] = ~layer2_out[16];
    assign layer3_out[137] = layer2_out[34] & layer2_out[35];
    assign layer3_out[138] = layer2_out[148] & layer2_out[149];
    assign layer3_out[139] = ~layer2_out[152];
    assign layer3_out[140] = ~(layer2_out[24] & layer2_out[25]);
    assign layer3_out[141] = layer2_out[107] & layer2_out[108];
    assign layer3_out[142] = layer2_out[140];
    assign layer3_out[143] = layer2_out[45];
    assign layer3_out[144] = ~layer2_out[160];
    assign layer3_out[145] = ~(layer2_out[27] | layer2_out[28]);
    assign layer3_out[146] = ~(layer2_out[137] | layer2_out[138]);
    assign layer3_out[147] = layer2_out[156] & layer2_out[157];
    assign layer3_out[148] = ~layer2_out[94];
    assign layer3_out[149] = layer2_out[178] & ~layer2_out[179];
    assign layer3_out[150] = ~(layer2_out[72] | layer2_out[73]);
    assign layer3_out[151] = ~layer2_out[88];
    assign layer3_out[152] = layer2_out[165];
    assign layer3_out[153] = layer2_out[26];
    assign layer3_out[154] = layer2_out[3] & layer2_out[4];
    assign layer3_out[155] = ~(layer2_out[128] ^ layer2_out[129]);
    assign layer3_out[156] = ~layer2_out[151] | layer2_out[150];
    assign layer3_out[157] = ~layer2_out[12];
    assign layer3_out[158] = layer2_out[152] & ~layer2_out[153];
    assign layer3_out[159] = ~layer2_out[146];
    assign layer3_out[160] = ~layer2_out[131];
    assign layer3_out[161] = layer2_out[162] ^ layer2_out[163];
    assign layer3_out[162] = ~layer2_out[135];
    assign layer3_out[163] = layer2_out[29];
    assign layer3_out[164] = layer2_out[54] & ~layer2_out[55];
    assign layer3_out[165] = ~(layer2_out[149] | layer2_out[150]);
    assign layer3_out[166] = layer2_out[108] & layer2_out[109];
    assign layer3_out[167] = ~layer2_out[110];
    assign layer3_out[168] = layer2_out[92];
    assign layer3_out[169] = layer2_out[62] & ~layer2_out[63];
    assign layer3_out[170] = ~layer2_out[26];
    assign layer3_out[171] = layer2_out[69] & ~layer2_out[70];
    assign layer3_out[172] = layer2_out[8];
    assign layer3_out[173] = layer2_out[16];
    assign layer3_out[174] = layer2_out[196] & layer2_out[197];
    assign layer3_out[175] = ~layer2_out[188];
    assign layer3_out[176] = layer2_out[104];
    assign layer3_out[177] = layer2_out[81];
    assign layer3_out[178] = layer2_out[196];
    assign layer3_out[179] = ~layer2_out[47] | layer2_out[46];
    assign layer3_out[180] = ~(layer2_out[45] | layer2_out[46]);
    assign layer3_out[181] = layer2_out[172];
    assign layer3_out[182] = ~(layer2_out[182] | layer2_out[183]);
    assign layer3_out[183] = layer2_out[134];
    assign layer3_out[184] = layer2_out[187];
    assign layer3_out[185] = ~layer2_out[85];
    assign layer3_out[186] = ~layer2_out[119];
    assign layer3_out[187] = ~layer2_out[80];
    assign layer3_out[188] = ~layer2_out[161];
    assign layer3_out[189] = ~(layer2_out[30] | layer2_out[31]);
    assign layer3_out[190] = layer2_out[134];
    assign layer3_out[191] = ~layer2_out[54];
    assign layer3_out[192] = ~layer2_out[74];
    assign layer3_out[193] = ~(layer2_out[82] | layer2_out[83]);
    assign layer3_out[194] = layer2_out[19];
    assign layer3_out[195] = layer2_out[139] & ~layer2_out[138];
    assign layer3_out[196] = layer2_out[7];
    assign layer3_out[197] = layer2_out[176];
    assign layer3_out[198] = ~layer2_out[124];
    assign layer3_out[199] = layer2_out[57] & layer2_out[58];
      wire [199:0] last_layer_output;
      assign last_layer_output = layer3_out;
      wire [4:0] res [9:0];

      assign res[0] = last_layer_output[0] + last_layer_output[1] + last_layer_output[2] + last_layer_output[3] + last_layer_output[4] + last_layer_output[5] + last_layer_output[6] + last_layer_output[7] + last_layer_output[8] + last_layer_output[9] + last_layer_output[10] + last_layer_output[11] + last_layer_output[12] + last_layer_output[13] + last_layer_output[14] + last_layer_output[15] + last_layer_output[16] + last_layer_output[17] + last_layer_output[18] + last_layer_output[19];
      assign res[1] = last_layer_output[20] + last_layer_output[21] + last_layer_output[22] + last_layer_output[23] + last_layer_output[24] + last_layer_output[25] + last_layer_output[26] + last_layer_output[27] + last_layer_output[28] + last_layer_output[29] + last_layer_output[30] + last_layer_output[31] + last_layer_output[32] + last_layer_output[33] + last_layer_output[34] + last_layer_output[35] + last_layer_output[36] + last_layer_output[37] + last_layer_output[38] + last_layer_output[39];
      assign res[2] = last_layer_output[40] + last_layer_output[41] + last_layer_output[42] + last_layer_output[43] + last_layer_output[44] + last_layer_output[45] + last_layer_output[46] + last_layer_output[47] + last_layer_output[48] + last_layer_output[49] + last_layer_output[50] + last_layer_output[51] + last_layer_output[52] + last_layer_output[53] + last_layer_output[54] + last_layer_output[55] + last_layer_output[56] + last_layer_output[57] + last_layer_output[58] + last_layer_output[59];
      assign res[3] = last_layer_output[60] + last_layer_output[61] + last_layer_output[62] + last_layer_output[63] + last_layer_output[64] + last_layer_output[65] + last_layer_output[66] + last_layer_output[67] + last_layer_output[68] + last_layer_output[69] + last_layer_output[70] + last_layer_output[71] + last_layer_output[72] + last_layer_output[73] + last_layer_output[74] + last_layer_output[75] + last_layer_output[76] + last_layer_output[77] + last_layer_output[78] + last_layer_output[79];
      assign res[4] = last_layer_output[80] + last_layer_output[81] + last_layer_output[82] + last_layer_output[83] + last_layer_output[84] + last_layer_output[85] + last_layer_output[86] + last_layer_output[87] + last_layer_output[88] + last_layer_output[89] + last_layer_output[90] + last_layer_output[91] + last_layer_output[92] + last_layer_output[93] + last_layer_output[94] + last_layer_output[95] + last_layer_output[96] + last_layer_output[97] + last_layer_output[98] + last_layer_output[99];
      assign res[5] = last_layer_output[100] + last_layer_output[101] + last_layer_output[102] + last_layer_output[103] + last_layer_output[104] + last_layer_output[105] + last_layer_output[106] + last_layer_output[107] + last_layer_output[108] + last_layer_output[109] + last_layer_output[110] + last_layer_output[111] + last_layer_output[112] + last_layer_output[113] + last_layer_output[114] + last_layer_output[115] + last_layer_output[116] + last_layer_output[117] + last_layer_output[118] + last_layer_output[119];
      assign res[6] = last_layer_output[120] + last_layer_output[121] + last_layer_output[122] + last_layer_output[123] + last_layer_output[124] + last_layer_output[125] + last_layer_output[126] + last_layer_output[127] + last_layer_output[128] + last_layer_output[129] + last_layer_output[130] + last_layer_output[131] + last_layer_output[132] + last_layer_output[133] + last_layer_output[134] + last_layer_output[135] + last_layer_output[136] + last_layer_output[137] + last_layer_output[138] + last_layer_output[139];
      assign res[7] = last_layer_output[140] + last_layer_output[141] + last_layer_output[142] + last_layer_output[143] + last_layer_output[144] + last_layer_output[145] + last_layer_output[146] + last_layer_output[147] + last_layer_output[148] + last_layer_output[149] + last_layer_output[150] + last_layer_output[151] + last_layer_output[152] + last_layer_output[153] + last_layer_output[154] + last_layer_output[155] + last_layer_output[156] + last_layer_output[157] + last_layer_output[158] + last_layer_output[159];
      assign res[8] = last_layer_output[160] + last_layer_output[161] + last_layer_output[162] + last_layer_output[163] + last_layer_output[164] + last_layer_output[165] + last_layer_output[166] + last_layer_output[167] + last_layer_output[168] + last_layer_output[169] + last_layer_output[170] + last_layer_output[171] + last_layer_output[172] + last_layer_output[173] + last_layer_output[174] + last_layer_output[175] + last_layer_output[176] + last_layer_output[177] + last_layer_output[178] + last_layer_output[179];
      assign res[9] = last_layer_output[180] + last_layer_output[181] + last_layer_output[182] + last_layer_output[183] + last_layer_output[184] + last_layer_output[185] + last_layer_output[186] + last_layer_output[187] + last_layer_output[188] + last_layer_output[189] + last_layer_output[190] + last_layer_output[191] + last_layer_output[192] + last_layer_output[193] + last_layer_output[194] + last_layer_output[195] + last_layer_output[196] + last_layer_output[197] + last_layer_output[198] + last_layer_output[199];
      assign y[49:45]=res[0];
      assign y[44:40]=res[1];
      assign y[39:35]=res[2];
      assign y[34:30]=res[3];
      assign y[29:25]=res[4];
      assign y[24:20]=res[5];
      assign y[19:15]=res[6];
      assign y[14:10]=res[7];
      assign y[9:5]=res[8];
      assign y[4:0]=res[9];
endmodule
