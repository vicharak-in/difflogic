module logic_network (    input wire [399:0] x,
    output wire [69:0] y
);
      wire [799:0] layer0_out;
      wire [799:0] layer1_out;
      wire [799:0] layer2_out;
      wire [799:0] layer3_out;
    assign layer0_out[0] = ~x[354];
    assign layer0_out[1] = ~(x[300] | x[302]);
    assign layer0_out[2] = ~(x[258] | x[259]);
    assign layer0_out[3] = x[6] | x[7];
    assign layer0_out[4] = ~(x[22] | x[24]);
    assign layer0_out[5] = ~x[41];
    assign layer0_out[6] = x[125] | x[127];
    assign layer0_out[7] = x[372] & x[374];
    assign layer0_out[8] = x[357];
    assign layer0_out[9] = ~x[7] | x[8];
    assign layer0_out[10] = 1'b1;
    assign layer0_out[11] = 1'b0;
    assign layer0_out[12] = ~(x[159] | x[161]);
    assign layer0_out[13] = ~x[73];
    assign layer0_out[14] = x[124] | x[125];
    assign layer0_out[15] = ~(x[304] | x[305]);
    assign layer0_out[16] = 1'b0;
    assign layer0_out[17] = ~x[163] | x[165];
    assign layer0_out[18] = ~x[313];
    assign layer0_out[19] = ~x[164] | x[165];
    assign layer0_out[20] = x[185] | x[187];
    assign layer0_out[21] = 1'b1;
    assign layer0_out[22] = ~x[252];
    assign layer0_out[23] = x[133] | x[134];
    assign layer0_out[24] = x[269] | x[270];
    assign layer0_out[25] = 1'b0;
    assign layer0_out[26] = x[285] | x[287];
    assign layer0_out[27] = x[166] & ~x[168];
    assign layer0_out[28] = x[172];
    assign layer0_out[29] = ~(x[148] | x[149]);
    assign layer0_out[30] = x[111] | x[113];
    assign layer0_out[31] = 1'b0;
    assign layer0_out[32] = x[311] | x[313];
    assign layer0_out[33] = ~(x[220] | x[222]);
    assign layer0_out[34] = 1'b1;
    assign layer0_out[35] = x[313] | x[315];
    assign layer0_out[36] = x[221] & ~x[223];
    assign layer0_out[37] = ~(x[270] | x[271]);
    assign layer0_out[38] = x[259] ^ x[261];
    assign layer0_out[39] = ~x[187];
    assign layer0_out[40] = x[89] ^ x[91];
    assign layer0_out[41] = ~(x[359] | x[361]);
    assign layer0_out[42] = x[360];
    assign layer0_out[43] = x[308];
    assign layer0_out[44] = x[221] | x[222];
    assign layer0_out[45] = ~x[300] | x[301];
    assign layer0_out[46] = x[73] | x[74];
    assign layer0_out[47] = x[208];
    assign layer0_out[48] = x[90];
    assign layer0_out[49] = x[10] | x[12];
    assign layer0_out[50] = ~(x[40] | x[42]);
    assign layer0_out[51] = 1'b0;
    assign layer0_out[52] = ~x[280] | x[279];
    assign layer0_out[53] = x[170];
    assign layer0_out[54] = ~(x[358] | x[359]);
    assign layer0_out[55] = ~x[51];
    assign layer0_out[56] = ~x[287] | x[289];
    assign layer0_out[57] = x[364];
    assign layer0_out[58] = x[177] | x[179];
    assign layer0_out[59] = ~(x[137] | x[139]);
    assign layer0_out[60] = 1'b1;
    assign layer0_out[61] = x[256] | x[258];
    assign layer0_out[62] = x[82] | x[84];
    assign layer0_out[63] = x[340] & ~x[339];
    assign layer0_out[64] = 1'b0;
    assign layer0_out[65] = ~x[395] | x[393];
    assign layer0_out[66] = x[287] | x[288];
    assign layer0_out[67] = x[179] & x[180];
    assign layer0_out[68] = x[394] | x[395];
    assign layer0_out[69] = x[323] | x[324];
    assign layer0_out[70] = x[264] | x[265];
    assign layer0_out[71] = ~(x[343] | x[344]);
    assign layer0_out[72] = ~(x[32] & x[34]);
    assign layer0_out[73] = ~x[229];
    assign layer0_out[74] = ~(x[20] & x[21]);
    assign layer0_out[75] = x[269] & ~x[268];
    assign layer0_out[76] = ~(x[242] | x[243]);
    assign layer0_out[77] = ~x[157] | x[156];
    assign layer0_out[78] = x[331];
    assign layer0_out[79] = ~(x[136] | x[138]);
    assign layer0_out[80] = ~(x[284] | x[285]);
    assign layer0_out[81] = 1'b0;
    assign layer0_out[82] = x[183] | x[184];
    assign layer0_out[83] = ~(x[152] | x[154]);
    assign layer0_out[84] = ~x[80];
    assign layer0_out[85] = ~(x[157] | x[158]);
    assign layer0_out[86] = ~x[91];
    assign layer0_out[87] = ~(x[199] | x[200]);
    assign layer0_out[88] = 1'b0;
    assign layer0_out[89] = ~(x[66] ^ x[68]);
    assign layer0_out[90] = 1'b1;
    assign layer0_out[91] = ~(x[47] | x[48]);
    assign layer0_out[92] = x[228];
    assign layer0_out[93] = ~x[201];
    assign layer0_out[94] = ~x[390];
    assign layer0_out[95] = x[186];
    assign layer0_out[96] = ~x[39];
    assign layer0_out[97] = x[333] | x[334];
    assign layer0_out[98] = ~x[248] | x[247];
    assign layer0_out[99] = ~(x[331] | x[332]);
    assign layer0_out[100] = x[112] | x[113];
    assign layer0_out[101] = 1'b0;
    assign layer0_out[102] = x[266] | x[268];
    assign layer0_out[103] = 1'b1;
    assign layer0_out[104] = ~x[176] | x[175];
    assign layer0_out[105] = 1'b0;
    assign layer0_out[106] = ~x[149];
    assign layer0_out[107] = ~x[25];
    assign layer0_out[108] = ~(x[248] | x[249]);
    assign layer0_out[109] = x[98] | x[99];
    assign layer0_out[110] = ~(x[188] & x[190]);
    assign layer0_out[111] = x[155] | x[156];
    assign layer0_out[112] = ~(x[143] | x[145]);
    assign layer0_out[113] = x[107] | x[108];
    assign layer0_out[114] = 1'b0;
    assign layer0_out[115] = ~(x[143] | x[144]);
    assign layer0_out[116] = x[388];
    assign layer0_out[117] = ~(x[274] | x[276]);
    assign layer0_out[118] = x[161];
    assign layer0_out[119] = x[243] | x[244];
    assign layer0_out[120] = ~x[333];
    assign layer0_out[121] = ~x[69] | x[71];
    assign layer0_out[122] = x[103] | x[104];
    assign layer0_out[123] = ~(x[116] | x[118]);
    assign layer0_out[124] = ~(x[229] | x[230]);
    assign layer0_out[125] = x[156] | x[158];
    assign layer0_out[126] = ~(x[51] & x[52]);
    assign layer0_out[127] = x[42] | x[44];
    assign layer0_out[128] = x[84] | x[86];
    assign layer0_out[129] = x[44] | x[45];
    assign layer0_out[130] = x[210] | x[211];
    assign layer0_out[131] = x[245];
    assign layer0_out[132] = ~x[241];
    assign layer0_out[133] = x[17] & ~x[15];
    assign layer0_out[134] = ~(x[305] | x[306]);
    assign layer0_out[135] = x[79] & ~x[78];
    assign layer0_out[136] = 1'b1;
    assign layer0_out[137] = x[1] & x[2];
    assign layer0_out[138] = x[209] | x[210];
    assign layer0_out[139] = ~x[152];
    assign layer0_out[140] = 1'b1;
    assign layer0_out[141] = x[115] | x[116];
    assign layer0_out[142] = ~x[46];
    assign layer0_out[143] = x[170] | x[171];
    assign layer0_out[144] = 1'b1;
    assign layer0_out[145] = x[171];
    assign layer0_out[146] = ~x[29] | x[30];
    assign layer0_out[147] = ~(x[204] | x[205]);
    assign layer0_out[148] = 1'b1;
    assign layer0_out[149] = x[389];
    assign layer0_out[150] = x[110];
    assign layer0_out[151] = ~x[178];
    assign layer0_out[152] = ~(x[255] | x[256]);
    assign layer0_out[153] = ~x[16] | x[14];
    assign layer0_out[154] = x[162] | x[163];
    assign layer0_out[155] = x[214];
    assign layer0_out[156] = ~x[187];
    assign layer0_out[157] = ~(x[317] | x[319]);
    assign layer0_out[158] = x[230];
    assign layer0_out[159] = x[381] & x[383];
    assign layer0_out[160] = 1'b0;
    assign layer0_out[161] = ~(x[342] & x[344]);
    assign layer0_out[162] = ~(x[307] & x[308]);
    assign layer0_out[163] = 1'b1;
    assign layer0_out[164] = ~(x[39] & x[41]);
    assign layer0_out[165] = ~(x[256] | x[257]);
    assign layer0_out[166] = ~(x[358] | x[360]);
    assign layer0_out[167] = 1'b0;
    assign layer0_out[168] = ~(x[284] | x[286]);
    assign layer0_out[169] = x[282] | x[284];
    assign layer0_out[170] = x[190] | x[191];
    assign layer0_out[171] = x[397] | x[399];
    assign layer0_out[172] = ~(x[283] | x[284]);
    assign layer0_out[173] = x[345] | x[347];
    assign layer0_out[174] = ~x[158];
    assign layer0_out[175] = ~(x[39] | x[40]);
    assign layer0_out[176] = x[348] | x[349];
    assign layer0_out[177] = 1'b0;
    assign layer0_out[178] = x[104] | x[106];
    assign layer0_out[179] = x[43];
    assign layer0_out[180] = x[303] | x[305];
    assign layer0_out[181] = ~x[56];
    assign layer0_out[182] = 1'b0;
    assign layer0_out[183] = x[100] & ~x[101];
    assign layer0_out[184] = ~(x[87] | x[88]);
    assign layer0_out[185] = 1'b1;
    assign layer0_out[186] = ~x[118];
    assign layer0_out[187] = ~x[278];
    assign layer0_out[188] = ~(x[254] | x[255]);
    assign layer0_out[189] = x[59] | x[61];
    assign layer0_out[190] = ~(x[124] | x[126]);
    assign layer0_out[191] = ~(x[347] & x[349]);
    assign layer0_out[192] = 1'b1;
    assign layer0_out[193] = ~(x[288] | x[289]);
    assign layer0_out[194] = ~(x[153] | x[155]);
    assign layer0_out[195] = x[373] & ~x[372];
    assign layer0_out[196] = ~(x[328] & x[330]);
    assign layer0_out[197] = x[356] | x[357];
    assign layer0_out[198] = x[132] | x[134];
    assign layer0_out[199] = x[126];
    assign layer0_out[200] = x[23] | x[24];
    assign layer0_out[201] = x[138] | x[139];
    assign layer0_out[202] = ~x[100] | x[102];
    assign layer0_out[203] = x[82];
    assign layer0_out[204] = ~x[329];
    assign layer0_out[205] = x[93] & x[95];
    assign layer0_out[206] = ~(x[115] | x[117]);
    assign layer0_out[207] = ~(x[5] | x[6]);
    assign layer0_out[208] = ~(x[71] ^ x[72]);
    assign layer0_out[209] = x[87];
    assign layer0_out[210] = ~(x[210] | x[212]);
    assign layer0_out[211] = ~(x[0] | x[1]);
    assign layer0_out[212] = x[23];
    assign layer0_out[213] = x[353] | x[354];
    assign layer0_out[214] = x[385] | x[387];
    assign layer0_out[215] = ~x[109];
    assign layer0_out[216] = ~x[218];
    assign layer0_out[217] = ~x[386];
    assign layer0_out[218] = ~x[141];
    assign layer0_out[219] = x[202] | x[204];
    assign layer0_out[220] = x[378];
    assign layer0_out[221] = ~x[397] | x[395];
    assign layer0_out[222] = x[64] ^ x[66];
    assign layer0_out[223] = ~(x[8] | x[10]);
    assign layer0_out[224] = ~(x[27] & x[29]);
    assign layer0_out[225] = ~(x[239] | x[240]);
    assign layer0_out[226] = x[31];
    assign layer0_out[227] = x[268] & x[270];
    assign layer0_out[228] = x[301] | x[302];
    assign layer0_out[229] = x[189];
    assign layer0_out[230] = 1'b0;
    assign layer0_out[231] = x[307];
    assign layer0_out[232] = 1'b1;
    assign layer0_out[233] = x[28];
    assign layer0_out[234] = x[244] | x[246];
    assign layer0_out[235] = ~(x[267] | x[269]);
    assign layer0_out[236] = 1'b1;
    assign layer0_out[237] = x[181] | x[182];
    assign layer0_out[238] = ~(x[53] & x[54]);
    assign layer0_out[239] = ~x[384];
    assign layer0_out[240] = ~(x[103] | x[105]);
    assign layer0_out[241] = ~(x[166] | x[167]);
    assign layer0_out[242] = x[359] & ~x[360];
    assign layer0_out[243] = ~(x[28] | x[29]);
    assign layer0_out[244] = ~(x[223] | x[224]);
    assign layer0_out[245] = ~(x[112] ^ x[114]);
    assign layer0_out[246] = x[241] | x[243];
    assign layer0_out[247] = ~(x[17] ^ x[18]);
    assign layer0_out[248] = ~x[92] | x[94];
    assign layer0_out[249] = ~(x[114] | x[116]);
    assign layer0_out[250] = x[117] | x[119];
    assign layer0_out[251] = x[203];
    assign layer0_out[252] = x[315] & x[317];
    assign layer0_out[253] = ~x[42];
    assign layer0_out[254] = ~(x[346] | x[348]);
    assign layer0_out[255] = 1'b0;
    assign layer0_out[256] = ~x[220];
    assign layer0_out[257] = x[75] | x[76];
    assign layer0_out[258] = x[182] | x[184];
    assign layer0_out[259] = 1'b0;
    assign layer0_out[260] = x[70] & ~x[71];
    assign layer0_out[261] = x[218] & ~x[216];
    assign layer0_out[262] = ~(x[152] | x[153]);
    assign layer0_out[263] = x[376] ^ x[378];
    assign layer0_out[264] = ~(x[324] | x[325]);
    assign layer0_out[265] = 1'b0;
    assign layer0_out[266] = x[334] | x[336];
    assign layer0_out[267] = ~x[273] | x[272];
    assign layer0_out[268] = ~(x[362] | x[363]);
    assign layer0_out[269] = ~x[52];
    assign layer0_out[270] = ~(x[206] | x[207]);
    assign layer0_out[271] = x[62] & x[63];
    assign layer0_out[272] = x[13] & ~x[15];
    assign layer0_out[273] = x[302] | x[303];
    assign layer0_out[274] = 1'b1;
    assign layer0_out[275] = 1'b0;
    assign layer0_out[276] = ~x[83];
    assign layer0_out[277] = ~(x[88] ^ x[90]);
    assign layer0_out[278] = ~x[49];
    assign layer0_out[279] = x[80];
    assign layer0_out[280] = x[379] & ~x[380];
    assign layer0_out[281] = x[204] | x[206];
    assign layer0_out[282] = x[165] | x[167];
    assign layer0_out[283] = 1'b0;
    assign layer0_out[284] = ~(x[389] | x[391]);
    assign layer0_out[285] = ~x[63];
    assign layer0_out[286] = ~(x[44] | x[46]);
    assign layer0_out[287] = ~(x[109] | x[111]);
    assign layer0_out[288] = ~(x[298] | x[300]);
    assign layer0_out[289] = x[253] & ~x[251];
    assign layer0_out[290] = ~(x[160] | x[162]);
    assign layer0_out[291] = x[76] & ~x[77];
    assign layer0_out[292] = x[311] | x[312];
    assign layer0_out[293] = x[192] & x[193];
    assign layer0_out[294] = ~(x[165] | x[166]);
    assign layer0_out[295] = x[232] | x[234];
    assign layer0_out[296] = x[133] | x[135];
    assign layer0_out[297] = x[94] & x[95];
    assign layer0_out[298] = x[147];
    assign layer0_out[299] = 1'b0;
    assign layer0_out[300] = ~x[208];
    assign layer0_out[301] = ~x[209];
    assign layer0_out[302] = x[379] ^ x[381];
    assign layer0_out[303] = x[35] | x[36];
    assign layer0_out[304] = ~(x[154] | x[155]);
    assign layer0_out[305] = ~x[147];
    assign layer0_out[306] = ~(x[367] | x[369]);
    assign layer0_out[307] = ~(x[352] | x[353]);
    assign layer0_out[308] = ~x[106];
    assign layer0_out[309] = x[110] | x[112];
    assign layer0_out[310] = x[309] ^ x[311];
    assign layer0_out[311] = x[90] | x[92];
    assign layer0_out[312] = x[364];
    assign layer0_out[313] = 1'b0;
    assign layer0_out[314] = ~(x[31] & x[32]);
    assign layer0_out[315] = ~(x[295] | x[296]);
    assign layer0_out[316] = x[262] | x[264];
    assign layer0_out[317] = 1'b1;
    assign layer0_out[318] = ~(x[140] | x[141]);
    assign layer0_out[319] = ~(x[45] | x[47]);
    assign layer0_out[320] = ~(x[16] | x[17]);
    assign layer0_out[321] = x[181] | x[183];
    assign layer0_out[322] = x[104];
    assign layer0_out[323] = 1'b0;
    assign layer0_out[324] = ~x[106] | x[105];
    assign layer0_out[325] = ~(x[324] | x[326]);
    assign layer0_out[326] = 1'b1;
    assign layer0_out[327] = 1'b1;
    assign layer0_out[328] = x[365] | x[366];
    assign layer0_out[329] = ~x[352];
    assign layer0_out[330] = x[179] & x[181];
    assign layer0_out[331] = ~x[328];
    assign layer0_out[332] = x[264] | x[266];
    assign layer0_out[333] = ~(x[202] | x[203]);
    assign layer0_out[334] = ~(x[198] | x[200]);
    assign layer0_out[335] = ~(x[195] | x[197]);
    assign layer0_out[336] = ~(x[385] | x[386]);
    assign layer0_out[337] = x[101] & x[103];
    assign layer0_out[338] = x[249] | x[251];
    assign layer0_out[339] = ~(x[81] | x[82]);
    assign layer0_out[340] = x[76] | x[78];
    assign layer0_out[341] = ~(x[318] ^ x[320]);
    assign layer0_out[342] = x[52] | x[54];
    assign layer0_out[343] = x[94] | x[96];
    assign layer0_out[344] = ~x[342] | x[343];
    assign layer0_out[345] = ~(x[96] | x[98]);
    assign layer0_out[346] = 1'b0;
    assign layer0_out[347] = ~(x[363] | x[364]);
    assign layer0_out[348] = x[240];
    assign layer0_out[349] = x[176] | x[177];
    assign layer0_out[350] = ~(x[334] | x[335]);
    assign layer0_out[351] = x[72];
    assign layer0_out[352] = 1'b1;
    assign layer0_out[353] = x[62] | x[64];
    assign layer0_out[354] = ~x[387];
    assign layer0_out[355] = ~(x[285] | x[286]);
    assign layer0_out[356] = ~x[360] | x[361];
    assign layer0_out[357] = ~(x[377] | x[378]);
    assign layer0_out[358] = x[164] | x[166];
    assign layer0_out[359] = x[344] | x[345];
    assign layer0_out[360] = x[180] & ~x[182];
    assign layer0_out[361] = ~(x[250] & x[251]);
    assign layer0_out[362] = x[51] & x[53];
    assign layer0_out[363] = x[277] | x[279];
    assign layer0_out[364] = x[254] | x[256];
    assign layer0_out[365] = ~x[120] | x[122];
    assign layer0_out[366] = ~x[13];
    assign layer0_out[367] = x[0] | x[3];
    assign layer0_out[368] = ~(x[95] | x[97]);
    assign layer0_out[369] = 1'b0;
    assign layer0_out[370] = ~x[282] | x[280];
    assign layer0_out[371] = ~(x[203] | x[204]);
    assign layer0_out[372] = ~(x[292] | x[293]);
    assign layer0_out[373] = ~(x[86] | x[87]);
    assign layer0_out[374] = x[142] | x[143];
    assign layer0_out[375] = x[58] & ~x[57];
    assign layer0_out[376] = x[255] | x[257];
    assign layer0_out[377] = ~(x[393] | x[394]);
    assign layer0_out[378] = 1'b1;
    assign layer0_out[379] = x[167] | x[169];
    assign layer0_out[380] = 1'b0;
    assign layer0_out[381] = 1'b0;
    assign layer0_out[382] = x[224] | x[225];
    assign layer0_out[383] = x[398];
    assign layer0_out[384] = ~(x[10] | x[11]);
    assign layer0_out[385] = ~(x[184] | x[186]);
    assign layer0_out[386] = ~x[148];
    assign layer0_out[387] = ~x[67];
    assign layer0_out[388] = x[12] & x[14];
    assign layer0_out[389] = x[68] & ~x[69];
    assign layer0_out[390] = x[35] & ~x[34];
    assign layer0_out[391] = x[18] | x[19];
    assign layer0_out[392] = x[283] | x[285];
    assign layer0_out[393] = x[126] | x[127];
    assign layer0_out[394] = ~(x[41] | x[42]);
    assign layer0_out[395] = ~x[80] | x[79];
    assign layer0_out[396] = 1'b0;
    assign layer0_out[397] = 1'b1;
    assign layer0_out[398] = x[212] | x[214];
    assign layer0_out[399] = x[63] | x[65];
    assign layer0_out[400] = 1'b1;
    assign layer0_out[401] = ~x[287];
    assign layer0_out[402] = ~(x[228] | x[229]);
    assign layer0_out[403] = x[104] | x[105];
    assign layer0_out[404] = ~x[278];
    assign layer0_out[405] = ~x[119] | x[118];
    assign layer0_out[406] = x[343] | x[345];
    assign layer0_out[407] = ~x[215];
    assign layer0_out[408] = ~(x[185] | x[186]);
    assign layer0_out[409] = ~x[120] | x[121];
    assign layer0_out[410] = ~(x[309] & x[310]);
    assign layer0_out[411] = x[263] | x[265];
    assign layer0_out[412] = ~x[192];
    assign layer0_out[413] = 1'b0;
    assign layer0_out[414] = ~x[290];
    assign layer0_out[415] = x[346] | x[347];
    assign layer0_out[416] = ~(x[45] & x[46]);
    assign layer0_out[417] = x[171] | x[172];
    assign layer0_out[418] = ~(x[318] & x[319]);
    assign layer0_out[419] = ~(x[49] | x[50]);
    assign layer0_out[420] = ~(x[167] | x[168]);
    assign layer0_out[421] = x[171];
    assign layer0_out[422] = 1'b1;
    assign layer0_out[423] = ~(x[388] | x[390]);
    assign layer0_out[424] = x[233];
    assign layer0_out[425] = 1'b1;
    assign layer0_out[426] = ~x[243];
    assign layer0_out[427] = ~(x[351] | x[353]);
    assign layer0_out[428] = 1'b1;
    assign layer0_out[429] = ~x[127];
    assign layer0_out[430] = ~(x[19] ^ x[20]);
    assign layer0_out[431] = ~(x[336] | x[338]);
    assign layer0_out[432] = ~x[59] | x[60];
    assign layer0_out[433] = ~(x[17] | x[19]);
    assign layer0_out[434] = ~(x[315] | x[316]);
    assign layer0_out[435] = x[259] | x[260];
    assign layer0_out[436] = ~x[136] | x[135];
    assign layer0_out[437] = ~(x[46] | x[48]);
    assign layer0_out[438] = 1'b0;
    assign layer0_out[439] = x[319] | x[320];
    assign layer0_out[440] = ~(x[333] | x[335]);
    assign layer0_out[441] = 1'b0;
    assign layer0_out[442] = x[387] | x[388];
    assign layer0_out[443] = x[341];
    assign layer0_out[444] = ~(x[226] | x[228]);
    assign layer0_out[445] = 1'b1;
    assign layer0_out[446] = ~(x[262] | x[263]);
    assign layer0_out[447] = x[85] & x[86];
    assign layer0_out[448] = ~(x[61] | x[62]);
    assign layer0_out[449] = ~(x[325] | x[326]);
    assign layer0_out[450] = ~x[351];
    assign layer0_out[451] = 1'b1;
    assign layer0_out[452] = ~(x[351] | x[352]);
    assign layer0_out[453] = x[263] | x[264];
    assign layer0_out[454] = x[361] & ~x[362];
    assign layer0_out[455] = ~(x[183] | x[185]);
    assign layer0_out[456] = ~(x[0] ^ x[2]);
    assign layer0_out[457] = ~x[90];
    assign layer0_out[458] = x[302] | x[304];
    assign layer0_out[459] = x[195];
    assign layer0_out[460] = ~x[233];
    assign layer0_out[461] = x[208] | x[209];
    assign layer0_out[462] = 1'b0;
    assign layer0_out[463] = x[53];
    assign layer0_out[464] = x[168];
    assign layer0_out[465] = ~x[66] | x[65];
    assign layer0_out[466] = x[121] | x[123];
    assign layer0_out[467] = x[299] ^ x[300];
    assign layer0_out[468] = ~(x[236] | x[238]);
    assign layer0_out[469] = x[381] & ~x[380];
    assign layer0_out[470] = ~(x[296] | x[298]);
    assign layer0_out[471] = ~(x[74] | x[75]);
    assign layer0_out[472] = 1'b0;
    assign layer0_out[473] = ~(x[345] | x[346]);
    assign layer0_out[474] = x[213] & ~x[215];
    assign layer0_out[475] = x[99] | x[100];
    assign layer0_out[476] = x[367];
    assign layer0_out[477] = x[56] | x[58];
    assign layer0_out[478] = 1'b0;
    assign layer0_out[479] = x[237] & ~x[236];
    assign layer0_out[480] = ~x[59];
    assign layer0_out[481] = x[136] | x[137];
    assign layer0_out[482] = ~x[38];
    assign layer0_out[483] = x[238] | x[239];
    assign layer0_out[484] = ~x[368];
    assign layer0_out[485] = ~(x[335] | x[337]);
    assign layer0_out[486] = x[155] | x[157];
    assign layer0_out[487] = 1'b0;
    assign layer0_out[488] = x[89] & ~x[88];
    assign layer0_out[489] = 1'b1;
    assign layer0_out[490] = x[193] ^ x[195];
    assign layer0_out[491] = x[2] ^ x[5];
    assign layer0_out[492] = ~x[340];
    assign layer0_out[493] = x[172];
    assign layer0_out[494] = x[276] | x[278];
    assign layer0_out[495] = x[316] | x[317];
    assign layer0_out[496] = ~x[117] | x[116];
    assign layer0_out[497] = ~(x[97] & x[99]);
    assign layer0_out[498] = x[368] | x[369];
    assign layer0_out[499] = ~(x[97] | x[98]);
    assign layer0_out[500] = ~(x[312] & x[314]);
    assign layer0_out[501] = ~(x[36] | x[38]);
    assign layer0_out[502] = x[213] & ~x[211];
    assign layer0_out[503] = x[349] & x[351];
    assign layer0_out[504] = ~(x[261] | x[263]);
    assign layer0_out[505] = x[150];
    assign layer0_out[506] = ~x[25];
    assign layer0_out[507] = ~(x[316] | x[318]);
    assign layer0_out[508] = x[225] & ~x[226];
    assign layer0_out[509] = ~(x[289] & x[291]);
    assign layer0_out[510] = x[149];
    assign layer0_out[511] = x[144] | x[145];
    assign layer0_out[512] = x[251] & ~x[252];
    assign layer0_out[513] = ~(x[257] | x[259]);
    assign layer0_out[514] = x[222] | x[223];
    assign layer0_out[515] = x[95] | x[96];
    assign layer0_out[516] = x[170] | x[172];
    assign layer0_out[517] = ~x[70] | x[69];
    assign layer0_out[518] = ~(x[261] | x[262]);
    assign layer0_out[519] = ~(x[18] | x[20]);
    assign layer0_out[520] = ~x[355];
    assign layer0_out[521] = ~(x[131] ^ x[132]);
    assign layer0_out[522] = x[140] & ~x[138];
    assign layer0_out[523] = 1'b1;
    assign layer0_out[524] = ~(x[266] | x[267]);
    assign layer0_out[525] = 1'b1;
    assign layer0_out[526] = ~x[367];
    assign layer0_out[527] = ~(x[119] ^ x[121]);
    assign layer0_out[528] = ~(x[274] | x[275]);
    assign layer0_out[529] = ~x[392] | x[390];
    assign layer0_out[530] = ~x[133] | x[131];
    assign layer0_out[531] = 1'b0;
    assign layer0_out[532] = 1'b0;
    assign layer0_out[533] = ~(x[361] | x[363]);
    assign layer0_out[534] = x[348];
    assign layer0_out[535] = ~x[170] | x[168];
    assign layer0_out[536] = 1'b0;
    assign layer0_out[537] = 1'b1;
    assign layer0_out[538] = x[150];
    assign layer0_out[539] = x[275] & ~x[273];
    assign layer0_out[540] = x[126];
    assign layer0_out[541] = 1'b1;
    assign layer0_out[542] = 1'b1;
    assign layer0_out[543] = x[161] | x[163];
    assign layer0_out[544] = x[161] | x[162];
    assign layer0_out[545] = 1'b0;
    assign layer0_out[546] = ~x[321];
    assign layer0_out[547] = x[8] | x[9];
    assign layer0_out[548] = 1'b1;
    assign layer0_out[549] = ~(x[75] | x[77]);
    assign layer0_out[550] = ~x[64] | x[65];
    assign layer0_out[551] = ~(x[218] | x[220]);
    assign layer0_out[552] = ~x[128];
    assign layer0_out[553] = 1'b0;
    assign layer0_out[554] = ~x[369];
    assign layer0_out[555] = ~(x[48] & x[50]);
    assign layer0_out[556] = ~(x[194] | x[196]);
    assign layer0_out[557] = x[322] | x[324];
    assign layer0_out[558] = ~(x[113] | x[115]);
    assign layer0_out[559] = x[325] | x[327];
    assign layer0_out[560] = x[24];
    assign layer0_out[561] = ~x[70];
    assign layer0_out[562] = x[114] | x[115];
    assign layer0_out[563] = 1'b1;
    assign layer0_out[564] = x[246] | x[247];
    assign layer0_out[565] = x[3] | x[5];
    assign layer0_out[566] = ~x[181];
    assign layer0_out[567] = x[105] | x[107];
    assign layer0_out[568] = ~x[299];
    assign layer0_out[569] = ~x[354];
    assign layer0_out[570] = x[11];
    assign layer0_out[571] = x[340] | x[342];
    assign layer0_out[572] = x[317] | x[318];
    assign layer0_out[573] = x[20] | x[22];
    assign layer0_out[574] = ~(x[220] | x[221]);
    assign layer0_out[575] = 1'b1;
    assign layer0_out[576] = x[73] | x[75];
    assign layer0_out[577] = x[346] & ~x[344];
    assign layer0_out[578] = ~x[311];
    assign layer0_out[579] = ~x[43];
    assign layer0_out[580] = ~x[271];
    assign layer0_out[581] = x[173] | x[174];
    assign layer0_out[582] = x[216] & ~x[214];
    assign layer0_out[583] = ~(x[147] | x[148]);
    assign layer0_out[584] = x[306] | x[307];
    assign layer0_out[585] = ~(x[154] | x[156]);
    assign layer0_out[586] = x[159] & ~x[158];
    assign layer0_out[587] = x[4] | x[6];
    assign layer0_out[588] = ~(x[25] | x[27]);
    assign layer0_out[589] = x[189];
    assign layer0_out[590] = ~(x[209] | x[211]);
    assign layer0_out[591] = x[2] | x[4];
    assign layer0_out[592] = x[240] & x[242];
    assign layer0_out[593] = x[367];
    assign layer0_out[594] = ~(x[275] | x[277]);
    assign layer0_out[595] = ~x[1];
    assign layer0_out[596] = ~(x[227] | x[229]);
    assign layer0_out[597] = x[122] | x[124];
    assign layer0_out[598] = 1'b1;
    assign layer0_out[599] = x[255] & ~x[253];
    assign layer0_out[600] = ~x[26];
    assign layer0_out[601] = x[21] & ~x[19];
    assign layer0_out[602] = x[341] & ~x[342];
    assign layer0_out[603] = ~x[213];
    assign layer0_out[604] = x[391];
    assign layer0_out[605] = ~x[122];
    assign layer0_out[606] = x[352] | x[354];
    assign layer0_out[607] = x[339];
    assign layer0_out[608] = x[223] | x[225];
    assign layer0_out[609] = ~(x[217] | x[219]);
    assign layer0_out[610] = x[129] | x[131];
    assign layer0_out[611] = ~x[97];
    assign layer0_out[612] = x[230] | x[232];
    assign layer0_out[613] = 1'b1;
    assign layer0_out[614] = 1'b0;
    assign layer0_out[615] = x[288] | x[290];
    assign layer0_out[616] = x[337] | x[339];
    assign layer0_out[617] = ~(x[14] | x[15]);
    assign layer0_out[618] = ~(x[175] | x[177]);
    assign layer0_out[619] = x[357] | x[358];
    assign layer0_out[620] = ~x[198];
    assign layer0_out[621] = ~(x[293] | x[294]);
    assign layer0_out[622] = ~(x[396] | x[397]);
    assign layer0_out[623] = x[86];
    assign layer0_out[624] = x[84];
    assign layer0_out[625] = ~x[370];
    assign layer0_out[626] = x[267] | x[268];
    assign layer0_out[627] = 1'b1;
    assign layer0_out[628] = ~(x[349] | x[350]);
    assign layer0_out[629] = ~(x[24] | x[26]);
    assign layer0_out[630] = ~x[274];
    assign layer0_out[631] = ~x[62];
    assign layer0_out[632] = ~(x[58] | x[59]);
    assign layer0_out[633] = ~(x[196] | x[197]);
    assign layer0_out[634] = ~x[378] | x[379];
    assign layer0_out[635] = ~(x[150] | x[151]);
    assign layer0_out[636] = ~(x[242] | x[244]);
    assign layer0_out[637] = x[159] & ~x[160];
    assign layer0_out[638] = ~x[379] | x[377];
    assign layer0_out[639] = ~(x[321] | x[323]);
    assign layer0_out[640] = x[218] | x[219];
    assign layer0_out[641] = x[163] | x[164];
    assign layer0_out[642] = x[234] | x[235];
    assign layer0_out[643] = x[91] ^ x[93];
    assign layer0_out[644] = x[134] | x[135];
    assign layer0_out[645] = x[60] | x[61];
    assign layer0_out[646] = x[308] | x[309];
    assign layer0_out[647] = x[140];
    assign layer0_out[648] = ~(x[26] | x[28]);
    assign layer0_out[649] = ~(x[193] | x[194]);
    assign layer0_out[650] = ~x[33];
    assign layer0_out[651] = x[224] | x[226];
    assign layer0_out[652] = x[338] | x[339];
    assign layer0_out[653] = x[265] | x[266];
    assign layer0_out[654] = x[364];
    assign layer0_out[655] = x[390];
    assign layer0_out[656] = ~(x[21] | x[22]);
    assign layer0_out[657] = ~x[77];
    assign layer0_out[658] = ~(x[332] & x[334]);
    assign layer0_out[659] = ~(x[203] | x[205]);
    assign layer0_out[660] = x[4] | x[5];
    assign layer0_out[661] = x[270] | x[272];
    assign layer0_out[662] = ~x[138];
    assign layer0_out[663] = x[200] | x[202];
    assign layer0_out[664] = x[192];
    assign layer0_out[665] = ~(x[235] | x[237]);
    assign layer0_out[666] = ~(x[198] | x[199]);
    assign layer0_out[667] = x[69];
    assign layer0_out[668] = x[391] & x[392];
    assign layer0_out[669] = x[276];
    assign layer0_out[670] = x[305] | x[307];
    assign layer0_out[671] = x[301] | x[303];
    assign layer0_out[672] = 1'b0;
    assign layer0_out[673] = 1'b0;
    assign layer0_out[674] = x[145] | x[147];
    assign layer0_out[675] = ~(x[222] | x[224]);
    assign layer0_out[676] = ~(x[151] | x[153]);
    assign layer0_out[677] = ~(x[3] | x[4]);
    assign layer0_out[678] = ~(x[238] & x[240]);
    assign layer0_out[679] = ~x[238];
    assign layer0_out[680] = x[30];
    assign layer0_out[681] = ~(x[93] | x[94]);
    assign layer0_out[682] = ~(x[233] | x[235]);
    assign layer0_out[683] = 1'b0;
    assign layer0_out[684] = ~(x[153] | x[154]);
    assign layer0_out[685] = 1'b0;
    assign layer0_out[686] = x[135] | x[137];
    assign layer0_out[687] = 1'b0;
    assign layer0_out[688] = ~(x[144] | x[146]);
    assign layer0_out[689] = ~(x[294] | x[295]);
    assign layer0_out[690] = x[267] & ~x[265];
    assign layer0_out[691] = ~x[252];
    assign layer0_out[692] = x[31];
    assign layer0_out[693] = 1'b0;
    assign layer0_out[694] = x[353] | x[355];
    assign layer0_out[695] = ~(x[282] | x[283]);
    assign layer0_out[696] = ~(x[355] | x[356]);
    assign layer0_out[697] = x[250] | x[252];
    assign layer0_out[698] = x[313] & ~x[314];
    assign layer0_out[699] = x[326];
    assign layer0_out[700] = ~x[30];
    assign layer0_out[701] = ~(x[328] | x[329]);
    assign layer0_out[702] = ~(x[132] & x[133]);
    assign layer0_out[703] = 1'b1;
    assign layer0_out[704] = ~x[250] | x[249];
    assign layer0_out[705] = ~(x[326] | x[328]);
    assign layer0_out[706] = x[205] | x[207];
    assign layer0_out[707] = ~(x[123] | x[124]);
    assign layer0_out[708] = ~(x[66] | x[67]);
    assign layer0_out[709] = x[50] & ~x[52];
    assign layer0_out[710] = ~(x[108] & x[109]);
    assign layer0_out[711] = ~(x[37] | x[39]);
    assign layer0_out[712] = ~(x[174] | x[176]);
    assign layer0_out[713] = ~(x[298] | x[299]);
    assign layer0_out[714] = 1'b0;
    assign layer0_out[715] = x[200] | x[201];
    assign layer0_out[716] = ~(x[341] | x[343]);
    assign layer0_out[717] = x[226] | x[227];
    assign layer0_out[718] = x[286] | x[288];
    assign layer0_out[719] = x[37] & ~x[35];
    assign layer0_out[720] = x[93] & ~x[92];
    assign layer0_out[721] = 1'b1;
    assign layer0_out[722] = ~x[65] | x[67];
    assign layer0_out[723] = x[1] & x[4];
    assign layer0_out[724] = x[381] & ~x[382];
    assign layer0_out[725] = x[189];
    assign layer0_out[726] = x[253] | x[254];
    assign layer0_out[727] = x[322] | x[323];
    assign layer0_out[728] = ~(x[258] | x[260]);
    assign layer0_out[729] = 1'b0;
    assign layer0_out[730] = x[201] & x[202];
    assign layer0_out[731] = 1'b1;
    assign layer0_out[732] = x[257];
    assign layer0_out[733] = 1'b1;
    assign layer0_out[734] = ~x[194] | x[192];
    assign layer0_out[735] = x[314] | x[315];
    assign layer0_out[736] = ~(x[215] | x[216]);
    assign layer0_out[737] = 1'b0;
    assign layer0_out[738] = x[80] & ~x[81];
    assign layer0_out[739] = 1'b0;
    assign layer0_out[740] = x[83] | x[85];
    assign layer0_out[741] = x[175] & ~x[174];
    assign layer0_out[742] = x[273];
    assign layer0_out[743] = x[314] | x[316];
    assign layer0_out[744] = ~(x[375] | x[377]);
    assign layer0_out[745] = ~x[193] | x[191];
    assign layer0_out[746] = ~(x[119] & x[120]);
    assign layer0_out[747] = ~x[130] | x[131];
    assign layer0_out[748] = ~x[208];
    assign layer0_out[749] = ~(x[376] | x[377]);
    assign layer0_out[750] = ~(x[241] | x[242]);
    assign layer0_out[751] = ~(x[74] | x[76]);
    assign layer0_out[752] = x[365];
    assign layer0_out[753] = ~(x[106] | x[107]);
    assign layer0_out[754] = x[145];
    assign layer0_out[755] = ~(x[304] | x[306]);
    assign layer0_out[756] = ~(x[107] | x[109]);
    assign layer0_out[757] = ~(x[176] ^ x[178]);
    assign layer0_out[758] = ~(x[182] | x[183]);
    assign layer0_out[759] = ~x[293];
    assign layer0_out[760] = ~(x[142] | x[144]);
    assign layer0_out[761] = x[312];
    assign layer0_out[762] = ~x[127];
    assign layer0_out[763] = x[61] & ~x[63];
    assign layer0_out[764] = ~(x[296] | x[297]);
    assign layer0_out[765] = x[323] | x[325];
    assign layer0_out[766] = ~x[296] | x[294];
    assign layer0_out[767] = 1'b1;
    assign layer0_out[768] = x[36];
    assign layer0_out[769] = x[30] & ~x[32];
    assign layer0_out[770] = ~(x[177] | x[178]);
    assign layer0_out[771] = 1'b0;
    assign layer0_out[772] = x[141] | x[143];
    assign layer0_out[773] = ~(x[248] | x[250]);
    assign layer0_out[774] = ~(x[375] | x[376]);
    assign layer0_out[775] = ~(x[134] | x[136]);
    assign layer0_out[776] = x[123] | x[125];
    assign layer0_out[777] = 1'b1;
    assign layer0_out[778] = ~(x[173] | x[175]);
    assign layer0_out[779] = x[54] & x[55];
    assign layer0_out[780] = ~x[396];
    assign layer0_out[781] = x[373] | x[375];
    assign layer0_out[782] = ~x[281] | x[280];
    assign layer0_out[783] = ~(x[245] | x[246]);
    assign layer0_out[784] = 1'b1;
    assign layer0_out[785] = 1'b1;
    assign layer0_out[786] = ~x[184];
    assign layer0_out[787] = 1'b0;
    assign layer0_out[788] = ~x[11];
    assign layer0_out[789] = x[292] & x[294];
    assign layer0_out[790] = ~(x[380] & x[382]);
    assign layer0_out[791] = x[260] | x[262];
    assign layer0_out[792] = x[225] & ~x[227];
    assign layer0_out[793] = 1'b1;
    assign layer0_out[794] = ~(x[113] | x[114]);
    assign layer0_out[795] = ~(x[247] | x[249]);
    assign layer0_out[796] = x[321] | x[322];
    assign layer0_out[797] = 1'b0;
    assign layer0_out[798] = 1'b1;
    assign layer0_out[799] = x[269];
    assign layer1_out[0] = layer0_out[320] & ~layer0_out[321];
    assign layer1_out[1] = 1'b1;
    assign layer1_out[2] = layer0_out[453];
    assign layer1_out[3] = layer0_out[321] | layer0_out[322];
    assign layer1_out[4] = ~layer0_out[716] | layer0_out[715];
    assign layer1_out[5] = layer0_out[275] & ~layer0_out[276];
    assign layer1_out[6] = ~layer0_out[190];
    assign layer1_out[7] = ~layer0_out[132] | layer0_out[131];
    assign layer1_out[8] = ~layer0_out[99];
    assign layer1_out[9] = layer0_out[713] & ~layer0_out[712];
    assign layer1_out[10] = layer0_out[632];
    assign layer1_out[11] = layer0_out[296];
    assign layer1_out[12] = ~layer0_out[265] | layer0_out[266];
    assign layer1_out[13] = layer0_out[744] & layer0_out[745];
    assign layer1_out[14] = ~(layer0_out[229] | layer0_out[230]);
    assign layer1_out[15] = layer0_out[616];
    assign layer1_out[16] = ~(layer0_out[747] & layer0_out[748]);
    assign layer1_out[17] = ~layer0_out[458] | layer0_out[459];
    assign layer1_out[18] = ~(layer0_out[202] ^ layer0_out[203]);
    assign layer1_out[19] = layer0_out[516];
    assign layer1_out[20] = ~layer0_out[657];
    assign layer1_out[21] = layer0_out[403] & ~layer0_out[402];
    assign layer1_out[22] = layer0_out[547] | layer0_out[548];
    assign layer1_out[23] = layer0_out[687] & ~layer0_out[686];
    assign layer1_out[24] = layer0_out[493];
    assign layer1_out[25] = ~(layer0_out[125] | layer0_out[126]);
    assign layer1_out[26] = ~(layer0_out[155] | layer0_out[156]);
    assign layer1_out[27] = ~layer0_out[714];
    assign layer1_out[28] = ~layer0_out[100] | layer0_out[101];
    assign layer1_out[29] = ~layer0_out[492] | layer0_out[493];
    assign layer1_out[30] = layer0_out[731] & layer0_out[732];
    assign layer1_out[31] = ~(layer0_out[570] | layer0_out[571]);
    assign layer1_out[32] = 1'b1;
    assign layer1_out[33] = layer0_out[359];
    assign layer1_out[34] = ~layer0_out[378] | layer0_out[377];
    assign layer1_out[35] = layer0_out[770] & ~layer0_out[771];
    assign layer1_out[36] = layer0_out[778];
    assign layer1_out[37] = layer0_out[716];
    assign layer1_out[38] = layer0_out[416] & layer0_out[417];
    assign layer1_out[39] = ~(layer0_out[541] | layer0_out[542]);
    assign layer1_out[40] = layer0_out[46] & ~layer0_out[47];
    assign layer1_out[41] = ~layer0_out[86];
    assign layer1_out[42] = layer0_out[269] & ~layer0_out[270];
    assign layer1_out[43] = ~layer0_out[692];
    assign layer1_out[44] = layer0_out[29];
    assign layer1_out[45] = layer0_out[613];
    assign layer1_out[46] = layer0_out[354] & ~layer0_out[353];
    assign layer1_out[47] = ~layer0_out[795];
    assign layer1_out[48] = 1'b1;
    assign layer1_out[49] = layer0_out[766];
    assign layer1_out[50] = layer0_out[316];
    assign layer1_out[51] = layer0_out[648] & ~layer0_out[647];
    assign layer1_out[52] = ~(layer0_out[534] | layer0_out[535]);
    assign layer1_out[53] = layer0_out[61];
    assign layer1_out[54] = layer0_out[138] & ~layer0_out[139];
    assign layer1_out[55] = ~(layer0_out[442] | layer0_out[443]);
    assign layer1_out[56] = 1'b0;
    assign layer1_out[57] = layer0_out[609] & layer0_out[610];
    assign layer1_out[58] = layer0_out[688] & layer0_out[689];
    assign layer1_out[59] = layer0_out[761] | layer0_out[762];
    assign layer1_out[60] = ~layer0_out[345] | layer0_out[344];
    assign layer1_out[61] = ~layer0_out[26];
    assign layer1_out[62] = layer0_out[734];
    assign layer1_out[63] = ~layer0_out[735];
    assign layer1_out[64] = 1'b0;
    assign layer1_out[65] = layer0_out[484];
    assign layer1_out[66] = ~layer0_out[725] | layer0_out[726];
    assign layer1_out[67] = layer0_out[580];
    assign layer1_out[68] = ~(layer0_out[175] & layer0_out[176]);
    assign layer1_out[69] = layer0_out[356] | layer0_out[357];
    assign layer1_out[70] = ~(layer0_out[14] & layer0_out[15]);
    assign layer1_out[71] = layer0_out[566] & ~layer0_out[567];
    assign layer1_out[72] = ~layer0_out[147];
    assign layer1_out[73] = layer0_out[8] & layer0_out[9];
    assign layer1_out[74] = layer0_out[473];
    assign layer1_out[75] = layer0_out[680];
    assign layer1_out[76] = layer0_out[603] & ~layer0_out[602];
    assign layer1_out[77] = ~layer0_out[728] | layer0_out[727];
    assign layer1_out[78] = layer0_out[368];
    assign layer1_out[79] = ~layer0_out[95] | layer0_out[96];
    assign layer1_out[80] = layer0_out[596];
    assign layer1_out[81] = ~layer0_out[606];
    assign layer1_out[82] = ~layer0_out[405];
    assign layer1_out[83] = layer0_out[598] | layer0_out[599];
    assign layer1_out[84] = ~layer0_out[169];
    assign layer1_out[85] = layer0_out[237];
    assign layer1_out[86] = ~layer0_out[511];
    assign layer1_out[87] = layer0_out[464];
    assign layer1_out[88] = layer0_out[274];
    assign layer1_out[89] = ~layer0_out[199];
    assign layer1_out[90] = ~(layer0_out[54] & layer0_out[55]);
    assign layer1_out[91] = ~layer0_out[65] | layer0_out[66];
    assign layer1_out[92] = layer0_out[512] & layer0_out[513];
    assign layer1_out[93] = ~(layer0_out[432] ^ layer0_out[433]);
    assign layer1_out[94] = ~(layer0_out[454] | layer0_out[455]);
    assign layer1_out[95] = layer0_out[490];
    assign layer1_out[96] = layer0_out[558] & layer0_out[559];
    assign layer1_out[97] = layer0_out[246] | layer0_out[247];
    assign layer1_out[98] = 1'b0;
    assign layer1_out[99] = layer0_out[319];
    assign layer1_out[100] = layer0_out[788];
    assign layer1_out[101] = layer0_out[728] & ~layer0_out[729];
    assign layer1_out[102] = ~layer0_out[708];
    assign layer1_out[103] = ~(layer0_out[702] ^ layer0_out[703]);
    assign layer1_out[104] = layer0_out[771];
    assign layer1_out[105] = ~layer0_out[362];
    assign layer1_out[106] = ~(layer0_out[314] & layer0_out[315]);
    assign layer1_out[107] = layer0_out[740];
    assign layer1_out[108] = layer0_out[382];
    assign layer1_out[109] = ~layer0_out[264] | layer0_out[263];
    assign layer1_out[110] = layer0_out[421];
    assign layer1_out[111] = layer0_out[610] & layer0_out[611];
    assign layer1_out[112] = 1'b1;
    assign layer1_out[113] = ~layer0_out[156];
    assign layer1_out[114] = layer0_out[301] & ~layer0_out[302];
    assign layer1_out[115] = 1'b1;
    assign layer1_out[116] = layer0_out[80];
    assign layer1_out[117] = 1'b0;
    assign layer1_out[118] = layer0_out[20];
    assign layer1_out[119] = ~(layer0_out[730] | layer0_out[731]);
    assign layer1_out[120] = layer0_out[640] | layer0_out[641];
    assign layer1_out[121] = ~layer0_out[237];
    assign layer1_out[122] = ~(layer0_out[328] & layer0_out[329]);
    assign layer1_out[123] = layer0_out[285] ^ layer0_out[286];
    assign layer1_out[124] = layer0_out[562];
    assign layer1_out[125] = layer0_out[673] | layer0_out[674];
    assign layer1_out[126] = layer0_out[363] | layer0_out[364];
    assign layer1_out[127] = ~layer0_out[510];
    assign layer1_out[128] = layer0_out[730];
    assign layer1_out[129] = ~layer0_out[529] | layer0_out[528];
    assign layer1_out[130] = ~layer0_out[480] | layer0_out[481];
    assign layer1_out[131] = layer0_out[605];
    assign layer1_out[132] = 1'b1;
    assign layer1_out[133] = layer0_out[434] & ~layer0_out[435];
    assign layer1_out[134] = layer0_out[379];
    assign layer1_out[135] = ~layer0_out[759] | layer0_out[760];
    assign layer1_out[136] = ~layer0_out[57];
    assign layer1_out[137] = layer0_out[284];
    assign layer1_out[138] = ~layer0_out[335];
    assign layer1_out[139] = layer0_out[576];
    assign layer1_out[140] = layer0_out[775];
    assign layer1_out[141] = 1'b0;
    assign layer1_out[142] = ~layer0_out[770] | layer0_out[769];
    assign layer1_out[143] = layer0_out[292] & ~layer0_out[291];
    assign layer1_out[144] = ~layer0_out[520] | layer0_out[519];
    assign layer1_out[145] = ~layer0_out[79];
    assign layer1_out[146] = ~(layer0_out[732] & layer0_out[733]);
    assign layer1_out[147] = layer0_out[187] & layer0_out[188];
    assign layer1_out[148] = layer0_out[337];
    assign layer1_out[149] = ~layer0_out[533];
    assign layer1_out[150] = layer0_out[278];
    assign layer1_out[151] = ~layer0_out[581];
    assign layer1_out[152] = layer0_out[145];
    assign layer1_out[153] = ~(layer0_out[755] & layer0_out[756]);
    assign layer1_out[154] = layer0_out[44];
    assign layer1_out[155] = layer0_out[491] & layer0_out[492];
    assign layer1_out[156] = layer0_out[188] & ~layer0_out[189];
    assign layer1_out[157] = layer0_out[200] | layer0_out[201];
    assign layer1_out[158] = ~layer0_out[322];
    assign layer1_out[159] = ~layer0_out[666] | layer0_out[667];
    assign layer1_out[160] = ~layer0_out[325];
    assign layer1_out[161] = layer0_out[590] & ~layer0_out[589];
    assign layer1_out[162] = ~layer0_out[327] | layer0_out[328];
    assign layer1_out[163] = ~(layer0_out[163] ^ layer0_out[164]);
    assign layer1_out[164] = layer0_out[425] & layer0_out[426];
    assign layer1_out[165] = ~(layer0_out[584] & layer0_out[585]);
    assign layer1_out[166] = ~(layer0_out[340] & layer0_out[341]);
    assign layer1_out[167] = layer0_out[484] & ~layer0_out[483];
    assign layer1_out[168] = layer0_out[569];
    assign layer1_out[169] = ~layer0_out[457] | layer0_out[458];
    assign layer1_out[170] = layer0_out[41];
    assign layer1_out[171] = layer0_out[430] & layer0_out[431];
    assign layer1_out[172] = layer0_out[441] & ~layer0_out[442];
    assign layer1_out[173] = ~(layer0_out[171] | layer0_out[172]);
    assign layer1_out[174] = layer0_out[736] & ~layer0_out[735];
    assign layer1_out[175] = layer0_out[675] & ~layer0_out[674];
    assign layer1_out[176] = ~(layer0_out[157] | layer0_out[158]);
    assign layer1_out[177] = ~(layer0_out[504] & layer0_out[505]);
    assign layer1_out[178] = ~layer0_out[13];
    assign layer1_out[179] = 1'b0;
    assign layer1_out[180] = layer0_out[37] | layer0_out[38];
    assign layer1_out[181] = layer0_out[69];
    assign layer1_out[182] = layer0_out[782] & layer0_out[783];
    assign layer1_out[183] = layer0_out[791] | layer0_out[792];
    assign layer1_out[184] = layer0_out[28];
    assign layer1_out[185] = layer0_out[280];
    assign layer1_out[186] = layer0_out[744] & ~layer0_out[743];
    assign layer1_out[187] = layer0_out[325];
    assign layer1_out[188] = ~(layer0_out[62] | layer0_out[63]);
    assign layer1_out[189] = layer0_out[130] & ~layer0_out[131];
    assign layer1_out[190] = ~layer0_out[97];
    assign layer1_out[191] = ~layer0_out[705];
    assign layer1_out[192] = ~(layer0_out[208] | layer0_out[209]);
    assign layer1_out[193] = layer0_out[562];
    assign layer1_out[194] = ~layer0_out[323];
    assign layer1_out[195] = ~(layer0_out[397] | layer0_out[398]);
    assign layer1_out[196] = layer0_out[615] & ~layer0_out[616];
    assign layer1_out[197] = layer0_out[86] & ~layer0_out[85];
    assign layer1_out[198] = ~layer0_out[251];
    assign layer1_out[199] = layer0_out[465] & ~layer0_out[466];
    assign layer1_out[200] = ~layer0_out[371];
    assign layer1_out[201] = layer0_out[552];
    assign layer1_out[202] = ~layer0_out[113];
    assign layer1_out[203] = layer0_out[752];
    assign layer1_out[204] = 1'b1;
    assign layer1_out[205] = ~(layer0_out[114] ^ layer0_out[115]);
    assign layer1_out[206] = layer0_out[762];
    assign layer1_out[207] = layer0_out[564] | layer0_out[565];
    assign layer1_out[208] = layer0_out[334];
    assign layer1_out[209] = layer0_out[308] & layer0_out[309];
    assign layer1_out[210] = layer0_out[254];
    assign layer1_out[211] = layer0_out[530];
    assign layer1_out[212] = 1'b0;
    assign layer1_out[213] = ~(layer0_out[401] & layer0_out[402]);
    assign layer1_out[214] = ~layer0_out[430];
    assign layer1_out[215] = layer0_out[235];
    assign layer1_out[216] = ~layer0_out[76];
    assign layer1_out[217] = layer0_out[161] & layer0_out[162];
    assign layer1_out[218] = ~layer0_out[233];
    assign layer1_out[219] = layer0_out[786];
    assign layer1_out[220] = layer0_out[678];
    assign layer1_out[221] = ~layer0_out[185] | layer0_out[184];
    assign layer1_out[222] = ~layer0_out[215] | layer0_out[214];
    assign layer1_out[223] = ~layer0_out[158] | layer0_out[159];
    assign layer1_out[224] = ~(layer0_out[240] & layer0_out[241]);
    assign layer1_out[225] = ~(layer0_out[533] ^ layer0_out[534]);
    assign layer1_out[226] = ~layer0_out[19] | layer0_out[20];
    assign layer1_out[227] = layer0_out[191];
    assign layer1_out[228] = ~layer0_out[684] | layer0_out[685];
    assign layer1_out[229] = layer0_out[538] | layer0_out[539];
    assign layer1_out[230] = layer0_out[348] | layer0_out[349];
    assign layer1_out[231] = layer0_out[609] & ~layer0_out[608];
    assign layer1_out[232] = layer0_out[677];
    assign layer1_out[233] = ~layer0_out[362] | layer0_out[363];
    assign layer1_out[234] = layer0_out[773] & ~layer0_out[772];
    assign layer1_out[235] = layer0_out[95];
    assign layer1_out[236] = layer0_out[9] | layer0_out[10];
    assign layer1_out[237] = ~(layer0_out[667] | layer0_out[668]);
    assign layer1_out[238] = ~(layer0_out[537] & layer0_out[538]);
    assign layer1_out[239] = layer0_out[404];
    assign layer1_out[240] = layer0_out[168] & ~layer0_out[169];
    assign layer1_out[241] = layer0_out[787] & ~layer0_out[786];
    assign layer1_out[242] = ~layer0_out[656];
    assign layer1_out[243] = layer0_out[556] & ~layer0_out[555];
    assign layer1_out[244] = layer0_out[262] & ~layer0_out[261];
    assign layer1_out[245] = layer0_out[58];
    assign layer1_out[246] = 1'b1;
    assign layer1_out[247] = ~(layer0_out[203] & layer0_out[204]);
    assign layer1_out[248] = ~(layer0_out[6] | layer0_out[7]);
    assign layer1_out[249] = ~layer0_out[486];
    assign layer1_out[250] = ~(layer0_out[317] | layer0_out[318]);
    assign layer1_out[251] = 1'b0;
    assign layer1_out[252] = layer0_out[503] & ~layer0_out[502];
    assign layer1_out[253] = layer0_out[557];
    assign layer1_out[254] = ~(layer0_out[452] | layer0_out[453]);
    assign layer1_out[255] = ~(layer0_out[206] & layer0_out[207]);
    assign layer1_out[256] = layer0_out[720];
    assign layer1_out[257] = ~(layer0_out[381] & layer0_out[382]);
    assign layer1_out[258] = layer0_out[7] | layer0_out[8];
    assign layer1_out[259] = 1'b0;
    assign layer1_out[260] = layer0_out[645] | layer0_out[646];
    assign layer1_out[261] = 1'b0;
    assign layer1_out[262] = layer0_out[50] & ~layer0_out[51];
    assign layer1_out[263] = 1'b1;
    assign layer1_out[264] = ~layer0_out[565];
    assign layer1_out[265] = ~layer0_out[212];
    assign layer1_out[266] = layer0_out[712];
    assign layer1_out[267] = layer0_out[278] & ~layer0_out[279];
    assign layer1_out[268] = layer0_out[448] & ~layer0_out[447];
    assign layer1_out[269] = ~layer0_out[39];
    assign layer1_out[270] = ~layer0_out[758] | layer0_out[757];
    assign layer1_out[271] = layer0_out[205] ^ layer0_out[206];
    assign layer1_out[272] = 1'b1;
    assign layer1_out[273] = layer0_out[615];
    assign layer1_out[274] = ~(layer0_out[74] | layer0_out[75]);
    assign layer1_out[275] = ~layer0_out[35];
    assign layer1_out[276] = ~layer0_out[428] | layer0_out[429];
    assign layer1_out[277] = ~layer0_out[245] | layer0_out[246];
    assign layer1_out[278] = layer0_out[374];
    assign layer1_out[279] = ~layer0_out[138];
    assign layer1_out[280] = 1'b1;
    assign layer1_out[281] = ~layer0_out[418] | layer0_out[419];
    assign layer1_out[282] = ~layer0_out[87];
    assign layer1_out[283] = layer0_out[74] & ~layer0_out[73];
    assign layer1_out[284] = ~layer0_out[788];
    assign layer1_out[285] = ~layer0_out[66];
    assign layer1_out[286] = layer0_out[33] & ~layer0_out[32];
    assign layer1_out[287] = layer0_out[373] & ~layer0_out[374];
    assign layer1_out[288] = layer0_out[341] & ~layer0_out[342];
    assign layer1_out[289] = ~layer0_out[612];
    assign layer1_out[290] = ~layer0_out[288];
    assign layer1_out[291] = ~layer0_out[587];
    assign layer1_out[292] = layer0_out[310];
    assign layer1_out[293] = layer0_out[216] & ~layer0_out[217];
    assign layer1_out[294] = ~layer0_out[524];
    assign layer1_out[295] = 1'b0;
    assign layer1_out[296] = ~layer0_out[26];
    assign layer1_out[297] = layer0_out[741] | layer0_out[742];
    assign layer1_out[298] = ~layer0_out[18];
    assign layer1_out[299] = layer0_out[665] & ~layer0_out[664];
    assign layer1_out[300] = layer0_out[218] & ~layer0_out[219];
    assign layer1_out[301] = ~layer0_out[559] | layer0_out[560];
    assign layer1_out[302] = 1'b0;
    assign layer1_out[303] = ~layer0_out[387];
    assign layer1_out[304] = ~layer0_out[794];
    assign layer1_out[305] = ~layer0_out[264];
    assign layer1_out[306] = ~layer0_out[691];
    assign layer1_out[307] = layer0_out[424];
    assign layer1_out[308] = layer0_out[76] & layer0_out[77];
    assign layer1_out[309] = layer0_out[127] & ~layer0_out[128];
    assign layer1_out[310] = layer0_out[795];
    assign layer1_out[311] = layer0_out[639];
    assign layer1_out[312] = ~layer0_out[626];
    assign layer1_out[313] = ~(layer0_out[648] & layer0_out[649]);
    assign layer1_out[314] = layer0_out[385] & layer0_out[386];
    assign layer1_out[315] = 1'b0;
    assign layer1_out[316] = ~layer0_out[586] | layer0_out[585];
    assign layer1_out[317] = ~(layer0_out[52] & layer0_out[53]);
    assign layer1_out[318] = layer0_out[59] & layer0_out[60];
    assign layer1_out[319] = ~layer0_out[196];
    assign layer1_out[320] = layer0_out[563] ^ layer0_out[564];
    assign layer1_out[321] = layer0_out[249] & ~layer0_out[250];
    assign layer1_out[322] = ~layer0_out[271] | layer0_out[272];
    assign layer1_out[323] = ~layer0_out[671];
    assign layer1_out[324] = ~layer0_out[546];
    assign layer1_out[325] = layer0_out[398] | layer0_out[399];
    assign layer1_out[326] = layer0_out[261];
    assign layer1_out[327] = ~layer0_out[72];
    assign layer1_out[328] = layer0_out[293] & ~layer0_out[292];
    assign layer1_out[329] = layer0_out[192] & layer0_out[193];
    assign layer1_out[330] = layer0_out[596] & ~layer0_out[597];
    assign layer1_out[331] = layer0_out[699] & ~layer0_out[700];
    assign layer1_out[332] = layer0_out[633] ^ layer0_out[634];
    assign layer1_out[333] = ~layer0_out[282];
    assign layer1_out[334] = layer0_out[1] & layer0_out[2];
    assign layer1_out[335] = layer0_out[55] | layer0_out[56];
    assign layer1_out[336] = layer0_out[69] | layer0_out[70];
    assign layer1_out[337] = layer0_out[569] & layer0_out[570];
    assign layer1_out[338] = ~layer0_out[407] | layer0_out[406];
    assign layer1_out[339] = layer0_out[391] & ~layer0_out[390];
    assign layer1_out[340] = ~layer0_out[366];
    assign layer1_out[341] = ~(layer0_out[669] | layer0_out[670]);
    assign layer1_out[342] = layer0_out[606];
    assign layer1_out[343] = layer0_out[707] & ~layer0_out[706];
    assign layer1_out[344] = layer0_out[498];
    assign layer1_out[345] = ~layer0_out[339] | layer0_out[340];
    assign layer1_out[346] = layer0_out[549];
    assign layer1_out[347] = ~layer0_out[288] | layer0_out[289];
    assign layer1_out[348] = layer0_out[182] & layer0_out[183];
    assign layer1_out[349] = ~layer0_out[28];
    assign layer1_out[350] = layer0_out[174];
    assign layer1_out[351] = layer0_out[242];
    assign layer1_out[352] = ~(layer0_out[510] | layer0_out[511]);
    assign layer1_out[353] = ~layer0_out[440] | layer0_out[439];
    assign layer1_out[354] = ~layer0_out[48];
    assign layer1_out[355] = ~(layer0_out[784] | layer0_out[785]);
    assign layer1_out[356] = layer0_out[422] ^ layer0_out[423];
    assign layer1_out[357] = layer0_out[631] & ~layer0_out[630];
    assign layer1_out[358] = layer0_out[352];
    assign layer1_out[359] = 1'b1;
    assign layer1_out[360] = 1'b1;
    assign layer1_out[361] = ~(layer0_out[0] & layer0_out[1]);
    assign layer1_out[362] = ~(layer0_out[527] & layer0_out[528]);
    assign layer1_out[363] = layer0_out[333] & ~layer0_out[332];
    assign layer1_out[364] = ~layer0_out[108] | layer0_out[107];
    assign layer1_out[365] = layer0_out[355] & ~layer0_out[354];
    assign layer1_out[366] = 1'b0;
    assign layer1_out[367] = layer0_out[85];
    assign layer1_out[368] = ~(layer0_out[724] ^ layer0_out[725]);
    assign layer1_out[369] = layer0_out[659] & ~layer0_out[658];
    assign layer1_out[370] = ~layer0_out[121] | layer0_out[122];
    assign layer1_out[371] = layer0_out[257];
    assign layer1_out[372] = ~(layer0_out[318] ^ layer0_out[319]);
    assign layer1_out[373] = ~(layer0_out[148] ^ layer0_out[149]);
    assign layer1_out[374] = layer0_out[796];
    assign layer1_out[375] = layer0_out[191];
    assign layer1_out[376] = layer0_out[501];
    assign layer1_out[377] = layer0_out[567] & layer0_out[568];
    assign layer1_out[378] = ~(layer0_out[679] & layer0_out[680]);
    assign layer1_out[379] = ~layer0_out[396] | layer0_out[397];
    assign layer1_out[380] = layer0_out[675];
    assign layer1_out[381] = 1'b0;
    assign layer1_out[382] = ~layer0_out[124];
    assign layer1_out[383] = layer0_out[636] & layer0_out[637];
    assign layer1_out[384] = ~(layer0_out[573] & layer0_out[574]);
    assign layer1_out[385] = layer0_out[22];
    assign layer1_out[386] = layer0_out[449] & ~layer0_out[448];
    assign layer1_out[387] = layer0_out[350] & ~layer0_out[349];
    assign layer1_out[388] = ~(layer0_out[4] | layer0_out[5]);
    assign layer1_out[389] = ~(layer0_out[300] & layer0_out[301]);
    assign layer1_out[390] = ~layer0_out[696];
    assign layer1_out[391] = ~layer0_out[515];
    assign layer1_out[392] = layer0_out[764];
    assign layer1_out[393] = ~layer0_out[764] | layer0_out[763];
    assign layer1_out[394] = layer0_out[115] & layer0_out[116];
    assign layer1_out[395] = layer0_out[516];
    assign layer1_out[396] = layer0_out[186];
    assign layer1_out[397] = ~layer0_out[315] | layer0_out[316];
    assign layer1_out[398] = ~layer0_out[177] | layer0_out[178];
    assign layer1_out[399] = layer0_out[497];
    assign layer1_out[400] = ~(layer0_out[242] | layer0_out[243]);
    assign layer1_out[401] = layer0_out[244] & ~layer0_out[243];
    assign layer1_out[402] = ~layer0_out[420] | layer0_out[419];
    assign layer1_out[403] = ~layer0_out[612];
    assign layer1_out[404] = ~layer0_out[93] | layer0_out[92];
    assign layer1_out[405] = ~(layer0_out[629] & layer0_out[630]);
    assign layer1_out[406] = layer0_out[141];
    assign layer1_out[407] = ~layer0_out[437];
    assign layer1_out[408] = ~layer0_out[97];
    assign layer1_out[409] = layer0_out[653] ^ layer0_out[654];
    assign layer1_out[410] = 1'b0;
    assign layer1_out[411] = layer0_out[401];
    assign layer1_out[412] = ~(layer0_out[603] & layer0_out[604]);
    assign layer1_out[413] = layer0_out[286] & ~layer0_out[287];
    assign layer1_out[414] = layer0_out[540];
    assign layer1_out[415] = layer0_out[710] & ~layer0_out[711];
    assign layer1_out[416] = ~layer0_out[311];
    assign layer1_out[417] = ~layer0_out[505];
    assign layer1_out[418] = layer0_out[207] | layer0_out[208];
    assign layer1_out[419] = layer0_out[102];
    assign layer1_out[420] = layer0_out[549];
    assign layer1_out[421] = layer0_out[255];
    assign layer1_out[422] = ~layer0_out[258];
    assign layer1_out[423] = layer0_out[226];
    assign layer1_out[424] = layer0_out[139];
    assign layer1_out[425] = layer0_out[145];
    assign layer1_out[426] = layer0_out[273];
    assign layer1_out[427] = ~layer0_out[91];
    assign layer1_out[428] = ~layer0_out[120] | layer0_out[119];
    assign layer1_out[429] = layer0_out[489];
    assign layer1_out[430] = layer0_out[776];
    assign layer1_out[431] = 1'b0;
    assign layer1_out[432] = layer0_out[682];
    assign layer1_out[433] = layer0_out[727];
    assign layer1_out[434] = ~layer0_out[437];
    assign layer1_out[435] = layer0_out[123] & ~layer0_out[122];
    assign layer1_out[436] = ~(layer0_out[507] | layer0_out[508]);
    assign layer1_out[437] = layer0_out[204] | layer0_out[205];
    assign layer1_out[438] = layer0_out[719];
    assign layer1_out[439] = ~layer0_out[211] | layer0_out[210];
    assign layer1_out[440] = layer0_out[513] | layer0_out[514];
    assign layer1_out[441] = layer0_out[520];
    assign layer1_out[442] = ~(layer0_out[789] & layer0_out[790]);
    assign layer1_out[443] = 1'b1;
    assign layer1_out[444] = ~layer0_out[49] | layer0_out[48];
    assign layer1_out[445] = layer0_out[5];
    assign layer1_out[446] = layer0_out[415];
    assign layer1_out[447] = layer0_out[506];
    assign layer1_out[448] = layer0_out[635];
    assign layer1_out[449] = ~layer0_out[707];
    assign layer1_out[450] = ~(layer0_out[560] | layer0_out[561]);
    assign layer1_out[451] = layer0_out[508] | layer0_out[509];
    assign layer1_out[452] = ~layer0_out[281];
    assign layer1_out[453] = layer0_out[395] & layer0_out[396];
    assign layer1_out[454] = layer0_out[653];
    assign layer1_out[455] = ~layer0_out[134];
    assign layer1_out[456] = ~layer0_out[78];
    assign layer1_out[457] = ~(layer0_out[517] & layer0_out[518]);
    assign layer1_out[458] = 1'b1;
    assign layer1_out[459] = layer0_out[357] & ~layer0_out[358];
    assign layer1_out[460] = layer0_out[353];
    assign layer1_out[461] = layer0_out[540];
    assign layer1_out[462] = ~(layer0_out[173] & layer0_out[174]);
    assign layer1_out[463] = layer0_out[39];
    assign layer1_out[464] = ~(layer0_out[165] ^ layer0_out[166]);
    assign layer1_out[465] = layer0_out[651];
    assign layer1_out[466] = layer0_out[306];
    assign layer1_out[467] = ~layer0_out[392];
    assign layer1_out[468] = ~layer0_out[142];
    assign layer1_out[469] = layer0_out[590] | layer0_out[591];
    assign layer1_out[470] = 1'b0;
    assign layer1_out[471] = 1'b0;
    assign layer1_out[472] = layer0_out[332];
    assign layer1_out[473] = layer0_out[93] ^ layer0_out[94];
    assign layer1_out[474] = ~(layer0_out[644] | layer0_out[645]);
    assign layer1_out[475] = ~layer0_out[408];
    assign layer1_out[476] = layer0_out[655];
    assign layer1_out[477] = layer0_out[421];
    assign layer1_out[478] = ~(layer0_out[233] | layer0_out[234]);
    assign layer1_out[479] = layer0_out[557];
    assign layer1_out[480] = layer0_out[781] & layer0_out[782];
    assign layer1_out[481] = ~layer0_out[106];
    assign layer1_out[482] = layer0_out[745];
    assign layer1_out[483] = layer0_out[672] | layer0_out[673];
    assign layer1_out[484] = ~(layer0_out[111] | layer0_out[112]);
    assign layer1_out[485] = ~layer0_out[600] | layer0_out[601];
    assign layer1_out[486] = layer0_out[42] & ~layer0_out[43];
    assign layer1_out[487] = ~layer0_out[194];
    assign layer1_out[488] = layer0_out[427] & layer0_out[428];
    assign layer1_out[489] = 1'b1;
    assign layer1_out[490] = layer0_out[399];
    assign layer1_out[491] = ~layer0_out[304];
    assign layer1_out[492] = ~layer0_out[414];
    assign layer1_out[493] = ~layer0_out[499];
    assign layer1_out[494] = layer0_out[227] & ~layer0_out[228];
    assign layer1_out[495] = layer0_out[760];
    assign layer1_out[496] = 1'b1;
    assign layer1_out[497] = layer0_out[15];
    assign layer1_out[498] = layer0_out[141];
    assign layer1_out[499] = ~(layer0_out[213] & layer0_out[214]);
    assign layer1_out[500] = ~(layer0_out[393] | layer0_out[394]);
    assign layer1_out[501] = ~(layer0_out[297] | layer0_out[298]);
    assign layer1_out[502] = layer0_out[463] & ~layer0_out[464];
    assign layer1_out[503] = layer0_out[112];
    assign layer1_out[504] = layer0_out[637] & ~layer0_out[638];
    assign layer1_out[505] = layer0_out[460];
    assign layer1_out[506] = ~layer0_out[244];
    assign layer1_out[507] = layer0_out[411] | layer0_out[412];
    assign layer1_out[508] = layer0_out[280] | layer0_out[281];
    assign layer1_out[509] = ~layer0_out[58];
    assign layer1_out[510] = ~layer0_out[490] | layer0_out[491];
    assign layer1_out[511] = layer0_out[128] | layer0_out[129];
    assign layer1_out[512] = ~layer0_out[677] | layer0_out[676];
    assign layer1_out[513] = layer0_out[588] | layer0_out[589];
    assign layer1_out[514] = ~(layer0_out[124] & layer0_out[125]);
    assign layer1_out[515] = ~(layer0_out[478] & layer0_out[479]);
    assign layer1_out[516] = layer0_out[476] & ~layer0_out[475];
    assign layer1_out[517] = layer0_out[636] & ~layer0_out[635];
    assign layer1_out[518] = ~layer0_out[163];
    assign layer1_out[519] = ~layer0_out[91];
    assign layer1_out[520] = ~layer0_out[183];
    assign layer1_out[521] = layer0_out[649] | layer0_out[650];
    assign layer1_out[522] = layer0_out[544] & layer0_out[545];
    assign layer1_out[523] = layer0_out[625] | layer0_out[626];
    assign layer1_out[524] = layer0_out[466];
    assign layer1_out[525] = ~layer0_out[221];
    assign layer1_out[526] = ~layer0_out[600];
    assign layer1_out[527] = layer0_out[172];
    assign layer1_out[528] = layer0_out[755];
    assign layer1_out[529] = ~layer0_out[444];
    assign layer1_out[530] = ~(layer0_out[758] & layer0_out[759]);
    assign layer1_out[531] = layer0_out[24] & ~layer0_out[23];
    assign layer1_out[532] = ~(layer0_out[546] & layer0_out[547]);
    assign layer1_out[533] = layer0_out[302];
    assign layer1_out[534] = layer0_out[226];
    assign layer1_out[535] = ~layer0_out[4] | layer0_out[3];
    assign layer1_out[536] = ~(layer0_out[749] & layer0_out[750]);
    assign layer1_out[537] = ~layer0_out[671];
    assign layer1_out[538] = layer0_out[355];
    assign layer1_out[539] = 1'b1;
    assign layer1_out[540] = layer0_out[592] & ~layer0_out[591];
    assign layer1_out[541] = layer0_out[379];
    assign layer1_out[542] = ~layer0_out[751] | layer0_out[750];
    assign layer1_out[543] = ~layer0_out[461];
    assign layer1_out[544] = layer0_out[551];
    assign layer1_out[545] = ~layer0_out[706];
    assign layer1_out[546] = ~layer0_out[659];
    assign layer1_out[547] = 1'b1;
    assign layer1_out[548] = layer0_out[774];
    assign layer1_out[549] = ~layer0_out[468];
    assign layer1_out[550] = ~layer0_out[519] | layer0_out[518];
    assign layer1_out[551] = layer0_out[268];
    assign layer1_out[552] = 1'b0;
    assign layer1_out[553] = layer0_out[647];
    assign layer1_out[554] = layer0_out[110];
    assign layer1_out[555] = layer0_out[572] | layer0_out[573];
    assign layer1_out[556] = layer0_out[715];
    assign layer1_out[557] = 1'b0;
    assign layer1_out[558] = 1'b1;
    assign layer1_out[559] = ~layer0_out[151];
    assign layer1_out[560] = layer0_out[773];
    assign layer1_out[561] = layer0_out[783] | layer0_out[784];
    assign layer1_out[562] = ~layer0_out[37];
    assign layer1_out[563] = layer0_out[435] & layer0_out[436];
    assign layer1_out[564] = 1'b0;
    assign layer1_out[565] = ~layer0_out[166];
    assign layer1_out[566] = layer0_out[219];
    assign layer1_out[567] = layer0_out[691];
    assign layer1_out[568] = layer0_out[181];
    assign layer1_out[569] = layer0_out[737] & layer0_out[738];
    assign layer1_out[570] = ~layer0_out[347] | layer0_out[346];
    assign layer1_out[571] = ~(layer0_out[748] & layer0_out[749]);
    assign layer1_out[572] = layer0_out[477] & layer0_out[478];
    assign layer1_out[573] = ~layer0_out[480] | layer0_out[479];
    assign layer1_out[574] = ~layer0_out[240];
    assign layer1_out[575] = layer0_out[236];
    assign layer1_out[576] = ~layer0_out[30];
    assign layer1_out[577] = ~layer0_out[597];
    assign layer1_out[578] = ~layer0_out[384];
    assign layer1_out[579] = layer0_out[594] ^ layer0_out[595];
    assign layer1_out[580] = layer0_out[338] & ~layer0_out[337];
    assign layer1_out[581] = ~layer0_out[522] | layer0_out[521];
    assign layer1_out[582] = layer0_out[471];
    assign layer1_out[583] = layer0_out[440];
    assign layer1_out[584] = ~layer0_out[660];
    assign layer1_out[585] = ~(layer0_out[43] | layer0_out[44]);
    assign layer1_out[586] = layer0_out[535] & ~layer0_out[536];
    assign layer1_out[587] = ~layer0_out[410] | layer0_out[411];
    assign layer1_out[588] = ~layer0_out[450];
    assign layer1_out[589] = layer0_out[644];
    assign layer1_out[590] = layer0_out[368] & ~layer0_out[367];
    assign layer1_out[591] = layer0_out[250] & ~layer0_out[251];
    assign layer1_out[592] = layer0_out[290];
    assign layer1_out[593] = ~(layer0_out[740] | layer0_out[741]);
    assign layer1_out[594] = layer0_out[619] & ~layer0_out[620];
    assign layer1_out[595] = layer0_out[621];
    assign layer1_out[596] = layer0_out[259] & layer0_out[260];
    assign layer1_out[597] = layer0_out[369];
    assign layer1_out[598] = layer0_out[82] | layer0_out[83];
    assign layer1_out[599] = ~(layer0_out[307] | layer0_out[308]);
    assign layer1_out[600] = layer0_out[178];
    assign layer1_out[601] = layer0_out[415] & layer0_out[416];
    assign layer1_out[602] = ~layer0_out[470] | layer0_out[471];
    assign layer1_out[603] = layer0_out[89] | layer0_out[90];
    assign layer1_out[604] = layer0_out[623] | layer0_out[624];
    assign layer1_out[605] = ~layer0_out[294];
    assign layer1_out[606] = layer0_out[643];
    assign layer1_out[607] = ~layer0_out[459];
    assign layer1_out[608] = ~(layer0_out[149] | layer0_out[150]);
    assign layer1_out[609] = layer0_out[201];
    assign layer1_out[610] = ~layer0_out[89] | layer0_out[88];
    assign layer1_out[611] = layer0_out[176];
    assign layer1_out[612] = layer0_out[799];
    assign layer1_out[613] = layer0_out[543];
    assign layer1_out[614] = ~layer0_out[277];
    assign layer1_out[615] = layer0_out[498];
    assign layer1_out[616] = ~layer0_out[446];
    assign layer1_out[617] = ~(layer0_out[61] | layer0_out[62]);
    assign layer1_out[618] = layer0_out[473];
    assign layer1_out[619] = layer0_out[130];
    assign layer1_out[620] = layer0_out[266] ^ layer0_out[267];
    assign layer1_out[621] = layer0_out[159];
    assign layer1_out[622] = layer0_out[164] & ~layer0_out[165];
    assign layer1_out[623] = ~layer0_out[168];
    assign layer1_out[624] = layer0_out[701] & ~layer0_out[700];
    assign layer1_out[625] = 1'b1;
    assign layer1_out[626] = layer0_out[151] & ~layer0_out[152];
    assign layer1_out[627] = 1'b0;
    assign layer1_out[628] = layer0_out[717];
    assign layer1_out[629] = layer0_out[450];
    assign layer1_out[630] = layer0_out[689];
    assign layer1_out[631] = layer0_out[257] | layer0_out[258];
    assign layer1_out[632] = 1'b0;
    assign layer1_out[633] = ~layer0_out[135] | layer0_out[136];
    assign layer1_out[634] = ~(layer0_out[407] & layer0_out[408]);
    assign layer1_out[635] = ~layer0_out[198] | layer0_out[197];
    assign layer1_out[636] = layer0_out[359];
    assign layer1_out[637] = ~layer0_out[756];
    assign layer1_out[638] = ~layer0_out[739];
    assign layer1_out[639] = 1'b0;
    assign layer1_out[640] = 1'b0;
    assign layer1_out[641] = layer0_out[627] & layer0_out[628];
    assign layer1_out[642] = ~(layer0_out[387] & layer0_out[388]);
    assign layer1_out[643] = ~layer0_out[100];
    assign layer1_out[644] = ~(layer0_out[694] | layer0_out[695]);
    assign layer1_out[645] = layer0_out[104] ^ layer0_out[105];
    assign layer1_out[646] = layer0_out[127];
    assign layer1_out[647] = ~layer0_out[588] | layer0_out[587];
    assign layer1_out[648] = layer0_out[217];
    assign layer1_out[649] = layer0_out[134] & ~layer0_out[133];
    assign layer1_out[650] = layer0_out[417] ^ layer0_out[418];
    assign layer1_out[651] = layer0_out[426] & ~layer0_out[427];
    assign layer1_out[652] = ~(layer0_out[703] | layer0_out[704]);
    assign layer1_out[653] = layer0_out[409] & layer0_out[410];
    assign layer1_out[654] = 1'b0;
    assign layer1_out[655] = layer0_out[143];
    assign layer1_out[656] = layer0_out[14] & ~layer0_out[13];
    assign layer1_out[657] = layer0_out[33];
    assign layer1_out[658] = layer0_out[117];
    assign layer1_out[659] = layer0_out[555] & ~layer0_out[554];
    assign layer1_out[660] = layer0_out[106];
    assign layer1_out[661] = ~layer0_out[82];
    assign layer1_out[662] = layer0_out[621] ^ layer0_out[622];
    assign layer1_out[663] = ~(layer0_out[571] | layer0_out[572]);
    assign layer1_out[664] = ~layer0_out[476] | layer0_out[477];
    assign layer1_out[665] = ~layer0_out[622];
    assign layer1_out[666] = ~layer0_out[110] | layer0_out[109];
    assign layer1_out[667] = ~layer0_out[229] | layer0_out[228];
    assign layer1_out[668] = ~layer0_out[765] | layer0_out[766];
    assign layer1_out[669] = layer0_out[23];
    assign layer1_out[670] = ~layer0_out[390];
    assign layer1_out[671] = ~(layer0_out[342] | layer0_out[343]);
    assign layer1_out[672] = ~layer0_out[133];
    assign layer1_out[673] = ~layer0_out[504];
    assign layer1_out[674] = ~layer0_out[312] | layer0_out[311];
    assign layer1_out[675] = ~layer0_out[632];
    assign layer1_out[676] = layer0_out[147] ^ layer0_out[148];
    assign layer1_out[677] = ~layer0_out[697];
    assign layer1_out[678] = ~layer0_out[526];
    assign layer1_out[679] = ~layer0_out[196] | layer0_out[197];
    assign layer1_out[680] = layer0_out[791] & ~layer0_out[790];
    assign layer1_out[681] = layer0_out[329] | layer0_out[330];
    assign layer1_out[682] = layer0_out[554];
    assign layer1_out[683] = ~(layer0_out[45] & layer0_out[46]);
    assign layer1_out[684] = layer0_out[343];
    assign layer1_out[685] = layer0_out[593];
    assign layer1_out[686] = layer0_out[495];
    assign layer1_out[687] = ~layer0_out[68] | layer0_out[67];
    assign layer1_out[688] = ~layer0_out[584];
    assign layer1_out[689] = ~layer0_out[686];
    assign layer1_out[690] = ~layer0_out[231];
    assign layer1_out[691] = layer0_out[618] & ~layer0_out[619];
    assign layer1_out[692] = layer0_out[194];
    assign layer1_out[693] = layer0_out[688];
    assign layer1_out[694] = ~(layer0_out[116] | layer0_out[117]);
    assign layer1_out[695] = 1'b0;
    assign layer1_out[696] = layer0_out[681];
    assign layer1_out[697] = layer0_out[24];
    assign layer1_out[698] = ~(layer0_out[299] | layer0_out[300]);
    assign layer1_out[699] = layer0_out[155] & ~layer0_out[154];
    assign layer1_out[700] = layer0_out[406];
    assign layer1_out[701] = 1'b0;
    assign layer1_out[702] = layer0_out[270];
    assign layer1_out[703] = layer0_out[530];
    assign layer1_out[704] = ~layer0_out[724] | layer0_out[723];
    assign layer1_out[705] = ~layer0_out[225] | layer0_out[224];
    assign layer1_out[706] = ~(layer0_out[601] & layer0_out[602]);
    assign layer1_out[707] = ~layer0_out[153] | layer0_out[154];
    assign layer1_out[708] = ~layer0_out[639] | layer0_out[640];
    assign layer1_out[709] = layer0_out[71] & ~layer0_out[70];
    assign layer1_out[710] = layer0_out[2] & ~layer0_out[0];
    assign layer1_out[711] = layer0_out[768];
    assign layer1_out[712] = layer0_out[593] & ~layer0_out[592];
    assign layer1_out[713] = 1'b1;
    assign layer1_out[714] = 1'b0;
    assign layer1_out[715] = layer0_out[102];
    assign layer1_out[716] = layer0_out[118] | layer0_out[119];
    assign layer1_out[717] = layer0_out[295];
    assign layer1_out[718] = layer0_out[451] ^ layer0_out[452];
    assign layer1_out[719] = ~layer0_out[423];
    assign layer1_out[720] = layer0_out[350] & ~layer0_out[351];
    assign layer1_out[721] = layer0_out[2] & layer0_out[3];
    assign layer1_out[722] = layer0_out[779] & layer0_out[780];
    assign layer1_out[723] = layer0_out[41] & ~layer0_out[42];
    assign layer1_out[724] = layer0_out[709];
    assign layer1_out[725] = ~layer0_out[662] | layer0_out[661];
    assign layer1_out[726] = layer0_out[262] & ~layer0_out[263];
    assign layer1_out[727] = layer0_out[483] & ~layer0_out[482];
    assign layer1_out[728] = layer0_out[641] | layer0_out[642];
    assign layer1_out[729] = ~(layer0_out[360] | layer0_out[361]);
    assign layer1_out[730] = layer0_out[578];
    assign layer1_out[731] = layer0_out[314] & ~layer0_out[313];
    assign layer1_out[732] = ~layer0_out[392] | layer0_out[391];
    assign layer1_out[733] = ~layer0_out[618];
    assign layer1_out[734] = layer0_out[72];
    assign layer1_out[735] = ~layer0_out[312];
    assign layer1_out[736] = ~layer0_out[339] | layer0_out[338];
    assign layer1_out[737] = layer0_out[684] & ~layer0_out[683];
    assign layer1_out[738] = layer0_out[482] & ~layer0_out[481];
    assign layer1_out[739] = layer0_out[215] ^ layer0_out[216];
    assign layer1_out[740] = ~layer0_out[152];
    assign layer1_out[741] = ~layer0_out[373];
    assign layer1_out[742] = ~(layer0_out[654] & layer0_out[655]);
    assign layer1_out[743] = ~layer0_out[625];
    assign layer1_out[744] = layer0_out[181] & ~layer0_out[180];
    assign layer1_out[745] = ~layer0_out[575] | layer0_out[574];
    assign layer1_out[746] = ~(layer0_out[170] | layer0_out[171]);
    assign layer1_out[747] = layer0_out[83] & layer0_out[84];
    assign layer1_out[748] = ~layer0_out[53];
    assign layer1_out[749] = ~(layer0_out[63] & layer0_out[64]);
    assign layer1_out[750] = layer0_out[80];
    assign layer1_out[751] = layer0_out[444];
    assign layer1_out[752] = ~layer0_out[252] | layer0_out[253];
    assign layer1_out[753] = layer0_out[469] | layer0_out[470];
    assign layer1_out[754] = layer0_out[376] & layer0_out[377];
    assign layer1_out[755] = ~(layer0_out[780] ^ layer0_out[781]);
    assign layer1_out[756] = ~(layer0_out[578] ^ layer0_out[579]);
    assign layer1_out[757] = 1'b1;
    assign layer1_out[758] = layer0_out[526];
    assign layer1_out[759] = ~layer0_out[697];
    assign layer1_out[760] = layer0_out[434];
    assign layer1_out[761] = ~layer0_out[663];
    assign layer1_out[762] = layer0_out[186] & layer0_out[187];
    assign layer1_out[763] = ~layer0_out[753] | layer0_out[752];
    assign layer1_out[764] = ~layer0_out[455] | layer0_out[456];
    assign layer1_out[765] = ~layer0_out[768] | layer0_out[767];
    assign layer1_out[766] = layer0_out[501];
    assign layer1_out[767] = ~layer0_out[551];
    assign layer1_out[768] = layer0_out[273];
    assign layer1_out[769] = 1'b0;
    assign layer1_out[770] = layer0_out[238] & ~layer0_out[239];
    assign layer1_out[771] = 1'b1;
    assign layer1_out[772] = ~(layer0_out[431] & layer0_out[432]);
    assign layer1_out[773] = layer0_out[651] | layer0_out[652];
    assign layer1_out[774] = layer0_out[737] & ~layer0_out[736];
    assign layer1_out[775] = ~layer0_out[747];
    assign layer1_out[776] = ~layer0_out[331] | layer0_out[330];
    assign layer1_out[777] = layer0_out[494] | layer0_out[495];
    assign layer1_out[778] = ~(layer0_out[364] & layer0_out[365]);
    assign layer1_out[779] = layer0_out[35];
    assign layer1_out[780] = layer0_out[742] | layer0_out[743];
    assign layer1_out[781] = ~(layer0_out[304] & layer0_out[305]);
    assign layer1_out[782] = layer0_out[608] & ~layer0_out[607];
    assign layer1_out[783] = layer0_out[120] & layer0_out[121];
    assign layer1_out[784] = 1'b0;
    assign layer1_out[785] = layer0_out[180];
    assign layer1_out[786] = layer0_out[446];
    assign layer1_out[787] = layer0_out[412];
    assign layer1_out[788] = ~layer0_out[753] | layer0_out[754];
    assign layer1_out[789] = ~(layer0_out[628] & layer0_out[629]);
    assign layer1_out[790] = ~layer0_out[210];
    assign layer1_out[791] = ~layer0_out[284];
    assign layer1_out[792] = ~(layer0_out[543] | layer0_out[544]);
    assign layer1_out[793] = 1'b0;
    assign layer1_out[794] = layer0_out[576];
    assign layer1_out[795] = layer0_out[524];
    assign layer1_out[796] = layer0_out[347];
    assign layer1_out[797] = layer0_out[583] & ~layer0_out[582];
    assign layer1_out[798] = ~(layer0_out[383] | layer0_out[384]);
    assign layer1_out[799] = ~layer0_out[722];
    assign layer2_out[0] = layer1_out[169];
    assign layer2_out[1] = layer1_out[521] | layer1_out[522];
    assign layer2_out[2] = layer1_out[523];
    assign layer2_out[3] = ~layer1_out[147];
    assign layer2_out[4] = ~layer1_out[13];
    assign layer2_out[5] = ~layer1_out[197];
    assign layer2_out[6] = layer1_out[303] & ~layer1_out[302];
    assign layer2_out[7] = ~layer1_out[35];
    assign layer2_out[8] = layer1_out[717] ^ layer1_out[718];
    assign layer2_out[9] = ~layer1_out[203];
    assign layer2_out[10] = layer1_out[763];
    assign layer2_out[11] = layer1_out[480] & ~layer1_out[481];
    assign layer2_out[12] = layer1_out[10] & ~layer1_out[9];
    assign layer2_out[13] = layer1_out[617];
    assign layer2_out[14] = layer1_out[561] & ~layer1_out[560];
    assign layer2_out[15] = layer1_out[621] | layer1_out[622];
    assign layer2_out[16] = layer1_out[574];
    assign layer2_out[17] = layer1_out[74];
    assign layer2_out[18] = layer1_out[578];
    assign layer2_out[19] = layer1_out[794] & layer1_out[795];
    assign layer2_out[20] = 1'b0;
    assign layer2_out[21] = layer1_out[253];
    assign layer2_out[22] = ~layer1_out[753] | layer1_out[754];
    assign layer2_out[23] = ~layer1_out[589];
    assign layer2_out[24] = layer1_out[11];
    assign layer2_out[25] = layer1_out[46];
    assign layer2_out[26] = ~layer1_out[386] | layer1_out[385];
    assign layer2_out[27] = layer1_out[455];
    assign layer2_out[28] = layer1_out[384] & ~layer1_out[385];
    assign layer2_out[29] = ~layer1_out[312];
    assign layer2_out[30] = ~layer1_out[649] | layer1_out[650];
    assign layer2_out[31] = ~layer1_out[523];
    assign layer2_out[32] = layer1_out[400] & ~layer1_out[399];
    assign layer2_out[33] = layer1_out[469];
    assign layer2_out[34] = ~(layer1_out[742] ^ layer1_out[743]);
    assign layer2_out[35] = ~layer1_out[357];
    assign layer2_out[36] = ~layer1_out[548] | layer1_out[549];
    assign layer2_out[37] = ~(layer1_out[574] | layer1_out[575]);
    assign layer2_out[38] = ~layer1_out[612] | layer1_out[613];
    assign layer2_out[39] = ~layer1_out[352];
    assign layer2_out[40] = layer1_out[583];
    assign layer2_out[41] = layer1_out[494];
    assign layer2_out[42] = ~layer1_out[519];
    assign layer2_out[43] = ~layer1_out[275];
    assign layer2_out[44] = ~layer1_out[610];
    assign layer2_out[45] = layer1_out[676] & ~layer1_out[677];
    assign layer2_out[46] = ~(layer1_out[125] | layer1_out[126]);
    assign layer2_out[47] = layer1_out[632];
    assign layer2_out[48] = ~layer1_out[668] | layer1_out[667];
    assign layer2_out[49] = layer1_out[42] & ~layer1_out[41];
    assign layer2_out[50] = 1'b0;
    assign layer2_out[51] = ~layer1_out[406];
    assign layer2_out[52] = layer1_out[28];
    assign layer2_out[53] = layer1_out[150] & ~layer1_out[149];
    assign layer2_out[54] = ~layer1_out[109];
    assign layer2_out[55] = layer1_out[777];
    assign layer2_out[56] = layer1_out[162];
    assign layer2_out[57] = ~layer1_out[539] | layer1_out[538];
    assign layer2_out[58] = ~layer1_out[408] | layer1_out[409];
    assign layer2_out[59] = ~layer1_out[722];
    assign layer2_out[60] = ~layer1_out[8] | layer1_out[9];
    assign layer2_out[61] = ~(layer1_out[531] & layer1_out[532]);
    assign layer2_out[62] = ~layer1_out[709];
    assign layer2_out[63] = layer1_out[546];
    assign layer2_out[64] = ~(layer1_out[572] & layer1_out[573]);
    assign layer2_out[65] = ~layer1_out[715];
    assign layer2_out[66] = layer1_out[788];
    assign layer2_out[67] = layer1_out[231] & layer1_out[232];
    assign layer2_out[68] = layer1_out[260] & layer1_out[261];
    assign layer2_out[69] = layer1_out[40];
    assign layer2_out[70] = ~layer1_out[655];
    assign layer2_out[71] = ~layer1_out[21];
    assign layer2_out[72] = ~layer1_out[454];
    assign layer2_out[73] = layer1_out[414];
    assign layer2_out[74] = layer1_out[298] & ~layer1_out[299];
    assign layer2_out[75] = layer1_out[265] & layer1_out[266];
    assign layer2_out[76] = ~layer1_out[101];
    assign layer2_out[77] = layer1_out[127] | layer1_out[128];
    assign layer2_out[78] = ~layer1_out[339] | layer1_out[338];
    assign layer2_out[79] = layer1_out[55] & ~layer1_out[56];
    assign layer2_out[80] = ~layer1_out[318] | layer1_out[319];
    assign layer2_out[81] = layer1_out[380];
    assign layer2_out[82] = layer1_out[772] | layer1_out[773];
    assign layer2_out[83] = ~layer1_out[262];
    assign layer2_out[84] = ~layer1_out[674] | layer1_out[673];
    assign layer2_out[85] = layer1_out[238];
    assign layer2_out[86] = ~(layer1_out[177] | layer1_out[178]);
    assign layer2_out[87] = ~layer1_out[704] | layer1_out[703];
    assign layer2_out[88] = ~layer1_out[158];
    assign layer2_out[89] = ~layer1_out[693];
    assign layer2_out[90] = layer1_out[62] & layer1_out[63];
    assign layer2_out[91] = layer1_out[51];
    assign layer2_out[92] = layer1_out[508];
    assign layer2_out[93] = ~(layer1_out[192] | layer1_out[193]);
    assign layer2_out[94] = layer1_out[561] & ~layer1_out[562];
    assign layer2_out[95] = ~layer1_out[99];
    assign layer2_out[96] = ~(layer1_out[359] | layer1_out[360]);
    assign layer2_out[97] = ~layer1_out[750];
    assign layer2_out[98] = ~(layer1_out[234] & layer1_out[235]);
    assign layer2_out[99] = ~(layer1_out[691] & layer1_out[692]);
    assign layer2_out[100] = ~layer1_out[307];
    assign layer2_out[101] = ~layer1_out[413] | layer1_out[414];
    assign layer2_out[102] = layer1_out[397];
    assign layer2_out[103] = layer1_out[552] & layer1_out[553];
    assign layer2_out[104] = layer1_out[203];
    assign layer2_out[105] = layer1_out[294] & layer1_out[295];
    assign layer2_out[106] = layer1_out[306];
    assign layer2_out[107] = layer1_out[726] ^ layer1_out[727];
    assign layer2_out[108] = ~(layer1_out[550] & layer1_out[551]);
    assign layer2_out[109] = layer1_out[237];
    assign layer2_out[110] = layer1_out[118];
    assign layer2_out[111] = ~layer1_out[410] | layer1_out[409];
    assign layer2_out[112] = layer1_out[408] & ~layer1_out[407];
    assign layer2_out[113] = ~layer1_out[576];
    assign layer2_out[114] = layer1_out[614] & layer1_out[615];
    assign layer2_out[115] = ~(layer1_out[227] | layer1_out[228]);
    assign layer2_out[116] = layer1_out[112] & layer1_out[113];
    assign layer2_out[117] = ~layer1_out[790];
    assign layer2_out[118] = ~(layer1_out[547] & layer1_out[548]);
    assign layer2_out[119] = ~(layer1_out[438] ^ layer1_out[439]);
    assign layer2_out[120] = 1'b1;
    assign layer2_out[121] = layer1_out[186] & layer1_out[187];
    assign layer2_out[122] = layer1_out[84];
    assign layer2_out[123] = layer1_out[244] ^ layer1_out[245];
    assign layer2_out[124] = ~layer1_out[646];
    assign layer2_out[125] = layer1_out[103];
    assign layer2_out[126] = layer1_out[382];
    assign layer2_out[127] = ~layer1_out[639] | layer1_out[638];
    assign layer2_out[128] = layer1_out[595] & ~layer1_out[596];
    assign layer2_out[129] = ~(layer1_out[637] ^ layer1_out[638]);
    assign layer2_out[130] = ~layer1_out[389] | layer1_out[388];
    assign layer2_out[131] = ~layer1_out[2];
    assign layer2_out[132] = layer1_out[329] & ~layer1_out[328];
    assign layer2_out[133] = ~layer1_out[71];
    assign layer2_out[134] = layer1_out[157];
    assign layer2_out[135] = ~layer1_out[663] | layer1_out[662];
    assign layer2_out[136] = layer1_out[792] & ~layer1_out[793];
    assign layer2_out[137] = ~layer1_out[401];
    assign layer2_out[138] = layer1_out[580];
    assign layer2_out[139] = layer1_out[748];
    assign layer2_out[140] = layer1_out[76] & ~layer1_out[77];
    assign layer2_out[141] = layer1_out[717];
    assign layer2_out[142] = layer1_out[697] | layer1_out[698];
    assign layer2_out[143] = ~(layer1_out[382] ^ layer1_out[383]);
    assign layer2_out[144] = layer1_out[204] & layer1_out[205];
    assign layer2_out[145] = ~(layer1_out[527] & layer1_out[528]);
    assign layer2_out[146] = ~layer1_out[725];
    assign layer2_out[147] = ~layer1_out[75] | layer1_out[74];
    assign layer2_out[148] = layer1_out[245];
    assign layer2_out[149] = ~(layer1_out[445] & layer1_out[446]);
    assign layer2_out[150] = layer1_out[377];
    assign layer2_out[151] = layer1_out[189] & layer1_out[190];
    assign layer2_out[152] = layer1_out[776];
    assign layer2_out[153] = ~layer1_out[685];
    assign layer2_out[154] = ~layer1_out[640] | layer1_out[639];
    assign layer2_out[155] = layer1_out[487] | layer1_out[488];
    assign layer2_out[156] = layer1_out[140] ^ layer1_out[141];
    assign layer2_out[157] = layer1_out[609];
    assign layer2_out[158] = layer1_out[349] & ~layer1_out[348];
    assign layer2_out[159] = ~layer1_out[175];
    assign layer2_out[160] = ~layer1_out[82];
    assign layer2_out[161] = ~layer1_out[528];
    assign layer2_out[162] = 1'b1;
    assign layer2_out[163] = 1'b0;
    assign layer2_out[164] = ~layer1_out[526];
    assign layer2_out[165] = ~layer1_out[154];
    assign layer2_out[166] = layer1_out[3];
    assign layer2_out[167] = ~layer1_out[513];
    assign layer2_out[168] = layer1_out[708];
    assign layer2_out[169] = layer1_out[161];
    assign layer2_out[170] = ~layer1_out[259] | layer1_out[258];
    assign layer2_out[171] = layer1_out[276] & ~layer1_out[277];
    assign layer2_out[172] = ~layer1_out[173];
    assign layer2_out[173] = ~layer1_out[416];
    assign layer2_out[174] = layer1_out[133];
    assign layer2_out[175] = ~layer1_out[86];
    assign layer2_out[176] = ~layer1_out[40];
    assign layer2_out[177] = ~layer1_out[425];
    assign layer2_out[178] = layer1_out[664];
    assign layer2_out[179] = layer1_out[351];
    assign layer2_out[180] = layer1_out[456] & ~layer1_out[457];
    assign layer2_out[181] = layer1_out[667];
    assign layer2_out[182] = ~layer1_out[576];
    assign layer2_out[183] = ~layer1_out[446];
    assign layer2_out[184] = ~layer1_out[257];
    assign layer2_out[185] = ~(layer1_out[235] & layer1_out[236]);
    assign layer2_out[186] = ~layer1_out[741];
    assign layer2_out[187] = layer1_out[174];
    assign layer2_out[188] = ~(layer1_out[755] & layer1_out[756]);
    assign layer2_out[189] = ~layer1_out[679];
    assign layer2_out[190] = layer1_out[160] & layer1_out[161];
    assign layer2_out[191] = ~layer1_out[321];
    assign layer2_out[192] = ~layer1_out[300];
    assign layer2_out[193] = layer1_out[788];
    assign layer2_out[194] = layer1_out[305];
    assign layer2_out[195] = ~layer1_out[482];
    assign layer2_out[196] = ~layer1_out[186] | layer1_out[185];
    assign layer2_out[197] = ~layer1_out[444];
    assign layer2_out[198] = layer1_out[241];
    assign layer2_out[199] = layer1_out[581] & ~layer1_out[582];
    assign layer2_out[200] = layer1_out[361] | layer1_out[362];
    assign layer2_out[201] = 1'b1;
    assign layer2_out[202] = layer1_out[534] ^ layer1_out[535];
    assign layer2_out[203] = layer1_out[95];
    assign layer2_out[204] = 1'b1;
    assign layer2_out[205] = ~layer1_out[226];
    assign layer2_out[206] = layer1_out[89];
    assign layer2_out[207] = ~layer1_out[419];
    assign layer2_out[208] = ~layer1_out[313];
    assign layer2_out[209] = layer1_out[375];
    assign layer2_out[210] = layer1_out[620];
    assign layer2_out[211] = ~layer1_out[179];
    assign layer2_out[212] = ~layer1_out[354];
    assign layer2_out[213] = layer1_out[371];
    assign layer2_out[214] = layer1_out[760] & layer1_out[761];
    assign layer2_out[215] = layer1_out[97] & layer1_out[98];
    assign layer2_out[216] = ~(layer1_out[148] | layer1_out[149]);
    assign layer2_out[217] = layer1_out[616];
    assign layer2_out[218] = layer1_out[570];
    assign layer2_out[219] = layer1_out[423] | layer1_out[424];
    assign layer2_out[220] = layer1_out[263] ^ layer1_out[264];
    assign layer2_out[221] = layer1_out[108];
    assign layer2_out[222] = layer1_out[560];
    assign layer2_out[223] = ~layer1_out[124];
    assign layer2_out[224] = ~layer1_out[363];
    assign layer2_out[225] = ~layer1_out[35];
    assign layer2_out[226] = layer1_out[80];
    assign layer2_out[227] = layer1_out[124];
    assign layer2_out[228] = ~(layer1_out[596] & layer1_out[597]);
    assign layer2_out[229] = ~layer1_out[199] | layer1_out[200];
    assign layer2_out[230] = ~layer1_out[15];
    assign layer2_out[231] = ~layer1_out[593];
    assign layer2_out[232] = layer1_out[249];
    assign layer2_out[233] = ~layer1_out[510] | layer1_out[511];
    assign layer2_out[234] = 1'b0;
    assign layer2_out[235] = ~layer1_out[37] | layer1_out[36];
    assign layer2_out[236] = layer1_out[61] & layer1_out[62];
    assign layer2_out[237] = ~layer1_out[111];
    assign layer2_out[238] = ~layer1_out[452];
    assign layer2_out[239] = layer1_out[689] & ~layer1_out[690];
    assign layer2_out[240] = layer1_out[262];
    assign layer2_out[241] = ~(layer1_out[663] ^ layer1_out[664]);
    assign layer2_out[242] = layer1_out[777];
    assign layer2_out[243] = layer1_out[697];
    assign layer2_out[244] = ~layer1_out[44];
    assign layer2_out[245] = ~layer1_out[679];
    assign layer2_out[246] = ~layer1_out[31];
    assign layer2_out[247] = ~layer1_out[620];
    assign layer2_out[248] = layer1_out[590] & ~layer1_out[591];
    assign layer2_out[249] = ~layer1_out[701];
    assign layer2_out[250] = layer1_out[787] & ~layer1_out[786];
    assign layer2_out[251] = ~layer1_out[94];
    assign layer2_out[252] = ~layer1_out[479] | layer1_out[480];
    assign layer2_out[253] = layer1_out[284];
    assign layer2_out[254] = layer1_out[299];
    assign layer2_out[255] = 1'b0;
    assign layer2_out[256] = ~layer1_out[81];
    assign layer2_out[257] = ~layer1_out[23] | layer1_out[22];
    assign layer2_out[258] = ~(layer1_out[201] & layer1_out[202]);
    assign layer2_out[259] = layer1_out[72];
    assign layer2_out[260] = ~layer1_out[333];
    assign layer2_out[261] = ~layer1_out[395];
    assign layer2_out[262] = ~layer1_out[491];
    assign layer2_out[263] = layer1_out[150] | layer1_out[151];
    assign layer2_out[264] = layer1_out[714] & ~layer1_out[713];
    assign layer2_out[265] = ~layer1_out[430];
    assign layer2_out[266] = ~layer1_out[540];
    assign layer2_out[267] = layer1_out[90];
    assign layer2_out[268] = layer1_out[563] ^ layer1_out[564];
    assign layer2_out[269] = layer1_out[272] & ~layer1_out[271];
    assign layer2_out[270] = ~layer1_out[402];
    assign layer2_out[271] = ~layer1_out[84];
    assign layer2_out[272] = ~layer1_out[635];
    assign layer2_out[273] = ~layer1_out[468];
    assign layer2_out[274] = ~layer1_out[63] | layer1_out[64];
    assign layer2_out[275] = layer1_out[457] & layer1_out[458];
    assign layer2_out[276] = ~layer1_out[696];
    assign layer2_out[277] = ~(layer1_out[6] | layer1_out[7]);
    assign layer2_out[278] = layer1_out[649];
    assign layer2_out[279] = ~layer1_out[402] | layer1_out[401];
    assign layer2_out[280] = layer1_out[658] & layer1_out[659];
    assign layer2_out[281] = layer1_out[136] & layer1_out[137];
    assign layer2_out[282] = ~(layer1_out[601] & layer1_out[602]);
    assign layer2_out[283] = layer1_out[66] ^ layer1_out[67];
    assign layer2_out[284] = 1'b0;
    assign layer2_out[285] = layer1_out[339] & ~layer1_out[340];
    assign layer2_out[286] = layer1_out[752] & ~layer1_out[751];
    assign layer2_out[287] = layer1_out[323] & layer1_out[324];
    assign layer2_out[288] = ~layer1_out[320];
    assign layer2_out[289] = layer1_out[228] & ~layer1_out[229];
    assign layer2_out[290] = ~layer1_out[145];
    assign layer2_out[291] = ~layer1_out[441];
    assign layer2_out[292] = layer1_out[129] & ~layer1_out[130];
    assign layer2_out[293] = layer1_out[50];
    assign layer2_out[294] = layer1_out[749] & layer1_out[750];
    assign layer2_out[295] = 1'b1;
    assign layer2_out[296] = ~layer1_out[747];
    assign layer2_out[297] = ~(layer1_out[360] ^ layer1_out[361]);
    assign layer2_out[298] = layer1_out[210];
    assign layer2_out[299] = layer1_out[108];
    assign layer2_out[300] = ~layer1_out[121];
    assign layer2_out[301] = ~layer1_out[541];
    assign layer2_out[302] = layer1_out[488] ^ layer1_out[489];
    assign layer2_out[303] = ~layer1_out[477];
    assign layer2_out[304] = layer1_out[213] | layer1_out[214];
    assign layer2_out[305] = layer1_out[466];
    assign layer2_out[306] = layer1_out[691];
    assign layer2_out[307] = ~layer1_out[587];
    assign layer2_out[308] = ~(layer1_out[60] & layer1_out[61]);
    assign layer2_out[309] = ~(layer1_out[10] | layer1_out[11]);
    assign layer2_out[310] = ~layer1_out[294];
    assign layer2_out[311] = ~layer1_out[551] | layer1_out[552];
    assign layer2_out[312] = ~(layer1_out[762] & layer1_out[763]);
    assign layer2_out[313] = layer1_out[75];
    assign layer2_out[314] = layer1_out[298];
    assign layer2_out[315] = ~layer1_out[380];
    assign layer2_out[316] = ~(layer1_out[699] | layer1_out[700]);
    assign layer2_out[317] = layer1_out[760];
    assign layer2_out[318] = 1'b0;
    assign layer2_out[319] = ~(layer1_out[494] & layer1_out[495]);
    assign layer2_out[320] = ~layer1_out[47];
    assign layer2_out[321] = ~layer1_out[641];
    assign layer2_out[322] = ~(layer1_out[774] & layer1_out[775]);
    assign layer2_out[323] = layer1_out[292];
    assign layer2_out[324] = layer1_out[378];
    assign layer2_out[325] = layer1_out[651] & ~layer1_out[652];
    assign layer2_out[326] = layer1_out[754];
    assign layer2_out[327] = ~layer1_out[419];
    assign layer2_out[328] = ~(layer1_out[246] | layer1_out[247]);
    assign layer2_out[329] = layer1_out[420] | layer1_out[421];
    assign layer2_out[330] = layer1_out[330];
    assign layer2_out[331] = 1'b1;
    assign layer2_out[332] = layer1_out[643] | layer1_out[644];
    assign layer2_out[333] = ~layer1_out[646];
    assign layer2_out[334] = ~layer1_out[226];
    assign layer2_out[335] = layer1_out[180];
    assign layer2_out[336] = ~layer1_out[747];
    assign layer2_out[337] = ~layer1_out[768] | layer1_out[769];
    assign layer2_out[338] = ~layer1_out[284];
    assign layer2_out[339] = layer1_out[467];
    assign layer2_out[340] = ~layer1_out[90];
    assign layer2_out[341] = ~(layer1_out[790] & layer1_out[791]);
    assign layer2_out[342] = layer1_out[16] & ~layer1_out[17];
    assign layer2_out[343] = ~layer1_out[297];
    assign layer2_out[344] = ~layer1_out[619];
    assign layer2_out[345] = layer1_out[524] ^ layer1_out[525];
    assign layer2_out[346] = layer1_out[252] | layer1_out[253];
    assign layer2_out[347] = ~layer1_out[492] | layer1_out[493];
    assign layer2_out[348] = ~layer1_out[593];
    assign layer2_out[349] = ~layer1_out[116] | layer1_out[117];
    assign layer2_out[350] = ~layer1_out[602];
    assign layer2_out[351] = ~layer1_out[782];
    assign layer2_out[352] = ~layer1_out[384];
    assign layer2_out[353] = layer1_out[222];
    assign layer2_out[354] = layer1_out[589];
    assign layer2_out[355] = layer1_out[442] & layer1_out[443];
    assign layer2_out[356] = ~layer1_out[13];
    assign layer2_out[357] = ~layer1_out[766];
    assign layer2_out[358] = layer1_out[753];
    assign layer2_out[359] = layer1_out[792];
    assign layer2_out[360] = layer1_out[734];
    assign layer2_out[361] = ~layer1_out[544] | layer1_out[543];
    assign layer2_out[362] = 1'b1;
    assign layer2_out[363] = layer1_out[310] & layer1_out[311];
    assign layer2_out[364] = ~layer1_out[240] | layer1_out[241];
    assign layer2_out[365] = layer1_out[28] ^ layer1_out[29];
    assign layer2_out[366] = layer1_out[629] ^ layer1_out[630];
    assign layer2_out[367] = layer1_out[144];
    assign layer2_out[368] = 1'b1;
    assign layer2_out[369] = ~(layer1_out[52] | layer1_out[53]);
    assign layer2_out[370] = layer1_out[411];
    assign layer2_out[371] = ~layer1_out[231] | layer1_out[230];
    assign layer2_out[372] = ~layer1_out[628];
    assign layer2_out[373] = layer1_out[734] & ~layer1_out[733];
    assign layer2_out[374] = ~layer1_out[398];
    assign layer2_out[375] = ~layer1_out[142];
    assign layer2_out[376] = ~(layer1_out[266] | layer1_out[267]);
    assign layer2_out[377] = layer1_out[222];
    assign layer2_out[378] = ~(layer1_out[448] | layer1_out[449]);
    assign layer2_out[379] = layer1_out[426] | layer1_out[427];
    assign layer2_out[380] = ~(layer1_out[264] & layer1_out[265]);
    assign layer2_out[381] = ~(layer1_out[295] ^ layer1_out[296]);
    assign layer2_out[382] = ~layer1_out[485];
    assign layer2_out[383] = ~layer1_out[623] | layer1_out[624];
    assign layer2_out[384] = layer1_out[530] | layer1_out[531];
    assign layer2_out[385] = ~layer1_out[234];
    assign layer2_out[386] = layer1_out[411] ^ layer1_out[412];
    assign layer2_out[387] = layer1_out[146] & layer1_out[147];
    assign layer2_out[388] = ~(layer1_out[490] | layer1_out[491]);
    assign layer2_out[389] = ~layer1_out[516] | layer1_out[517];
    assign layer2_out[390] = ~layer1_out[721];
    assign layer2_out[391] = layer1_out[489] & layer1_out[490];
    assign layer2_out[392] = ~(layer1_out[314] ^ layer1_out[315]);
    assign layer2_out[393] = layer1_out[343];
    assign layer2_out[394] = ~layer1_out[196];
    assign layer2_out[395] = layer1_out[344];
    assign layer2_out[396] = ~layer1_out[287];
    assign layer2_out[397] = layer1_out[770] & ~layer1_out[771];
    assign layer2_out[398] = layer1_out[24];
    assign layer2_out[399] = ~layer1_out[687] | layer1_out[686];
    assign layer2_out[400] = ~layer1_out[669];
    assign layer2_out[401] = layer1_out[29] & ~layer1_out[30];
    assign layer2_out[402] = ~layer1_out[200];
    assign layer2_out[403] = layer1_out[137];
    assign layer2_out[404] = layer1_out[693];
    assign layer2_out[405] = layer1_out[683] & ~layer1_out[684];
    assign layer2_out[406] = ~layer1_out[217] | layer1_out[216];
    assign layer2_out[407] = layer1_out[675] | layer1_out[676];
    assign layer2_out[408] = layer1_out[440];
    assign layer2_out[409] = layer1_out[277];
    assign layer2_out[410] = layer1_out[595];
    assign layer2_out[411] = layer1_out[331] | layer1_out[332];
    assign layer2_out[412] = ~layer1_out[310] | layer1_out[309];
    assign layer2_out[413] = ~(layer1_out[415] | layer1_out[416]);
    assign layer2_out[414] = layer1_out[212] ^ layer1_out[213];
    assign layer2_out[415] = ~layer1_out[181];
    assign layer2_out[416] = ~layer1_out[159];
    assign layer2_out[417] = ~layer1_out[303] | layer1_out[304];
    assign layer2_out[418] = ~layer1_out[6];
    assign layer2_out[419] = layer1_out[131] | layer1_out[132];
    assign layer2_out[420] = layer1_out[238];
    assign layer2_out[421] = layer1_out[346];
    assign layer2_out[422] = ~layer1_out[629];
    assign layer2_out[423] = ~layer1_out[727] | layer1_out[728];
    assign layer2_out[424] = layer1_out[497];
    assign layer2_out[425] = layer1_out[270];
    assign layer2_out[426] = ~layer1_out[7];
    assign layer2_out[427] = ~layer1_out[642] | layer1_out[641];
    assign layer2_out[428] = layer1_out[58];
    assign layer2_out[429] = ~layer1_out[519];
    assign layer2_out[430] = ~layer1_out[534];
    assign layer2_out[431] = layer1_out[329] | layer1_out[330];
    assign layer2_out[432] = layer1_out[726];
    assign layer2_out[433] = ~(layer1_out[362] & layer1_out[363]);
    assign layer2_out[434] = layer1_out[229];
    assign layer2_out[435] = ~(layer1_out[390] | layer1_out[391]);
    assign layer2_out[436] = layer1_out[343];
    assign layer2_out[437] = ~layer1_out[406];
    assign layer2_out[438] = ~layer1_out[25] | layer1_out[26];
    assign layer2_out[439] = ~layer1_out[538];
    assign layer2_out[440] = ~layer1_out[508];
    assign layer2_out[441] = layer1_out[553];
    assign layer2_out[442] = ~layer1_out[671];
    assign layer2_out[443] = layer1_out[501];
    assign layer2_out[444] = ~layer1_out[737];
    assign layer2_out[445] = ~(layer1_out[657] ^ layer1_out[658]);
    assign layer2_out[446] = layer1_out[504] ^ layer1_out[505];
    assign layer2_out[447] = ~layer1_out[437] | layer1_out[436];
    assign layer2_out[448] = layer1_out[332];
    assign layer2_out[449] = ~layer1_out[433];
    assign layer2_out[450] = layer1_out[163] | layer1_out[164];
    assign layer2_out[451] = ~(layer1_out[43] | layer1_out[44]);
    assign layer2_out[452] = ~layer1_out[661];
    assign layer2_out[453] = ~(layer1_out[356] | layer1_out[357]);
    assign layer2_out[454] = ~layer1_out[273];
    assign layer2_out[455] = layer1_out[554];
    assign layer2_out[456] = layer1_out[556];
    assign layer2_out[457] = ~(layer1_out[656] & layer1_out[657]);
    assign layer2_out[458] = layer1_out[249];
    assign layer2_out[459] = layer1_out[68];
    assign layer2_out[460] = ~layer1_out[283] | layer1_out[282];
    assign layer2_out[461] = ~layer1_out[460];
    assign layer2_out[462] = ~(layer1_out[665] ^ layer1_out[666]);
    assign layer2_out[463] = layer1_out[432] | layer1_out[433];
    assign layer2_out[464] = ~layer1_out[293] | layer1_out[292];
    assign layer2_out[465] = 1'b1;
    assign layer2_out[466] = ~layer1_out[138];
    assign layer2_out[467] = layer1_out[723] & ~layer1_out[724];
    assign layer2_out[468] = ~layer1_out[316];
    assign layer2_out[469] = layer1_out[218];
    assign layer2_out[470] = layer1_out[707];
    assign layer2_out[471] = layer1_out[106] & ~layer1_out[107];
    assign layer2_out[472] = layer1_out[68];
    assign layer2_out[473] = ~layer1_out[38];
    assign layer2_out[474] = ~layer1_out[140];
    assign layer2_out[475] = ~layer1_out[223] | layer1_out[224];
    assign layer2_out[476] = layer1_out[197];
    assign layer2_out[477] = layer1_out[606];
    assign layer2_out[478] = layer1_out[688];
    assign layer2_out[479] = layer1_out[737];
    assign layer2_out[480] = layer1_out[514];
    assign layer2_out[481] = ~layer1_out[732];
    assign layer2_out[482] = 1'b0;
    assign layer2_out[483] = layer1_out[454] | layer1_out[455];
    assign layer2_out[484] = ~(layer1_out[535] | layer1_out[536]);
    assign layer2_out[485] = layer1_out[761];
    assign layer2_out[486] = layer1_out[64] ^ layer1_out[65];
    assign layer2_out[487] = layer1_out[606];
    assign layer2_out[488] = ~layer1_out[17] | layer1_out[18];
    assign layer2_out[489] = ~layer1_out[387] | layer1_out[388];
    assign layer2_out[490] = layer1_out[260];
    assign layer2_out[491] = ~(layer1_out[472] | layer1_out[473]);
    assign layer2_out[492] = ~(layer1_out[624] | layer1_out[625]);
    assign layer2_out[493] = ~layer1_out[732] | layer1_out[731];
    assign layer2_out[494] = ~(layer1_out[568] & layer1_out[569]);
    assign layer2_out[495] = ~layer1_out[325];
    assign layer2_out[496] = layer1_out[757] & ~layer1_out[756];
    assign layer2_out[497] = ~layer1_out[256] | layer1_out[257];
    assign layer2_out[498] = layer1_out[481];
    assign layer2_out[499] = ~layer1_out[367] | layer1_out[366];
    assign layer2_out[500] = layer1_out[705];
    assign layer2_out[501] = layer1_out[187] & layer1_out[188];
    assign layer2_out[502] = layer1_out[118];
    assign layer2_out[503] = ~layer1_out[559];
    assign layer2_out[504] = layer1_out[2];
    assign layer2_out[505] = layer1_out[623];
    assign layer2_out[506] = layer1_out[466] | layer1_out[467];
    assign layer2_out[507] = layer1_out[633];
    assign layer2_out[508] = ~layer1_out[86];
    assign layer2_out[509] = ~(layer1_out[544] & layer1_out[545]);
    assign layer2_out[510] = layer1_out[171] ^ layer1_out[172];
    assign layer2_out[511] = ~layer1_out[169];
    assign layer2_out[512] = ~layer1_out[182];
    assign layer2_out[513] = layer1_out[744];
    assign layer2_out[514] = layer1_out[70];
    assign layer2_out[515] = layer1_out[336];
    assign layer2_out[516] = layer1_out[678] & ~layer1_out[677];
    assign layer2_out[517] = ~layer1_out[405];
    assign layer2_out[518] = layer1_out[317];
    assign layer2_out[519] = layer1_out[214] & layer1_out[215];
    assign layer2_out[520] = ~layer1_out[364] | layer1_out[365];
    assign layer2_out[521] = layer1_out[479] & ~layer1_out[478];
    assign layer2_out[522] = layer1_out[212] & ~layer1_out[211];
    assign layer2_out[523] = layer1_out[126] | layer1_out[127];
    assign layer2_out[524] = layer1_out[571];
    assign layer2_out[525] = ~layer1_out[289];
    assign layer2_out[526] = layer1_out[275];
    assign layer2_out[527] = ~layer1_out[474];
    assign layer2_out[528] = layer1_out[255] | layer1_out[256];
    assign layer2_out[529] = layer1_out[704] & ~layer1_out[705];
    assign layer2_out[530] = ~(layer1_out[142] ^ layer1_out[143]);
    assign layer2_out[531] = layer1_out[105] & ~layer1_out[106];
    assign layer2_out[532] = layer1_out[604];
    assign layer2_out[533] = layer1_out[386] | layer1_out[387];
    assign layer2_out[534] = layer1_out[476];
    assign layer2_out[535] = ~layer1_out[555] | layer1_out[556];
    assign layer2_out[536] = layer1_out[741] & ~layer1_out[740];
    assign layer2_out[537] = layer1_out[453];
    assign layer2_out[538] = ~(layer1_out[767] ^ layer1_out[768]);
    assign layer2_out[539] = layer1_out[499] & ~layer1_out[500];
    assign layer2_out[540] = ~(layer1_out[701] ^ layer1_out[702]);
    assign layer2_out[541] = ~layer1_out[568];
    assign layer2_out[542] = layer1_out[321] & ~layer1_out[320];
    assign layer2_out[543] = ~layer1_out[653];
    assign layer2_out[544] = ~layer1_out[199];
    assign layer2_out[545] = ~layer1_out[778] | layer1_out[779];
    assign layer2_out[546] = ~layer1_out[33];
    assign layer2_out[547] = ~layer1_out[122];
    assign layer2_out[548] = layer1_out[393] | layer1_out[394];
    assign layer2_out[549] = layer1_out[119] & ~layer1_out[120];
    assign layer2_out[550] = layer1_out[758];
    assign layer2_out[551] = layer1_out[647];
    assign layer2_out[552] = ~layer1_out[49] | layer1_out[50];
    assign layer2_out[553] = layer1_out[267];
    assign layer2_out[554] = ~layer1_out[435] | layer1_out[436];
    assign layer2_out[555] = layer1_out[207];
    assign layer2_out[556] = layer1_out[375] & ~layer1_out[374];
    assign layer2_out[557] = layer1_out[14] | layer1_out[15];
    assign layer2_out[558] = ~layer1_out[33];
    assign layer2_out[559] = layer1_out[473];
    assign layer2_out[560] = layer1_out[243] | layer1_out[244];
    assign layer2_out[561] = ~layer1_out[96];
    assign layer2_out[562] = layer1_out[26] & layer1_out[27];
    assign layer2_out[563] = ~(layer1_out[373] | layer1_out[374]);
    assign layer2_out[564] = layer1_out[171];
    assign layer2_out[565] = ~layer1_out[517];
    assign layer2_out[566] = layer1_out[133];
    assign layer2_out[567] = ~layer1_out[428];
    assign layer2_out[568] = layer1_out[643];
    assign layer2_out[569] = layer1_out[671];
    assign layer2_out[570] = ~layer1_out[287];
    assign layer2_out[571] = ~layer1_out[4];
    assign layer2_out[572] = layer1_out[680] | layer1_out[681];
    assign layer2_out[573] = 1'b0;
    assign layer2_out[574] = layer1_out[254];
    assign layer2_out[575] = layer1_out[87] | layer1_out[88];
    assign layer2_out[576] = ~layer1_out[685] | layer1_out[684];
    assign layer2_out[577] = layer1_out[598];
    assign layer2_out[578] = layer1_out[120];
    assign layer2_out[579] = layer1_out[191] & ~layer1_out[190];
    assign layer2_out[580] = layer1_out[308];
    assign layer2_out[581] = ~layer1_out[506];
    assign layer2_out[582] = layer1_out[437] & layer1_out[438];
    assign layer2_out[583] = layer1_out[772];
    assign layer2_out[584] = layer1_out[48] & ~layer1_out[47];
    assign layer2_out[585] = layer1_out[215] & layer1_out[216];
    assign layer2_out[586] = layer1_out[654] ^ layer1_out[655];
    assign layer2_out[587] = ~layer1_out[55];
    assign layer2_out[588] = ~layer1_out[325] | layer1_out[326];
    assign layer2_out[589] = layer1_out[219] & layer1_out[220];
    assign layer2_out[590] = layer1_out[464] & ~layer1_out[463];
    assign layer2_out[591] = layer1_out[720];
    assign layer2_out[592] = ~(layer1_out[417] & layer1_out[418]);
    assign layer2_out[593] = ~layer1_out[281];
    assign layer2_out[594] = layer1_out[529] | layer1_out[530];
    assign layer2_out[595] = layer1_out[765] | layer1_out[766];
    assign layer2_out[596] = layer1_out[521];
    assign layer2_out[597] = ~(layer1_out[184] ^ layer1_out[185]);
    assign layer2_out[598] = layer1_out[434];
    assign layer2_out[599] = ~(layer1_out[506] & layer1_out[507]);
    assign layer2_out[600] = ~layer1_out[308];
    assign layer2_out[601] = ~(layer1_out[709] | layer1_out[710]);
    assign layer2_out[602] = layer1_out[396] & ~layer1_out[395];
    assign layer2_out[603] = ~layer1_out[314] | layer1_out[313];
    assign layer2_out[604] = ~(layer1_out[353] | layer1_out[354]);
    assign layer2_out[605] = ~(layer1_out[422] | layer1_out[423]);
    assign layer2_out[606] = ~layer1_out[19];
    assign layer2_out[607] = layer1_out[515] ^ layer1_out[516];
    assign layer2_out[608] = layer1_out[248];
    assign layer2_out[609] = layer1_out[358] | layer1_out[359];
    assign layer2_out[610] = layer1_out[786] & ~layer1_out[785];
    assign layer2_out[611] = layer1_out[567];
    assign layer2_out[612] = ~layer1_out[472];
    assign layer2_out[613] = ~layer1_out[630] | layer1_out[631];
    assign layer2_out[614] = ~layer1_out[674] | layer1_out[675];
    assign layer2_out[615] = layer1_out[347] ^ layer1_out[348];
    assign layer2_out[616] = layer1_out[798];
    assign layer2_out[617] = layer1_out[368];
    assign layer2_out[618] = layer1_out[351];
    assign layer2_out[619] = ~layer1_out[153] | layer1_out[152];
    assign layer2_out[620] = layer1_out[626];
    assign layer2_out[621] = ~layer1_out[430];
    assign layer2_out[622] = layer1_out[115] | layer1_out[116];
    assign layer2_out[623] = ~layer1_out[376];
    assign layer2_out[624] = layer1_out[644];
    assign layer2_out[625] = layer1_out[584] & layer1_out[585];
    assign layer2_out[626] = ~layer1_out[156] | layer1_out[155];
    assign layer2_out[627] = ~(layer1_out[42] | layer1_out[43]);
    assign layer2_out[628] = ~layer1_out[672] | layer1_out[673];
    assign layer2_out[629] = ~layer1_out[165];
    assign layer2_out[630] = layer1_out[206] & ~layer1_out[205];
    assign layer2_out[631] = layer1_out[565] | layer1_out[566];
    assign layer2_out[632] = layer1_out[695];
    assign layer2_out[633] = layer1_out[440];
    assign layer2_out[634] = ~layer1_out[167];
    assign layer2_out[635] = layer1_out[209];
    assign layer2_out[636] = ~layer1_out[502] | layer1_out[503];
    assign layer2_out[637] = ~layer1_out[659];
    assign layer2_out[638] = ~layer1_out[422];
    assign layer2_out[639] = layer1_out[81];
    assign layer2_out[640] = ~layer1_out[731];
    assign layer2_out[641] = ~layer1_out[546];
    assign layer2_out[642] = ~(layer1_out[94] | layer1_out[95]);
    assign layer2_out[643] = layer1_out[65] & layer1_out[66];
    assign layer2_out[644] = ~layer1_out[22];
    assign layer2_out[645] = layer1_out[740];
    assign layer2_out[646] = layer1_out[650] | layer1_out[651];
    assign layer2_out[647] = layer1_out[718];
    assign layer2_out[648] = layer1_out[779] | layer1_out[780];
    assign layer2_out[649] = ~layer1_out[349];
    assign layer2_out[650] = layer1_out[532];
    assign layer2_out[651] = layer1_out[633] ^ layer1_out[634];
    assign layer2_out[652] = ~(layer1_out[176] | layer1_out[177]);
    assign layer2_out[653] = ~layer1_out[154];
    assign layer2_out[654] = ~layer1_out[501];
    assign layer2_out[655] = layer1_out[450];
    assign layer2_out[656] = ~layer1_out[611] | layer1_out[612];
    assign layer2_out[657] = ~layer1_out[688];
    assign layer2_out[658] = layer1_out[412] & ~layer1_out[413];
    assign layer2_out[659] = ~layer1_out[728] | layer1_out[729];
    assign layer2_out[660] = ~(layer1_out[250] & layer1_out[251]);
    assign layer2_out[661] = ~layer1_out[785];
    assign layer2_out[662] = ~layer1_out[240];
    assign layer2_out[663] = ~layer1_out[114];
    assign layer2_out[664] = ~layer1_out[290];
    assign layer2_out[665] = layer1_out[372];
    assign layer2_out[666] = ~layer1_out[77];
    assign layer2_out[667] = 1'b1;
    assign layer2_out[668] = ~layer1_out[404] | layer1_out[403];
    assign layer2_out[669] = layer1_out[463];
    assign layer2_out[670] = layer1_out[562];
    assign layer2_out[671] = ~(layer1_out[322] & layer1_out[323]);
    assign layer2_out[672] = ~layer1_out[2];
    assign layer2_out[673] = layer1_out[37] & layer1_out[38];
    assign layer2_out[674] = layer1_out[337];
    assign layer2_out[675] = ~(layer1_out[58] & layer1_out[59]);
    assign layer2_out[676] = ~layer1_out[795];
    assign layer2_out[677] = ~(layer1_out[316] ^ layer1_out[317]);
    assign layer2_out[678] = ~(layer1_out[232] & layer1_out[233]);
    assign layer2_out[679] = ~layer1_out[511];
    assign layer2_out[680] = ~layer1_out[782] | layer1_out[783];
    assign layer2_out[681] = layer1_out[208] & ~layer1_out[207];
    assign layer2_out[682] = ~layer1_out[334];
    assign layer2_out[683] = layer1_out[591];
    assign layer2_out[684] = ~layer1_out[286];
    assign layer2_out[685] = ~layer1_out[543];
    assign layer2_out[686] = layer1_out[24];
    assign layer2_out[687] = ~layer1_out[537] | layer1_out[536];
    assign layer2_out[688] = ~(layer1_out[135] & layer1_out[136]);
    assign layer2_out[689] = ~layer1_out[570];
    assign layer2_out[690] = layer1_out[653];
    assign layer2_out[691] = layer1_out[145];
    assign layer2_out[692] = layer1_out[503];
    assign layer2_out[693] = layer1_out[134];
    assign layer2_out[694] = ~layer1_out[290];
    assign layer2_out[695] = ~layer1_out[613];
    assign layer2_out[696] = ~layer1_out[72];
    assign layer2_out[697] = layer1_out[798] & ~layer1_out[797];
    assign layer2_out[698] = ~layer1_out[131];
    assign layer2_out[699] = layer1_out[91] | layer1_out[92];
    assign layer2_out[700] = layer1_out[495];
    assign layer2_out[701] = ~layer1_out[425] | layer1_out[424];
    assign layer2_out[702] = layer1_out[191];
    assign layer2_out[703] = layer1_out[765];
    assign layer2_out[704] = ~layer1_out[342] | layer1_out[341];
    assign layer2_out[705] = ~layer1_out[188];
    assign layer2_out[706] = ~layer1_out[744];
    assign layer2_out[707] = layer1_out[781];
    assign layer2_out[708] = layer1_out[736] & ~layer1_out[735];
    assign layer2_out[709] = ~(layer1_out[242] ^ layer1_out[243]);
    assign layer2_out[710] = layer1_out[165] & ~layer1_out[166];
    assign layer2_out[711] = ~layer1_out[56];
    assign layer2_out[712] = ~layer1_out[193];
    assign layer2_out[713] = ~layer1_out[475];
    assign layer2_out[714] = layer1_out[783] ^ layer1_out[784];
    assign layer2_out[715] = layer1_out[484];
    assign layer2_out[716] = layer1_out[103];
    assign layer2_out[717] = layer1_out[715] | layer1_out[716];
    assign layer2_out[718] = layer1_out[345];
    assign layer2_out[719] = ~layer1_out[512];
    assign layer2_out[720] = ~layer1_out[391];
    assign layer2_out[721] = ~layer1_out[184] | layer1_out[183];
    assign layer2_out[722] = layer1_out[151] | layer1_out[152];
    assign layer2_out[723] = ~layer1_out[712];
    assign layer2_out[724] = ~layer1_out[156] | layer1_out[157];
    assign layer2_out[725] = layer1_out[278] & ~layer1_out[279];
    assign layer2_out[726] = layer1_out[599] | layer1_out[600];
    assign layer2_out[727] = ~layer1_out[712];
    assign layer2_out[728] = layer1_out[273] | layer1_out[274];
    assign layer2_out[729] = layer1_out[509] & layer1_out[510];
    assign layer2_out[730] = layer1_out[796];
    assign layer2_out[731] = layer1_out[100];
    assign layer2_out[732] = ~layer1_out[195] | layer1_out[194];
    assign layer2_out[733] = layer1_out[600];
    assign layer2_out[734] = layer1_out[451];
    assign layer2_out[735] = ~layer1_out[0];
    assign layer2_out[736] = ~layer1_out[48];
    assign layer2_out[737] = layer1_out[183];
    assign layer2_out[738] = layer1_out[462];
    assign layer2_out[739] = layer1_out[746];
    assign layer2_out[740] = layer1_out[588];
    assign layer2_out[741] = ~layer1_out[341] | layer1_out[340];
    assign layer2_out[742] = layer1_out[662] & ~layer1_out[661];
    assign layer2_out[743] = layer1_out[636];
    assign layer2_out[744] = layer1_out[759] & ~layer1_out[758];
    assign layer2_out[745] = ~layer1_out[730] | layer1_out[729];
    assign layer2_out[746] = layer1_out[371] & ~layer1_out[372];
    assign layer2_out[747] = ~layer1_out[392] | layer1_out[393];
    assign layer2_out[748] = ~layer1_out[698];
    assign layer2_out[749] = ~layer1_out[269];
    assign layer2_out[750] = 1'b0;
    assign layer2_out[751] = ~layer1_out[110];
    assign layer2_out[752] = ~layer1_out[269];
    assign layer2_out[753] = layer1_out[550] & ~layer1_out[549];
    assign layer2_out[754] = layer1_out[458] & ~layer1_out[459];
    assign layer2_out[755] = layer1_out[738] & layer1_out[739];
    assign layer2_out[756] = ~(layer1_out[217] & layer1_out[218]);
    assign layer2_out[757] = ~layer1_out[487];
    assign layer2_out[758] = layer1_out[93];
    assign layer2_out[759] = ~(layer1_out[604] | layer1_out[605]);
    assign layer2_out[760] = ~(layer1_out[365] & layer1_out[366]);
    assign layer2_out[761] = layer1_out[208] & ~layer1_out[209];
    assign layer2_out[762] = layer1_out[668] & layer1_out[669];
    assign layer2_out[763] = ~layer1_out[128];
    assign layer2_out[764] = layer1_out[20];
    assign layer2_out[765] = layer1_out[607] & ~layer1_out[608];
    assign layer2_out[766] = ~(layer1_out[578] | layer1_out[579]);
    assign layer2_out[767] = ~layer1_out[356];
    assign layer2_out[768] = layer1_out[586];
    assign layer2_out[769] = layer1_out[448];
    assign layer2_out[770] = layer1_out[390];
    assign layer2_out[771] = layer1_out[397];
    assign layer2_out[772] = layer1_out[626] & ~layer1_out[625];
    assign layer2_out[773] = layer1_out[681] | layer1_out[682];
    assign layer2_out[774] = layer1_out[101];
    assign layer2_out[775] = ~(layer1_out[443] | layer1_out[444]);
    assign layer2_out[776] = ~layer1_out[682];
    assign layer2_out[777] = layer1_out[336];
    assign layer2_out[778] = layer1_out[30];
    assign layer2_out[779] = ~layer1_out[78];
    assign layer2_out[780] = layer1_out[173];
    assign layer2_out[781] = layer1_out[498];
    assign layer2_out[782] = ~layer1_out[221] | layer1_out[220];
    assign layer2_out[783] = ~layer1_out[635];
    assign layer2_out[784] = ~(layer1_out[557] | layer1_out[558]);
    assign layer2_out[785] = layer1_out[224];
    assign layer2_out[786] = ~(layer1_out[104] & layer1_out[105]);
    assign layer2_out[787] = ~layer1_out[432];
    assign layer2_out[788] = layer1_out[497];
    assign layer2_out[789] = ~layer1_out[54];
    assign layer2_out[790] = ~layer1_out[580];
    assign layer2_out[791] = ~layer1_out[711];
    assign layer2_out[792] = layer1_out[598];
    assign layer2_out[793] = ~layer1_out[370];
    assign layer2_out[794] = ~layer1_out[428];
    assign layer2_out[795] = layer1_out[793] & ~layer1_out[794];
    assign layer2_out[796] = ~layer1_out[461];
    assign layer2_out[797] = ~(layer1_out[525] | layer1_out[526]);
    assign layer2_out[798] = ~(layer1_out[59] ^ layer1_out[60]);
    assign layer2_out[799] = layer1_out[281] & ~layer1_out[282];
    assign layer3_out[0] = layer2_out[495];
    assign layer3_out[1] = layer2_out[124];
    assign layer3_out[2] = layer2_out[115] & ~layer2_out[116];
    assign layer3_out[3] = layer2_out[737];
    assign layer3_out[4] = layer2_out[344];
    assign layer3_out[5] = layer2_out[203];
    assign layer3_out[6] = layer2_out[7];
    assign layer3_out[7] = ~layer2_out[649];
    assign layer3_out[8] = layer2_out[76];
    assign layer3_out[9] = ~(layer2_out[685] | layer2_out[686]);
    assign layer3_out[10] = layer2_out[564] & layer2_out[565];
    assign layer3_out[11] = ~layer2_out[663];
    assign layer3_out[12] = layer2_out[169];
    assign layer3_out[13] = ~layer2_out[75] | layer2_out[76];
    assign layer3_out[14] = ~layer2_out[533];
    assign layer3_out[15] = layer2_out[21] & layer2_out[22];
    assign layer3_out[16] = ~layer2_out[126];
    assign layer3_out[17] = layer2_out[395];
    assign layer3_out[18] = layer2_out[276] & ~layer2_out[277];
    assign layer3_out[19] = ~layer2_out[283];
    assign layer3_out[20] = layer2_out[117];
    assign layer3_out[21] = layer2_out[777] | layer2_out[778];
    assign layer3_out[22] = ~layer2_out[252];
    assign layer3_out[23] = layer2_out[250];
    assign layer3_out[24] = layer2_out[597];
    assign layer3_out[25] = layer2_out[515];
    assign layer3_out[26] = layer2_out[70];
    assign layer3_out[27] = layer2_out[584];
    assign layer3_out[28] = layer2_out[320];
    assign layer3_out[29] = layer2_out[739];
    assign layer3_out[30] = layer2_out[655];
    assign layer3_out[31] = ~(layer2_out[728] | layer2_out[729]);
    assign layer3_out[32] = ~layer2_out[81];
    assign layer3_out[33] = ~layer2_out[503] | layer2_out[504];
    assign layer3_out[34] = layer2_out[159];
    assign layer3_out[35] = ~(layer2_out[549] | layer2_out[550]);
    assign layer3_out[36] = layer2_out[303];
    assign layer3_out[37] = ~layer2_out[466];
    assign layer3_out[38] = ~layer2_out[661];
    assign layer3_out[39] = ~layer2_out[304];
    assign layer3_out[40] = layer2_out[742];
    assign layer3_out[41] = ~layer2_out[51];
    assign layer3_out[42] = layer2_out[585];
    assign layer3_out[43] = ~layer2_out[351];
    assign layer3_out[44] = ~layer2_out[359];
    assign layer3_out[45] = ~layer2_out[109] | layer2_out[110];
    assign layer3_out[46] = layer2_out[192];
    assign layer3_out[47] = ~layer2_out[294];
    assign layer3_out[48] = layer2_out[601];
    assign layer3_out[49] = layer2_out[615];
    assign layer3_out[50] = ~layer2_out[599] | layer2_out[600];
    assign layer3_out[51] = ~(layer2_out[507] ^ layer2_out[508]);
    assign layer3_out[52] = layer2_out[62];
    assign layer3_out[53] = ~layer2_out[524];
    assign layer3_out[54] = layer2_out[779];
    assign layer3_out[55] = layer2_out[148];
    assign layer3_out[56] = layer2_out[780];
    assign layer3_out[57] = ~(layer2_out[415] | layer2_out[416]);
    assign layer3_out[58] = ~layer2_out[656];
    assign layer3_out[59] = ~layer2_out[176];
    assign layer3_out[60] = ~(layer2_out[524] | layer2_out[525]);
    assign layer3_out[61] = layer2_out[792];
    assign layer3_out[62] = ~layer2_out[799];
    assign layer3_out[63] = layer2_out[315];
    assign layer3_out[64] = layer2_out[726] & ~layer2_out[725];
    assign layer3_out[65] = layer2_out[411];
    assign layer3_out[66] = layer2_out[190];
    assign layer3_out[67] = ~layer2_out[653];
    assign layer3_out[68] = ~layer2_out[480];
    assign layer3_out[69] = layer2_out[547] ^ layer2_out[548];
    assign layer3_out[70] = ~layer2_out[142];
    assign layer3_out[71] = layer2_out[293] & ~layer2_out[292];
    assign layer3_out[72] = ~layer2_out[356];
    assign layer3_out[73] = ~(layer2_out[436] | layer2_out[437]);
    assign layer3_out[74] = layer2_out[3];
    assign layer3_out[75] = layer2_out[346];
    assign layer3_out[76] = ~layer2_out[580];
    assign layer3_out[77] = layer2_out[212];
    assign layer3_out[78] = ~layer2_out[490];
    assign layer3_out[79] = ~layer2_out[653];
    assign layer3_out[80] = layer2_out[174];
    assign layer3_out[81] = layer2_out[408] & ~layer2_out[407];
    assign layer3_out[82] = layer2_out[553] & ~layer2_out[554];
    assign layer3_out[83] = layer2_out[186] & layer2_out[187];
    assign layer3_out[84] = layer2_out[215] & layer2_out[216];
    assign layer3_out[85] = layer2_out[100] & ~layer2_out[101];
    assign layer3_out[86] = layer2_out[171];
    assign layer3_out[87] = layer2_out[86] & layer2_out[87];
    assign layer3_out[88] = layer2_out[67] & ~layer2_out[66];
    assign layer3_out[89] = layer2_out[98] ^ layer2_out[99];
    assign layer3_out[90] = layer2_out[753] & ~layer2_out[754];
    assign layer3_out[91] = layer2_out[12] & ~layer2_out[11];
    assign layer3_out[92] = ~(layer2_out[84] | layer2_out[85]);
    assign layer3_out[93] = layer2_out[641] & ~layer2_out[640];
    assign layer3_out[94] = ~layer2_out[509];
    assign layer3_out[95] = layer2_out[343];
    assign layer3_out[96] = layer2_out[13] & layer2_out[14];
    assign layer3_out[97] = ~(layer2_out[768] | layer2_out[769]);
    assign layer3_out[98] = layer2_out[495];
    assign layer3_out[99] = layer2_out[185] & layer2_out[186];
    assign layer3_out[100] = layer2_out[119] & ~layer2_out[118];
    assign layer3_out[101] = ~layer2_out[21];
    assign layer3_out[102] = layer2_out[121] & layer2_out[122];
    assign layer3_out[103] = ~layer2_out[95];
    assign layer3_out[104] = ~layer2_out[299];
    assign layer3_out[105] = ~layer2_out[787];
    assign layer3_out[106] = layer2_out[533] & ~layer2_out[532];
    assign layer3_out[107] = ~layer2_out[58];
    assign layer3_out[108] = layer2_out[100] & ~layer2_out[99];
    assign layer3_out[109] = layer2_out[696];
    assign layer3_out[110] = ~(layer2_out[200] & layer2_out[201]);
    assign layer3_out[111] = layer2_out[635];
    assign layer3_out[112] = ~(layer2_out[527] | layer2_out[528]);
    assign layer3_out[113] = layer2_out[360] & ~layer2_out[361];
    assign layer3_out[114] = layer2_out[651] & layer2_out[652];
    assign layer3_out[115] = ~(layer2_out[379] | layer2_out[380]);
    assign layer3_out[116] = layer2_out[428] & layer2_out[429];
    assign layer3_out[117] = layer2_out[410] & ~layer2_out[411];
    assign layer3_out[118] = ~layer2_out[354];
    assign layer3_out[119] = ~(layer2_out[441] | layer2_out[442]);
    assign layer3_out[120] = layer2_out[642];
    assign layer3_out[121] = layer2_out[163] ^ layer2_out[164];
    assign layer3_out[122] = ~layer2_out[489];
    assign layer3_out[123] = layer2_out[759] & layer2_out[760];
    assign layer3_out[124] = ~(layer2_out[237] | layer2_out[238]);
    assign layer3_out[125] = layer2_out[248] & ~layer2_out[247];
    assign layer3_out[126] = layer2_out[385] & layer2_out[386];
    assign layer3_out[127] = layer2_out[417] & layer2_out[418];
    assign layer3_out[128] = layer2_out[151];
    assign layer3_out[129] = ~layer2_out[48];
    assign layer3_out[130] = layer2_out[679];
    assign layer3_out[131] = layer2_out[621];
    assign layer3_out[132] = layer2_out[428];
    assign layer3_out[133] = ~(layer2_out[270] | layer2_out[271]);
    assign layer3_out[134] = ~layer2_out[371];
    assign layer3_out[135] = ~(layer2_out[518] ^ layer2_out[519]);
    assign layer3_out[136] = layer2_out[91] & ~layer2_out[92];
    assign layer3_out[137] = layer2_out[112] & layer2_out[113];
    assign layer3_out[138] = layer2_out[284] ^ layer2_out[285];
    assign layer3_out[139] = ~layer2_out[48];
    assign layer3_out[140] = ~layer2_out[613];
    assign layer3_out[141] = layer2_out[25] & layer2_out[26];
    assign layer3_out[142] = layer2_out[513] & ~layer2_out[512];
    assign layer3_out[143] = layer2_out[531];
    assign layer3_out[144] = layer2_out[292];
    assign layer3_out[145] = layer2_out[517] & ~layer2_out[518];
    assign layer3_out[146] = layer2_out[663] & ~layer2_out[662];
    assign layer3_out[147] = layer2_out[484];
    assign layer3_out[148] = layer2_out[112];
    assign layer3_out[149] = layer2_out[151] & ~layer2_out[150];
    assign layer3_out[150] = ~layer2_out[613];
    assign layer3_out[151] = ~layer2_out[396];
    assign layer3_out[152] = layer2_out[752];
    assign layer3_out[153] = ~layer2_out[675];
    assign layer3_out[154] = layer2_out[607] & layer2_out[608];
    assign layer3_out[155] = ~(layer2_out[746] | layer2_out[747]);
    assign layer3_out[156] = ~layer2_out[38];
    assign layer3_out[157] = ~(layer2_out[226] | layer2_out[227]);
    assign layer3_out[158] = layer2_out[393] & ~layer2_out[394];
    assign layer3_out[159] = ~layer2_out[603] | layer2_out[604];
    assign layer3_out[160] = layer2_out[267];
    assign layer3_out[161] = ~layer2_out[370];
    assign layer3_out[162] = layer2_out[609] ^ layer2_out[610];
    assign layer3_out[163] = ~(layer2_out[425] & layer2_out[426]);
    assign layer3_out[164] = layer2_out[206] & ~layer2_out[207];
    assign layer3_out[165] = ~layer2_out[65];
    assign layer3_out[166] = ~layer2_out[94];
    assign layer3_out[167] = ~layer2_out[94];
    assign layer3_out[168] = ~layer2_out[535];
    assign layer3_out[169] = ~layer2_out[467] | layer2_out[468];
    assign layer3_out[170] = ~layer2_out[260];
    assign layer3_out[171] = ~layer2_out[498];
    assign layer3_out[172] = layer2_out[521];
    assign layer3_out[173] = layer2_out[366];
    assign layer3_out[174] = layer2_out[706];
    assign layer3_out[175] = ~layer2_out[785];
    assign layer3_out[176] = ~layer2_out[392];
    assign layer3_out[177] = ~layer2_out[794];
    assign layer3_out[178] = layer2_out[671];
    assign layer3_out[179] = ~layer2_out[272];
    assign layer3_out[180] = layer2_out[447];
    assign layer3_out[181] = layer2_out[145] & ~layer2_out[144];
    assign layer3_out[182] = layer2_out[288];
    assign layer3_out[183] = layer2_out[471];
    assign layer3_out[184] = layer2_out[505];
    assign layer3_out[185] = ~(layer2_out[604] | layer2_out[605]);
    assign layer3_out[186] = ~(layer2_out[123] & layer2_out[124]);
    assign layer3_out[187] = ~(layer2_out[89] | layer2_out[90]);
    assign layer3_out[188] = ~layer2_out[210];
    assign layer3_out[189] = layer2_out[233];
    assign layer3_out[190] = layer2_out[543];
    assign layer3_out[191] = ~layer2_out[294];
    assign layer3_out[192] = ~layer2_out[65];
    assign layer3_out[193] = layer2_out[0];
    assign layer3_out[194] = layer2_out[59];
    assign layer3_out[195] = ~layer2_out[245];
    assign layer3_out[196] = ~(layer2_out[697] ^ layer2_out[698]);
    assign layer3_out[197] = layer2_out[708];
    assign layer3_out[198] = layer2_out[669];
    assign layer3_out[199] = layer2_out[456] ^ layer2_out[457];
    assign layer3_out[200] = ~layer2_out[383];
    assign layer3_out[201] = ~layer2_out[26] | layer2_out[27];
    assign layer3_out[202] = layer2_out[687];
    assign layer3_out[203] = ~layer2_out[128];
    assign layer3_out[204] = ~layer2_out[664];
    assign layer3_out[205] = ~layer2_out[735];
    assign layer3_out[206] = layer2_out[659];
    assign layer3_out[207] = layer2_out[745] & ~layer2_out[746];
    assign layer3_out[208] = ~layer2_out[735];
    assign layer3_out[209] = layer2_out[708];
    assign layer3_out[210] = layer2_out[270];
    assign layer3_out[211] = layer2_out[387] ^ layer2_out[388];
    assign layer3_out[212] = layer2_out[194];
    assign layer3_out[213] = layer2_out[55];
    assign layer3_out[214] = layer2_out[85];
    assign layer3_out[215] = layer2_out[212];
    assign layer3_out[216] = layer2_out[399];
    assign layer3_out[217] = layer2_out[80] & layer2_out[81];
    assign layer3_out[218] = ~layer2_out[216];
    assign layer3_out[219] = layer2_out[403];
    assign layer3_out[220] = layer2_out[481] | layer2_out[482];
    assign layer3_out[221] = ~layer2_out[722];
    assign layer3_out[222] = ~layer2_out[166];
    assign layer3_out[223] = layer2_out[560];
    assign layer3_out[224] = layer2_out[8];
    assign layer3_out[225] = layer2_out[557];
    assign layer3_out[226] = layer2_out[127] ^ layer2_out[128];
    assign layer3_out[227] = ~layer2_out[236];
    assign layer3_out[228] = layer2_out[669] & layer2_out[670];
    assign layer3_out[229] = layer2_out[334];
    assign layer3_out[230] = ~layer2_out[470];
    assign layer3_out[231] = ~layer2_out[5] | layer2_out[4];
    assign layer3_out[232] = ~layer2_out[39];
    assign layer3_out[233] = layer2_out[329];
    assign layer3_out[234] = ~(layer2_out[674] | layer2_out[675]);
    assign layer3_out[235] = ~(layer2_out[693] & layer2_out[694]);
    assign layer3_out[236] = ~layer2_out[230];
    assign layer3_out[237] = ~layer2_out[690];
    assign layer3_out[238] = layer2_out[443];
    assign layer3_out[239] = layer2_out[743] ^ layer2_out[744];
    assign layer3_out[240] = ~layer2_out[475];
    assign layer3_out[241] = ~layer2_out[166];
    assign layer3_out[242] = ~(layer2_out[183] | layer2_out[184]);
    assign layer3_out[243] = ~layer2_out[35] | layer2_out[36];
    assign layer3_out[244] = ~(layer2_out[702] & layer2_out[703]);
    assign layer3_out[245] = ~(layer2_out[315] | layer2_out[316]);
    assign layer3_out[246] = layer2_out[641];
    assign layer3_out[247] = layer2_out[378];
    assign layer3_out[248] = layer2_out[146];
    assign layer3_out[249] = ~layer2_out[243];
    assign layer3_out[250] = layer2_out[424];
    assign layer3_out[251] = layer2_out[72] & ~layer2_out[73];
    assign layer3_out[252] = ~(layer2_out[628] | layer2_out[629]);
    assign layer3_out[253] = layer2_out[496] & ~layer2_out[497];
    assign layer3_out[254] = ~layer2_out[723];
    assign layer3_out[255] = layer2_out[398];
    assign layer3_out[256] = ~layer2_out[181];
    assign layer3_out[257] = layer2_out[589];
    assign layer3_out[258] = ~layer2_out[323];
    assign layer3_out[259] = ~(layer2_out[308] ^ layer2_out[309]);
    assign layer3_out[260] = ~layer2_out[348];
    assign layer3_out[261] = layer2_out[136] & ~layer2_out[137];
    assign layer3_out[262] = layer2_out[619];
    assign layer3_out[263] = layer2_out[444];
    assign layer3_out[264] = layer2_out[71] & ~layer2_out[70];
    assign layer3_out[265] = ~layer2_out[73];
    assign layer3_out[266] = ~(layer2_out[228] & layer2_out[229]);
    assign layer3_out[267] = layer2_out[454];
    assign layer3_out[268] = ~layer2_out[385];
    assign layer3_out[269] = layer2_out[464] ^ layer2_out[465];
    assign layer3_out[270] = ~layer2_out[29];
    assign layer3_out[271] = ~layer2_out[364];
    assign layer3_out[272] = ~layer2_out[769];
    assign layer3_out[273] = ~layer2_out[558];
    assign layer3_out[274] = ~(layer2_out[56] ^ layer2_out[57]);
    assign layer3_out[275] = ~layer2_out[332];
    assign layer3_out[276] = ~layer2_out[774];
    assign layer3_out[277] = layer2_out[583];
    assign layer3_out[278] = ~(layer2_out[258] | layer2_out[259]);
    assign layer3_out[279] = layer2_out[431] & ~layer2_out[432];
    assign layer3_out[280] = layer2_out[520];
    assign layer3_out[281] = ~(layer2_out[750] ^ layer2_out[751]);
    assign layer3_out[282] = layer2_out[325] & ~layer2_out[324];
    assign layer3_out[283] = layer2_out[330] & layer2_out[331];
    assign layer3_out[284] = layer2_out[274];
    assign layer3_out[285] = ~(layer2_out[139] | layer2_out[140]);
    assign layer3_out[286] = ~layer2_out[773];
    assign layer3_out[287] = layer2_out[434];
    assign layer3_out[288] = layer2_out[574];
    assign layer3_out[289] = ~layer2_out[633];
    assign layer3_out[290] = layer2_out[793];
    assign layer3_out[291] = layer2_out[545] & ~layer2_out[546];
    assign layer3_out[292] = layer2_out[770] | layer2_out[771];
    assign layer3_out[293] = layer2_out[422];
    assign layer3_out[294] = ~(layer2_out[698] | layer2_out[699]);
    assign layer3_out[295] = ~(layer2_out[676] | layer2_out[677]);
    assign layer3_out[296] = layer2_out[787];
    assign layer3_out[297] = ~(layer2_out[52] | layer2_out[53]);
    assign layer3_out[298] = layer2_out[31];
    assign layer3_out[299] = ~layer2_out[231];
    assign layer3_out[300] = layer2_out[103] ^ layer2_out[104];
    assign layer3_out[301] = ~layer2_out[445];
    assign layer3_out[302] = ~layer2_out[486];
    assign layer3_out[303] = layer2_out[640] & ~layer2_out[639];
    assign layer3_out[304] = layer2_out[398];
    assign layer3_out[305] = layer2_out[146];
    assign layer3_out[306] = ~layer2_out[572];
    assign layer3_out[307] = ~layer2_out[299];
    assign layer3_out[308] = layer2_out[372] & ~layer2_out[371];
    assign layer3_out[309] = ~layer2_out[169];
    assign layer3_out[310] = ~layer2_out[597];
    assign layer3_out[311] = ~(layer2_out[285] | layer2_out[286]);
    assign layer3_out[312] = ~layer2_out[387];
    assign layer3_out[313] = layer2_out[251] & ~layer2_out[250];
    assign layer3_out[314] = layer2_out[31] | layer2_out[32];
    assign layer3_out[315] = layer2_out[645];
    assign layer3_out[316] = ~layer2_out[717];
    assign layer3_out[317] = ~layer2_out[317];
    assign layer3_out[318] = ~layer2_out[542];
    assign layer3_out[319] = layer2_out[199];
    assign layer3_out[320] = layer2_out[172];
    assign layer3_out[321] = ~(layer2_out[378] | layer2_out[379]);
    assign layer3_out[322] = layer2_out[357];
    assign layer3_out[323] = layer2_out[605];
    assign layer3_out[324] = layer2_out[138];
    assign layer3_out[325] = layer2_out[730] & layer2_out[731];
    assign layer3_out[326] = ~layer2_out[235];
    assign layer3_out[327] = ~(layer2_out[262] & layer2_out[263]);
    assign layer3_out[328] = ~layer2_out[71];
    assign layer3_out[329] = ~(layer2_out[246] | layer2_out[247]);
    assign layer3_out[330] = layer2_out[594] & ~layer2_out[593];
    assign layer3_out[331] = layer2_out[643];
    assign layer3_out[332] = layer2_out[153];
    assign layer3_out[333] = layer2_out[109] & ~layer2_out[108];
    assign layer3_out[334] = layer2_out[49];
    assign layer3_out[335] = ~layer2_out[700];
    assign layer3_out[336] = ~layer2_out[621];
    assign layer3_out[337] = layer2_out[63];
    assign layer3_out[338] = ~layer2_out[741];
    assign layer3_out[339] = ~layer2_out[463];
    assign layer3_out[340] = ~layer2_out[440];
    assign layer3_out[341] = ~layer2_out[696];
    assign layer3_out[342] = layer2_out[590] | layer2_out[591];
    assign layer3_out[343] = layer2_out[221];
    assign layer3_out[344] = layer2_out[690];
    assign layer3_out[345] = layer2_out[53];
    assign layer3_out[346] = layer2_out[408] & layer2_out[409];
    assign layer3_out[347] = layer2_out[298];
    assign layer3_out[348] = layer2_out[338];
    assign layer3_out[349] = layer2_out[694] & ~layer2_out[695];
    assign layer3_out[350] = ~layer2_out[308];
    assign layer3_out[351] = layer2_out[656];
    assign layer3_out[352] = ~layer2_out[514];
    assign layer3_out[353] = layer2_out[121];
    assign layer3_out[354] = layer2_out[45];
    assign layer3_out[355] = layer2_out[133] & ~layer2_out[134];
    assign layer3_out[356] = layer2_out[773];
    assign layer3_out[357] = ~layer2_out[321];
    assign layer3_out[358] = ~(layer2_out[763] & layer2_out[764]);
    assign layer3_out[359] = layer2_out[126];
    assign layer3_out[360] = layer2_out[469];
    assign layer3_out[361] = layer2_out[142];
    assign layer3_out[362] = ~layer2_out[756];
    assign layer3_out[363] = ~(layer2_out[264] ^ layer2_out[265]);
    assign layer3_out[364] = layer2_out[414];
    assign layer3_out[365] = ~layer2_out[418];
    assign layer3_out[366] = ~layer2_out[446];
    assign layer3_out[367] = layer2_out[788];
    assign layer3_out[368] = layer2_out[2] & ~layer2_out[0];
    assign layer3_out[369] = ~layer2_out[325];
    assign layer3_out[370] = layer2_out[340];
    assign layer3_out[371] = ~layer2_out[488];
    assign layer3_out[372] = ~layer2_out[413];
    assign layer3_out[373] = layer2_out[506];
    assign layer3_out[374] = layer2_out[289];
    assign layer3_out[375] = ~layer2_out[700];
    assign layer3_out[376] = layer2_out[280] | layer2_out[281];
    assign layer3_out[377] = ~layer2_out[23];
    assign layer3_out[378] = layer2_out[40] | layer2_out[41];
    assign layer3_out[379] = ~layer2_out[181];
    assign layer3_out[380] = layer2_out[155];
    assign layer3_out[381] = ~layer2_out[668];
    assign layer3_out[382] = layer2_out[367] ^ layer2_out[368];
    assign layer3_out[383] = layer2_out[766] & ~layer2_out[765];
    assign layer3_out[384] = layer2_out[762];
    assign layer3_out[385] = layer2_out[209];
    assign layer3_out[386] = layer2_out[224] & ~layer2_out[223];
    assign layer3_out[387] = layer2_out[666];
    assign layer3_out[388] = ~layer2_out[279];
    assign layer3_out[389] = layer2_out[415];
    assign layer3_out[390] = ~layer2_out[313];
    assign layer3_out[391] = layer2_out[730];
    assign layer3_out[392] = layer2_out[241];
    assign layer3_out[393] = ~(layer2_out[629] | layer2_out[630]);
    assign layer3_out[394] = ~layer2_out[344];
    assign layer3_out[395] = ~layer2_out[713];
    assign layer3_out[396] = ~layer2_out[97];
    assign layer3_out[397] = layer2_out[472] & ~layer2_out[473];
    assign layer3_out[398] = ~layer2_out[581];
    assign layer3_out[399] = layer2_out[452];
    assign layer3_out[400] = ~(layer2_out[257] ^ layer2_out[258]);
    assign layer3_out[401] = ~layer2_out[781];
    assign layer3_out[402] = ~layer2_out[528];
    assign layer3_out[403] = layer2_out[309];
    assign layer3_out[404] = layer2_out[235];
    assign layer3_out[405] = ~layer2_out[499];
    assign layer3_out[406] = layer2_out[254] ^ layer2_out[255];
    assign layer3_out[407] = layer2_out[156];
    assign layer3_out[408] = ~layer2_out[449];
    assign layer3_out[409] = ~layer2_out[359];
    assign layer3_out[410] = ~(layer2_out[691] | layer2_out[692]);
    assign layer3_out[411] = ~layer2_out[474];
    assign layer3_out[412] = layer2_out[42] ^ layer2_out[43];
    assign layer3_out[413] = layer2_out[711] & ~layer2_out[710];
    assign layer3_out[414] = layer2_out[318] & ~layer2_out[319];
    assign layer3_out[415] = layer2_out[375];
    assign layer3_out[416] = ~layer2_out[409];
    assign layer3_out[417] = ~layer2_out[301];
    assign layer3_out[418] = ~(layer2_out[736] ^ layer2_out[737]);
    assign layer3_out[419] = layer2_out[544];
    assign layer3_out[420] = layer2_out[133];
    assign layer3_out[421] = layer2_out[574];
    assign layer3_out[422] = layer2_out[502] & layer2_out[503];
    assign layer3_out[423] = layer2_out[584] ^ layer2_out[585];
    assign layer3_out[424] = layer2_out[590] & ~layer2_out[589];
    assign layer3_out[425] = ~layer2_out[796];
    assign layer3_out[426] = layer2_out[93];
    assign layer3_out[427] = layer2_out[204] ^ layer2_out[205];
    assign layer3_out[428] = ~(layer2_out[727] | layer2_out[728]);
    assign layer3_out[429] = layer2_out[568];
    assign layer3_out[430] = ~layer2_out[791];
    assign layer3_out[431] = ~(layer2_out[448] | layer2_out[449]);
    assign layer3_out[432] = layer2_out[789] & layer2_out[790];
    assign layer3_out[433] = ~(layer2_out[537] | layer2_out[538]);
    assign layer3_out[434] = layer2_out[538] ^ layer2_out[539];
    assign layer3_out[435] = ~layer2_out[798];
    assign layer3_out[436] = layer2_out[357];
    assign layer3_out[437] = layer2_out[601] | layer2_out[602];
    assign layer3_out[438] = ~layer2_out[555];
    assign layer3_out[439] = layer2_out[19] & ~layer2_out[18];
    assign layer3_out[440] = layer2_out[432];
    assign layer3_out[441] = layer2_out[715];
    assign layer3_out[442] = ~layer2_out[283];
    assign layer3_out[443] = ~(layer2_out[749] | layer2_out[750]);
    assign layer3_out[444] = layer2_out[712];
    assign layer3_out[445] = ~layer2_out[185] | layer2_out[184];
    assign layer3_out[446] = layer2_out[731];
    assign layer3_out[447] = ~layer2_out[571];
    assign layer3_out[448] = layer2_out[219];
    assign layer3_out[449] = ~layer2_out[783];
    assign layer3_out[450] = ~layer2_out[296];
    assign layer3_out[451] = ~layer2_out[576];
    assign layer3_out[452] = ~layer2_out[102];
    assign layer3_out[453] = layer2_out[110];
    assign layer3_out[454] = layer2_out[493] ^ layer2_out[494];
    assign layer3_out[455] = layer2_out[646];
    assign layer3_out[456] = layer2_out[248] & layer2_out[249];
    assign layer3_out[457] = ~(layer2_out[275] ^ layer2_out[276]);
    assign layer3_out[458] = ~layer2_out[417];
    assign layer3_out[459] = layer2_out[502];
    assign layer3_out[460] = ~layer2_out[659];
    assign layer3_out[461] = layer2_out[587] ^ layer2_out[588];
    assign layer3_out[462] = ~layer2_out[202];
    assign layer3_out[463] = layer2_out[122] & layer2_out[123];
    assign layer3_out[464] = layer2_out[614] | layer2_out[615];
    assign layer3_out[465] = layer2_out[761];
    assign layer3_out[466] = layer2_out[332];
    assign layer3_out[467] = ~layer2_out[288] | layer2_out[287];
    assign layer3_out[468] = layer2_out[311] & ~layer2_out[312];
    assign layer3_out[469] = ~layer2_out[487];
    assign layer3_out[470] = layer2_out[310];
    assign layer3_out[471] = layer2_out[452];
    assign layer3_out[472] = ~layer2_out[608];
    assign layer3_out[473] = ~layer2_out[34] | layer2_out[33];
    assign layer3_out[474] = ~(layer2_out[648] ^ layer2_out[649]);
    assign layer3_out[475] = layer2_out[479] & layer2_out[480];
    assign layer3_out[476] = layer2_out[51];
    assign layer3_out[477] = layer2_out[375];
    assign layer3_out[478] = layer2_out[785] & layer2_out[786];
    assign layer3_out[479] = layer2_out[116] | layer2_out[117];
    assign layer3_out[480] = layer2_out[420] & layer2_out[421];
    assign layer3_out[481] = ~layer2_out[474];
    assign layer3_out[482] = layer2_out[555];
    assign layer3_out[483] = layer2_out[200] & ~layer2_out[199];
    assign layer3_out[484] = layer2_out[115];
    assign layer3_out[485] = layer2_out[647];
    assign layer3_out[486] = layer2_out[364];
    assign layer3_out[487] = layer2_out[717] & ~layer2_out[718];
    assign layer3_out[488] = ~layer2_out[313];
    assign layer3_out[489] = ~layer2_out[17];
    assign layer3_out[490] = layer2_out[381] & ~layer2_out[380];
    assign layer3_out[491] = layer2_out[388] & ~layer2_out[389];
    assign layer3_out[492] = ~layer2_out[627];
    assign layer3_out[493] = layer2_out[516];
    assign layer3_out[494] = ~layer2_out[251];
    assign layer3_out[495] = ~(layer2_out[350] | layer2_out[351]);
    assign layer3_out[496] = layer2_out[238] | layer2_out[239];
    assign layer3_out[497] = ~layer2_out[532];
    assign layer3_out[498] = ~layer2_out[603] | layer2_out[602];
    assign layer3_out[499] = layer2_out[373];
    assign layer3_out[500] = ~layer2_out[178];
    assign layer3_out[501] = layer2_out[548] | layer2_out[549];
    assign layer3_out[502] = ~layer2_out[767];
    assign layer3_out[503] = ~layer2_out[612];
    assign layer3_out[504] = layer2_out[405];
    assign layer3_out[505] = layer2_out[1];
    assign layer3_out[506] = ~layer2_out[267];
    assign layer3_out[507] = ~layer2_out[389];
    assign layer3_out[508] = layer2_out[560] & ~layer2_out[561];
    assign layer3_out[509] = layer2_out[232] & ~layer2_out[233];
    assign layer3_out[510] = ~layer2_out[459];
    assign layer3_out[511] = layer2_out[512];
    assign layer3_out[512] = layer2_out[458] & ~layer2_out[459];
    assign layer3_out[513] = layer2_out[290];
    assign layer3_out[514] = ~layer2_out[279];
    assign layer3_out[515] = layer2_out[421];
    assign layer3_out[516] = layer2_out[400] & ~layer2_out[401];
    assign layer3_out[517] = layer2_out[579];
    assign layer3_out[518] = ~layer2_out[567];
    assign layer3_out[519] = ~(layer2_out[711] ^ layer2_out[712]);
    assign layer3_out[520] = layer2_out[43];
    assign layer3_out[521] = layer2_out[104] ^ layer2_out[105];
    assign layer3_out[522] = ~layer2_out[637];
    assign layer3_out[523] = ~layer2_out[79];
    assign layer3_out[524] = ~layer2_out[506];
    assign layer3_out[525] = ~layer2_out[576];
    assign layer3_out[526] = ~layer2_out[446];
    assign layer3_out[527] = layer2_out[437] & layer2_out[438];
    assign layer3_out[528] = layer2_out[721] & ~layer2_out[720];
    assign layer3_out[529] = ~layer2_out[155];
    assign layer3_out[530] = layer2_out[461] & layer2_out[462];
    assign layer3_out[531] = ~layer2_out[282];
    assign layer3_out[532] = ~(layer2_out[46] ^ layer2_out[47]);
    assign layer3_out[533] = layer2_out[273] & ~layer2_out[272];
    assign layer3_out[534] = layer2_out[542];
    assign layer3_out[535] = ~layer2_out[336];
    assign layer3_out[536] = layer2_out[96] ^ layer2_out[97];
    assign layer3_out[537] = layer2_out[797];
    assign layer3_out[538] = ~layer2_out[680];
    assign layer3_out[539] = layer2_out[106];
    assign layer3_out[540] = ~layer2_out[727];
    assign layer3_out[541] = ~layer2_out[69];
    assign layer3_out[542] = ~layer2_out[245];
    assign layer3_out[543] = ~layer2_out[401];
    assign layer3_out[544] = layer2_out[606];
    assign layer3_out[545] = ~layer2_out[738];
    assign layer3_out[546] = layer2_out[568];
    assign layer3_out[547] = ~(layer2_out[526] | layer2_out[527]);
    assign layer3_out[548] = layer2_out[569];
    assign layer3_out[549] = ~layer2_out[783];
    assign layer3_out[550] = ~layer2_out[704];
    assign layer3_out[551] = ~layer2_out[639];
    assign layer3_out[552] = layer2_out[457] & layer2_out[458];
    assign layer3_out[553] = ~layer2_out[348];
    assign layer3_out[554] = layer2_out[161];
    assign layer3_out[555] = ~layer2_out[581];
    assign layer3_out[556] = layer2_out[499] ^ layer2_out[500];
    assign layer3_out[557] = ~layer2_out[172];
    assign layer3_out[558] = ~layer2_out[24];
    assign layer3_out[559] = ~layer2_out[149];
    assign layer3_out[560] = layer2_out[637] & ~layer2_out[638];
    assign layer3_out[561] = ~layer2_out[792];
    assign layer3_out[562] = layer2_out[350] & ~layer2_out[349];
    assign layer3_out[563] = layer2_out[563];
    assign layer3_out[564] = ~layer2_out[102];
    assign layer3_out[565] = layer2_out[189] & ~layer2_out[190];
    assign layer3_out[566] = layer2_out[334];
    assign layer3_out[567] = layer2_out[453];
    assign layer3_out[568] = layer2_out[565] & layer2_out[566];
    assign layer3_out[569] = layer2_out[491];
    assign layer3_out[570] = ~layer2_out[709] | layer2_out[710];
    assign layer3_out[571] = layer2_out[153] & ~layer2_out[152];
    assign layer3_out[572] = ~(layer2_out[78] ^ layer2_out[79]);
    assign layer3_out[573] = ~layer2_out[75];
    assign layer3_out[574] = layer2_out[205] & layer2_out[206];
    assign layer3_out[575] = ~layer2_out[553];
    assign layer3_out[576] = ~(layer2_out[263] ^ layer2_out[264]);
    assign layer3_out[577] = layer2_out[327];
    assign layer3_out[578] = layer2_out[556];
    assign layer3_out[579] = layer2_out[723] & ~layer2_out[722];
    assign layer3_out[580] = layer2_out[301];
    assign layer3_out[581] = layer2_out[767];
    assign layer3_out[582] = ~layer2_out[631];
    assign layer3_out[583] = layer2_out[6];
    assign layer3_out[584] = layer2_out[440];
    assign layer3_out[585] = ~layer2_out[384];
    assign layer3_out[586] = layer2_out[165] & ~layer2_out[164];
    assign layer3_out[587] = ~layer2_out[161];
    assign layer3_out[588] = layer2_out[130];
    assign layer3_out[589] = layer2_out[541] & ~layer2_out[540];
    assign layer3_out[590] = layer2_out[136] & ~layer2_out[135];
    assign layer3_out[591] = ~layer2_out[535] | layer2_out[536];
    assign layer3_out[592] = layer2_out[678];
    assign layer3_out[593] = ~layer2_out[137];
    assign layer3_out[594] = layer2_out[619] & ~layer2_out[620];
    assign layer3_out[595] = ~layer2_out[244];
    assign layer3_out[596] = ~layer2_out[10];
    assign layer3_out[597] = layer2_out[704];
    assign layer3_out[598] = layer2_out[571] & layer2_out[572];
    assign layer3_out[599] = layer2_out[134];
    assign layer3_out[600] = ~layer2_out[329] | layer2_out[328];
    assign layer3_out[601] = ~layer2_out[390] | layer2_out[391];
    assign layer3_out[602] = ~layer2_out[771];
    assign layer3_out[603] = layer2_out[764] & ~layer2_out[765];
    assign layer3_out[604] = layer2_out[404];
    assign layer3_out[605] = ~(layer2_out[419] ^ layer2_out[420]);
    assign layer3_out[606] = ~layer2_out[382];
    assign layer3_out[607] = ~layer2_out[82] | layer2_out[83];
    assign layer3_out[608] = ~layer2_out[776];
    assign layer3_out[609] = ~layer2_out[693];
    assign layer3_out[610] = ~layer2_out[55];
    assign layer3_out[611] = ~layer2_out[777];
    assign layer3_out[612] = layer2_out[317];
    assign layer3_out[613] = ~layer2_out[392];
    assign layer3_out[614] = layer2_out[256] ^ layer2_out[257];
    assign layer3_out[615] = ~layer2_out[23];
    assign layer3_out[616] = layer2_out[19];
    assign layer3_out[617] = layer2_out[435];
    assign layer3_out[618] = ~layer2_out[196];
    assign layer3_out[619] = ~layer2_out[12];
    assign layer3_out[620] = layer2_out[623];
    assign layer3_out[621] = ~layer2_out[645];
    assign layer3_out[622] = layer2_out[167];
    assign layer3_out[623] = ~(layer2_out[36] | layer2_out[37]);
    assign layer3_out[624] = layer2_out[14] & ~layer2_out[15];
    assign layer3_out[625] = layer2_out[666] & ~layer2_out[665];
    assign layer3_out[626] = layer2_out[551] & ~layer2_out[552];
    assign layer3_out[627] = layer2_out[672] & ~layer2_out[673];
    assign layer3_out[628] = ~layer2_out[273];
    assign layer3_out[629] = ~layer2_out[754];
    assign layer3_out[630] = layer2_out[689];
    assign layer3_out[631] = ~layer2_out[159];
    assign layer3_out[632] = ~layer2_out[684] | layer2_out[683];
    assign layer3_out[633] = layer2_out[227];
    assign layer3_out[634] = layer2_out[230] & layer2_out[231];
    assign layer3_out[635] = layer2_out[426] & layer2_out[427];
    assign layer3_out[636] = layer2_out[352];
    assign layer3_out[637] = layer2_out[60] & layer2_out[61];
    assign layer3_out[638] = ~layer2_out[84];
    assign layer3_out[639] = ~layer2_out[59];
    assign layer3_out[640] = layer2_out[685];
    assign layer3_out[641] = ~layer2_out[324];
    assign layer3_out[642] = layer2_out[369];
    assign layer3_out[643] = layer2_out[488];
    assign layer3_out[644] = layer2_out[758] & ~layer2_out[757];
    assign layer3_out[645] = layer2_out[219];
    assign layer3_out[646] = layer2_out[224] ^ layer2_out[225];
    assign layer3_out[647] = layer2_out[150];
    assign layer3_out[648] = layer2_out[213];
    assign layer3_out[649] = ~layer2_out[130];
    assign layer3_out[650] = ~(layer2_out[406] ^ layer2_out[407]);
    assign layer3_out[651] = layer2_out[435];
    assign layer3_out[652] = layer2_out[187];
    assign layer3_out[653] = layer2_out[259] ^ layer2_out[260];
    assign layer3_out[654] = layer2_out[439];
    assign layer3_out[655] = ~layer2_out[8];
    assign layer3_out[656] = layer2_out[269];
    assign layer3_out[657] = ~(layer2_out[630] | layer2_out[631]);
    assign layer3_out[658] = ~layer2_out[469];
    assign layer3_out[659] = layer2_out[176];
    assign layer3_out[660] = ~layer2_out[33];
    assign layer3_out[661] = layer2_out[254];
    assign layer3_out[662] = layer2_out[191] & ~layer2_out[192];
    assign layer3_out[663] = ~layer2_out[241];
    assign layer3_out[664] = layer2_out[10] ^ layer2_out[11];
    assign layer3_out[665] = layer2_out[562];
    assign layer3_out[666] = ~layer2_out[341];
    assign layer3_out[667] = ~layer2_out[759];
    assign layer3_out[668] = layer2_out[266] & ~layer2_out[265];
    assign layer3_out[669] = ~layer2_out[261];
    assign layer3_out[670] = ~layer2_out[113] | layer2_out[114];
    assign layer3_out[671] = layer2_out[342];
    assign layer3_out[672] = layer2_out[743] & ~layer2_out[742];
    assign layer3_out[673] = ~layer2_out[617];
    assign layer3_out[674] = layer2_out[547];
    assign layer3_out[675] = layer2_out[563] ^ layer2_out[564];
    assign layer3_out[676] = layer2_out[193];
    assign layer3_out[677] = layer2_out[483];
    assign layer3_out[678] = ~layer2_out[430];
    assign layer3_out[679] = ~layer2_out[757];
    assign layer3_out[680] = layer2_out[732] & layer2_out[733];
    assign layer3_out[681] = layer2_out[119] & layer2_out[120];
    assign layer3_out[682] = layer2_out[593];
    assign layer3_out[683] = layer2_out[240] & ~layer2_out[239];
    assign layer3_out[684] = ~(layer2_out[222] | layer2_out[223]);
    assign layer3_out[685] = ~layer2_out[372];
    assign layer3_out[686] = ~(layer2_out[140] ^ layer2_out[141]);
    assign layer3_out[687] = layer2_out[525] ^ layer2_out[526];
    assign layer3_out[688] = ~(layer2_out[3] | layer2_out[4]);
    assign layer3_out[689] = ~layer2_out[365];
    assign layer3_out[690] = layer2_out[591] | layer2_out[592];
    assign layer3_out[691] = layer2_out[336];
    assign layer3_out[692] = ~layer2_out[610];
    assign layer3_out[693] = layer2_out[77] ^ layer2_out[78];
    assign layer3_out[694] = ~layer2_out[577];
    assign layer3_out[695] = ~layer2_out[277];
    assign layer3_out[696] = layer2_out[34];
    assign layer3_out[697] = ~layer2_out[226];
    assign layer3_out[698] = ~layer2_out[748];
    assign layer3_out[699] = ~layer2_out[460];
    assign layer3_out[700] = ~layer2_out[595] | layer2_out[594];
    assign layer3_out[701] = ~(layer2_out[687] ^ layer2_out[688]);
    assign layer3_out[702] = ~layer2_out[131];
    assign layer3_out[703] = layer2_out[27];
    assign layer3_out[704] = ~layer2_out[550];
    assign layer3_out[705] = ~layer2_out[188] | layer2_out[189];
    assign layer3_out[706] = layer2_out[395];
    assign layer3_out[707] = layer2_out[197];
    assign layer3_out[708] = layer2_out[306] & ~layer2_out[305];
    assign layer3_out[709] = layer2_out[214] ^ layer2_out[215];
    assign layer3_out[710] = layer2_out[286];
    assign layer3_out[711] = ~layer2_out[617];
    assign layer3_out[712] = layer2_out[624];
    assign layer3_out[713] = ~(layer2_out[361] & layer2_out[362]);
    assign layer3_out[714] = ~layer2_out[455];
    assign layer3_out[715] = layer2_out[451];
    assign layer3_out[716] = layer2_out[90] & ~layer2_out[91];
    assign layer3_out[717] = ~layer2_out[177];
    assign layer3_out[718] = ~layer2_out[748];
    assign layer3_out[719] = ~layer2_out[752];
    assign layer3_out[720] = layer2_out[207] & ~layer2_out[208];
    assign layer3_out[721] = layer2_out[67];
    assign layer3_out[722] = ~(layer2_out[634] | layer2_out[635]);
    assign layer3_out[723] = ~layer2_out[218];
    assign layer3_out[724] = ~layer2_out[523] | layer2_out[522];
    assign layer3_out[725] = layer2_out[322] & ~layer2_out[321];
    assign layer3_out[726] = ~layer2_out[701];
    assign layer3_out[727] = ~layer2_out[303];
    assign layer3_out[728] = layer2_out[707] & ~layer2_out[706];
    assign layer3_out[729] = ~(layer2_out[203] ^ layer2_out[204]);
    assign layer3_out[730] = ~(layer2_out[482] | layer2_out[483]);
    assign layer3_out[731] = ~layer2_out[220];
    assign layer3_out[732] = ~layer2_out[346];
    assign layer3_out[733] = ~(layer2_out[63] ^ layer2_out[64]);
    assign layer3_out[734] = layer2_out[39] & layer2_out[40];
    assign layer3_out[735] = layer2_out[633] & ~layer2_out[634];
    assign layer3_out[736] = layer2_out[339] & ~layer2_out[338];
    assign layer3_out[737] = ~layer2_out[662];
    assign layer3_out[738] = ~(layer2_out[520] | layer2_out[521]);
    assign layer3_out[739] = layer2_out[197];
    assign layer3_out[740] = layer2_out[719];
    assign layer3_out[741] = ~layer2_out[626];
    assign layer3_out[742] = ~layer2_out[596];
    assign layer3_out[743] = layer2_out[296] & ~layer2_out[297];
    assign layer3_out[744] = ~(layer2_out[107] | layer2_out[108]);
    assign layer3_out[745] = layer2_out[477] & ~layer2_out[476];
    assign layer3_out[746] = ~layer2_out[44] | layer2_out[45];
    assign layer3_out[747] = layer2_out[586] & ~layer2_out[587];
    assign layer3_out[748] = ~(layer2_out[255] ^ layer2_out[256]);
    assign layer3_out[749] = layer2_out[16];
    assign layer3_out[750] = ~(layer2_out[500] ^ layer2_out[501]);
    assign layer3_out[751] = ~(layer2_out[162] ^ layer2_out[163]);
    assign layer3_out[752] = layer2_out[681];
    assign layer3_out[753] = layer2_out[180];
    assign layer3_out[754] = layer2_out[88];
    assign layer3_out[755] = ~layer2_out[423] | layer2_out[424];
    assign layer3_out[756] = layer2_out[478];
    assign layer3_out[757] = ~layer2_out[724] | layer2_out[725];
    assign layer3_out[758] = layer2_out[183];
    assign layer3_out[759] = ~layer2_out[682];
    assign layer3_out[760] = ~layer2_out[158];
    assign layer3_out[761] = layer2_out[88];
    assign layer3_out[762] = layer2_out[762];
    assign layer3_out[763] = layer2_out[354];
    assign layer3_out[764] = layer2_out[536];
    assign layer3_out[765] = layer2_out[175];
    assign layer3_out[766] = ~layer2_out[430];
    assign layer3_out[767] = ~layer2_out[515];
    assign layer3_out[768] = layer2_out[598] & layer2_out[599];
    assign layer3_out[769] = layer2_out[781] & ~layer2_out[780];
    assign layer3_out[770] = ~layer2_out[716];
    assign layer3_out[771] = ~layer2_out[479];
    assign layer3_out[772] = layer2_out[733] & layer2_out[734];
    assign layer3_out[773] = layer2_out[307];
    assign layer3_out[774] = layer2_out[144];
    assign layer3_out[775] = ~layer2_out[651];
    assign layer3_out[776] = layer2_out[672] & ~layer2_out[671];
    assign layer3_out[777] = layer2_out[658] & ~layer2_out[657];
    assign layer3_out[778] = layer2_out[376] & ~layer2_out[377];
    assign layer3_out[779] = ~layer2_out[404];
    assign layer3_out[780] = layer2_out[464] & ~layer2_out[463];
    assign layer3_out[781] = layer2_out[210] & layer2_out[211];
    assign layer3_out[782] = layer2_out[674];
    assign layer3_out[783] = layer2_out[625];
    assign layer3_out[784] = layer2_out[17] & layer2_out[18];
    assign layer3_out[785] = ~(layer2_out[29] | layer2_out[30]);
    assign layer3_out[786] = ~layer2_out[493];
    assign layer3_out[787] = ~layer2_out[107];
    assign layer3_out[788] = layer2_out[467];
    assign layer3_out[789] = layer2_out[719];
    assign layer3_out[790] = layer2_out[508];
    assign layer3_out[791] = layer2_out[511];
    assign layer3_out[792] = layer2_out[681] & ~layer2_out[682];
    assign layer3_out[793] = ~layer2_out[744];
    assign layer3_out[794] = layer2_out[627] & ~layer2_out[628];
    assign layer3_out[795] = ~layer2_out[42];
    assign layer3_out[796] = layer2_out[539] & layer2_out[540];
    assign layer3_out[797] = layer2_out[529] | layer2_out[530];
    assign layer3_out[798] = layer2_out[363];
    assign layer3_out[799] = layer2_out[327];
      wire [799:0] last_layer_output;
      assign last_layer_output = layer3_out;
      wire [6:0] result [9:0];

      assign result[0] = last_layer_output[0] + last_layer_output[1] + last_layer_output[2] + last_layer_output[3] + last_layer_output[4] + last_layer_output[5] + last_layer_output[6] + last_layer_output[7] + last_layer_output[8] + last_layer_output[9] + last_layer_output[10] + last_layer_output[11] + last_layer_output[12] + last_layer_output[13] + last_layer_output[14] + last_layer_output[15] + last_layer_output[16] + last_layer_output[17] + last_layer_output[18] + last_layer_output[19] + last_layer_output[20] + last_layer_output[21] + last_layer_output[22] + last_layer_output[23] + last_layer_output[24] + last_layer_output[25] + last_layer_output[26] + last_layer_output[27] + last_layer_output[28] + last_layer_output[29] + last_layer_output[30] + last_layer_output[31] + last_layer_output[32] + last_layer_output[33] + last_layer_output[34] + last_layer_output[35] + last_layer_output[36] + last_layer_output[37] + last_layer_output[38] + last_layer_output[39] + last_layer_output[40] + last_layer_output[41] + last_layer_output[42] + last_layer_output[43] + last_layer_output[44] + last_layer_output[45] + last_layer_output[46] + last_layer_output[47] + last_layer_output[48] + last_layer_output[49] + last_layer_output[50] + last_layer_output[51] + last_layer_output[52] + last_layer_output[53] + last_layer_output[54] + last_layer_output[55] + last_layer_output[56] + last_layer_output[57] + last_layer_output[58] + last_layer_output[59] + last_layer_output[60] + last_layer_output[61] + last_layer_output[62] + last_layer_output[63] + last_layer_output[64] + last_layer_output[65] + last_layer_output[66] + last_layer_output[67] + last_layer_output[68] + last_layer_output[69] + last_layer_output[70] + last_layer_output[71] + last_layer_output[72] + last_layer_output[73] + last_layer_output[74] + last_layer_output[75] + last_layer_output[76] + last_layer_output[77] + last_layer_output[78] + last_layer_output[79];
      assign result[1] = last_layer_output[80] + last_layer_output[81] + last_layer_output[82] + last_layer_output[83] + last_layer_output[84] + last_layer_output[85] + last_layer_output[86] + last_layer_output[87] + last_layer_output[88] + last_layer_output[89] + last_layer_output[90] + last_layer_output[91] + last_layer_output[92] + last_layer_output[93] + last_layer_output[94] + last_layer_output[95] + last_layer_output[96] + last_layer_output[97] + last_layer_output[98] + last_layer_output[99] + last_layer_output[100] + last_layer_output[101] + last_layer_output[102] + last_layer_output[103] + last_layer_output[104] + last_layer_output[105] + last_layer_output[106] + last_layer_output[107] + last_layer_output[108] + last_layer_output[109] + last_layer_output[110] + last_layer_output[111] + last_layer_output[112] + last_layer_output[113] + last_layer_output[114] + last_layer_output[115] + last_layer_output[116] + last_layer_output[117] + last_layer_output[118] + last_layer_output[119] + last_layer_output[120] + last_layer_output[121] + last_layer_output[122] + last_layer_output[123] + last_layer_output[124] + last_layer_output[125] + last_layer_output[126] + last_layer_output[127] + last_layer_output[128] + last_layer_output[129] + last_layer_output[130] + last_layer_output[131] + last_layer_output[132] + last_layer_output[133] + last_layer_output[134] + last_layer_output[135] + last_layer_output[136] + last_layer_output[137] + last_layer_output[138] + last_layer_output[139] + last_layer_output[140] + last_layer_output[141] + last_layer_output[142] + last_layer_output[143] + last_layer_output[144] + last_layer_output[145] + last_layer_output[146] + last_layer_output[147] + last_layer_output[148] + last_layer_output[149] + last_layer_output[150] + last_layer_output[151] + last_layer_output[152] + last_layer_output[153] + last_layer_output[154] + last_layer_output[155] + last_layer_output[156] + last_layer_output[157] + last_layer_output[158] + last_layer_output[159];
      assign result[2] = last_layer_output[160] + last_layer_output[161] + last_layer_output[162] + last_layer_output[163] + last_layer_output[164] + last_layer_output[165] + last_layer_output[166] + last_layer_output[167] + last_layer_output[168] + last_layer_output[169] + last_layer_output[170] + last_layer_output[171] + last_layer_output[172] + last_layer_output[173] + last_layer_output[174] + last_layer_output[175] + last_layer_output[176] + last_layer_output[177] + last_layer_output[178] + last_layer_output[179] + last_layer_output[180] + last_layer_output[181] + last_layer_output[182] + last_layer_output[183] + last_layer_output[184] + last_layer_output[185] + last_layer_output[186] + last_layer_output[187] + last_layer_output[188] + last_layer_output[189] + last_layer_output[190] + last_layer_output[191] + last_layer_output[192] + last_layer_output[193] + last_layer_output[194] + last_layer_output[195] + last_layer_output[196] + last_layer_output[197] + last_layer_output[198] + last_layer_output[199] + last_layer_output[200] + last_layer_output[201] + last_layer_output[202] + last_layer_output[203] + last_layer_output[204] + last_layer_output[205] + last_layer_output[206] + last_layer_output[207] + last_layer_output[208] + last_layer_output[209] + last_layer_output[210] + last_layer_output[211] + last_layer_output[212] + last_layer_output[213] + last_layer_output[214] + last_layer_output[215] + last_layer_output[216] + last_layer_output[217] + last_layer_output[218] + last_layer_output[219] + last_layer_output[220] + last_layer_output[221] + last_layer_output[222] + last_layer_output[223] + last_layer_output[224] + last_layer_output[225] + last_layer_output[226] + last_layer_output[227] + last_layer_output[228] + last_layer_output[229] + last_layer_output[230] + last_layer_output[231] + last_layer_output[232] + last_layer_output[233] + last_layer_output[234] + last_layer_output[235] + last_layer_output[236] + last_layer_output[237] + last_layer_output[238] + last_layer_output[239];
      assign result[3] = last_layer_output[240] + last_layer_output[241] + last_layer_output[242] + last_layer_output[243] + last_layer_output[244] + last_layer_output[245] + last_layer_output[246] + last_layer_output[247] + last_layer_output[248] + last_layer_output[249] + last_layer_output[250] + last_layer_output[251] + last_layer_output[252] + last_layer_output[253] + last_layer_output[254] + last_layer_output[255] + last_layer_output[256] + last_layer_output[257] + last_layer_output[258] + last_layer_output[259] + last_layer_output[260] + last_layer_output[261] + last_layer_output[262] + last_layer_output[263] + last_layer_output[264] + last_layer_output[265] + last_layer_output[266] + last_layer_output[267] + last_layer_output[268] + last_layer_output[269] + last_layer_output[270] + last_layer_output[271] + last_layer_output[272] + last_layer_output[273] + last_layer_output[274] + last_layer_output[275] + last_layer_output[276] + last_layer_output[277] + last_layer_output[278] + last_layer_output[279] + last_layer_output[280] + last_layer_output[281] + last_layer_output[282] + last_layer_output[283] + last_layer_output[284] + last_layer_output[285] + last_layer_output[286] + last_layer_output[287] + last_layer_output[288] + last_layer_output[289] + last_layer_output[290] + last_layer_output[291] + last_layer_output[292] + last_layer_output[293] + last_layer_output[294] + last_layer_output[295] + last_layer_output[296] + last_layer_output[297] + last_layer_output[298] + last_layer_output[299] + last_layer_output[300] + last_layer_output[301] + last_layer_output[302] + last_layer_output[303] + last_layer_output[304] + last_layer_output[305] + last_layer_output[306] + last_layer_output[307] + last_layer_output[308] + last_layer_output[309] + last_layer_output[310] + last_layer_output[311] + last_layer_output[312] + last_layer_output[313] + last_layer_output[314] + last_layer_output[315] + last_layer_output[316] + last_layer_output[317] + last_layer_output[318] + last_layer_output[319];
      assign result[4] = last_layer_output[320] + last_layer_output[321] + last_layer_output[322] + last_layer_output[323] + last_layer_output[324] + last_layer_output[325] + last_layer_output[326] + last_layer_output[327] + last_layer_output[328] + last_layer_output[329] + last_layer_output[330] + last_layer_output[331] + last_layer_output[332] + last_layer_output[333] + last_layer_output[334] + last_layer_output[335] + last_layer_output[336] + last_layer_output[337] + last_layer_output[338] + last_layer_output[339] + last_layer_output[340] + last_layer_output[341] + last_layer_output[342] + last_layer_output[343] + last_layer_output[344] + last_layer_output[345] + last_layer_output[346] + last_layer_output[347] + last_layer_output[348] + last_layer_output[349] + last_layer_output[350] + last_layer_output[351] + last_layer_output[352] + last_layer_output[353] + last_layer_output[354] + last_layer_output[355] + last_layer_output[356] + last_layer_output[357] + last_layer_output[358] + last_layer_output[359] + last_layer_output[360] + last_layer_output[361] + last_layer_output[362] + last_layer_output[363] + last_layer_output[364] + last_layer_output[365] + last_layer_output[366] + last_layer_output[367] + last_layer_output[368] + last_layer_output[369] + last_layer_output[370] + last_layer_output[371] + last_layer_output[372] + last_layer_output[373] + last_layer_output[374] + last_layer_output[375] + last_layer_output[376] + last_layer_output[377] + last_layer_output[378] + last_layer_output[379] + last_layer_output[380] + last_layer_output[381] + last_layer_output[382] + last_layer_output[383] + last_layer_output[384] + last_layer_output[385] + last_layer_output[386] + last_layer_output[387] + last_layer_output[388] + last_layer_output[389] + last_layer_output[390] + last_layer_output[391] + last_layer_output[392] + last_layer_output[393] + last_layer_output[394] + last_layer_output[395] + last_layer_output[396] + last_layer_output[397] + last_layer_output[398] + last_layer_output[399];
      assign result[5] = last_layer_output[400] + last_layer_output[401] + last_layer_output[402] + last_layer_output[403] + last_layer_output[404] + last_layer_output[405] + last_layer_output[406] + last_layer_output[407] + last_layer_output[408] + last_layer_output[409] + last_layer_output[410] + last_layer_output[411] + last_layer_output[412] + last_layer_output[413] + last_layer_output[414] + last_layer_output[415] + last_layer_output[416] + last_layer_output[417] + last_layer_output[418] + last_layer_output[419] + last_layer_output[420] + last_layer_output[421] + last_layer_output[422] + last_layer_output[423] + last_layer_output[424] + last_layer_output[425] + last_layer_output[426] + last_layer_output[427] + last_layer_output[428] + last_layer_output[429] + last_layer_output[430] + last_layer_output[431] + last_layer_output[432] + last_layer_output[433] + last_layer_output[434] + last_layer_output[435] + last_layer_output[436] + last_layer_output[437] + last_layer_output[438] + last_layer_output[439] + last_layer_output[440] + last_layer_output[441] + last_layer_output[442] + last_layer_output[443] + last_layer_output[444] + last_layer_output[445] + last_layer_output[446] + last_layer_output[447] + last_layer_output[448] + last_layer_output[449] + last_layer_output[450] + last_layer_output[451] + last_layer_output[452] + last_layer_output[453] + last_layer_output[454] + last_layer_output[455] + last_layer_output[456] + last_layer_output[457] + last_layer_output[458] + last_layer_output[459] + last_layer_output[460] + last_layer_output[461] + last_layer_output[462] + last_layer_output[463] + last_layer_output[464] + last_layer_output[465] + last_layer_output[466] + last_layer_output[467] + last_layer_output[468] + last_layer_output[469] + last_layer_output[470] + last_layer_output[471] + last_layer_output[472] + last_layer_output[473] + last_layer_output[474] + last_layer_output[475] + last_layer_output[476] + last_layer_output[477] + last_layer_output[478] + last_layer_output[479];
      assign result[6] = last_layer_output[480] + last_layer_output[481] + last_layer_output[482] + last_layer_output[483] + last_layer_output[484] + last_layer_output[485] + last_layer_output[486] + last_layer_output[487] + last_layer_output[488] + last_layer_output[489] + last_layer_output[490] + last_layer_output[491] + last_layer_output[492] + last_layer_output[493] + last_layer_output[494] + last_layer_output[495] + last_layer_output[496] + last_layer_output[497] + last_layer_output[498] + last_layer_output[499] + last_layer_output[500] + last_layer_output[501] + last_layer_output[502] + last_layer_output[503] + last_layer_output[504] + last_layer_output[505] + last_layer_output[506] + last_layer_output[507] + last_layer_output[508] + last_layer_output[509] + last_layer_output[510] + last_layer_output[511] + last_layer_output[512] + last_layer_output[513] + last_layer_output[514] + last_layer_output[515] + last_layer_output[516] + last_layer_output[517] + last_layer_output[518] + last_layer_output[519] + last_layer_output[520] + last_layer_output[521] + last_layer_output[522] + last_layer_output[523] + last_layer_output[524] + last_layer_output[525] + last_layer_output[526] + last_layer_output[527] + last_layer_output[528] + last_layer_output[529] + last_layer_output[530] + last_layer_output[531] + last_layer_output[532] + last_layer_output[533] + last_layer_output[534] + last_layer_output[535] + last_layer_output[536] + last_layer_output[537] + last_layer_output[538] + last_layer_output[539] + last_layer_output[540] + last_layer_output[541] + last_layer_output[542] + last_layer_output[543] + last_layer_output[544] + last_layer_output[545] + last_layer_output[546] + last_layer_output[547] + last_layer_output[548] + last_layer_output[549] + last_layer_output[550] + last_layer_output[551] + last_layer_output[552] + last_layer_output[553] + last_layer_output[554] + last_layer_output[555] + last_layer_output[556] + last_layer_output[557] + last_layer_output[558] + last_layer_output[559];
      assign result[7] = last_layer_output[560] + last_layer_output[561] + last_layer_output[562] + last_layer_output[563] + last_layer_output[564] + last_layer_output[565] + last_layer_output[566] + last_layer_output[567] + last_layer_output[568] + last_layer_output[569] + last_layer_output[570] + last_layer_output[571] + last_layer_output[572] + last_layer_output[573] + last_layer_output[574] + last_layer_output[575] + last_layer_output[576] + last_layer_output[577] + last_layer_output[578] + last_layer_output[579] + last_layer_output[580] + last_layer_output[581] + last_layer_output[582] + last_layer_output[583] + last_layer_output[584] + last_layer_output[585] + last_layer_output[586] + last_layer_output[587] + last_layer_output[588] + last_layer_output[589] + last_layer_output[590] + last_layer_output[591] + last_layer_output[592] + last_layer_output[593] + last_layer_output[594] + last_layer_output[595] + last_layer_output[596] + last_layer_output[597] + last_layer_output[598] + last_layer_output[599] + last_layer_output[600] + last_layer_output[601] + last_layer_output[602] + last_layer_output[603] + last_layer_output[604] + last_layer_output[605] + last_layer_output[606] + last_layer_output[607] + last_layer_output[608] + last_layer_output[609] + last_layer_output[610] + last_layer_output[611] + last_layer_output[612] + last_layer_output[613] + last_layer_output[614] + last_layer_output[615] + last_layer_output[616] + last_layer_output[617] + last_layer_output[618] + last_layer_output[619] + last_layer_output[620] + last_layer_output[621] + last_layer_output[622] + last_layer_output[623] + last_layer_output[624] + last_layer_output[625] + last_layer_output[626] + last_layer_output[627] + last_layer_output[628] + last_layer_output[629] + last_layer_output[630] + last_layer_output[631] + last_layer_output[632] + last_layer_output[633] + last_layer_output[634] + last_layer_output[635] + last_layer_output[636] + last_layer_output[637] + last_layer_output[638] + last_layer_output[639];
      assign result[8] = last_layer_output[640] + last_layer_output[641] + last_layer_output[642] + last_layer_output[643] + last_layer_output[644] + last_layer_output[645] + last_layer_output[646] + last_layer_output[647] + last_layer_output[648] + last_layer_output[649] + last_layer_output[650] + last_layer_output[651] + last_layer_output[652] + last_layer_output[653] + last_layer_output[654] + last_layer_output[655] + last_layer_output[656] + last_layer_output[657] + last_layer_output[658] + last_layer_output[659] + last_layer_output[660] + last_layer_output[661] + last_layer_output[662] + last_layer_output[663] + last_layer_output[664] + last_layer_output[665] + last_layer_output[666] + last_layer_output[667] + last_layer_output[668] + last_layer_output[669] + last_layer_output[670] + last_layer_output[671] + last_layer_output[672] + last_layer_output[673] + last_layer_output[674] + last_layer_output[675] + last_layer_output[676] + last_layer_output[677] + last_layer_output[678] + last_layer_output[679] + last_layer_output[680] + last_layer_output[681] + last_layer_output[682] + last_layer_output[683] + last_layer_output[684] + last_layer_output[685] + last_layer_output[686] + last_layer_output[687] + last_layer_output[688] + last_layer_output[689] + last_layer_output[690] + last_layer_output[691] + last_layer_output[692] + last_layer_output[693] + last_layer_output[694] + last_layer_output[695] + last_layer_output[696] + last_layer_output[697] + last_layer_output[698] + last_layer_output[699] + last_layer_output[700] + last_layer_output[701] + last_layer_output[702] + last_layer_output[703] + last_layer_output[704] + last_layer_output[705] + last_layer_output[706] + last_layer_output[707] + last_layer_output[708] + last_layer_output[709] + last_layer_output[710] + last_layer_output[711] + last_layer_output[712] + last_layer_output[713] + last_layer_output[714] + last_layer_output[715] + last_layer_output[716] + last_layer_output[717] + last_layer_output[718] + last_layer_output[719];
      assign result[9] = last_layer_output[720] + last_layer_output[721] + last_layer_output[722] + last_layer_output[723] + last_layer_output[724] + last_layer_output[725] + last_layer_output[726] + last_layer_output[727] + last_layer_output[728] + last_layer_output[729] + last_layer_output[730] + last_layer_output[731] + last_layer_output[732] + last_layer_output[733] + last_layer_output[734] + last_layer_output[735] + last_layer_output[736] + last_layer_output[737] + last_layer_output[738] + last_layer_output[739] + last_layer_output[740] + last_layer_output[741] + last_layer_output[742] + last_layer_output[743] + last_layer_output[744] + last_layer_output[745] + last_layer_output[746] + last_layer_output[747] + last_layer_output[748] + last_layer_output[749] + last_layer_output[750] + last_layer_output[751] + last_layer_output[752] + last_layer_output[753] + last_layer_output[754] + last_layer_output[755] + last_layer_output[756] + last_layer_output[757] + last_layer_output[758] + last_layer_output[759] + last_layer_output[760] + last_layer_output[761] + last_layer_output[762] + last_layer_output[763] + last_layer_output[764] + last_layer_output[765] + last_layer_output[766] + last_layer_output[767] + last_layer_output[768] + last_layer_output[769] + last_layer_output[770] + last_layer_output[771] + last_layer_output[772] + last_layer_output[773] + last_layer_output[774] + last_layer_output[775] + last_layer_output[776] + last_layer_output[777] + last_layer_output[778] + last_layer_output[779] + last_layer_output[780] + last_layer_output[781] + last_layer_output[782] + last_layer_output[783] + last_layer_output[784] + last_layer_output[785] + last_layer_output[786] + last_layer_output[787] + last_layer_output[788] + last_layer_output[789] + last_layer_output[790] + last_layer_output[791] + last_layer_output[792] + last_layer_output[793] + last_layer_output[794] + last_layer_output[795] + last_layer_output[796] + last_layer_output[797] + last_layer_output[798] + last_layer_output[799];
      assign y[69:63]=result[0];
      assign y[62:56]=result[1];
      assign y[55:49]=result[2];
      assign y[48:42]=result[3];
      assign y[41:35]=result[4];
      assign y[34:28]=result[5];
      assign y[27:21]=result[6];
      assign y[20:14]=result[7];
      assign y[13:7]=result[8];
      assign y[6:0]=result[9];
endmodule
